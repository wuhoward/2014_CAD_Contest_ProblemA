module top (out,n3,n21,n26,n28,n29,n31,n35,n38,n44
        ,n62,n76,n77,n78,n79,n80,n81,n82,n83,n87
        ,n88,n89,n93,n95,n97,n134,n136,n137,n138,n149
        ,n150,n151,n152,n164,n165,n166,n167,n180,n181,n182
        ,n183,n189,n191,n192,n195,n197,n200,n202,n203,n204
        ,n284,n390,n393,n395,n549,n551,n552,n555,n558,n559
        ,n560,n561,n564,n566,n570,n581,n582,n599,n602,n604
        ,n605,n607,n611,n617,n620,n622,n624,n628,n631,n633
        ,n635,n639,n642,n644,n646,n648,n656,n659,n661,n663
        ,n667,n670,n672,n674,n678,n681,n683,n685,n689,n692
        ,n694,n696,n704,n707,n709,n711,n715,n718,n720,n722
        ,n726,n729,n731,n733,n737,n740,n742,n744,n752,n755
        ,n757,n759,n776,n779,n781,n783,n792,n795,n797,n799
        ,n808,n811,n813,n815,n824,n827,n829,n831,n840,n843
        ,n845,n847,n855,n858,n860,n862,n935,n938,n940,n942
        ,n946,n949,n951,n953,n957,n960,n962,n964,n968,n971
        ,n973,n975,n984,n987,n989,n991,n995,n998,n1000,n1002
        ,n1006,n1009,n1011,n1013,n1017,n1020,n1022,n1024,n1032,n1035
        ,n1037,n1039,n1043,n1046,n1048,n1050,n1054,n1057,n1059,n1061
        ,n1065,n1068,n1070,n1072,n1248,n1251,n1253,n1255,n1264,n1267
        ,n1269,n1271,n1280,n1283,n1285,n1287,n1296,n1299,n1301,n1303
        ,n1312,n1315,n1317,n1319,n1328,n1331,n1333,n1335,n1344,n1347
        ,n1349,n1351,n1359,n1362,n1364,n1366,n1689,n1692,n1694,n1696
        ,n1705,n1708,n1710,n1712,n1724,n1727,n1729,n1731,n1750,n1753
        ,n1755,n1757,n1766,n1769,n1771,n1773,n1787,n1790,n1792,n1794
        ,n1817,n1820,n1822,n1824,n1840,n1843,n1845,n1847,n2084,n2087
        ,n2089,n2091,n2100,n2103,n2105,n2107,n2116,n2119,n2121,n2123
        ,n2132,n2135,n2137,n2139,n2148,n2151,n2153,n2155,n2164,n2167
        ,n2169,n2171,n2181,n2184,n2186,n2188,n2196,n2199,n2201,n2203
        ,n2711,n2713,n2715,n2717,n2723,n2725,n2727,n2729,n2735,n2737
        ,n2739,n2741,n2747,n2749,n2890,n2901,n2928,n2954,n2962,n2971
        ,n2982,n2985,n2988,n2991,n2996,n2999,n3002,n3005,n3010,n3013
        ,n3023,n3024,n3038,n3039,n3057,n3058,n3061,n3062,n3065,n3066
        ,n3069,n3070,n3075,n3076,n3079,n3080,n3083,n3084,n3087,n3088
        ,n3093,n3094,n3097,n3098,n3101,n3102,n3105,n3106,n3111,n3112
        ,n3115,n3116,n3126,n3127,n3141,n3142,n3160,n3161,n3164,n3165
        ,n3168,n3169,n3172,n3173,n3178,n3179,n3182,n3183,n3186,n3187
        ,n3190,n3191,n3196,n3197,n3200,n3201,n3204,n3205,n3208,n3209
        ,n3214,n3215,n3218,n3219,n3229,n3230,n3244,n3245,n3263,n3264
        ,n3267,n3268,n3271,n3272,n3275,n3276,n3281,n3282,n3285,n3286
        ,n3289,n3290,n3293,n3294,n3299,n3300,n3303,n3304,n3307,n3308
        ,n3311,n3312,n3317,n3318,n3321,n3322,n3332,n3333,n3347,n3348
        ,n3366,n3367,n3370,n3371,n3374,n3375,n3378,n3379,n3384,n3385
        ,n3388,n3389,n3392,n3393,n3396,n3397,n3402,n3403,n3406,n3407
        ,n3410,n3411,n3414,n3415,n3420,n3421,n3424,n3425,n3435,n3436
        ,n3450,n3451,n3469,n3470,n3473,n3474,n3477,n3478,n3481,n3482
        ,n3487,n3488,n3491,n3492,n3495,n3496,n3499,n3500,n3505,n3506
        ,n3509,n3510,n3513,n3514,n3517,n3518,n3523,n3524,n3527,n3528
        ,n3538,n3539,n3553,n3554,n3572,n3573,n3576,n3577,n3580,n3581
        ,n3584,n3585,n3590,n3591,n3594,n3595,n3598,n3599,n3602,n3603
        ,n3608,n3609,n3612,n3613,n3616,n3617,n3620,n3621,n3626,n3627
        ,n3630,n3631,n3641,n3642,n3656,n3657,n3674,n3675,n3678,n3679
        ,n3682,n3683,n3686,n3687,n3692,n3693,n3696,n3697,n3700,n3701
        ,n3704,n3705,n3710,n3711,n3714,n3715,n3718,n3719,n3722,n3723
        ,n3728,n3729,n3732,n3733,n3743,n3744,n3758,n3759,n3800,n3801
        ,n3820,n3821,n3835,n3836,n3863,n3864,n3883,n3884,n3898,n3899
        ,n3926,n3927,n3946,n3947,n3961,n3962,n3989,n3990,n4009,n4010
        ,n4024,n4025,n4052,n4053,n4072,n4073,n4087,n4088,n4115,n4116
        ,n4135,n4136,n4150,n4151,n4178,n4179,n4198,n4199,n4213,n4214
        ,n4240,n4241,n4260,n4261,n4275,n4276,n4393,n4394,n4408,n4409
        ,n4418,n4419,n4436,n4437,n4451,n4452,n4461,n4462,n4479,n4480
        ,n4494,n4495,n4504,n4505,n4522,n4523,n4537,n4538,n4547,n4548
        ,n4565,n4566,n4580,n4581,n4590,n4591,n4608,n4609,n4623,n4624
        ,n4633,n4634,n4651,n4652,n4666,n4667,n4676,n4677,n4693,n4694
        ,n4708,n4709,n4718,n4719,n4965,n4975,n4979,n4981,n4986,n4988
        ,n4993,n4995,n5000,n5002,n5012,n5013,n5027,n5032,n5037,n5044
        ,n5047,n5050,n5053,n5058,n5059,n5062,n5065,n5068,n5073,n5076
        ,n5081,n5088,n5089,n5092,n5095,n5098,n5103,n5106,n5109,n5112
        ,n5117,n5118,n5121,n5124,n5127,n5132,n5135,n5138,n5141,n5142
        ,n5152,n5153,n5156,n5159,n5162,n5167,n5170,n5173,n5176,n5181
        ,n5182,n5185,n5188,n5191,n5196,n5199,n5204,n5211,n5212,n5215
        ,n5218,n5221,n5226,n5229,n5232,n5235,n5240,n5241,n5244,n5247
        ,n5250,n5255,n5258,n5261,n5264,n5265,n5275,n5276,n5279,n5282
        ,n5285,n5290,n5293,n5296,n5299,n5304,n5305,n5308,n5311,n5314
        ,n5319,n5322,n5327,n5334,n5335,n5338,n5341,n5344,n5349,n5352
        ,n5355,n5358,n5363,n5364,n5367,n5370,n5373,n5378,n5381,n5384
        ,n5387,n5388,n5398,n5399,n5402,n5405,n5408,n5413,n5416,n5419
        ,n5422,n5427,n5428,n5431,n5434,n5437,n5442,n5445,n5450,n5457
        ,n5458,n5461,n5464,n5467,n5472,n5475,n5478,n5481,n5486,n5487
        ,n5490,n5493,n5496,n5501,n5504,n5507,n5510,n5511,n5521,n5522
        ,n5525,n5528,n5531,n5536,n5539,n5542,n5545,n5550,n5551,n5554
        ,n5557,n5560,n5565,n5568,n5573,n5580,n5581,n5584,n5587,n5590
        ,n5595,n5598,n5601,n5604,n5609,n5610,n5613,n5616,n5619,n5624
        ,n5627,n5630,n5633,n5634,n5644,n5645,n5648,n5651,n5654,n5659
        ,n5662,n5665,n5668,n5673,n5674,n5677,n5680,n5683,n5688,n5691
        ,n5696,n5703,n5704,n5707,n5710,n5713,n5718,n5721,n5724,n5727
        ,n5732,n5733,n5736,n5739,n5742,n5747,n5750,n5753,n5756,n5757
        ,n5767,n5768,n5771,n5774,n5777,n5782,n5785,n5788,n5791,n5796
        ,n5797,n5800,n5803,n5806,n5811,n5814,n5819,n5826,n5827,n5830
        ,n5833,n5836,n5841,n5844,n5847,n5850,n5855,n5856,n5859,n5862
        ,n5865,n5870,n5873,n5876,n5879,n5880,n5889,n5890,n5893,n5896
        ,n5899,n5904,n5907,n5910,n5913,n5918,n5919,n5922,n5925,n5928
        ,n5933,n5936,n5941,n5948,n5949,n5952,n5955,n5958,n5963,n5966
        ,n5969,n5972,n5977,n5978,n5981,n5984,n5987,n5992,n5995,n5998
        ,n6001,n6002,n6020,n6022,n6026,n6028,n6033,n6035,n6081,n6124
        ,n6170,n6213,n6259,n6302,n6348,n6391,n6437,n6480,n6526,n6569
        ,n6615,n6658,n6703,n6746,n6760,n6762,n6766,n6768,n6773,n6775
        ,n6780,n6782,n6787,n6789,n6801,n6802,n6805,n6808,n6811,n6816
        ,n6819,n6824,n6831,n6832,n6835,n6838,n6841,n6846,n6849,n6852
        ,n6855,n6858,n6870,n6871,n6874,n6877,n6880,n6885,n6888,n6893
        ,n6900,n6901,n6904,n6907,n6910,n6915,n6918,n6921,n6924,n6927
        ,n6939,n6940,n6943,n6946,n6949,n6954,n6957,n6962,n6969,n6970
        ,n6973,n6976,n6979,n6984,n6987,n6990,n6993,n6996,n7008,n7009
        ,n7012,n7015,n7018,n7023,n7026,n7031,n7038,n7039,n7042,n7045
        ,n7048,n7053,n7056,n7059,n7062,n7065,n7077,n7078,n7081,n7084
        ,n7087,n7092,n7095,n7100,n7107,n7108,n7111,n7114,n7117,n7122
        ,n7125,n7128,n7131,n7134,n7146,n7147,n7150,n7153,n7156,n7161
        ,n7164,n7169,n7176,n7177,n7180,n7183,n7186,n7191,n7194,n7197
        ,n7200,n7203,n7215,n7216,n7219,n7222,n7225,n7230,n7233,n7238
        ,n7245,n7246,n7249,n7252,n7255,n7260,n7263,n7266,n7269,n7272
        ,n7283,n7284,n7287,n7290,n7293,n7298,n7301,n7306,n7313,n7314
        ,n7317,n7320,n7323,n7328,n7331,n7334,n7337,n7340,n7644,n7646
        ,n7653,n7655,n7669,n7671,n7678,n7680,n7685,n7687,n7692,n7694
        ,n7708,n7710,n7717,n7719,n7885,n7888,n7997,n8000,n8109,n8112
        ,n8221,n8224,n8329,n8332,n8437,n8440,n8544,n8547,n9092,n9106
        ,n9120,n9142,n9166,n9189,n9215,n9231,n9405,n9417,n9429,n9441
        ,n9453,n9465,n9477,n9488,n9941,n9944,n10553,n10554,n10568,n10574
        ,n10575,n10589,n10590,n10617,n10618,n10632,n10638,n10639,n10653,n10654
        ,n10681,n10682,n10696,n10702,n10703,n10717,n10718,n10745,n10746,n10760
        ,n10766,n10767,n10781,n10782,n10810,n10811,n10825,n10831,n10832,n10847
        ,n10848,n10877,n10878,n10893,n10899,n10900,n10914,n10915,n10942,n10943
        ,n10957,n10963,n10964,n10978,n10979,n11006,n11007,n11022,n11028,n11029
        ,n11044,n11045,n11163,n11164,n11174,n11180,n11181,n11191,n11192,n11210
        ,n11211,n11221,n11227,n11228,n11238,n11239,n11257,n11258,n11268,n11274
        ,n11275,n11285,n11286,n11304,n11305,n11315,n11321,n11322,n11332,n11333
        ,n11351,n11352,n11362,n11368,n11369,n11378,n11379,n11396,n11397,n11407
        ,n11413,n11414,n11424,n11425,n11443,n11444,n11454,n11460,n11461,n11471
        ,n11472,n11489,n11490,n11500,n11506,n11507,n11517,n11518,n11747,n11751
        ,n11756,n11761,n11766,n11776,n11777,n11780,n11783,n11786,n11791,n11794
        ,n11797,n11800,n11803,n11813,n11814,n11817,n11820,n11823,n11828,n11831
        ,n11834,n11837,n11840,n11850,n11851,n11854,n11857,n11860,n11865,n11868
        ,n11871,n11874,n11877,n11887,n11888,n11891,n11894,n11897,n11902,n11905
        ,n11908,n11911,n11914,n11924,n11925,n11928,n11931,n11934,n11939,n11942
        ,n11945,n11948,n11951,n11961,n11962,n11965,n11968,n11971,n11976,n11979
        ,n11982,n11985,n11988,n11998,n11999,n12002,n12005,n12008,n12013,n12016
        ,n12019,n12022,n12025,n12034,n12035,n12038,n12041,n12044,n12049,n12052
        ,n12055,n12058,n12061,n12124,n12127,n12131,n12134,n12144,n12145,n12148
        ,n12151,n12154,n12159,n12162,n12165,n12168,n12171,n12181,n12182,n12185
        ,n12188,n12191,n12196,n12199,n12202,n12205,n12208,n12218,n12219,n12222
        ,n12225,n12228,n12233,n12236,n12239,n12242,n12245,n12255,n12256,n12259
        ,n12262,n12265,n12270,n12273,n12276,n12279,n12282,n12292,n12293,n12296
        ,n12299,n12302,n12307,n12310,n12313,n12316,n12319,n12329,n12330,n12333
        ,n12336,n12339,n12344,n12347,n12350,n12353,n12356,n12366,n12367,n12370
        ,n12373,n12376,n12381,n12384,n12387,n12390,n12393,n12402,n12403,n12406
        ,n12409,n12412,n12417,n12420,n12423,n12426,n12429,n12455,n12824,n12831
        ,n12874,n12877,n13067,n13070,n13179,n13182,n13291,n13294,n13403,n13406
        ,n13511,n13514,n13619,n13622,n13726,n13729,n13888,n13890,n13892,n13894
        ,n13896,n13899,n13906,n13908,n13909,n13912,n13919,n13922,n13927,n13934
        ,n13954,n13956,n13958,n13960,n13962,n13964,n13966,n13968,n13970,n13972
        ,n13974,n13976,n13978,n13980,n13982,n13984,n13989,n13997,n14002,n14008
        ,n14010,n14012,n14014,n14016,n14018,n14020,n14022,n14024,n14026,n14028
        ,n14030,n14032,n14034,n14036,n14038,n14043,n14045,n14047,n14049,n14051
        ,n14053,n14055,n14057,n14059,n14061,n14063,n14065,n14067,n14069,n14071
        ,n14073,n14077,n14079,n14081,n14083,n14085,n14087,n14089,n14091,n14093
        ,n14095,n14097,n14099,n14101,n14103,n14105,n14107,n14114,n14115,n14121
        ,n14122,n14127,n14128,n14129,n14130,n14146,n14155,n14170,n14175,n14198
        ,n14202,n14204,n14209,n14213,n14214,n14215,n14216,n14219,n14220,n14222
        ,n14223,n14240,n14253,n14285,n14287,n14290,n14292,n14302,n14304,n14307
        ,n14309,n14314,n14320,n14323,n14341,n14351,n14354,n14357,n14360,n14373
        ,n14392,n14411,n14420,n14428,n14436,n14441,n14461,n14463,n14465,n14467
        ,n14471,n14474,n14480,n14486,n14507,n14510,n14524,n14526,n14528,n14530
        ,n14534,n14541,n14547,n14556,n14557,n14562,n14582,n14584,n14586,n14588
        ,n14592,n14595,n14601,n14607,n14618,n14642,n14645,n14648,n14650,n14660
        ,n14662,n14665,n14667,n14676,n14678,n14681,n14683,n14692,n14694,n14697
        ,n14699,n14708,n14710,n14713,n14715,n14725,n14727,n14729,n14731,n14735
        ,n14738,n14744,n14750,n14760,n14767,n14780,n14787,n14789,n14796,n14798
        ,n14800,n14802,n14806,n14813,n14819,n14826,n14828,n14830,n14832,n14836
        ,n14839,n14845,n14851,n14855,n14857,n14859,n14865,n14868,n14870,n14872
        ,n14874,n14876,n14880,n14881,n14891,n14893,n14904,n14909,n14925,n14927
        ,n14929,n14931,n14935,n14938,n14944,n14950,n14961,n14978,n14980,n14982
        ,n14988,n14991,n14993,n14995,n14997,n14999,n15003,n15004,n15017,n15019
        ,n15022,n15024,n15031,n15034,n15036,n15044,n15046,n15049,n15051,n15061
        ,n15063,n15066,n15068,n15077,n15079,n15082,n15084,n15097,n15100,n15107
        ,n15111,n15113,n15117,n15124,n15126,n15128,n15130,n15134,n15137,n15143
        ,n15149,n15156,n15158,n15160,n15162,n15166,n15169,n15175,n15181,n15185
        ,n15188,n15196,n15198,n15200,n15202,n15206,n15213,n15219,n15228,n15233
        ,n15249,n15251,n15253,n15255,n15259,n15262,n15268,n15274,n15285,n15306
        ,n15309,n15312,n15314,n15324,n15326,n15329,n15331,n15340,n15342,n15345
        ,n15347,n15356,n15358,n15361,n15363,n15372,n15374,n15377,n15379,n15388
        ,n15390,n15392,n15394,n15398,n15401,n15407,n15413,n15423,n15430,n15443
        ,n15450,n15452,n15459,n15461,n15463,n15465,n15469,n15476,n15482,n15489
        ,n15491,n15493,n15495,n15499,n15502,n15508,n15514,n15519,n15521,n15523
        ,n15529,n15532,n15534,n15536,n15538,n15540,n15544,n15545,n15555,n15557
        ,n15568,n15573,n15589,n15591,n15593,n15595,n15599,n15602,n15608,n15614
        ,n15625,n15645,n15648,n15651,n15653,n15663,n15665,n15668,n15670,n15679
        ,n15681,n15684,n15686,n15695,n15697,n15700,n15702,n15711,n15713,n15716
        ,n15718,n15727,n15729,n15731,n15733,n15737,n15740,n15746,n15752,n15762
        ,n15769,n15782,n15789,n15791,n15798,n15800,n15802,n15804,n15808,n15815
        ,n15821,n15828,n15830,n15832,n15834,n15838,n15841,n15847,n15853,n15858
        ,n15860,n15862,n15868,n15871,n15873,n15875,n15877,n15879,n15883,n15884
        ,n15894,n15896,n15907,n15912,n15928,n15930,n15932,n15934,n15938,n15941
        ,n15947,n15953,n15964,n15985,n15988,n15991,n15993,n16003,n16005,n16008
        ,n16010,n16019,n16021,n16024,n16026,n16035,n16037,n16040,n16042,n16051
        ,n16053,n16056,n16058,n16067,n16069,n16071,n16073,n16077,n16080,n16086
        ,n16092,n16102,n16109,n16122,n16129,n16131,n16138,n16140,n16142,n16144
        ,n16148,n16155,n16161,n16168,n16170,n16172,n16174,n16178,n16181,n16187
        ,n16193,n16198,n16200,n16202,n16208,n16211,n16213,n16215,n16217,n16219
        ,n16223,n16224,n16234,n16236,n16247,n16252,n16268,n16270,n16272,n16274
        ,n16278,n16281,n16287,n16293,n16304,n16325,n16328,n16331,n16333,n16343
        ,n16345,n16348,n16350,n16359,n16361,n16364,n16366,n16375,n16377,n16380
        ,n16382,n16391,n16393,n16396,n16398,n16407,n16409,n16411,n16413,n16417
        ,n16420,n16426,n16432,n16442,n16449,n16462,n16469,n16471,n16478,n16480
        ,n16482,n16484,n16488,n16495,n16501,n16508,n16510,n16512,n16514,n16518
        ,n16521,n16527,n16533,n16538,n16540,n16542,n16548,n16551,n16553,n16555
        ,n16557,n16559,n16563,n16564,n16574,n16576,n16587,n16592,n16610,n16611
        ,n16612,n16622,n16623,n16624,n16631,n16636,n16675,n16693,n16696,n16699
        ,n16701,n16711,n16713,n16716,n16718,n16727,n16729,n16732,n16734,n16743
        ,n16745,n16748,n16750,n16759,n16761,n16764,n16766,n16775,n16777,n16779
        ,n16781,n16785,n16788,n16794,n16800,n16810,n16817,n16830,n16837,n16839
        ,n16846,n16848,n16850,n16852,n16856,n16863,n16869,n16876,n16878,n16880
        ,n16882,n16886,n16889,n16895,n16901,n16906,n16908,n16910,n16916,n16919
        ,n16921,n16923,n16925,n16927,n16931,n16932,n16942,n16944,n16955,n16975
        ,n16977,n16979,n16981,n16985,n16988,n16994,n17000,n17011,n17400,n17404
        ,n17407,n17409,n17416,n17417,n17453,n17457,n17460,n17462,n17469,n17470
        ,n17499,n17503,n17506,n17508,n17515,n17516,n17546,n17550,n17553,n17555
        ,n17562,n17563,n17592,n17596,n17599,n17601,n17634,n17638,n17641,n17643
        ,n17665,n17669,n17672,n17674,n17695,n17699,n17702,n17704,n17743,n17761
        ,n17789,n17791,n17888,n17898,n17919,n17921,n17923,n18002,n18018,n18042
        ,n18044,n18046,n18125,n18135,n18156,n18158,n18160,n18239,n18249,n18270
        ,n18272,n18274,n18353,n18363,n18384,n18386,n18388,n18467,n18477,n18498
        ,n18500,n18502,n18580,n18590,n18611,n18613,n18615,n18746,n18788,n18831
        ,n18874,n18917,n18960,n19003,n19045,n19208,n19215,n19259,n19288,n19295
        ,n19338,n19361,n19368,n19411,n19445,n19452,n19492,n19515,n19522,n19562
        ,n19586,n19593,n19633,n19656,n19663,n19703,n19740,n19747,n19787);
output out;
input n3;
input n21;
input n26;
input n28;
input n29;
input n31;
input n35;
input n38;
input n44;
input n62;
input n76;
input n77;
input n78;
input n79;
input n80;
input n81;
input n82;
input n83;
input n87;
input n88;
input n89;
input n93;
input n95;
input n97;
input n134;
input n136;
input n137;
input n138;
input n149;
input n150;
input n151;
input n152;
input n164;
input n165;
input n166;
input n167;
input n180;
input n181;
input n182;
input n183;
input n189;
input n191;
input n192;
input n195;
input n197;
input n200;
input n202;
input n203;
input n204;
input n284;
input n390;
input n393;
input n395;
input n549;
input n551;
input n552;
input n555;
input n558;
input n559;
input n560;
input n561;
input n564;
input n566;
input n570;
input n581;
input n582;
input n599;
input n602;
input n604;
input n605;
input n607;
input n611;
input n617;
input n620;
input n622;
input n624;
input n628;
input n631;
input n633;
input n635;
input n639;
input n642;
input n644;
input n646;
input n648;
input n656;
input n659;
input n661;
input n663;
input n667;
input n670;
input n672;
input n674;
input n678;
input n681;
input n683;
input n685;
input n689;
input n692;
input n694;
input n696;
input n704;
input n707;
input n709;
input n711;
input n715;
input n718;
input n720;
input n722;
input n726;
input n729;
input n731;
input n733;
input n737;
input n740;
input n742;
input n744;
input n752;
input n755;
input n757;
input n759;
input n776;
input n779;
input n781;
input n783;
input n792;
input n795;
input n797;
input n799;
input n808;
input n811;
input n813;
input n815;
input n824;
input n827;
input n829;
input n831;
input n840;
input n843;
input n845;
input n847;
input n855;
input n858;
input n860;
input n862;
input n935;
input n938;
input n940;
input n942;
input n946;
input n949;
input n951;
input n953;
input n957;
input n960;
input n962;
input n964;
input n968;
input n971;
input n973;
input n975;
input n984;
input n987;
input n989;
input n991;
input n995;
input n998;
input n1000;
input n1002;
input n1006;
input n1009;
input n1011;
input n1013;
input n1017;
input n1020;
input n1022;
input n1024;
input n1032;
input n1035;
input n1037;
input n1039;
input n1043;
input n1046;
input n1048;
input n1050;
input n1054;
input n1057;
input n1059;
input n1061;
input n1065;
input n1068;
input n1070;
input n1072;
input n1248;
input n1251;
input n1253;
input n1255;
input n1264;
input n1267;
input n1269;
input n1271;
input n1280;
input n1283;
input n1285;
input n1287;
input n1296;
input n1299;
input n1301;
input n1303;
input n1312;
input n1315;
input n1317;
input n1319;
input n1328;
input n1331;
input n1333;
input n1335;
input n1344;
input n1347;
input n1349;
input n1351;
input n1359;
input n1362;
input n1364;
input n1366;
input n1689;
input n1692;
input n1694;
input n1696;
input n1705;
input n1708;
input n1710;
input n1712;
input n1724;
input n1727;
input n1729;
input n1731;
input n1750;
input n1753;
input n1755;
input n1757;
input n1766;
input n1769;
input n1771;
input n1773;
input n1787;
input n1790;
input n1792;
input n1794;
input n1817;
input n1820;
input n1822;
input n1824;
input n1840;
input n1843;
input n1845;
input n1847;
input n2084;
input n2087;
input n2089;
input n2091;
input n2100;
input n2103;
input n2105;
input n2107;
input n2116;
input n2119;
input n2121;
input n2123;
input n2132;
input n2135;
input n2137;
input n2139;
input n2148;
input n2151;
input n2153;
input n2155;
input n2164;
input n2167;
input n2169;
input n2171;
input n2181;
input n2184;
input n2186;
input n2188;
input n2196;
input n2199;
input n2201;
input n2203;
input n2711;
input n2713;
input n2715;
input n2717;
input n2723;
input n2725;
input n2727;
input n2729;
input n2735;
input n2737;
input n2739;
input n2741;
input n2747;
input n2749;
input n2890;
input n2901;
input n2928;
input n2954;
input n2962;
input n2971;
input n2982;
input n2985;
input n2988;
input n2991;
input n2996;
input n2999;
input n3002;
input n3005;
input n3010;
input n3013;
input n3023;
input n3024;
input n3038;
input n3039;
input n3057;
input n3058;
input n3061;
input n3062;
input n3065;
input n3066;
input n3069;
input n3070;
input n3075;
input n3076;
input n3079;
input n3080;
input n3083;
input n3084;
input n3087;
input n3088;
input n3093;
input n3094;
input n3097;
input n3098;
input n3101;
input n3102;
input n3105;
input n3106;
input n3111;
input n3112;
input n3115;
input n3116;
input n3126;
input n3127;
input n3141;
input n3142;
input n3160;
input n3161;
input n3164;
input n3165;
input n3168;
input n3169;
input n3172;
input n3173;
input n3178;
input n3179;
input n3182;
input n3183;
input n3186;
input n3187;
input n3190;
input n3191;
input n3196;
input n3197;
input n3200;
input n3201;
input n3204;
input n3205;
input n3208;
input n3209;
input n3214;
input n3215;
input n3218;
input n3219;
input n3229;
input n3230;
input n3244;
input n3245;
input n3263;
input n3264;
input n3267;
input n3268;
input n3271;
input n3272;
input n3275;
input n3276;
input n3281;
input n3282;
input n3285;
input n3286;
input n3289;
input n3290;
input n3293;
input n3294;
input n3299;
input n3300;
input n3303;
input n3304;
input n3307;
input n3308;
input n3311;
input n3312;
input n3317;
input n3318;
input n3321;
input n3322;
input n3332;
input n3333;
input n3347;
input n3348;
input n3366;
input n3367;
input n3370;
input n3371;
input n3374;
input n3375;
input n3378;
input n3379;
input n3384;
input n3385;
input n3388;
input n3389;
input n3392;
input n3393;
input n3396;
input n3397;
input n3402;
input n3403;
input n3406;
input n3407;
input n3410;
input n3411;
input n3414;
input n3415;
input n3420;
input n3421;
input n3424;
input n3425;
input n3435;
input n3436;
input n3450;
input n3451;
input n3469;
input n3470;
input n3473;
input n3474;
input n3477;
input n3478;
input n3481;
input n3482;
input n3487;
input n3488;
input n3491;
input n3492;
input n3495;
input n3496;
input n3499;
input n3500;
input n3505;
input n3506;
input n3509;
input n3510;
input n3513;
input n3514;
input n3517;
input n3518;
input n3523;
input n3524;
input n3527;
input n3528;
input n3538;
input n3539;
input n3553;
input n3554;
input n3572;
input n3573;
input n3576;
input n3577;
input n3580;
input n3581;
input n3584;
input n3585;
input n3590;
input n3591;
input n3594;
input n3595;
input n3598;
input n3599;
input n3602;
input n3603;
input n3608;
input n3609;
input n3612;
input n3613;
input n3616;
input n3617;
input n3620;
input n3621;
input n3626;
input n3627;
input n3630;
input n3631;
input n3641;
input n3642;
input n3656;
input n3657;
input n3674;
input n3675;
input n3678;
input n3679;
input n3682;
input n3683;
input n3686;
input n3687;
input n3692;
input n3693;
input n3696;
input n3697;
input n3700;
input n3701;
input n3704;
input n3705;
input n3710;
input n3711;
input n3714;
input n3715;
input n3718;
input n3719;
input n3722;
input n3723;
input n3728;
input n3729;
input n3732;
input n3733;
input n3743;
input n3744;
input n3758;
input n3759;
input n3800;
input n3801;
input n3820;
input n3821;
input n3835;
input n3836;
input n3863;
input n3864;
input n3883;
input n3884;
input n3898;
input n3899;
input n3926;
input n3927;
input n3946;
input n3947;
input n3961;
input n3962;
input n3989;
input n3990;
input n4009;
input n4010;
input n4024;
input n4025;
input n4052;
input n4053;
input n4072;
input n4073;
input n4087;
input n4088;
input n4115;
input n4116;
input n4135;
input n4136;
input n4150;
input n4151;
input n4178;
input n4179;
input n4198;
input n4199;
input n4213;
input n4214;
input n4240;
input n4241;
input n4260;
input n4261;
input n4275;
input n4276;
input n4393;
input n4394;
input n4408;
input n4409;
input n4418;
input n4419;
input n4436;
input n4437;
input n4451;
input n4452;
input n4461;
input n4462;
input n4479;
input n4480;
input n4494;
input n4495;
input n4504;
input n4505;
input n4522;
input n4523;
input n4537;
input n4538;
input n4547;
input n4548;
input n4565;
input n4566;
input n4580;
input n4581;
input n4590;
input n4591;
input n4608;
input n4609;
input n4623;
input n4624;
input n4633;
input n4634;
input n4651;
input n4652;
input n4666;
input n4667;
input n4676;
input n4677;
input n4693;
input n4694;
input n4708;
input n4709;
input n4718;
input n4719;
input n4965;
input n4975;
input n4979;
input n4981;
input n4986;
input n4988;
input n4993;
input n4995;
input n5000;
input n5002;
input n5012;
input n5013;
input n5027;
input n5032;
input n5037;
input n5044;
input n5047;
input n5050;
input n5053;
input n5058;
input n5059;
input n5062;
input n5065;
input n5068;
input n5073;
input n5076;
input n5081;
input n5088;
input n5089;
input n5092;
input n5095;
input n5098;
input n5103;
input n5106;
input n5109;
input n5112;
input n5117;
input n5118;
input n5121;
input n5124;
input n5127;
input n5132;
input n5135;
input n5138;
input n5141;
input n5142;
input n5152;
input n5153;
input n5156;
input n5159;
input n5162;
input n5167;
input n5170;
input n5173;
input n5176;
input n5181;
input n5182;
input n5185;
input n5188;
input n5191;
input n5196;
input n5199;
input n5204;
input n5211;
input n5212;
input n5215;
input n5218;
input n5221;
input n5226;
input n5229;
input n5232;
input n5235;
input n5240;
input n5241;
input n5244;
input n5247;
input n5250;
input n5255;
input n5258;
input n5261;
input n5264;
input n5265;
input n5275;
input n5276;
input n5279;
input n5282;
input n5285;
input n5290;
input n5293;
input n5296;
input n5299;
input n5304;
input n5305;
input n5308;
input n5311;
input n5314;
input n5319;
input n5322;
input n5327;
input n5334;
input n5335;
input n5338;
input n5341;
input n5344;
input n5349;
input n5352;
input n5355;
input n5358;
input n5363;
input n5364;
input n5367;
input n5370;
input n5373;
input n5378;
input n5381;
input n5384;
input n5387;
input n5388;
input n5398;
input n5399;
input n5402;
input n5405;
input n5408;
input n5413;
input n5416;
input n5419;
input n5422;
input n5427;
input n5428;
input n5431;
input n5434;
input n5437;
input n5442;
input n5445;
input n5450;
input n5457;
input n5458;
input n5461;
input n5464;
input n5467;
input n5472;
input n5475;
input n5478;
input n5481;
input n5486;
input n5487;
input n5490;
input n5493;
input n5496;
input n5501;
input n5504;
input n5507;
input n5510;
input n5511;
input n5521;
input n5522;
input n5525;
input n5528;
input n5531;
input n5536;
input n5539;
input n5542;
input n5545;
input n5550;
input n5551;
input n5554;
input n5557;
input n5560;
input n5565;
input n5568;
input n5573;
input n5580;
input n5581;
input n5584;
input n5587;
input n5590;
input n5595;
input n5598;
input n5601;
input n5604;
input n5609;
input n5610;
input n5613;
input n5616;
input n5619;
input n5624;
input n5627;
input n5630;
input n5633;
input n5634;
input n5644;
input n5645;
input n5648;
input n5651;
input n5654;
input n5659;
input n5662;
input n5665;
input n5668;
input n5673;
input n5674;
input n5677;
input n5680;
input n5683;
input n5688;
input n5691;
input n5696;
input n5703;
input n5704;
input n5707;
input n5710;
input n5713;
input n5718;
input n5721;
input n5724;
input n5727;
input n5732;
input n5733;
input n5736;
input n5739;
input n5742;
input n5747;
input n5750;
input n5753;
input n5756;
input n5757;
input n5767;
input n5768;
input n5771;
input n5774;
input n5777;
input n5782;
input n5785;
input n5788;
input n5791;
input n5796;
input n5797;
input n5800;
input n5803;
input n5806;
input n5811;
input n5814;
input n5819;
input n5826;
input n5827;
input n5830;
input n5833;
input n5836;
input n5841;
input n5844;
input n5847;
input n5850;
input n5855;
input n5856;
input n5859;
input n5862;
input n5865;
input n5870;
input n5873;
input n5876;
input n5879;
input n5880;
input n5889;
input n5890;
input n5893;
input n5896;
input n5899;
input n5904;
input n5907;
input n5910;
input n5913;
input n5918;
input n5919;
input n5922;
input n5925;
input n5928;
input n5933;
input n5936;
input n5941;
input n5948;
input n5949;
input n5952;
input n5955;
input n5958;
input n5963;
input n5966;
input n5969;
input n5972;
input n5977;
input n5978;
input n5981;
input n5984;
input n5987;
input n5992;
input n5995;
input n5998;
input n6001;
input n6002;
input n6020;
input n6022;
input n6026;
input n6028;
input n6033;
input n6035;
input n6081;
input n6124;
input n6170;
input n6213;
input n6259;
input n6302;
input n6348;
input n6391;
input n6437;
input n6480;
input n6526;
input n6569;
input n6615;
input n6658;
input n6703;
input n6746;
input n6760;
input n6762;
input n6766;
input n6768;
input n6773;
input n6775;
input n6780;
input n6782;
input n6787;
input n6789;
input n6801;
input n6802;
input n6805;
input n6808;
input n6811;
input n6816;
input n6819;
input n6824;
input n6831;
input n6832;
input n6835;
input n6838;
input n6841;
input n6846;
input n6849;
input n6852;
input n6855;
input n6858;
input n6870;
input n6871;
input n6874;
input n6877;
input n6880;
input n6885;
input n6888;
input n6893;
input n6900;
input n6901;
input n6904;
input n6907;
input n6910;
input n6915;
input n6918;
input n6921;
input n6924;
input n6927;
input n6939;
input n6940;
input n6943;
input n6946;
input n6949;
input n6954;
input n6957;
input n6962;
input n6969;
input n6970;
input n6973;
input n6976;
input n6979;
input n6984;
input n6987;
input n6990;
input n6993;
input n6996;
input n7008;
input n7009;
input n7012;
input n7015;
input n7018;
input n7023;
input n7026;
input n7031;
input n7038;
input n7039;
input n7042;
input n7045;
input n7048;
input n7053;
input n7056;
input n7059;
input n7062;
input n7065;
input n7077;
input n7078;
input n7081;
input n7084;
input n7087;
input n7092;
input n7095;
input n7100;
input n7107;
input n7108;
input n7111;
input n7114;
input n7117;
input n7122;
input n7125;
input n7128;
input n7131;
input n7134;
input n7146;
input n7147;
input n7150;
input n7153;
input n7156;
input n7161;
input n7164;
input n7169;
input n7176;
input n7177;
input n7180;
input n7183;
input n7186;
input n7191;
input n7194;
input n7197;
input n7200;
input n7203;
input n7215;
input n7216;
input n7219;
input n7222;
input n7225;
input n7230;
input n7233;
input n7238;
input n7245;
input n7246;
input n7249;
input n7252;
input n7255;
input n7260;
input n7263;
input n7266;
input n7269;
input n7272;
input n7283;
input n7284;
input n7287;
input n7290;
input n7293;
input n7298;
input n7301;
input n7306;
input n7313;
input n7314;
input n7317;
input n7320;
input n7323;
input n7328;
input n7331;
input n7334;
input n7337;
input n7340;
input n7644;
input n7646;
input n7653;
input n7655;
input n7669;
input n7671;
input n7678;
input n7680;
input n7685;
input n7687;
input n7692;
input n7694;
input n7708;
input n7710;
input n7717;
input n7719;
input n7885;
input n7888;
input n7997;
input n8000;
input n8109;
input n8112;
input n8221;
input n8224;
input n8329;
input n8332;
input n8437;
input n8440;
input n8544;
input n8547;
input n9092;
input n9106;
input n9120;
input n9142;
input n9166;
input n9189;
input n9215;
input n9231;
input n9405;
input n9417;
input n9429;
input n9441;
input n9453;
input n9465;
input n9477;
input n9488;
input n9941;
input n9944;
input n10553;
input n10554;
input n10568;
input n10574;
input n10575;
input n10589;
input n10590;
input n10617;
input n10618;
input n10632;
input n10638;
input n10639;
input n10653;
input n10654;
input n10681;
input n10682;
input n10696;
input n10702;
input n10703;
input n10717;
input n10718;
input n10745;
input n10746;
input n10760;
input n10766;
input n10767;
input n10781;
input n10782;
input n10810;
input n10811;
input n10825;
input n10831;
input n10832;
input n10847;
input n10848;
input n10877;
input n10878;
input n10893;
input n10899;
input n10900;
input n10914;
input n10915;
input n10942;
input n10943;
input n10957;
input n10963;
input n10964;
input n10978;
input n10979;
input n11006;
input n11007;
input n11022;
input n11028;
input n11029;
input n11044;
input n11045;
input n11163;
input n11164;
input n11174;
input n11180;
input n11181;
input n11191;
input n11192;
input n11210;
input n11211;
input n11221;
input n11227;
input n11228;
input n11238;
input n11239;
input n11257;
input n11258;
input n11268;
input n11274;
input n11275;
input n11285;
input n11286;
input n11304;
input n11305;
input n11315;
input n11321;
input n11322;
input n11332;
input n11333;
input n11351;
input n11352;
input n11362;
input n11368;
input n11369;
input n11378;
input n11379;
input n11396;
input n11397;
input n11407;
input n11413;
input n11414;
input n11424;
input n11425;
input n11443;
input n11444;
input n11454;
input n11460;
input n11461;
input n11471;
input n11472;
input n11489;
input n11490;
input n11500;
input n11506;
input n11507;
input n11517;
input n11518;
input n11747;
input n11751;
input n11756;
input n11761;
input n11766;
input n11776;
input n11777;
input n11780;
input n11783;
input n11786;
input n11791;
input n11794;
input n11797;
input n11800;
input n11803;
input n11813;
input n11814;
input n11817;
input n11820;
input n11823;
input n11828;
input n11831;
input n11834;
input n11837;
input n11840;
input n11850;
input n11851;
input n11854;
input n11857;
input n11860;
input n11865;
input n11868;
input n11871;
input n11874;
input n11877;
input n11887;
input n11888;
input n11891;
input n11894;
input n11897;
input n11902;
input n11905;
input n11908;
input n11911;
input n11914;
input n11924;
input n11925;
input n11928;
input n11931;
input n11934;
input n11939;
input n11942;
input n11945;
input n11948;
input n11951;
input n11961;
input n11962;
input n11965;
input n11968;
input n11971;
input n11976;
input n11979;
input n11982;
input n11985;
input n11988;
input n11998;
input n11999;
input n12002;
input n12005;
input n12008;
input n12013;
input n12016;
input n12019;
input n12022;
input n12025;
input n12034;
input n12035;
input n12038;
input n12041;
input n12044;
input n12049;
input n12052;
input n12055;
input n12058;
input n12061;
input n12124;
input n12127;
input n12131;
input n12134;
input n12144;
input n12145;
input n12148;
input n12151;
input n12154;
input n12159;
input n12162;
input n12165;
input n12168;
input n12171;
input n12181;
input n12182;
input n12185;
input n12188;
input n12191;
input n12196;
input n12199;
input n12202;
input n12205;
input n12208;
input n12218;
input n12219;
input n12222;
input n12225;
input n12228;
input n12233;
input n12236;
input n12239;
input n12242;
input n12245;
input n12255;
input n12256;
input n12259;
input n12262;
input n12265;
input n12270;
input n12273;
input n12276;
input n12279;
input n12282;
input n12292;
input n12293;
input n12296;
input n12299;
input n12302;
input n12307;
input n12310;
input n12313;
input n12316;
input n12319;
input n12329;
input n12330;
input n12333;
input n12336;
input n12339;
input n12344;
input n12347;
input n12350;
input n12353;
input n12356;
input n12366;
input n12367;
input n12370;
input n12373;
input n12376;
input n12381;
input n12384;
input n12387;
input n12390;
input n12393;
input n12402;
input n12403;
input n12406;
input n12409;
input n12412;
input n12417;
input n12420;
input n12423;
input n12426;
input n12429;
input n12455;
input n12824;
input n12831;
input n12874;
input n12877;
input n13067;
input n13070;
input n13179;
input n13182;
input n13291;
input n13294;
input n13403;
input n13406;
input n13511;
input n13514;
input n13619;
input n13622;
input n13726;
input n13729;
input n13888;
input n13890;
input n13892;
input n13894;
input n13896;
input n13899;
input n13906;
input n13908;
input n13909;
input n13912;
input n13919;
input n13922;
input n13927;
input n13934;
input n13954;
input n13956;
input n13958;
input n13960;
input n13962;
input n13964;
input n13966;
input n13968;
input n13970;
input n13972;
input n13974;
input n13976;
input n13978;
input n13980;
input n13982;
input n13984;
input n13989;
input n13997;
input n14002;
input n14008;
input n14010;
input n14012;
input n14014;
input n14016;
input n14018;
input n14020;
input n14022;
input n14024;
input n14026;
input n14028;
input n14030;
input n14032;
input n14034;
input n14036;
input n14038;
input n14043;
input n14045;
input n14047;
input n14049;
input n14051;
input n14053;
input n14055;
input n14057;
input n14059;
input n14061;
input n14063;
input n14065;
input n14067;
input n14069;
input n14071;
input n14073;
input n14077;
input n14079;
input n14081;
input n14083;
input n14085;
input n14087;
input n14089;
input n14091;
input n14093;
input n14095;
input n14097;
input n14099;
input n14101;
input n14103;
input n14105;
input n14107;
input n14114;
input n14115;
input n14121;
input n14122;
input n14127;
input n14128;
input n14129;
input n14130;
input n14146;
input n14155;
input n14170;
input n14175;
input n14198;
input n14202;
input n14204;
input n14209;
input n14213;
input n14214;
input n14215;
input n14216;
input n14219;
input n14220;
input n14222;
input n14223;
input n14240;
input n14253;
input n14285;
input n14287;
input n14290;
input n14292;
input n14302;
input n14304;
input n14307;
input n14309;
input n14314;
input n14320;
input n14323;
input n14341;
input n14351;
input n14354;
input n14357;
input n14360;
input n14373;
input n14392;
input n14411;
input n14420;
input n14428;
input n14436;
input n14441;
input n14461;
input n14463;
input n14465;
input n14467;
input n14471;
input n14474;
input n14480;
input n14486;
input n14507;
input n14510;
input n14524;
input n14526;
input n14528;
input n14530;
input n14534;
input n14541;
input n14547;
input n14556;
input n14557;
input n14562;
input n14582;
input n14584;
input n14586;
input n14588;
input n14592;
input n14595;
input n14601;
input n14607;
input n14618;
input n14642;
input n14645;
input n14648;
input n14650;
input n14660;
input n14662;
input n14665;
input n14667;
input n14676;
input n14678;
input n14681;
input n14683;
input n14692;
input n14694;
input n14697;
input n14699;
input n14708;
input n14710;
input n14713;
input n14715;
input n14725;
input n14727;
input n14729;
input n14731;
input n14735;
input n14738;
input n14744;
input n14750;
input n14760;
input n14767;
input n14780;
input n14787;
input n14789;
input n14796;
input n14798;
input n14800;
input n14802;
input n14806;
input n14813;
input n14819;
input n14826;
input n14828;
input n14830;
input n14832;
input n14836;
input n14839;
input n14845;
input n14851;
input n14855;
input n14857;
input n14859;
input n14865;
input n14868;
input n14870;
input n14872;
input n14874;
input n14876;
input n14880;
input n14881;
input n14891;
input n14893;
input n14904;
input n14909;
input n14925;
input n14927;
input n14929;
input n14931;
input n14935;
input n14938;
input n14944;
input n14950;
input n14961;
input n14978;
input n14980;
input n14982;
input n14988;
input n14991;
input n14993;
input n14995;
input n14997;
input n14999;
input n15003;
input n15004;
input n15017;
input n15019;
input n15022;
input n15024;
input n15031;
input n15034;
input n15036;
input n15044;
input n15046;
input n15049;
input n15051;
input n15061;
input n15063;
input n15066;
input n15068;
input n15077;
input n15079;
input n15082;
input n15084;
input n15097;
input n15100;
input n15107;
input n15111;
input n15113;
input n15117;
input n15124;
input n15126;
input n15128;
input n15130;
input n15134;
input n15137;
input n15143;
input n15149;
input n15156;
input n15158;
input n15160;
input n15162;
input n15166;
input n15169;
input n15175;
input n15181;
input n15185;
input n15188;
input n15196;
input n15198;
input n15200;
input n15202;
input n15206;
input n15213;
input n15219;
input n15228;
input n15233;
input n15249;
input n15251;
input n15253;
input n15255;
input n15259;
input n15262;
input n15268;
input n15274;
input n15285;
input n15306;
input n15309;
input n15312;
input n15314;
input n15324;
input n15326;
input n15329;
input n15331;
input n15340;
input n15342;
input n15345;
input n15347;
input n15356;
input n15358;
input n15361;
input n15363;
input n15372;
input n15374;
input n15377;
input n15379;
input n15388;
input n15390;
input n15392;
input n15394;
input n15398;
input n15401;
input n15407;
input n15413;
input n15423;
input n15430;
input n15443;
input n15450;
input n15452;
input n15459;
input n15461;
input n15463;
input n15465;
input n15469;
input n15476;
input n15482;
input n15489;
input n15491;
input n15493;
input n15495;
input n15499;
input n15502;
input n15508;
input n15514;
input n15519;
input n15521;
input n15523;
input n15529;
input n15532;
input n15534;
input n15536;
input n15538;
input n15540;
input n15544;
input n15545;
input n15555;
input n15557;
input n15568;
input n15573;
input n15589;
input n15591;
input n15593;
input n15595;
input n15599;
input n15602;
input n15608;
input n15614;
input n15625;
input n15645;
input n15648;
input n15651;
input n15653;
input n15663;
input n15665;
input n15668;
input n15670;
input n15679;
input n15681;
input n15684;
input n15686;
input n15695;
input n15697;
input n15700;
input n15702;
input n15711;
input n15713;
input n15716;
input n15718;
input n15727;
input n15729;
input n15731;
input n15733;
input n15737;
input n15740;
input n15746;
input n15752;
input n15762;
input n15769;
input n15782;
input n15789;
input n15791;
input n15798;
input n15800;
input n15802;
input n15804;
input n15808;
input n15815;
input n15821;
input n15828;
input n15830;
input n15832;
input n15834;
input n15838;
input n15841;
input n15847;
input n15853;
input n15858;
input n15860;
input n15862;
input n15868;
input n15871;
input n15873;
input n15875;
input n15877;
input n15879;
input n15883;
input n15884;
input n15894;
input n15896;
input n15907;
input n15912;
input n15928;
input n15930;
input n15932;
input n15934;
input n15938;
input n15941;
input n15947;
input n15953;
input n15964;
input n15985;
input n15988;
input n15991;
input n15993;
input n16003;
input n16005;
input n16008;
input n16010;
input n16019;
input n16021;
input n16024;
input n16026;
input n16035;
input n16037;
input n16040;
input n16042;
input n16051;
input n16053;
input n16056;
input n16058;
input n16067;
input n16069;
input n16071;
input n16073;
input n16077;
input n16080;
input n16086;
input n16092;
input n16102;
input n16109;
input n16122;
input n16129;
input n16131;
input n16138;
input n16140;
input n16142;
input n16144;
input n16148;
input n16155;
input n16161;
input n16168;
input n16170;
input n16172;
input n16174;
input n16178;
input n16181;
input n16187;
input n16193;
input n16198;
input n16200;
input n16202;
input n16208;
input n16211;
input n16213;
input n16215;
input n16217;
input n16219;
input n16223;
input n16224;
input n16234;
input n16236;
input n16247;
input n16252;
input n16268;
input n16270;
input n16272;
input n16274;
input n16278;
input n16281;
input n16287;
input n16293;
input n16304;
input n16325;
input n16328;
input n16331;
input n16333;
input n16343;
input n16345;
input n16348;
input n16350;
input n16359;
input n16361;
input n16364;
input n16366;
input n16375;
input n16377;
input n16380;
input n16382;
input n16391;
input n16393;
input n16396;
input n16398;
input n16407;
input n16409;
input n16411;
input n16413;
input n16417;
input n16420;
input n16426;
input n16432;
input n16442;
input n16449;
input n16462;
input n16469;
input n16471;
input n16478;
input n16480;
input n16482;
input n16484;
input n16488;
input n16495;
input n16501;
input n16508;
input n16510;
input n16512;
input n16514;
input n16518;
input n16521;
input n16527;
input n16533;
input n16538;
input n16540;
input n16542;
input n16548;
input n16551;
input n16553;
input n16555;
input n16557;
input n16559;
input n16563;
input n16564;
input n16574;
input n16576;
input n16587;
input n16592;
input n16610;
input n16611;
input n16612;
input n16622;
input n16623;
input n16624;
input n16631;
input n16636;
input n16675;
input n16693;
input n16696;
input n16699;
input n16701;
input n16711;
input n16713;
input n16716;
input n16718;
input n16727;
input n16729;
input n16732;
input n16734;
input n16743;
input n16745;
input n16748;
input n16750;
input n16759;
input n16761;
input n16764;
input n16766;
input n16775;
input n16777;
input n16779;
input n16781;
input n16785;
input n16788;
input n16794;
input n16800;
input n16810;
input n16817;
input n16830;
input n16837;
input n16839;
input n16846;
input n16848;
input n16850;
input n16852;
input n16856;
input n16863;
input n16869;
input n16876;
input n16878;
input n16880;
input n16882;
input n16886;
input n16889;
input n16895;
input n16901;
input n16906;
input n16908;
input n16910;
input n16916;
input n16919;
input n16921;
input n16923;
input n16925;
input n16927;
input n16931;
input n16932;
input n16942;
input n16944;
input n16955;
input n16975;
input n16977;
input n16979;
input n16981;
input n16985;
input n16988;
input n16994;
input n17000;
input n17011;
input n17400;
input n17404;
input n17407;
input n17409;
input n17416;
input n17417;
input n17453;
input n17457;
input n17460;
input n17462;
input n17469;
input n17470;
input n17499;
input n17503;
input n17506;
input n17508;
input n17515;
input n17516;
input n17546;
input n17550;
input n17553;
input n17555;
input n17562;
input n17563;
input n17592;
input n17596;
input n17599;
input n17601;
input n17634;
input n17638;
input n17641;
input n17643;
input n17665;
input n17669;
input n17672;
input n17674;
input n17695;
input n17699;
input n17702;
input n17704;
input n17743;
input n17761;
input n17789;
input n17791;
input n17888;
input n17898;
input n17919;
input n17921;
input n17923;
input n18002;
input n18018;
input n18042;
input n18044;
input n18046;
input n18125;
input n18135;
input n18156;
input n18158;
input n18160;
input n18239;
input n18249;
input n18270;
input n18272;
input n18274;
input n18353;
input n18363;
input n18384;
input n18386;
input n18388;
input n18467;
input n18477;
input n18498;
input n18500;
input n18502;
input n18580;
input n18590;
input n18611;
input n18613;
input n18615;
input n18746;
input n18788;
input n18831;
input n18874;
input n18917;
input n18960;
input n19003;
input n19045;
input n19208;
input n19215;
input n19259;
input n19288;
input n19295;
input n19338;
input n19361;
input n19368;
input n19411;
input n19445;
input n19452;
input n19492;
input n19515;
input n19522;
input n19562;
input n19586;
input n19593;
input n19633;
input n19656;
input n19663;
input n19703;
input n19740;
input n19747;
input n19787;
wire n0;
wire n1;
wire n2;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n17;
wire n18;
wire n19;
wire n20;
wire n22;
wire n23;
wire n24;
wire n25;
wire n27;
wire n30;
wire n32;
wire n33;
wire n34;
wire n36;
wire n37;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n84;
wire n85;
wire n86;
wire n90;
wire n91;
wire n92;
wire n94;
wire n96;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n135;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n190;
wire n193;
wire n194;
wire n196;
wire n198;
wire n199;
wire n201;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n391;
wire n392;
wire n394;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n550;
wire n553;
wire n554;
wire n556;
wire n557;
wire n562;
wire n563;
wire n565;
wire n567;
wire n568;
wire n569;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n600;
wire n601;
wire n603;
wire n606;
wire n608;
wire n609;
wire n610;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n618;
wire n619;
wire n621;
wire n623;
wire n625;
wire n626;
wire n627;
wire n629;
wire n630;
wire n632;
wire n634;
wire n636;
wire n637;
wire n638;
wire n640;
wire n641;
wire n643;
wire n645;
wire n647;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n657;
wire n658;
wire n660;
wire n662;
wire n664;
wire n665;
wire n666;
wire n668;
wire n669;
wire n671;
wire n673;
wire n675;
wire n676;
wire n677;
wire n679;
wire n680;
wire n682;
wire n684;
wire n686;
wire n687;
wire n688;
wire n690;
wire n691;
wire n693;
wire n695;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n705;
wire n706;
wire n708;
wire n710;
wire n712;
wire n713;
wire n714;
wire n716;
wire n717;
wire n719;
wire n721;
wire n723;
wire n724;
wire n725;
wire n727;
wire n728;
wire n730;
wire n732;
wire n734;
wire n735;
wire n736;
wire n738;
wire n739;
wire n741;
wire n743;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n753;
wire n754;
wire n756;
wire n758;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n777;
wire n778;
wire n780;
wire n782;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n793;
wire n794;
wire n796;
wire n798;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n809;
wire n810;
wire n812;
wire n814;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n825;
wire n826;
wire n828;
wire n830;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n841;
wire n842;
wire n844;
wire n846;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n856;
wire n857;
wire n859;
wire n861;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n936;
wire n937;
wire n939;
wire n941;
wire n943;
wire n944;
wire n945;
wire n947;
wire n948;
wire n950;
wire n952;
wire n954;
wire n955;
wire n956;
wire n958;
wire n959;
wire n961;
wire n963;
wire n965;
wire n966;
wire n967;
wire n969;
wire n970;
wire n972;
wire n974;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n985;
wire n986;
wire n988;
wire n990;
wire n992;
wire n993;
wire n994;
wire n996;
wire n997;
wire n999;
wire n1001;
wire n1003;
wire n1004;
wire n1005;
wire n1007;
wire n1008;
wire n1010;
wire n1012;
wire n1014;
wire n1015;
wire n1016;
wire n1018;
wire n1019;
wire n1021;
wire n1023;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1033;
wire n1034;
wire n1036;
wire n1038;
wire n1040;
wire n1041;
wire n1042;
wire n1044;
wire n1045;
wire n1047;
wire n1049;
wire n1051;
wire n1052;
wire n1053;
wire n1055;
wire n1056;
wire n1058;
wire n1060;
wire n1062;
wire n1063;
wire n1064;
wire n1066;
wire n1067;
wire n1069;
wire n1071;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1249;
wire n1250;
wire n1252;
wire n1254;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1265;
wire n1266;
wire n1268;
wire n1270;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1281;
wire n1282;
wire n1284;
wire n1286;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1297;
wire n1298;
wire n1300;
wire n1302;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1313;
wire n1314;
wire n1316;
wire n1318;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1329;
wire n1330;
wire n1332;
wire n1334;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1345;
wire n1346;
wire n1348;
wire n1350;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1360;
wire n1361;
wire n1363;
wire n1365;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1690;
wire n1691;
wire n1693;
wire n1695;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1706;
wire n1707;
wire n1709;
wire n1711;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1725;
wire n1726;
wire n1728;
wire n1730;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1751;
wire n1752;
wire n1754;
wire n1756;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1767;
wire n1768;
wire n1770;
wire n1772;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1788;
wire n1789;
wire n1791;
wire n1793;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1818;
wire n1819;
wire n1821;
wire n1823;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1841;
wire n1842;
wire n1844;
wire n1846;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2085;
wire n2086;
wire n2088;
wire n2090;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2101;
wire n2102;
wire n2104;
wire n2106;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2117;
wire n2118;
wire n2120;
wire n2122;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2133;
wire n2134;
wire n2136;
wire n2138;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2149;
wire n2150;
wire n2152;
wire n2154;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2165;
wire n2166;
wire n2168;
wire n2170;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2182;
wire n2183;
wire n2185;
wire n2187;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2197;
wire n2198;
wire n2200;
wire n2202;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2712;
wire n2714;
wire n2716;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2724;
wire n2726;
wire n2728;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2736;
wire n2738;
wire n2740;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2748;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2983;
wire n2984;
wire n2986;
wire n2987;
wire n2989;
wire n2990;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2997;
wire n2998;
wire n3000;
wire n3001;
wire n3003;
wire n3004;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3011;
wire n3012;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
wire n3056;
wire n3059;
wire n3060;
wire n3063;
wire n3064;
wire n3067;
wire n3068;
wire n3071;
wire n3072;
wire n3073;
wire n3074;
wire n3077;
wire n3078;
wire n3081;
wire n3082;
wire n3085;
wire n3086;
wire n3089;
wire n3090;
wire n3091;
wire n3092;
wire n3095;
wire n3096;
wire n3099;
wire n3100;
wire n3103;
wire n3104;
wire n3107;
wire n3108;
wire n3109;
wire n3110;
wire n3113;
wire n3114;
wire n3117;
wire n3118;
wire n3119;
wire n3120;
wire n3121;
wire n3122;
wire n3123;
wire n3124;
wire n3125;
wire n3128;
wire n3129;
wire n3130;
wire n3131;
wire n3132;
wire n3133;
wire n3134;
wire n3135;
wire n3136;
wire n3137;
wire n3138;
wire n3139;
wire n3140;
wire n3143;
wire n3144;
wire n3145;
wire n3146;
wire n3147;
wire n3148;
wire n3149;
wire n3150;
wire n3151;
wire n3152;
wire n3153;
wire n3154;
wire n3155;
wire n3156;
wire n3157;
wire n3158;
wire n3159;
wire n3162;
wire n3163;
wire n3166;
wire n3167;
wire n3170;
wire n3171;
wire n3174;
wire n3175;
wire n3176;
wire n3177;
wire n3180;
wire n3181;
wire n3184;
wire n3185;
wire n3188;
wire n3189;
wire n3192;
wire n3193;
wire n3194;
wire n3195;
wire n3198;
wire n3199;
wire n3202;
wire n3203;
wire n3206;
wire n3207;
wire n3210;
wire n3211;
wire n3212;
wire n3213;
wire n3216;
wire n3217;
wire n3220;
wire n3221;
wire n3222;
wire n3223;
wire n3224;
wire n3225;
wire n3226;
wire n3227;
wire n3228;
wire n3231;
wire n3232;
wire n3233;
wire n3234;
wire n3235;
wire n3236;
wire n3237;
wire n3238;
wire n3239;
wire n3240;
wire n3241;
wire n3242;
wire n3243;
wire n3246;
wire n3247;
wire n3248;
wire n3249;
wire n3250;
wire n3251;
wire n3252;
wire n3253;
wire n3254;
wire n3255;
wire n3256;
wire n3257;
wire n3258;
wire n3259;
wire n3260;
wire n3261;
wire n3262;
wire n3265;
wire n3266;
wire n3269;
wire n3270;
wire n3273;
wire n3274;
wire n3277;
wire n3278;
wire n3279;
wire n3280;
wire n3283;
wire n3284;
wire n3287;
wire n3288;
wire n3291;
wire n3292;
wire n3295;
wire n3296;
wire n3297;
wire n3298;
wire n3301;
wire n3302;
wire n3305;
wire n3306;
wire n3309;
wire n3310;
wire n3313;
wire n3314;
wire n3315;
wire n3316;
wire n3319;
wire n3320;
wire n3323;
wire n3324;
wire n3325;
wire n3326;
wire n3327;
wire n3328;
wire n3329;
wire n3330;
wire n3331;
wire n3334;
wire n3335;
wire n3336;
wire n3337;
wire n3338;
wire n3339;
wire n3340;
wire n3341;
wire n3342;
wire n3343;
wire n3344;
wire n3345;
wire n3346;
wire n3349;
wire n3350;
wire n3351;
wire n3352;
wire n3353;
wire n3354;
wire n3355;
wire n3356;
wire n3357;
wire n3358;
wire n3359;
wire n3360;
wire n3361;
wire n3362;
wire n3363;
wire n3364;
wire n3365;
wire n3368;
wire n3369;
wire n3372;
wire n3373;
wire n3376;
wire n3377;
wire n3380;
wire n3381;
wire n3382;
wire n3383;
wire n3386;
wire n3387;
wire n3390;
wire n3391;
wire n3394;
wire n3395;
wire n3398;
wire n3399;
wire n3400;
wire n3401;
wire n3404;
wire n3405;
wire n3408;
wire n3409;
wire n3412;
wire n3413;
wire n3416;
wire n3417;
wire n3418;
wire n3419;
wire n3422;
wire n3423;
wire n3426;
wire n3427;
wire n3428;
wire n3429;
wire n3430;
wire n3431;
wire n3432;
wire n3433;
wire n3434;
wire n3437;
wire n3438;
wire n3439;
wire n3440;
wire n3441;
wire n3442;
wire n3443;
wire n3444;
wire n3445;
wire n3446;
wire n3447;
wire n3448;
wire n3449;
wire n3452;
wire n3453;
wire n3454;
wire n3455;
wire n3456;
wire n3457;
wire n3458;
wire n3459;
wire n3460;
wire n3461;
wire n3462;
wire n3463;
wire n3464;
wire n3465;
wire n3466;
wire n3467;
wire n3468;
wire n3471;
wire n3472;
wire n3475;
wire n3476;
wire n3479;
wire n3480;
wire n3483;
wire n3484;
wire n3485;
wire n3486;
wire n3489;
wire n3490;
wire n3493;
wire n3494;
wire n3497;
wire n3498;
wire n3501;
wire n3502;
wire n3503;
wire n3504;
wire n3507;
wire n3508;
wire n3511;
wire n3512;
wire n3515;
wire n3516;
wire n3519;
wire n3520;
wire n3521;
wire n3522;
wire n3525;
wire n3526;
wire n3529;
wire n3530;
wire n3531;
wire n3532;
wire n3533;
wire n3534;
wire n3535;
wire n3536;
wire n3537;
wire n3540;
wire n3541;
wire n3542;
wire n3543;
wire n3544;
wire n3545;
wire n3546;
wire n3547;
wire n3548;
wire n3549;
wire n3550;
wire n3551;
wire n3552;
wire n3555;
wire n3556;
wire n3557;
wire n3558;
wire n3559;
wire n3560;
wire n3561;
wire n3562;
wire n3563;
wire n3564;
wire n3565;
wire n3566;
wire n3567;
wire n3568;
wire n3569;
wire n3570;
wire n3571;
wire n3574;
wire n3575;
wire n3578;
wire n3579;
wire n3582;
wire n3583;
wire n3586;
wire n3587;
wire n3588;
wire n3589;
wire n3592;
wire n3593;
wire n3596;
wire n3597;
wire n3600;
wire n3601;
wire n3604;
wire n3605;
wire n3606;
wire n3607;
wire n3610;
wire n3611;
wire n3614;
wire n3615;
wire n3618;
wire n3619;
wire n3622;
wire n3623;
wire n3624;
wire n3625;
wire n3628;
wire n3629;
wire n3632;
wire n3633;
wire n3634;
wire n3635;
wire n3636;
wire n3637;
wire n3638;
wire n3639;
wire n3640;
wire n3643;
wire n3644;
wire n3645;
wire n3646;
wire n3647;
wire n3648;
wire n3649;
wire n3650;
wire n3651;
wire n3652;
wire n3653;
wire n3654;
wire n3655;
wire n3658;
wire n3659;
wire n3660;
wire n3661;
wire n3662;
wire n3663;
wire n3664;
wire n3665;
wire n3666;
wire n3667;
wire n3668;
wire n3669;
wire n3670;
wire n3671;
wire n3672;
wire n3673;
wire n3676;
wire n3677;
wire n3680;
wire n3681;
wire n3684;
wire n3685;
wire n3688;
wire n3689;
wire n3690;
wire n3691;
wire n3694;
wire n3695;
wire n3698;
wire n3699;
wire n3702;
wire n3703;
wire n3706;
wire n3707;
wire n3708;
wire n3709;
wire n3712;
wire n3713;
wire n3716;
wire n3717;
wire n3720;
wire n3721;
wire n3724;
wire n3725;
wire n3726;
wire n3727;
wire n3730;
wire n3731;
wire n3734;
wire n3735;
wire n3736;
wire n3737;
wire n3738;
wire n3739;
wire n3740;
wire n3741;
wire n3742;
wire n3745;
wire n3746;
wire n3747;
wire n3748;
wire n3749;
wire n3750;
wire n3751;
wire n3752;
wire n3753;
wire n3754;
wire n3755;
wire n3756;
wire n3757;
wire n3760;
wire n3761;
wire n3762;
wire n3763;
wire n3764;
wire n3765;
wire n3766;
wire n3767;
wire n3768;
wire n3769;
wire n3770;
wire n3771;
wire n3772;
wire n3773;
wire n3774;
wire n3775;
wire n3776;
wire n3777;
wire n3778;
wire n3779;
wire n3780;
wire n3781;
wire n3782;
wire n3783;
wire n3784;
wire n3785;
wire n3786;
wire n3787;
wire n3788;
wire n3789;
wire n3790;
wire n3791;
wire n3792;
wire n3793;
wire n3794;
wire n3795;
wire n3796;
wire n3797;
wire n3798;
wire n3799;
wire n3802;
wire n3803;
wire n3804;
wire n3805;
wire n3806;
wire n3807;
wire n3808;
wire n3809;
wire n3810;
wire n3811;
wire n3812;
wire n3813;
wire n3814;
wire n3815;
wire n3816;
wire n3817;
wire n3818;
wire n3819;
wire n3822;
wire n3823;
wire n3824;
wire n3825;
wire n3826;
wire n3827;
wire n3828;
wire n3829;
wire n3830;
wire n3831;
wire n3832;
wire n3833;
wire n3834;
wire n3837;
wire n3838;
wire n3839;
wire n3840;
wire n3841;
wire n3842;
wire n3843;
wire n3844;
wire n3845;
wire n3846;
wire n3847;
wire n3848;
wire n3849;
wire n3850;
wire n3851;
wire n3852;
wire n3853;
wire n3854;
wire n3855;
wire n3856;
wire n3857;
wire n3858;
wire n3859;
wire n3860;
wire n3861;
wire n3862;
wire n3865;
wire n3866;
wire n3867;
wire n3868;
wire n3869;
wire n3870;
wire n3871;
wire n3872;
wire n3873;
wire n3874;
wire n3875;
wire n3876;
wire n3877;
wire n3878;
wire n3879;
wire n3880;
wire n3881;
wire n3882;
wire n3885;
wire n3886;
wire n3887;
wire n3888;
wire n3889;
wire n3890;
wire n3891;
wire n3892;
wire n3893;
wire n3894;
wire n3895;
wire n3896;
wire n3897;
wire n3900;
wire n3901;
wire n3902;
wire n3903;
wire n3904;
wire n3905;
wire n3906;
wire n3907;
wire n3908;
wire n3909;
wire n3910;
wire n3911;
wire n3912;
wire n3913;
wire n3914;
wire n3915;
wire n3916;
wire n3917;
wire n3918;
wire n3919;
wire n3920;
wire n3921;
wire n3922;
wire n3923;
wire n3924;
wire n3925;
wire n3928;
wire n3929;
wire n3930;
wire n3931;
wire n3932;
wire n3933;
wire n3934;
wire n3935;
wire n3936;
wire n3937;
wire n3938;
wire n3939;
wire n3940;
wire n3941;
wire n3942;
wire n3943;
wire n3944;
wire n3945;
wire n3948;
wire n3949;
wire n3950;
wire n3951;
wire n3952;
wire n3953;
wire n3954;
wire n3955;
wire n3956;
wire n3957;
wire n3958;
wire n3959;
wire n3960;
wire n3963;
wire n3964;
wire n3965;
wire n3966;
wire n3967;
wire n3968;
wire n3969;
wire n3970;
wire n3971;
wire n3972;
wire n3973;
wire n3974;
wire n3975;
wire n3976;
wire n3977;
wire n3978;
wire n3979;
wire n3980;
wire n3981;
wire n3982;
wire n3983;
wire n3984;
wire n3985;
wire n3986;
wire n3987;
wire n3988;
wire n3991;
wire n3992;
wire n3993;
wire n3994;
wire n3995;
wire n3996;
wire n3997;
wire n3998;
wire n3999;
wire n4000;
wire n4001;
wire n4002;
wire n4003;
wire n4004;
wire n4005;
wire n4006;
wire n4007;
wire n4008;
wire n4011;
wire n4012;
wire n4013;
wire n4014;
wire n4015;
wire n4016;
wire n4017;
wire n4018;
wire n4019;
wire n4020;
wire n4021;
wire n4022;
wire n4023;
wire n4026;
wire n4027;
wire n4028;
wire n4029;
wire n4030;
wire n4031;
wire n4032;
wire n4033;
wire n4034;
wire n4035;
wire n4036;
wire n4037;
wire n4038;
wire n4039;
wire n4040;
wire n4041;
wire n4042;
wire n4043;
wire n4044;
wire n4045;
wire n4046;
wire n4047;
wire n4048;
wire n4049;
wire n4050;
wire n4051;
wire n4054;
wire n4055;
wire n4056;
wire n4057;
wire n4058;
wire n4059;
wire n4060;
wire n4061;
wire n4062;
wire n4063;
wire n4064;
wire n4065;
wire n4066;
wire n4067;
wire n4068;
wire n4069;
wire n4070;
wire n4071;
wire n4074;
wire n4075;
wire n4076;
wire n4077;
wire n4078;
wire n4079;
wire n4080;
wire n4081;
wire n4082;
wire n4083;
wire n4084;
wire n4085;
wire n4086;
wire n4089;
wire n4090;
wire n4091;
wire n4092;
wire n4093;
wire n4094;
wire n4095;
wire n4096;
wire n4097;
wire n4098;
wire n4099;
wire n4100;
wire n4101;
wire n4102;
wire n4103;
wire n4104;
wire n4105;
wire n4106;
wire n4107;
wire n4108;
wire n4109;
wire n4110;
wire n4111;
wire n4112;
wire n4113;
wire n4114;
wire n4117;
wire n4118;
wire n4119;
wire n4120;
wire n4121;
wire n4122;
wire n4123;
wire n4124;
wire n4125;
wire n4126;
wire n4127;
wire n4128;
wire n4129;
wire n4130;
wire n4131;
wire n4132;
wire n4133;
wire n4134;
wire n4137;
wire n4138;
wire n4139;
wire n4140;
wire n4141;
wire n4142;
wire n4143;
wire n4144;
wire n4145;
wire n4146;
wire n4147;
wire n4148;
wire n4149;
wire n4152;
wire n4153;
wire n4154;
wire n4155;
wire n4156;
wire n4157;
wire n4158;
wire n4159;
wire n4160;
wire n4161;
wire n4162;
wire n4163;
wire n4164;
wire n4165;
wire n4166;
wire n4167;
wire n4168;
wire n4169;
wire n4170;
wire n4171;
wire n4172;
wire n4173;
wire n4174;
wire n4175;
wire n4176;
wire n4177;
wire n4180;
wire n4181;
wire n4182;
wire n4183;
wire n4184;
wire n4185;
wire n4186;
wire n4187;
wire n4188;
wire n4189;
wire n4190;
wire n4191;
wire n4192;
wire n4193;
wire n4194;
wire n4195;
wire n4196;
wire n4197;
wire n4200;
wire n4201;
wire n4202;
wire n4203;
wire n4204;
wire n4205;
wire n4206;
wire n4207;
wire n4208;
wire n4209;
wire n4210;
wire n4211;
wire n4212;
wire n4215;
wire n4216;
wire n4217;
wire n4218;
wire n4219;
wire n4220;
wire n4221;
wire n4222;
wire n4223;
wire n4224;
wire n4225;
wire n4226;
wire n4227;
wire n4228;
wire n4229;
wire n4230;
wire n4231;
wire n4232;
wire n4233;
wire n4234;
wire n4235;
wire n4236;
wire n4237;
wire n4238;
wire n4239;
wire n4242;
wire n4243;
wire n4244;
wire n4245;
wire n4246;
wire n4247;
wire n4248;
wire n4249;
wire n4250;
wire n4251;
wire n4252;
wire n4253;
wire n4254;
wire n4255;
wire n4256;
wire n4257;
wire n4258;
wire n4259;
wire n4262;
wire n4263;
wire n4264;
wire n4265;
wire n4266;
wire n4267;
wire n4268;
wire n4269;
wire n4270;
wire n4271;
wire n4272;
wire n4273;
wire n4274;
wire n4277;
wire n4278;
wire n4279;
wire n4280;
wire n4281;
wire n4282;
wire n4283;
wire n4284;
wire n4285;
wire n4286;
wire n4287;
wire n4288;
wire n4289;
wire n4290;
wire n4291;
wire n4292;
wire n4293;
wire n4294;
wire n4295;
wire n4296;
wire n4297;
wire n4298;
wire n4299;
wire n4300;
wire n4301;
wire n4302;
wire n4303;
wire n4304;
wire n4305;
wire n4306;
wire n4307;
wire n4308;
wire n4309;
wire n4310;
wire n4311;
wire n4312;
wire n4313;
wire n4314;
wire n4315;
wire n4316;
wire n4317;
wire n4318;
wire n4319;
wire n4320;
wire n4321;
wire n4322;
wire n4323;
wire n4324;
wire n4325;
wire n4326;
wire n4327;
wire n4328;
wire n4329;
wire n4330;
wire n4331;
wire n4332;
wire n4333;
wire n4334;
wire n4335;
wire n4336;
wire n4337;
wire n4338;
wire n4339;
wire n4340;
wire n4341;
wire n4342;
wire n4343;
wire n4344;
wire n4345;
wire n4346;
wire n4347;
wire n4348;
wire n4349;
wire n4350;
wire n4351;
wire n4352;
wire n4353;
wire n4354;
wire n4355;
wire n4356;
wire n4357;
wire n4358;
wire n4359;
wire n4360;
wire n4361;
wire n4362;
wire n4363;
wire n4364;
wire n4365;
wire n4366;
wire n4367;
wire n4368;
wire n4369;
wire n4370;
wire n4371;
wire n4372;
wire n4373;
wire n4374;
wire n4375;
wire n4376;
wire n4377;
wire n4378;
wire n4379;
wire n4380;
wire n4381;
wire n4382;
wire n4383;
wire n4384;
wire n4385;
wire n4386;
wire n4387;
wire n4388;
wire n4389;
wire n4390;
wire n4391;
wire n4392;
wire n4395;
wire n4396;
wire n4397;
wire n4398;
wire n4399;
wire n4400;
wire n4401;
wire n4402;
wire n4403;
wire n4404;
wire n4405;
wire n4406;
wire n4407;
wire n4410;
wire n4411;
wire n4412;
wire n4413;
wire n4414;
wire n4415;
wire n4416;
wire n4417;
wire n4420;
wire n4421;
wire n4422;
wire n4423;
wire n4424;
wire n4425;
wire n4426;
wire n4427;
wire n4428;
wire n4429;
wire n4430;
wire n4431;
wire n4432;
wire n4433;
wire n4434;
wire n4435;
wire n4438;
wire n4439;
wire n4440;
wire n4441;
wire n4442;
wire n4443;
wire n4444;
wire n4445;
wire n4446;
wire n4447;
wire n4448;
wire n4449;
wire n4450;
wire n4453;
wire n4454;
wire n4455;
wire n4456;
wire n4457;
wire n4458;
wire n4459;
wire n4460;
wire n4463;
wire n4464;
wire n4465;
wire n4466;
wire n4467;
wire n4468;
wire n4469;
wire n4470;
wire n4471;
wire n4472;
wire n4473;
wire n4474;
wire n4475;
wire n4476;
wire n4477;
wire n4478;
wire n4481;
wire n4482;
wire n4483;
wire n4484;
wire n4485;
wire n4486;
wire n4487;
wire n4488;
wire n4489;
wire n4490;
wire n4491;
wire n4492;
wire n4493;
wire n4496;
wire n4497;
wire n4498;
wire n4499;
wire n4500;
wire n4501;
wire n4502;
wire n4503;
wire n4506;
wire n4507;
wire n4508;
wire n4509;
wire n4510;
wire n4511;
wire n4512;
wire n4513;
wire n4514;
wire n4515;
wire n4516;
wire n4517;
wire n4518;
wire n4519;
wire n4520;
wire n4521;
wire n4524;
wire n4525;
wire n4526;
wire n4527;
wire n4528;
wire n4529;
wire n4530;
wire n4531;
wire n4532;
wire n4533;
wire n4534;
wire n4535;
wire n4536;
wire n4539;
wire n4540;
wire n4541;
wire n4542;
wire n4543;
wire n4544;
wire n4545;
wire n4546;
wire n4549;
wire n4550;
wire n4551;
wire n4552;
wire n4553;
wire n4554;
wire n4555;
wire n4556;
wire n4557;
wire n4558;
wire n4559;
wire n4560;
wire n4561;
wire n4562;
wire n4563;
wire n4564;
wire n4567;
wire n4568;
wire n4569;
wire n4570;
wire n4571;
wire n4572;
wire n4573;
wire n4574;
wire n4575;
wire n4576;
wire n4577;
wire n4578;
wire n4579;
wire n4582;
wire n4583;
wire n4584;
wire n4585;
wire n4586;
wire n4587;
wire n4588;
wire n4589;
wire n4592;
wire n4593;
wire n4594;
wire n4595;
wire n4596;
wire n4597;
wire n4598;
wire n4599;
wire n4600;
wire n4601;
wire n4602;
wire n4603;
wire n4604;
wire n4605;
wire n4606;
wire n4607;
wire n4610;
wire n4611;
wire n4612;
wire n4613;
wire n4614;
wire n4615;
wire n4616;
wire n4617;
wire n4618;
wire n4619;
wire n4620;
wire n4621;
wire n4622;
wire n4625;
wire n4626;
wire n4627;
wire n4628;
wire n4629;
wire n4630;
wire n4631;
wire n4632;
wire n4635;
wire n4636;
wire n4637;
wire n4638;
wire n4639;
wire n4640;
wire n4641;
wire n4642;
wire n4643;
wire n4644;
wire n4645;
wire n4646;
wire n4647;
wire n4648;
wire n4649;
wire n4650;
wire n4653;
wire n4654;
wire n4655;
wire n4656;
wire n4657;
wire n4658;
wire n4659;
wire n4660;
wire n4661;
wire n4662;
wire n4663;
wire n4664;
wire n4665;
wire n4668;
wire n4669;
wire n4670;
wire n4671;
wire n4672;
wire n4673;
wire n4674;
wire n4675;
wire n4678;
wire n4679;
wire n4680;
wire n4681;
wire n4682;
wire n4683;
wire n4684;
wire n4685;
wire n4686;
wire n4687;
wire n4688;
wire n4689;
wire n4690;
wire n4691;
wire n4692;
wire n4695;
wire n4696;
wire n4697;
wire n4698;
wire n4699;
wire n4700;
wire n4701;
wire n4702;
wire n4703;
wire n4704;
wire n4705;
wire n4706;
wire n4707;
wire n4710;
wire n4711;
wire n4712;
wire n4713;
wire n4714;
wire n4715;
wire n4716;
wire n4717;
wire n4720;
wire n4721;
wire n4722;
wire n4723;
wire n4724;
wire n4725;
wire n4726;
wire n4727;
wire n4728;
wire n4729;
wire n4730;
wire n4731;
wire n4732;
wire n4733;
wire n4734;
wire n4735;
wire n4736;
wire n4737;
wire n4738;
wire n4739;
wire n4740;
wire n4741;
wire n4742;
wire n4743;
wire n4744;
wire n4745;
wire n4746;
wire n4747;
wire n4748;
wire n4749;
wire n4750;
wire n4751;
wire n4752;
wire n4753;
wire n4754;
wire n4755;
wire n4756;
wire n4757;
wire n4758;
wire n4759;
wire n4760;
wire n4761;
wire n4762;
wire n4763;
wire n4764;
wire n4765;
wire n4766;
wire n4767;
wire n4768;
wire n4769;
wire n4770;
wire n4771;
wire n4772;
wire n4773;
wire n4774;
wire n4775;
wire n4776;
wire n4777;
wire n4778;
wire n4779;
wire n4780;
wire n4781;
wire n4782;
wire n4783;
wire n4784;
wire n4785;
wire n4786;
wire n4787;
wire n4788;
wire n4789;
wire n4790;
wire n4791;
wire n4792;
wire n4793;
wire n4794;
wire n4795;
wire n4796;
wire n4797;
wire n4798;
wire n4799;
wire n4800;
wire n4801;
wire n4802;
wire n4803;
wire n4804;
wire n4805;
wire n4806;
wire n4807;
wire n4808;
wire n4809;
wire n4810;
wire n4811;
wire n4812;
wire n4813;
wire n4814;
wire n4815;
wire n4816;
wire n4817;
wire n4818;
wire n4819;
wire n4820;
wire n4821;
wire n4822;
wire n4823;
wire n4824;
wire n4825;
wire n4826;
wire n4827;
wire n4828;
wire n4829;
wire n4830;
wire n4831;
wire n4832;
wire n4833;
wire n4834;
wire n4835;
wire n4836;
wire n4837;
wire n4838;
wire n4839;
wire n4840;
wire n4841;
wire n4842;
wire n4843;
wire n4844;
wire n4845;
wire n4846;
wire n4847;
wire n4848;
wire n4849;
wire n4850;
wire n4851;
wire n4852;
wire n4853;
wire n4854;
wire n4855;
wire n4856;
wire n4857;
wire n4858;
wire n4859;
wire n4860;
wire n4861;
wire n4862;
wire n4863;
wire n4864;
wire n4865;
wire n4866;
wire n4867;
wire n4868;
wire n4869;
wire n4870;
wire n4871;
wire n4872;
wire n4873;
wire n4874;
wire n4875;
wire n4876;
wire n4877;
wire n4878;
wire n4879;
wire n4880;
wire n4881;
wire n4882;
wire n4883;
wire n4884;
wire n4885;
wire n4886;
wire n4887;
wire n4888;
wire n4889;
wire n4890;
wire n4891;
wire n4892;
wire n4893;
wire n4894;
wire n4895;
wire n4896;
wire n4897;
wire n4898;
wire n4899;
wire n4900;
wire n4901;
wire n4902;
wire n4903;
wire n4904;
wire n4905;
wire n4906;
wire n4907;
wire n4908;
wire n4909;
wire n4910;
wire n4911;
wire n4912;
wire n4913;
wire n4914;
wire n4915;
wire n4916;
wire n4917;
wire n4918;
wire n4919;
wire n4920;
wire n4921;
wire n4922;
wire n4923;
wire n4924;
wire n4925;
wire n4926;
wire n4927;
wire n4928;
wire n4929;
wire n4930;
wire n4931;
wire n4932;
wire n4933;
wire n4934;
wire n4935;
wire n4936;
wire n4937;
wire n4938;
wire n4939;
wire n4940;
wire n4941;
wire n4942;
wire n4943;
wire n4944;
wire n4945;
wire n4946;
wire n4947;
wire n4948;
wire n4949;
wire n4950;
wire n4951;
wire n4952;
wire n4953;
wire n4954;
wire n4955;
wire n4956;
wire n4957;
wire n4958;
wire n4959;
wire n4960;
wire n4961;
wire n4962;
wire n4963;
wire n4964;
wire n4966;
wire n4967;
wire n4968;
wire n4969;
wire n4970;
wire n4971;
wire n4972;
wire n4973;
wire n4974;
wire n4976;
wire n4977;
wire n4978;
wire n4980;
wire n4982;
wire n4983;
wire n4984;
wire n4985;
wire n4987;
wire n4989;
wire n4990;
wire n4991;
wire n4992;
wire n4994;
wire n4996;
wire n4997;
wire n4998;
wire n4999;
wire n5001;
wire n5003;
wire n5004;
wire n5005;
wire n5006;
wire n5007;
wire n5008;
wire n5009;
wire n5010;
wire n5011;
wire n5014;
wire n5015;
wire n5016;
wire n5017;
wire n5018;
wire n5019;
wire n5020;
wire n5021;
wire n5022;
wire n5023;
wire n5024;
wire n5025;
wire n5026;
wire n5028;
wire n5029;
wire n5030;
wire n5031;
wire n5033;
wire n5034;
wire n5035;
wire n5036;
wire n5038;
wire n5039;
wire n5040;
wire n5041;
wire n5042;
wire n5043;
wire n5045;
wire n5046;
wire n5048;
wire n5049;
wire n5051;
wire n5052;
wire n5054;
wire n5055;
wire n5056;
wire n5057;
wire n5060;
wire n5061;
wire n5063;
wire n5064;
wire n5066;
wire n5067;
wire n5069;
wire n5070;
wire n5071;
wire n5072;
wire n5074;
wire n5075;
wire n5077;
wire n5078;
wire n5079;
wire n5080;
wire n5082;
wire n5083;
wire n5084;
wire n5085;
wire n5086;
wire n5087;
wire n5090;
wire n5091;
wire n5093;
wire n5094;
wire n5096;
wire n5097;
wire n5099;
wire n5100;
wire n5101;
wire n5102;
wire n5104;
wire n5105;
wire n5107;
wire n5108;
wire n5110;
wire n5111;
wire n5113;
wire n5114;
wire n5115;
wire n5116;
wire n5119;
wire n5120;
wire n5122;
wire n5123;
wire n5125;
wire n5126;
wire n5128;
wire n5129;
wire n5130;
wire n5131;
wire n5133;
wire n5134;
wire n5136;
wire n5137;
wire n5139;
wire n5140;
wire n5143;
wire n5144;
wire n5145;
wire n5146;
wire n5147;
wire n5148;
wire n5149;
wire n5150;
wire n5151;
wire n5154;
wire n5155;
wire n5157;
wire n5158;
wire n5160;
wire n5161;
wire n5163;
wire n5164;
wire n5165;
wire n5166;
wire n5168;
wire n5169;
wire n5171;
wire n5172;
wire n5174;
wire n5175;
wire n5177;
wire n5178;
wire n5179;
wire n5180;
wire n5183;
wire n5184;
wire n5186;
wire n5187;
wire n5189;
wire n5190;
wire n5192;
wire n5193;
wire n5194;
wire n5195;
wire n5197;
wire n5198;
wire n5200;
wire n5201;
wire n5202;
wire n5203;
wire n5205;
wire n5206;
wire n5207;
wire n5208;
wire n5209;
wire n5210;
wire n5213;
wire n5214;
wire n5216;
wire n5217;
wire n5219;
wire n5220;
wire n5222;
wire n5223;
wire n5224;
wire n5225;
wire n5227;
wire n5228;
wire n5230;
wire n5231;
wire n5233;
wire n5234;
wire n5236;
wire n5237;
wire n5238;
wire n5239;
wire n5242;
wire n5243;
wire n5245;
wire n5246;
wire n5248;
wire n5249;
wire n5251;
wire n5252;
wire n5253;
wire n5254;
wire n5256;
wire n5257;
wire n5259;
wire n5260;
wire n5262;
wire n5263;
wire n5266;
wire n5267;
wire n5268;
wire n5269;
wire n5270;
wire n5271;
wire n5272;
wire n5273;
wire n5274;
wire n5277;
wire n5278;
wire n5280;
wire n5281;
wire n5283;
wire n5284;
wire n5286;
wire n5287;
wire n5288;
wire n5289;
wire n5291;
wire n5292;
wire n5294;
wire n5295;
wire n5297;
wire n5298;
wire n5300;
wire n5301;
wire n5302;
wire n5303;
wire n5306;
wire n5307;
wire n5309;
wire n5310;
wire n5312;
wire n5313;
wire n5315;
wire n5316;
wire n5317;
wire n5318;
wire n5320;
wire n5321;
wire n5323;
wire n5324;
wire n5325;
wire n5326;
wire n5328;
wire n5329;
wire n5330;
wire n5331;
wire n5332;
wire n5333;
wire n5336;
wire n5337;
wire n5339;
wire n5340;
wire n5342;
wire n5343;
wire n5345;
wire n5346;
wire n5347;
wire n5348;
wire n5350;
wire n5351;
wire n5353;
wire n5354;
wire n5356;
wire n5357;
wire n5359;
wire n5360;
wire n5361;
wire n5362;
wire n5365;
wire n5366;
wire n5368;
wire n5369;
wire n5371;
wire n5372;
wire n5374;
wire n5375;
wire n5376;
wire n5377;
wire n5379;
wire n5380;
wire n5382;
wire n5383;
wire n5385;
wire n5386;
wire n5389;
wire n5390;
wire n5391;
wire n5392;
wire n5393;
wire n5394;
wire n5395;
wire n5396;
wire n5397;
wire n5400;
wire n5401;
wire n5403;
wire n5404;
wire n5406;
wire n5407;
wire n5409;
wire n5410;
wire n5411;
wire n5412;
wire n5414;
wire n5415;
wire n5417;
wire n5418;
wire n5420;
wire n5421;
wire n5423;
wire n5424;
wire n5425;
wire n5426;
wire n5429;
wire n5430;
wire n5432;
wire n5433;
wire n5435;
wire n5436;
wire n5438;
wire n5439;
wire n5440;
wire n5441;
wire n5443;
wire n5444;
wire n5446;
wire n5447;
wire n5448;
wire n5449;
wire n5451;
wire n5452;
wire n5453;
wire n5454;
wire n5455;
wire n5456;
wire n5459;
wire n5460;
wire n5462;
wire n5463;
wire n5465;
wire n5466;
wire n5468;
wire n5469;
wire n5470;
wire n5471;
wire n5473;
wire n5474;
wire n5476;
wire n5477;
wire n5479;
wire n5480;
wire n5482;
wire n5483;
wire n5484;
wire n5485;
wire n5488;
wire n5489;
wire n5491;
wire n5492;
wire n5494;
wire n5495;
wire n5497;
wire n5498;
wire n5499;
wire n5500;
wire n5502;
wire n5503;
wire n5505;
wire n5506;
wire n5508;
wire n5509;
wire n5512;
wire n5513;
wire n5514;
wire n5515;
wire n5516;
wire n5517;
wire n5518;
wire n5519;
wire n5520;
wire n5523;
wire n5524;
wire n5526;
wire n5527;
wire n5529;
wire n5530;
wire n5532;
wire n5533;
wire n5534;
wire n5535;
wire n5537;
wire n5538;
wire n5540;
wire n5541;
wire n5543;
wire n5544;
wire n5546;
wire n5547;
wire n5548;
wire n5549;
wire n5552;
wire n5553;
wire n5555;
wire n5556;
wire n5558;
wire n5559;
wire n5561;
wire n5562;
wire n5563;
wire n5564;
wire n5566;
wire n5567;
wire n5569;
wire n5570;
wire n5571;
wire n5572;
wire n5574;
wire n5575;
wire n5576;
wire n5577;
wire n5578;
wire n5579;
wire n5582;
wire n5583;
wire n5585;
wire n5586;
wire n5588;
wire n5589;
wire n5591;
wire n5592;
wire n5593;
wire n5594;
wire n5596;
wire n5597;
wire n5599;
wire n5600;
wire n5602;
wire n5603;
wire n5605;
wire n5606;
wire n5607;
wire n5608;
wire n5611;
wire n5612;
wire n5614;
wire n5615;
wire n5617;
wire n5618;
wire n5620;
wire n5621;
wire n5622;
wire n5623;
wire n5625;
wire n5626;
wire n5628;
wire n5629;
wire n5631;
wire n5632;
wire n5635;
wire n5636;
wire n5637;
wire n5638;
wire n5639;
wire n5640;
wire n5641;
wire n5642;
wire n5643;
wire n5646;
wire n5647;
wire n5649;
wire n5650;
wire n5652;
wire n5653;
wire n5655;
wire n5656;
wire n5657;
wire n5658;
wire n5660;
wire n5661;
wire n5663;
wire n5664;
wire n5666;
wire n5667;
wire n5669;
wire n5670;
wire n5671;
wire n5672;
wire n5675;
wire n5676;
wire n5678;
wire n5679;
wire n5681;
wire n5682;
wire n5684;
wire n5685;
wire n5686;
wire n5687;
wire n5689;
wire n5690;
wire n5692;
wire n5693;
wire n5694;
wire n5695;
wire n5697;
wire n5698;
wire n5699;
wire n5700;
wire n5701;
wire n5702;
wire n5705;
wire n5706;
wire n5708;
wire n5709;
wire n5711;
wire n5712;
wire n5714;
wire n5715;
wire n5716;
wire n5717;
wire n5719;
wire n5720;
wire n5722;
wire n5723;
wire n5725;
wire n5726;
wire n5728;
wire n5729;
wire n5730;
wire n5731;
wire n5734;
wire n5735;
wire n5737;
wire n5738;
wire n5740;
wire n5741;
wire n5743;
wire n5744;
wire n5745;
wire n5746;
wire n5748;
wire n5749;
wire n5751;
wire n5752;
wire n5754;
wire n5755;
wire n5758;
wire n5759;
wire n5760;
wire n5761;
wire n5762;
wire n5763;
wire n5764;
wire n5765;
wire n5766;
wire n5769;
wire n5770;
wire n5772;
wire n5773;
wire n5775;
wire n5776;
wire n5778;
wire n5779;
wire n5780;
wire n5781;
wire n5783;
wire n5784;
wire n5786;
wire n5787;
wire n5789;
wire n5790;
wire n5792;
wire n5793;
wire n5794;
wire n5795;
wire n5798;
wire n5799;
wire n5801;
wire n5802;
wire n5804;
wire n5805;
wire n5807;
wire n5808;
wire n5809;
wire n5810;
wire n5812;
wire n5813;
wire n5815;
wire n5816;
wire n5817;
wire n5818;
wire n5820;
wire n5821;
wire n5822;
wire n5823;
wire n5824;
wire n5825;
wire n5828;
wire n5829;
wire n5831;
wire n5832;
wire n5834;
wire n5835;
wire n5837;
wire n5838;
wire n5839;
wire n5840;
wire n5842;
wire n5843;
wire n5845;
wire n5846;
wire n5848;
wire n5849;
wire n5851;
wire n5852;
wire n5853;
wire n5854;
wire n5857;
wire n5858;
wire n5860;
wire n5861;
wire n5863;
wire n5864;
wire n5866;
wire n5867;
wire n5868;
wire n5869;
wire n5871;
wire n5872;
wire n5874;
wire n5875;
wire n5877;
wire n5878;
wire n5881;
wire n5882;
wire n5883;
wire n5884;
wire n5885;
wire n5886;
wire n5887;
wire n5888;
wire n5891;
wire n5892;
wire n5894;
wire n5895;
wire n5897;
wire n5898;
wire n5900;
wire n5901;
wire n5902;
wire n5903;
wire n5905;
wire n5906;
wire n5908;
wire n5909;
wire n5911;
wire n5912;
wire n5914;
wire n5915;
wire n5916;
wire n5917;
wire n5920;
wire n5921;
wire n5923;
wire n5924;
wire n5926;
wire n5927;
wire n5929;
wire n5930;
wire n5931;
wire n5932;
wire n5934;
wire n5935;
wire n5937;
wire n5938;
wire n5939;
wire n5940;
wire n5942;
wire n5943;
wire n5944;
wire n5945;
wire n5946;
wire n5947;
wire n5950;
wire n5951;
wire n5953;
wire n5954;
wire n5956;
wire n5957;
wire n5959;
wire n5960;
wire n5961;
wire n5962;
wire n5964;
wire n5965;
wire n5967;
wire n5968;
wire n5970;
wire n5971;
wire n5973;
wire n5974;
wire n5975;
wire n5976;
wire n5979;
wire n5980;
wire n5982;
wire n5983;
wire n5985;
wire n5986;
wire n5988;
wire n5989;
wire n5990;
wire n5991;
wire n5993;
wire n5994;
wire n5996;
wire n5997;
wire n5999;
wire n6000;
wire n6003;
wire n6004;
wire n6005;
wire n6006;
wire n6007;
wire n6008;
wire n6009;
wire n6010;
wire n6011;
wire n6012;
wire n6013;
wire n6014;
wire n6015;
wire n6016;
wire n6017;
wire n6018;
wire n6019;
wire n6021;
wire n6023;
wire n6024;
wire n6025;
wire n6027;
wire n6029;
wire n6030;
wire n6031;
wire n6032;
wire n6034;
wire n6036;
wire n6037;
wire n6038;
wire n6039;
wire n6040;
wire n6041;
wire n6042;
wire n6043;
wire n6044;
wire n6045;
wire n6046;
wire n6047;
wire n6048;
wire n6049;
wire n6050;
wire n6051;
wire n6052;
wire n6053;
wire n6054;
wire n6055;
wire n6056;
wire n6057;
wire n6058;
wire n6059;
wire n6060;
wire n6061;
wire n6062;
wire n6063;
wire n6064;
wire n6065;
wire n6066;
wire n6067;
wire n6068;
wire n6069;
wire n6070;
wire n6071;
wire n6072;
wire n6073;
wire n6074;
wire n6075;
wire n6076;
wire n6077;
wire n6078;
wire n6079;
wire n6080;
wire n6082;
wire n6083;
wire n6084;
wire n6085;
wire n6086;
wire n6087;
wire n6088;
wire n6089;
wire n6090;
wire n6091;
wire n6092;
wire n6093;
wire n6094;
wire n6095;
wire n6096;
wire n6097;
wire n6098;
wire n6099;
wire n6100;
wire n6101;
wire n6102;
wire n6103;
wire n6104;
wire n6105;
wire n6106;
wire n6107;
wire n6108;
wire n6109;
wire n6110;
wire n6111;
wire n6112;
wire n6113;
wire n6114;
wire n6115;
wire n6116;
wire n6117;
wire n6118;
wire n6119;
wire n6120;
wire n6121;
wire n6122;
wire n6123;
wire n6125;
wire n6126;
wire n6127;
wire n6128;
wire n6129;
wire n6130;
wire n6131;
wire n6132;
wire n6133;
wire n6134;
wire n6135;
wire n6136;
wire n6137;
wire n6138;
wire n6139;
wire n6140;
wire n6141;
wire n6142;
wire n6143;
wire n6144;
wire n6145;
wire n6146;
wire n6147;
wire n6148;
wire n6149;
wire n6150;
wire n6151;
wire n6152;
wire n6153;
wire n6154;
wire n6155;
wire n6156;
wire n6157;
wire n6158;
wire n6159;
wire n6160;
wire n6161;
wire n6162;
wire n6163;
wire n6164;
wire n6165;
wire n6166;
wire n6167;
wire n6168;
wire n6169;
wire n6171;
wire n6172;
wire n6173;
wire n6174;
wire n6175;
wire n6176;
wire n6177;
wire n6178;
wire n6179;
wire n6180;
wire n6181;
wire n6182;
wire n6183;
wire n6184;
wire n6185;
wire n6186;
wire n6187;
wire n6188;
wire n6189;
wire n6190;
wire n6191;
wire n6192;
wire n6193;
wire n6194;
wire n6195;
wire n6196;
wire n6197;
wire n6198;
wire n6199;
wire n6200;
wire n6201;
wire n6202;
wire n6203;
wire n6204;
wire n6205;
wire n6206;
wire n6207;
wire n6208;
wire n6209;
wire n6210;
wire n6211;
wire n6212;
wire n6214;
wire n6215;
wire n6216;
wire n6217;
wire n6218;
wire n6219;
wire n6220;
wire n6221;
wire n6222;
wire n6223;
wire n6224;
wire n6225;
wire n6226;
wire n6227;
wire n6228;
wire n6229;
wire n6230;
wire n6231;
wire n6232;
wire n6233;
wire n6234;
wire n6235;
wire n6236;
wire n6237;
wire n6238;
wire n6239;
wire n6240;
wire n6241;
wire n6242;
wire n6243;
wire n6244;
wire n6245;
wire n6246;
wire n6247;
wire n6248;
wire n6249;
wire n6250;
wire n6251;
wire n6252;
wire n6253;
wire n6254;
wire n6255;
wire n6256;
wire n6257;
wire n6258;
wire n6260;
wire n6261;
wire n6262;
wire n6263;
wire n6264;
wire n6265;
wire n6266;
wire n6267;
wire n6268;
wire n6269;
wire n6270;
wire n6271;
wire n6272;
wire n6273;
wire n6274;
wire n6275;
wire n6276;
wire n6277;
wire n6278;
wire n6279;
wire n6280;
wire n6281;
wire n6282;
wire n6283;
wire n6284;
wire n6285;
wire n6286;
wire n6287;
wire n6288;
wire n6289;
wire n6290;
wire n6291;
wire n6292;
wire n6293;
wire n6294;
wire n6295;
wire n6296;
wire n6297;
wire n6298;
wire n6299;
wire n6300;
wire n6301;
wire n6303;
wire n6304;
wire n6305;
wire n6306;
wire n6307;
wire n6308;
wire n6309;
wire n6310;
wire n6311;
wire n6312;
wire n6313;
wire n6314;
wire n6315;
wire n6316;
wire n6317;
wire n6318;
wire n6319;
wire n6320;
wire n6321;
wire n6322;
wire n6323;
wire n6324;
wire n6325;
wire n6326;
wire n6327;
wire n6328;
wire n6329;
wire n6330;
wire n6331;
wire n6332;
wire n6333;
wire n6334;
wire n6335;
wire n6336;
wire n6337;
wire n6338;
wire n6339;
wire n6340;
wire n6341;
wire n6342;
wire n6343;
wire n6344;
wire n6345;
wire n6346;
wire n6347;
wire n6349;
wire n6350;
wire n6351;
wire n6352;
wire n6353;
wire n6354;
wire n6355;
wire n6356;
wire n6357;
wire n6358;
wire n6359;
wire n6360;
wire n6361;
wire n6362;
wire n6363;
wire n6364;
wire n6365;
wire n6366;
wire n6367;
wire n6368;
wire n6369;
wire n6370;
wire n6371;
wire n6372;
wire n6373;
wire n6374;
wire n6375;
wire n6376;
wire n6377;
wire n6378;
wire n6379;
wire n6380;
wire n6381;
wire n6382;
wire n6383;
wire n6384;
wire n6385;
wire n6386;
wire n6387;
wire n6388;
wire n6389;
wire n6390;
wire n6392;
wire n6393;
wire n6394;
wire n6395;
wire n6396;
wire n6397;
wire n6398;
wire n6399;
wire n6400;
wire n6401;
wire n6402;
wire n6403;
wire n6404;
wire n6405;
wire n6406;
wire n6407;
wire n6408;
wire n6409;
wire n6410;
wire n6411;
wire n6412;
wire n6413;
wire n6414;
wire n6415;
wire n6416;
wire n6417;
wire n6418;
wire n6419;
wire n6420;
wire n6421;
wire n6422;
wire n6423;
wire n6424;
wire n6425;
wire n6426;
wire n6427;
wire n6428;
wire n6429;
wire n6430;
wire n6431;
wire n6432;
wire n6433;
wire n6434;
wire n6435;
wire n6436;
wire n6438;
wire n6439;
wire n6440;
wire n6441;
wire n6442;
wire n6443;
wire n6444;
wire n6445;
wire n6446;
wire n6447;
wire n6448;
wire n6449;
wire n6450;
wire n6451;
wire n6452;
wire n6453;
wire n6454;
wire n6455;
wire n6456;
wire n6457;
wire n6458;
wire n6459;
wire n6460;
wire n6461;
wire n6462;
wire n6463;
wire n6464;
wire n6465;
wire n6466;
wire n6467;
wire n6468;
wire n6469;
wire n6470;
wire n6471;
wire n6472;
wire n6473;
wire n6474;
wire n6475;
wire n6476;
wire n6477;
wire n6478;
wire n6479;
wire n6481;
wire n6482;
wire n6483;
wire n6484;
wire n6485;
wire n6486;
wire n6487;
wire n6488;
wire n6489;
wire n6490;
wire n6491;
wire n6492;
wire n6493;
wire n6494;
wire n6495;
wire n6496;
wire n6497;
wire n6498;
wire n6499;
wire n6500;
wire n6501;
wire n6502;
wire n6503;
wire n6504;
wire n6505;
wire n6506;
wire n6507;
wire n6508;
wire n6509;
wire n6510;
wire n6511;
wire n6512;
wire n6513;
wire n6514;
wire n6515;
wire n6516;
wire n6517;
wire n6518;
wire n6519;
wire n6520;
wire n6521;
wire n6522;
wire n6523;
wire n6524;
wire n6525;
wire n6527;
wire n6528;
wire n6529;
wire n6530;
wire n6531;
wire n6532;
wire n6533;
wire n6534;
wire n6535;
wire n6536;
wire n6537;
wire n6538;
wire n6539;
wire n6540;
wire n6541;
wire n6542;
wire n6543;
wire n6544;
wire n6545;
wire n6546;
wire n6547;
wire n6548;
wire n6549;
wire n6550;
wire n6551;
wire n6552;
wire n6553;
wire n6554;
wire n6555;
wire n6556;
wire n6557;
wire n6558;
wire n6559;
wire n6560;
wire n6561;
wire n6562;
wire n6563;
wire n6564;
wire n6565;
wire n6566;
wire n6567;
wire n6568;
wire n6570;
wire n6571;
wire n6572;
wire n6573;
wire n6574;
wire n6575;
wire n6576;
wire n6577;
wire n6578;
wire n6579;
wire n6580;
wire n6581;
wire n6582;
wire n6583;
wire n6584;
wire n6585;
wire n6586;
wire n6587;
wire n6588;
wire n6589;
wire n6590;
wire n6591;
wire n6592;
wire n6593;
wire n6594;
wire n6595;
wire n6596;
wire n6597;
wire n6598;
wire n6599;
wire n6600;
wire n6601;
wire n6602;
wire n6603;
wire n6604;
wire n6605;
wire n6606;
wire n6607;
wire n6608;
wire n6609;
wire n6610;
wire n6611;
wire n6612;
wire n6613;
wire n6614;
wire n6616;
wire n6617;
wire n6618;
wire n6619;
wire n6620;
wire n6621;
wire n6622;
wire n6623;
wire n6624;
wire n6625;
wire n6626;
wire n6627;
wire n6628;
wire n6629;
wire n6630;
wire n6631;
wire n6632;
wire n6633;
wire n6634;
wire n6635;
wire n6636;
wire n6637;
wire n6638;
wire n6639;
wire n6640;
wire n6641;
wire n6642;
wire n6643;
wire n6644;
wire n6645;
wire n6646;
wire n6647;
wire n6648;
wire n6649;
wire n6650;
wire n6651;
wire n6652;
wire n6653;
wire n6654;
wire n6655;
wire n6656;
wire n6657;
wire n6659;
wire n6660;
wire n6661;
wire n6662;
wire n6663;
wire n6664;
wire n6665;
wire n6666;
wire n6667;
wire n6668;
wire n6669;
wire n6670;
wire n6671;
wire n6672;
wire n6673;
wire n6674;
wire n6675;
wire n6676;
wire n6677;
wire n6678;
wire n6679;
wire n6680;
wire n6681;
wire n6682;
wire n6683;
wire n6684;
wire n6685;
wire n6686;
wire n6687;
wire n6688;
wire n6689;
wire n6690;
wire n6691;
wire n6692;
wire n6693;
wire n6694;
wire n6695;
wire n6696;
wire n6697;
wire n6698;
wire n6699;
wire n6700;
wire n6701;
wire n6702;
wire n6704;
wire n6705;
wire n6706;
wire n6707;
wire n6708;
wire n6709;
wire n6710;
wire n6711;
wire n6712;
wire n6713;
wire n6714;
wire n6715;
wire n6716;
wire n6717;
wire n6718;
wire n6719;
wire n6720;
wire n6721;
wire n6722;
wire n6723;
wire n6724;
wire n6725;
wire n6726;
wire n6727;
wire n6728;
wire n6729;
wire n6730;
wire n6731;
wire n6732;
wire n6733;
wire n6734;
wire n6735;
wire n6736;
wire n6737;
wire n6738;
wire n6739;
wire n6740;
wire n6741;
wire n6742;
wire n6743;
wire n6744;
wire n6745;
wire n6747;
wire n6748;
wire n6749;
wire n6750;
wire n6751;
wire n6752;
wire n6753;
wire n6754;
wire n6755;
wire n6756;
wire n6757;
wire n6758;
wire n6759;
wire n6761;
wire n6763;
wire n6764;
wire n6765;
wire n6767;
wire n6769;
wire n6770;
wire n6771;
wire n6772;
wire n6774;
wire n6776;
wire n6777;
wire n6778;
wire n6779;
wire n6781;
wire n6783;
wire n6784;
wire n6785;
wire n6786;
wire n6788;
wire n6790;
wire n6791;
wire n6792;
wire n6793;
wire n6794;
wire n6795;
wire n6796;
wire n6797;
wire n6798;
wire n6799;
wire n6800;
wire n6803;
wire n6804;
wire n6806;
wire n6807;
wire n6809;
wire n6810;
wire n6812;
wire n6813;
wire n6814;
wire n6815;
wire n6817;
wire n6818;
wire n6820;
wire n6821;
wire n6822;
wire n6823;
wire n6825;
wire n6826;
wire n6827;
wire n6828;
wire n6829;
wire n6830;
wire n6833;
wire n6834;
wire n6836;
wire n6837;
wire n6839;
wire n6840;
wire n6842;
wire n6843;
wire n6844;
wire n6845;
wire n6847;
wire n6848;
wire n6850;
wire n6851;
wire n6853;
wire n6854;
wire n6856;
wire n6857;
wire n6859;
wire n6860;
wire n6861;
wire n6862;
wire n6863;
wire n6864;
wire n6865;
wire n6866;
wire n6867;
wire n6868;
wire n6869;
wire n6872;
wire n6873;
wire n6875;
wire n6876;
wire n6878;
wire n6879;
wire n6881;
wire n6882;
wire n6883;
wire n6884;
wire n6886;
wire n6887;
wire n6889;
wire n6890;
wire n6891;
wire n6892;
wire n6894;
wire n6895;
wire n6896;
wire n6897;
wire n6898;
wire n6899;
wire n6902;
wire n6903;
wire n6905;
wire n6906;
wire n6908;
wire n6909;
wire n6911;
wire n6912;
wire n6913;
wire n6914;
wire n6916;
wire n6917;
wire n6919;
wire n6920;
wire n6922;
wire n6923;
wire n6925;
wire n6926;
wire n6928;
wire n6929;
wire n6930;
wire n6931;
wire n6932;
wire n6933;
wire n6934;
wire n6935;
wire n6936;
wire n6937;
wire n6938;
wire n6941;
wire n6942;
wire n6944;
wire n6945;
wire n6947;
wire n6948;
wire n6950;
wire n6951;
wire n6952;
wire n6953;
wire n6955;
wire n6956;
wire n6958;
wire n6959;
wire n6960;
wire n6961;
wire n6963;
wire n6964;
wire n6965;
wire n6966;
wire n6967;
wire n6968;
wire n6971;
wire n6972;
wire n6974;
wire n6975;
wire n6977;
wire n6978;
wire n6980;
wire n6981;
wire n6982;
wire n6983;
wire n6985;
wire n6986;
wire n6988;
wire n6989;
wire n6991;
wire n6992;
wire n6994;
wire n6995;
wire n6997;
wire n6998;
wire n6999;
wire n7000;
wire n7001;
wire n7002;
wire n7003;
wire n7004;
wire n7005;
wire n7006;
wire n7007;
wire n7010;
wire n7011;
wire n7013;
wire n7014;
wire n7016;
wire n7017;
wire n7019;
wire n7020;
wire n7021;
wire n7022;
wire n7024;
wire n7025;
wire n7027;
wire n7028;
wire n7029;
wire n7030;
wire n7032;
wire n7033;
wire n7034;
wire n7035;
wire n7036;
wire n7037;
wire n7040;
wire n7041;
wire n7043;
wire n7044;
wire n7046;
wire n7047;
wire n7049;
wire n7050;
wire n7051;
wire n7052;
wire n7054;
wire n7055;
wire n7057;
wire n7058;
wire n7060;
wire n7061;
wire n7063;
wire n7064;
wire n7066;
wire n7067;
wire n7068;
wire n7069;
wire n7070;
wire n7071;
wire n7072;
wire n7073;
wire n7074;
wire n7075;
wire n7076;
wire n7079;
wire n7080;
wire n7082;
wire n7083;
wire n7085;
wire n7086;
wire n7088;
wire n7089;
wire n7090;
wire n7091;
wire n7093;
wire n7094;
wire n7096;
wire n7097;
wire n7098;
wire n7099;
wire n7101;
wire n7102;
wire n7103;
wire n7104;
wire n7105;
wire n7106;
wire n7109;
wire n7110;
wire n7112;
wire n7113;
wire n7115;
wire n7116;
wire n7118;
wire n7119;
wire n7120;
wire n7121;
wire n7123;
wire n7124;
wire n7126;
wire n7127;
wire n7129;
wire n7130;
wire n7132;
wire n7133;
wire n7135;
wire n7136;
wire n7137;
wire n7138;
wire n7139;
wire n7140;
wire n7141;
wire n7142;
wire n7143;
wire n7144;
wire n7145;
wire n7148;
wire n7149;
wire n7151;
wire n7152;
wire n7154;
wire n7155;
wire n7157;
wire n7158;
wire n7159;
wire n7160;
wire n7162;
wire n7163;
wire n7165;
wire n7166;
wire n7167;
wire n7168;
wire n7170;
wire n7171;
wire n7172;
wire n7173;
wire n7174;
wire n7175;
wire n7178;
wire n7179;
wire n7181;
wire n7182;
wire n7184;
wire n7185;
wire n7187;
wire n7188;
wire n7189;
wire n7190;
wire n7192;
wire n7193;
wire n7195;
wire n7196;
wire n7198;
wire n7199;
wire n7201;
wire n7202;
wire n7204;
wire n7205;
wire n7206;
wire n7207;
wire n7208;
wire n7209;
wire n7210;
wire n7211;
wire n7212;
wire n7213;
wire n7214;
wire n7217;
wire n7218;
wire n7220;
wire n7221;
wire n7223;
wire n7224;
wire n7226;
wire n7227;
wire n7228;
wire n7229;
wire n7231;
wire n7232;
wire n7234;
wire n7235;
wire n7236;
wire n7237;
wire n7239;
wire n7240;
wire n7241;
wire n7242;
wire n7243;
wire n7244;
wire n7247;
wire n7248;
wire n7250;
wire n7251;
wire n7253;
wire n7254;
wire n7256;
wire n7257;
wire n7258;
wire n7259;
wire n7261;
wire n7262;
wire n7264;
wire n7265;
wire n7267;
wire n7268;
wire n7270;
wire n7271;
wire n7273;
wire n7274;
wire n7275;
wire n7276;
wire n7277;
wire n7278;
wire n7279;
wire n7280;
wire n7281;
wire n7282;
wire n7285;
wire n7286;
wire n7288;
wire n7289;
wire n7291;
wire n7292;
wire n7294;
wire n7295;
wire n7296;
wire n7297;
wire n7299;
wire n7300;
wire n7302;
wire n7303;
wire n7304;
wire n7305;
wire n7307;
wire n7308;
wire n7309;
wire n7310;
wire n7311;
wire n7312;
wire n7315;
wire n7316;
wire n7318;
wire n7319;
wire n7321;
wire n7322;
wire n7324;
wire n7325;
wire n7326;
wire n7327;
wire n7329;
wire n7330;
wire n7332;
wire n7333;
wire n7335;
wire n7336;
wire n7338;
wire n7339;
wire n7341;
wire n7342;
wire n7343;
wire n7344;
wire n7345;
wire n7346;
wire n7347;
wire n7348;
wire n7349;
wire n7350;
wire n7351;
wire n7352;
wire n7353;
wire n7354;
wire n7355;
wire n7356;
wire n7357;
wire n7358;
wire n7359;
wire n7360;
wire n7361;
wire n7362;
wire n7363;
wire n7364;
wire n7365;
wire n7366;
wire n7367;
wire n7368;
wire n7369;
wire n7370;
wire n7371;
wire n7372;
wire n7373;
wire n7374;
wire n7375;
wire n7376;
wire n7377;
wire n7378;
wire n7379;
wire n7380;
wire n7381;
wire n7382;
wire n7383;
wire n7384;
wire n7385;
wire n7386;
wire n7387;
wire n7388;
wire n7389;
wire n7390;
wire n7391;
wire n7392;
wire n7393;
wire n7394;
wire n7395;
wire n7396;
wire n7397;
wire n7398;
wire n7399;
wire n7400;
wire n7401;
wire n7402;
wire n7403;
wire n7404;
wire n7405;
wire n7406;
wire n7407;
wire n7408;
wire n7409;
wire n7410;
wire n7411;
wire n7412;
wire n7413;
wire n7414;
wire n7415;
wire n7416;
wire n7417;
wire n7418;
wire n7419;
wire n7420;
wire n7421;
wire n7422;
wire n7423;
wire n7424;
wire n7425;
wire n7426;
wire n7427;
wire n7428;
wire n7429;
wire n7430;
wire n7431;
wire n7432;
wire n7433;
wire n7434;
wire n7435;
wire n7436;
wire n7437;
wire n7438;
wire n7439;
wire n7440;
wire n7441;
wire n7442;
wire n7443;
wire n7444;
wire n7445;
wire n7446;
wire n7447;
wire n7448;
wire n7449;
wire n7450;
wire n7451;
wire n7452;
wire n7453;
wire n7454;
wire n7455;
wire n7456;
wire n7457;
wire n7458;
wire n7459;
wire n7460;
wire n7461;
wire n7462;
wire n7463;
wire n7464;
wire n7465;
wire n7466;
wire n7467;
wire n7468;
wire n7469;
wire n7470;
wire n7471;
wire n7472;
wire n7473;
wire n7474;
wire n7475;
wire n7476;
wire n7477;
wire n7478;
wire n7479;
wire n7480;
wire n7481;
wire n7482;
wire n7483;
wire n7484;
wire n7485;
wire n7486;
wire n7487;
wire n7488;
wire n7489;
wire n7490;
wire n7491;
wire n7492;
wire n7493;
wire n7494;
wire n7495;
wire n7496;
wire n7497;
wire n7498;
wire n7499;
wire n7500;
wire n7501;
wire n7502;
wire n7503;
wire n7504;
wire n7505;
wire n7506;
wire n7507;
wire n7508;
wire n7509;
wire n7510;
wire n7511;
wire n7512;
wire n7513;
wire n7514;
wire n7515;
wire n7516;
wire n7517;
wire n7518;
wire n7519;
wire n7520;
wire n7521;
wire n7522;
wire n7523;
wire n7524;
wire n7525;
wire n7526;
wire n7527;
wire n7528;
wire n7529;
wire n7530;
wire n7531;
wire n7532;
wire n7533;
wire n7534;
wire n7535;
wire n7536;
wire n7537;
wire n7538;
wire n7539;
wire n7540;
wire n7541;
wire n7542;
wire n7543;
wire n7544;
wire n7545;
wire n7546;
wire n7547;
wire n7548;
wire n7549;
wire n7550;
wire n7551;
wire n7552;
wire n7553;
wire n7554;
wire n7555;
wire n7556;
wire n7557;
wire n7558;
wire n7559;
wire n7560;
wire n7561;
wire n7562;
wire n7563;
wire n7564;
wire n7565;
wire n7566;
wire n7567;
wire n7568;
wire n7569;
wire n7570;
wire n7571;
wire n7572;
wire n7573;
wire n7574;
wire n7575;
wire n7576;
wire n7577;
wire n7578;
wire n7579;
wire n7580;
wire n7581;
wire n7582;
wire n7583;
wire n7584;
wire n7585;
wire n7586;
wire n7587;
wire n7588;
wire n7589;
wire n7590;
wire n7591;
wire n7592;
wire n7593;
wire n7594;
wire n7595;
wire n7596;
wire n7597;
wire n7598;
wire n7599;
wire n7600;
wire n7601;
wire n7602;
wire n7603;
wire n7604;
wire n7605;
wire n7606;
wire n7607;
wire n7608;
wire n7609;
wire n7610;
wire n7611;
wire n7612;
wire n7613;
wire n7614;
wire n7615;
wire n7616;
wire n7617;
wire n7618;
wire n7619;
wire n7620;
wire n7621;
wire n7622;
wire n7623;
wire n7624;
wire n7625;
wire n7626;
wire n7627;
wire n7628;
wire n7629;
wire n7630;
wire n7631;
wire n7632;
wire n7633;
wire n7634;
wire n7635;
wire n7636;
wire n7637;
wire n7638;
wire n7639;
wire n7640;
wire n7641;
wire n7642;
wire n7643;
wire n7645;
wire n7647;
wire n7648;
wire n7649;
wire n7650;
wire n7651;
wire n7652;
wire n7654;
wire n7656;
wire n7657;
wire n7658;
wire n7659;
wire n7660;
wire n7661;
wire n7662;
wire n7663;
wire n7664;
wire n7665;
wire n7666;
wire n7667;
wire n7668;
wire n7670;
wire n7672;
wire n7673;
wire n7674;
wire n7675;
wire n7676;
wire n7677;
wire n7679;
wire n7681;
wire n7682;
wire n7683;
wire n7684;
wire n7686;
wire n7688;
wire n7689;
wire n7690;
wire n7691;
wire n7693;
wire n7695;
wire n7696;
wire n7697;
wire n7698;
wire n7699;
wire n7700;
wire n7701;
wire n7702;
wire n7703;
wire n7704;
wire n7705;
wire n7706;
wire n7707;
wire n7709;
wire n7711;
wire n7712;
wire n7713;
wire n7714;
wire n7715;
wire n7716;
wire n7718;
wire n7720;
wire n7721;
wire n7722;
wire n7723;
wire n7724;
wire n7725;
wire n7726;
wire n7727;
wire n7728;
wire n7729;
wire n7730;
wire n7731;
wire n7732;
wire n7733;
wire n7734;
wire n7735;
wire n7736;
wire n7737;
wire n7738;
wire n7739;
wire n7740;
wire n7741;
wire n7742;
wire n7743;
wire n7744;
wire n7745;
wire n7746;
wire n7747;
wire n7748;
wire n7749;
wire n7750;
wire n7751;
wire n7752;
wire n7753;
wire n7754;
wire n7755;
wire n7756;
wire n7757;
wire n7758;
wire n7759;
wire n7760;
wire n7761;
wire n7762;
wire n7763;
wire n7764;
wire n7765;
wire n7766;
wire n7767;
wire n7768;
wire n7769;
wire n7770;
wire n7771;
wire n7772;
wire n7773;
wire n7774;
wire n7775;
wire n7776;
wire n7777;
wire n7778;
wire n7779;
wire n7780;
wire n7781;
wire n7782;
wire n7783;
wire n7784;
wire n7785;
wire n7786;
wire n7787;
wire n7788;
wire n7789;
wire n7790;
wire n7791;
wire n7792;
wire n7793;
wire n7794;
wire n7795;
wire n7796;
wire n7797;
wire n7798;
wire n7799;
wire n7800;
wire n7801;
wire n7802;
wire n7803;
wire n7804;
wire n7805;
wire n7806;
wire n7807;
wire n7808;
wire n7809;
wire n7810;
wire n7811;
wire n7812;
wire n7813;
wire n7814;
wire n7815;
wire n7816;
wire n7817;
wire n7818;
wire n7819;
wire n7820;
wire n7821;
wire n7822;
wire n7823;
wire n7824;
wire n7825;
wire n7826;
wire n7827;
wire n7828;
wire n7829;
wire n7830;
wire n7831;
wire n7832;
wire n7833;
wire n7834;
wire n7835;
wire n7836;
wire n7837;
wire n7838;
wire n7839;
wire n7840;
wire n7841;
wire n7842;
wire n7843;
wire n7844;
wire n7845;
wire n7846;
wire n7847;
wire n7848;
wire n7849;
wire n7850;
wire n7851;
wire n7852;
wire n7853;
wire n7854;
wire n7855;
wire n7856;
wire n7857;
wire n7858;
wire n7859;
wire n7860;
wire n7861;
wire n7862;
wire n7863;
wire n7864;
wire n7865;
wire n7866;
wire n7867;
wire n7868;
wire n7869;
wire n7870;
wire n7871;
wire n7872;
wire n7873;
wire n7874;
wire n7875;
wire n7876;
wire n7877;
wire n7878;
wire n7879;
wire n7880;
wire n7881;
wire n7882;
wire n7883;
wire n7884;
wire n7886;
wire n7887;
wire n7889;
wire n7890;
wire n7891;
wire n7892;
wire n7893;
wire n7894;
wire n7895;
wire n7896;
wire n7897;
wire n7898;
wire n7899;
wire n7900;
wire n7901;
wire n7902;
wire n7903;
wire n7904;
wire n7905;
wire n7906;
wire n7907;
wire n7908;
wire n7909;
wire n7910;
wire n7911;
wire n7912;
wire n7913;
wire n7914;
wire n7915;
wire n7916;
wire n7917;
wire n7918;
wire n7919;
wire n7920;
wire n7921;
wire n7922;
wire n7923;
wire n7924;
wire n7925;
wire n7926;
wire n7927;
wire n7928;
wire n7929;
wire n7930;
wire n7931;
wire n7932;
wire n7933;
wire n7934;
wire n7935;
wire n7936;
wire n7937;
wire n7938;
wire n7939;
wire n7940;
wire n7941;
wire n7942;
wire n7943;
wire n7944;
wire n7945;
wire n7946;
wire n7947;
wire n7948;
wire n7949;
wire n7950;
wire n7951;
wire n7952;
wire n7953;
wire n7954;
wire n7955;
wire n7956;
wire n7957;
wire n7958;
wire n7959;
wire n7960;
wire n7961;
wire n7962;
wire n7963;
wire n7964;
wire n7965;
wire n7966;
wire n7967;
wire n7968;
wire n7969;
wire n7970;
wire n7971;
wire n7972;
wire n7973;
wire n7974;
wire n7975;
wire n7976;
wire n7977;
wire n7978;
wire n7979;
wire n7980;
wire n7981;
wire n7982;
wire n7983;
wire n7984;
wire n7985;
wire n7986;
wire n7987;
wire n7988;
wire n7989;
wire n7990;
wire n7991;
wire n7992;
wire n7993;
wire n7994;
wire n7995;
wire n7996;
wire n7998;
wire n7999;
wire n8001;
wire n8002;
wire n8003;
wire n8004;
wire n8005;
wire n8006;
wire n8007;
wire n8008;
wire n8009;
wire n8010;
wire n8011;
wire n8012;
wire n8013;
wire n8014;
wire n8015;
wire n8016;
wire n8017;
wire n8018;
wire n8019;
wire n8020;
wire n8021;
wire n8022;
wire n8023;
wire n8024;
wire n8025;
wire n8026;
wire n8027;
wire n8028;
wire n8029;
wire n8030;
wire n8031;
wire n8032;
wire n8033;
wire n8034;
wire n8035;
wire n8036;
wire n8037;
wire n8038;
wire n8039;
wire n8040;
wire n8041;
wire n8042;
wire n8043;
wire n8044;
wire n8045;
wire n8046;
wire n8047;
wire n8048;
wire n8049;
wire n8050;
wire n8051;
wire n8052;
wire n8053;
wire n8054;
wire n8055;
wire n8056;
wire n8057;
wire n8058;
wire n8059;
wire n8060;
wire n8061;
wire n8062;
wire n8063;
wire n8064;
wire n8065;
wire n8066;
wire n8067;
wire n8068;
wire n8069;
wire n8070;
wire n8071;
wire n8072;
wire n8073;
wire n8074;
wire n8075;
wire n8076;
wire n8077;
wire n8078;
wire n8079;
wire n8080;
wire n8081;
wire n8082;
wire n8083;
wire n8084;
wire n8085;
wire n8086;
wire n8087;
wire n8088;
wire n8089;
wire n8090;
wire n8091;
wire n8092;
wire n8093;
wire n8094;
wire n8095;
wire n8096;
wire n8097;
wire n8098;
wire n8099;
wire n8100;
wire n8101;
wire n8102;
wire n8103;
wire n8104;
wire n8105;
wire n8106;
wire n8107;
wire n8108;
wire n8110;
wire n8111;
wire n8113;
wire n8114;
wire n8115;
wire n8116;
wire n8117;
wire n8118;
wire n8119;
wire n8120;
wire n8121;
wire n8122;
wire n8123;
wire n8124;
wire n8125;
wire n8126;
wire n8127;
wire n8128;
wire n8129;
wire n8130;
wire n8131;
wire n8132;
wire n8133;
wire n8134;
wire n8135;
wire n8136;
wire n8137;
wire n8138;
wire n8139;
wire n8140;
wire n8141;
wire n8142;
wire n8143;
wire n8144;
wire n8145;
wire n8146;
wire n8147;
wire n8148;
wire n8149;
wire n8150;
wire n8151;
wire n8152;
wire n8153;
wire n8154;
wire n8155;
wire n8156;
wire n8157;
wire n8158;
wire n8159;
wire n8160;
wire n8161;
wire n8162;
wire n8163;
wire n8164;
wire n8165;
wire n8166;
wire n8167;
wire n8168;
wire n8169;
wire n8170;
wire n8171;
wire n8172;
wire n8173;
wire n8174;
wire n8175;
wire n8176;
wire n8177;
wire n8178;
wire n8179;
wire n8180;
wire n8181;
wire n8182;
wire n8183;
wire n8184;
wire n8185;
wire n8186;
wire n8187;
wire n8188;
wire n8189;
wire n8190;
wire n8191;
wire n8192;
wire n8193;
wire n8194;
wire n8195;
wire n8196;
wire n8197;
wire n8198;
wire n8199;
wire n8200;
wire n8201;
wire n8202;
wire n8203;
wire n8204;
wire n8205;
wire n8206;
wire n8207;
wire n8208;
wire n8209;
wire n8210;
wire n8211;
wire n8212;
wire n8213;
wire n8214;
wire n8215;
wire n8216;
wire n8217;
wire n8218;
wire n8219;
wire n8220;
wire n8222;
wire n8223;
wire n8225;
wire n8226;
wire n8227;
wire n8228;
wire n8229;
wire n8230;
wire n8231;
wire n8232;
wire n8233;
wire n8234;
wire n8235;
wire n8236;
wire n8237;
wire n8238;
wire n8239;
wire n8240;
wire n8241;
wire n8242;
wire n8243;
wire n8244;
wire n8245;
wire n8246;
wire n8247;
wire n8248;
wire n8249;
wire n8250;
wire n8251;
wire n8252;
wire n8253;
wire n8254;
wire n8255;
wire n8256;
wire n8257;
wire n8258;
wire n8259;
wire n8260;
wire n8261;
wire n8262;
wire n8263;
wire n8264;
wire n8265;
wire n8266;
wire n8267;
wire n8268;
wire n8269;
wire n8270;
wire n8271;
wire n8272;
wire n8273;
wire n8274;
wire n8275;
wire n8276;
wire n8277;
wire n8278;
wire n8279;
wire n8280;
wire n8281;
wire n8282;
wire n8283;
wire n8284;
wire n8285;
wire n8286;
wire n8287;
wire n8288;
wire n8289;
wire n8290;
wire n8291;
wire n8292;
wire n8293;
wire n8294;
wire n8295;
wire n8296;
wire n8297;
wire n8298;
wire n8299;
wire n8300;
wire n8301;
wire n8302;
wire n8303;
wire n8304;
wire n8305;
wire n8306;
wire n8307;
wire n8308;
wire n8309;
wire n8310;
wire n8311;
wire n8312;
wire n8313;
wire n8314;
wire n8315;
wire n8316;
wire n8317;
wire n8318;
wire n8319;
wire n8320;
wire n8321;
wire n8322;
wire n8323;
wire n8324;
wire n8325;
wire n8326;
wire n8327;
wire n8328;
wire n8330;
wire n8331;
wire n8333;
wire n8334;
wire n8335;
wire n8336;
wire n8337;
wire n8338;
wire n8339;
wire n8340;
wire n8341;
wire n8342;
wire n8343;
wire n8344;
wire n8345;
wire n8346;
wire n8347;
wire n8348;
wire n8349;
wire n8350;
wire n8351;
wire n8352;
wire n8353;
wire n8354;
wire n8355;
wire n8356;
wire n8357;
wire n8358;
wire n8359;
wire n8360;
wire n8361;
wire n8362;
wire n8363;
wire n8364;
wire n8365;
wire n8366;
wire n8367;
wire n8368;
wire n8369;
wire n8370;
wire n8371;
wire n8372;
wire n8373;
wire n8374;
wire n8375;
wire n8376;
wire n8377;
wire n8378;
wire n8379;
wire n8380;
wire n8381;
wire n8382;
wire n8383;
wire n8384;
wire n8385;
wire n8386;
wire n8387;
wire n8388;
wire n8389;
wire n8390;
wire n8391;
wire n8392;
wire n8393;
wire n8394;
wire n8395;
wire n8396;
wire n8397;
wire n8398;
wire n8399;
wire n8400;
wire n8401;
wire n8402;
wire n8403;
wire n8404;
wire n8405;
wire n8406;
wire n8407;
wire n8408;
wire n8409;
wire n8410;
wire n8411;
wire n8412;
wire n8413;
wire n8414;
wire n8415;
wire n8416;
wire n8417;
wire n8418;
wire n8419;
wire n8420;
wire n8421;
wire n8422;
wire n8423;
wire n8424;
wire n8425;
wire n8426;
wire n8427;
wire n8428;
wire n8429;
wire n8430;
wire n8431;
wire n8432;
wire n8433;
wire n8434;
wire n8435;
wire n8436;
wire n8438;
wire n8439;
wire n8441;
wire n8442;
wire n8443;
wire n8444;
wire n8445;
wire n8446;
wire n8447;
wire n8448;
wire n8449;
wire n8450;
wire n8451;
wire n8452;
wire n8453;
wire n8454;
wire n8455;
wire n8456;
wire n8457;
wire n8458;
wire n8459;
wire n8460;
wire n8461;
wire n8462;
wire n8463;
wire n8464;
wire n8465;
wire n8466;
wire n8467;
wire n8468;
wire n8469;
wire n8470;
wire n8471;
wire n8472;
wire n8473;
wire n8474;
wire n8475;
wire n8476;
wire n8477;
wire n8478;
wire n8479;
wire n8480;
wire n8481;
wire n8482;
wire n8483;
wire n8484;
wire n8485;
wire n8486;
wire n8487;
wire n8488;
wire n8489;
wire n8490;
wire n8491;
wire n8492;
wire n8493;
wire n8494;
wire n8495;
wire n8496;
wire n8497;
wire n8498;
wire n8499;
wire n8500;
wire n8501;
wire n8502;
wire n8503;
wire n8504;
wire n8505;
wire n8506;
wire n8507;
wire n8508;
wire n8509;
wire n8510;
wire n8511;
wire n8512;
wire n8513;
wire n8514;
wire n8515;
wire n8516;
wire n8517;
wire n8518;
wire n8519;
wire n8520;
wire n8521;
wire n8522;
wire n8523;
wire n8524;
wire n8525;
wire n8526;
wire n8527;
wire n8528;
wire n8529;
wire n8530;
wire n8531;
wire n8532;
wire n8533;
wire n8534;
wire n8535;
wire n8536;
wire n8537;
wire n8538;
wire n8539;
wire n8540;
wire n8541;
wire n8542;
wire n8543;
wire n8545;
wire n8546;
wire n8548;
wire n8549;
wire n8550;
wire n8551;
wire n8552;
wire n8553;
wire n8554;
wire n8555;
wire n8556;
wire n8557;
wire n8558;
wire n8559;
wire n8560;
wire n8561;
wire n8562;
wire n8563;
wire n8564;
wire n8565;
wire n8566;
wire n8567;
wire n8568;
wire n8569;
wire n8570;
wire n8571;
wire n8572;
wire n8573;
wire n8574;
wire n8575;
wire n8576;
wire n8577;
wire n8578;
wire n8579;
wire n8580;
wire n8581;
wire n8582;
wire n8583;
wire n8584;
wire n8585;
wire n8586;
wire n8587;
wire n8588;
wire n8589;
wire n8590;
wire n8591;
wire n8592;
wire n8593;
wire n8594;
wire n8595;
wire n8596;
wire n8597;
wire n8598;
wire n8599;
wire n8600;
wire n8601;
wire n8602;
wire n8603;
wire n8604;
wire n8605;
wire n8606;
wire n8607;
wire n8608;
wire n8609;
wire n8610;
wire n8611;
wire n8612;
wire n8613;
wire n8614;
wire n8615;
wire n8616;
wire n8617;
wire n8618;
wire n8619;
wire n8620;
wire n8621;
wire n8622;
wire n8623;
wire n8624;
wire n8625;
wire n8626;
wire n8627;
wire n8628;
wire n8629;
wire n8630;
wire n8631;
wire n8632;
wire n8633;
wire n8634;
wire n8635;
wire n8636;
wire n8637;
wire n8638;
wire n8639;
wire n8640;
wire n8641;
wire n8642;
wire n8643;
wire n8644;
wire n8645;
wire n8646;
wire n8647;
wire n8648;
wire n8649;
wire n8650;
wire n8651;
wire n8652;
wire n8653;
wire n8654;
wire n8655;
wire n8656;
wire n8657;
wire n8658;
wire n8659;
wire n8660;
wire n8661;
wire n8662;
wire n8663;
wire n8664;
wire n8665;
wire n8666;
wire n8667;
wire n8668;
wire n8669;
wire n8670;
wire n8671;
wire n8672;
wire n8673;
wire n8674;
wire n8675;
wire n8676;
wire n8677;
wire n8678;
wire n8679;
wire n8680;
wire n8681;
wire n8682;
wire n8683;
wire n8684;
wire n8685;
wire n8686;
wire n8687;
wire n8688;
wire n8689;
wire n8690;
wire n8691;
wire n8692;
wire n8693;
wire n8694;
wire n8695;
wire n8696;
wire n8697;
wire n8698;
wire n8699;
wire n8700;
wire n8701;
wire n8702;
wire n8703;
wire n8704;
wire n8705;
wire n8706;
wire n8707;
wire n8708;
wire n8709;
wire n8710;
wire n8711;
wire n8712;
wire n8713;
wire n8714;
wire n8715;
wire n8716;
wire n8717;
wire n8718;
wire n8719;
wire n8720;
wire n8721;
wire n8722;
wire n8723;
wire n8724;
wire n8725;
wire n8726;
wire n8727;
wire n8728;
wire n8729;
wire n8730;
wire n8731;
wire n8732;
wire n8733;
wire n8734;
wire n8735;
wire n8736;
wire n8737;
wire n8738;
wire n8739;
wire n8740;
wire n8741;
wire n8742;
wire n8743;
wire n8744;
wire n8745;
wire n8746;
wire n8747;
wire n8748;
wire n8749;
wire n8750;
wire n8751;
wire n8752;
wire n8753;
wire n8754;
wire n8755;
wire n8756;
wire n8757;
wire n8758;
wire n8759;
wire n8760;
wire n8761;
wire n8762;
wire n8763;
wire n8764;
wire n8765;
wire n8766;
wire n8767;
wire n8768;
wire n8769;
wire n8770;
wire n8771;
wire n8772;
wire n8773;
wire n8774;
wire n8775;
wire n8776;
wire n8777;
wire n8778;
wire n8779;
wire n8780;
wire n8781;
wire n8782;
wire n8783;
wire n8784;
wire n8785;
wire n8786;
wire n8787;
wire n8788;
wire n8789;
wire n8790;
wire n8791;
wire n8792;
wire n8793;
wire n8794;
wire n8795;
wire n8796;
wire n8797;
wire n8798;
wire n8799;
wire n8800;
wire n8801;
wire n8802;
wire n8803;
wire n8804;
wire n8805;
wire n8806;
wire n8807;
wire n8808;
wire n8809;
wire n8810;
wire n8811;
wire n8812;
wire n8813;
wire n8814;
wire n8815;
wire n8816;
wire n8817;
wire n8818;
wire n8819;
wire n8820;
wire n8821;
wire n8822;
wire n8823;
wire n8824;
wire n8825;
wire n8826;
wire n8827;
wire n8828;
wire n8829;
wire n8830;
wire n8831;
wire n8832;
wire n8833;
wire n8834;
wire n8835;
wire n8836;
wire n8837;
wire n8838;
wire n8839;
wire n8840;
wire n8841;
wire n8842;
wire n8843;
wire n8844;
wire n8845;
wire n8846;
wire n8847;
wire n8848;
wire n8849;
wire n8850;
wire n8851;
wire n8852;
wire n8853;
wire n8854;
wire n8855;
wire n8856;
wire n8857;
wire n8858;
wire n8859;
wire n8860;
wire n8861;
wire n8862;
wire n8863;
wire n8864;
wire n8865;
wire n8866;
wire n8867;
wire n8868;
wire n8869;
wire n8870;
wire n8871;
wire n8872;
wire n8873;
wire n8874;
wire n8875;
wire n8876;
wire n8877;
wire n8878;
wire n8879;
wire n8880;
wire n8881;
wire n8882;
wire n8883;
wire n8884;
wire n8885;
wire n8886;
wire n8887;
wire n8888;
wire n8889;
wire n8890;
wire n8891;
wire n8892;
wire n8893;
wire n8894;
wire n8895;
wire n8896;
wire n8897;
wire n8898;
wire n8899;
wire n8900;
wire n8901;
wire n8902;
wire n8903;
wire n8904;
wire n8905;
wire n8906;
wire n8907;
wire n8908;
wire n8909;
wire n8910;
wire n8911;
wire n8912;
wire n8913;
wire n8914;
wire n8915;
wire n8916;
wire n8917;
wire n8918;
wire n8919;
wire n8920;
wire n8921;
wire n8922;
wire n8923;
wire n8924;
wire n8925;
wire n8926;
wire n8927;
wire n8928;
wire n8929;
wire n8930;
wire n8931;
wire n8932;
wire n8933;
wire n8934;
wire n8935;
wire n8936;
wire n8937;
wire n8938;
wire n8939;
wire n8940;
wire n8941;
wire n8942;
wire n8943;
wire n8944;
wire n8945;
wire n8946;
wire n8947;
wire n8948;
wire n8949;
wire n8950;
wire n8951;
wire n8952;
wire n8953;
wire n8954;
wire n8955;
wire n8956;
wire n8957;
wire n8958;
wire n8959;
wire n8960;
wire n8961;
wire n8962;
wire n8963;
wire n8964;
wire n8965;
wire n8966;
wire n8967;
wire n8968;
wire n8969;
wire n8970;
wire n8971;
wire n8972;
wire n8973;
wire n8974;
wire n8975;
wire n8976;
wire n8977;
wire n8978;
wire n8979;
wire n8980;
wire n8981;
wire n8982;
wire n8983;
wire n8984;
wire n8985;
wire n8986;
wire n8987;
wire n8988;
wire n8989;
wire n8990;
wire n8991;
wire n8992;
wire n8993;
wire n8994;
wire n8995;
wire n8996;
wire n8997;
wire n8998;
wire n8999;
wire n9000;
wire n9001;
wire n9002;
wire n9003;
wire n9004;
wire n9005;
wire n9006;
wire n9007;
wire n9008;
wire n9009;
wire n9010;
wire n9011;
wire n9012;
wire n9013;
wire n9014;
wire n9015;
wire n9016;
wire n9017;
wire n9018;
wire n9019;
wire n9020;
wire n9021;
wire n9022;
wire n9023;
wire n9024;
wire n9025;
wire n9026;
wire n9027;
wire n9028;
wire n9029;
wire n9030;
wire n9031;
wire n9032;
wire n9033;
wire n9034;
wire n9035;
wire n9036;
wire n9037;
wire n9038;
wire n9039;
wire n9040;
wire n9041;
wire n9042;
wire n9043;
wire n9044;
wire n9045;
wire n9046;
wire n9047;
wire n9048;
wire n9049;
wire n9050;
wire n9051;
wire n9052;
wire n9053;
wire n9054;
wire n9055;
wire n9056;
wire n9057;
wire n9058;
wire n9059;
wire n9060;
wire n9061;
wire n9062;
wire n9063;
wire n9064;
wire n9065;
wire n9066;
wire n9067;
wire n9068;
wire n9069;
wire n9070;
wire n9071;
wire n9072;
wire n9073;
wire n9074;
wire n9075;
wire n9076;
wire n9077;
wire n9078;
wire n9079;
wire n9080;
wire n9081;
wire n9082;
wire n9083;
wire n9084;
wire n9085;
wire n9086;
wire n9087;
wire n9088;
wire n9089;
wire n9090;
wire n9091;
wire n9093;
wire n9094;
wire n9095;
wire n9096;
wire n9097;
wire n9098;
wire n9099;
wire n9100;
wire n9101;
wire n9102;
wire n9103;
wire n9104;
wire n9105;
wire n9107;
wire n9108;
wire n9109;
wire n9110;
wire n9111;
wire n9112;
wire n9113;
wire n9114;
wire n9115;
wire n9116;
wire n9117;
wire n9118;
wire n9119;
wire n9121;
wire n9122;
wire n9123;
wire n9124;
wire n9125;
wire n9126;
wire n9127;
wire n9128;
wire n9129;
wire n9130;
wire n9131;
wire n9132;
wire n9133;
wire n9134;
wire n9135;
wire n9136;
wire n9137;
wire n9138;
wire n9139;
wire n9140;
wire n9141;
wire n9143;
wire n9144;
wire n9145;
wire n9146;
wire n9147;
wire n9148;
wire n9149;
wire n9150;
wire n9151;
wire n9152;
wire n9153;
wire n9154;
wire n9155;
wire n9156;
wire n9157;
wire n9158;
wire n9159;
wire n9160;
wire n9161;
wire n9162;
wire n9163;
wire n9164;
wire n9165;
wire n9167;
wire n9168;
wire n9169;
wire n9170;
wire n9171;
wire n9172;
wire n9173;
wire n9174;
wire n9175;
wire n9176;
wire n9177;
wire n9178;
wire n9179;
wire n9180;
wire n9181;
wire n9182;
wire n9183;
wire n9184;
wire n9185;
wire n9186;
wire n9187;
wire n9188;
wire n9190;
wire n9191;
wire n9192;
wire n9193;
wire n9194;
wire n9195;
wire n9196;
wire n9197;
wire n9198;
wire n9199;
wire n9200;
wire n9201;
wire n9202;
wire n9203;
wire n9204;
wire n9205;
wire n9206;
wire n9207;
wire n9208;
wire n9209;
wire n9210;
wire n9211;
wire n9212;
wire n9213;
wire n9214;
wire n9216;
wire n9217;
wire n9218;
wire n9219;
wire n9220;
wire n9221;
wire n9222;
wire n9223;
wire n9224;
wire n9225;
wire n9226;
wire n9227;
wire n9228;
wire n9229;
wire n9230;
wire n9232;
wire n9233;
wire n9234;
wire n9235;
wire n9236;
wire n9237;
wire n9238;
wire n9239;
wire n9240;
wire n9241;
wire n9242;
wire n9243;
wire n9244;
wire n9245;
wire n9246;
wire n9247;
wire n9248;
wire n9249;
wire n9250;
wire n9251;
wire n9252;
wire n9253;
wire n9254;
wire n9255;
wire n9256;
wire n9257;
wire n9258;
wire n9259;
wire n9260;
wire n9261;
wire n9262;
wire n9263;
wire n9264;
wire n9265;
wire n9266;
wire n9267;
wire n9268;
wire n9269;
wire n9270;
wire n9271;
wire n9272;
wire n9273;
wire n9274;
wire n9275;
wire n9276;
wire n9277;
wire n9278;
wire n9279;
wire n9280;
wire n9281;
wire n9282;
wire n9283;
wire n9284;
wire n9285;
wire n9286;
wire n9287;
wire n9288;
wire n9289;
wire n9290;
wire n9291;
wire n9292;
wire n9293;
wire n9294;
wire n9295;
wire n9296;
wire n9297;
wire n9298;
wire n9299;
wire n9300;
wire n9301;
wire n9302;
wire n9303;
wire n9304;
wire n9305;
wire n9306;
wire n9307;
wire n9308;
wire n9309;
wire n9310;
wire n9311;
wire n9312;
wire n9313;
wire n9314;
wire n9315;
wire n9316;
wire n9317;
wire n9318;
wire n9319;
wire n9320;
wire n9321;
wire n9322;
wire n9323;
wire n9324;
wire n9325;
wire n9326;
wire n9327;
wire n9328;
wire n9329;
wire n9330;
wire n9331;
wire n9332;
wire n9333;
wire n9334;
wire n9335;
wire n9336;
wire n9337;
wire n9338;
wire n9339;
wire n9340;
wire n9341;
wire n9342;
wire n9343;
wire n9344;
wire n9345;
wire n9346;
wire n9347;
wire n9348;
wire n9349;
wire n9350;
wire n9351;
wire n9352;
wire n9353;
wire n9354;
wire n9355;
wire n9356;
wire n9357;
wire n9358;
wire n9359;
wire n9360;
wire n9361;
wire n9362;
wire n9363;
wire n9364;
wire n9365;
wire n9366;
wire n9367;
wire n9368;
wire n9369;
wire n9370;
wire n9371;
wire n9372;
wire n9373;
wire n9374;
wire n9375;
wire n9376;
wire n9377;
wire n9378;
wire n9379;
wire n9380;
wire n9381;
wire n9382;
wire n9383;
wire n9384;
wire n9385;
wire n9386;
wire n9387;
wire n9388;
wire n9389;
wire n9390;
wire n9391;
wire n9392;
wire n9393;
wire n9394;
wire n9395;
wire n9396;
wire n9397;
wire n9398;
wire n9399;
wire n9400;
wire n9401;
wire n9402;
wire n9403;
wire n9404;
wire n9406;
wire n9407;
wire n9408;
wire n9409;
wire n9410;
wire n9411;
wire n9412;
wire n9413;
wire n9414;
wire n9415;
wire n9416;
wire n9418;
wire n9419;
wire n9420;
wire n9421;
wire n9422;
wire n9423;
wire n9424;
wire n9425;
wire n9426;
wire n9427;
wire n9428;
wire n9430;
wire n9431;
wire n9432;
wire n9433;
wire n9434;
wire n9435;
wire n9436;
wire n9437;
wire n9438;
wire n9439;
wire n9440;
wire n9442;
wire n9443;
wire n9444;
wire n9445;
wire n9446;
wire n9447;
wire n9448;
wire n9449;
wire n9450;
wire n9451;
wire n9452;
wire n9454;
wire n9455;
wire n9456;
wire n9457;
wire n9458;
wire n9459;
wire n9460;
wire n9461;
wire n9462;
wire n9463;
wire n9464;
wire n9466;
wire n9467;
wire n9468;
wire n9469;
wire n9470;
wire n9471;
wire n9472;
wire n9473;
wire n9474;
wire n9475;
wire n9476;
wire n9478;
wire n9479;
wire n9480;
wire n9481;
wire n9482;
wire n9483;
wire n9484;
wire n9485;
wire n9486;
wire n9487;
wire n9489;
wire n9490;
wire n9491;
wire n9492;
wire n9493;
wire n9494;
wire n9495;
wire n9496;
wire n9497;
wire n9498;
wire n9499;
wire n9500;
wire n9501;
wire n9502;
wire n9503;
wire n9504;
wire n9505;
wire n9506;
wire n9507;
wire n9508;
wire n9509;
wire n9510;
wire n9511;
wire n9512;
wire n9513;
wire n9514;
wire n9515;
wire n9516;
wire n9517;
wire n9518;
wire n9519;
wire n9520;
wire n9521;
wire n9522;
wire n9523;
wire n9524;
wire n9525;
wire n9526;
wire n9527;
wire n9528;
wire n9529;
wire n9530;
wire n9531;
wire n9532;
wire n9533;
wire n9534;
wire n9535;
wire n9536;
wire n9537;
wire n9538;
wire n9539;
wire n9540;
wire n9541;
wire n9542;
wire n9543;
wire n9544;
wire n9545;
wire n9546;
wire n9547;
wire n9548;
wire n9549;
wire n9550;
wire n9551;
wire n9552;
wire n9553;
wire n9554;
wire n9555;
wire n9556;
wire n9557;
wire n9558;
wire n9559;
wire n9560;
wire n9561;
wire n9562;
wire n9563;
wire n9564;
wire n9565;
wire n9566;
wire n9567;
wire n9568;
wire n9569;
wire n9570;
wire n9571;
wire n9572;
wire n9573;
wire n9574;
wire n9575;
wire n9576;
wire n9577;
wire n9578;
wire n9579;
wire n9580;
wire n9581;
wire n9582;
wire n9583;
wire n9584;
wire n9585;
wire n9586;
wire n9587;
wire n9588;
wire n9589;
wire n9590;
wire n9591;
wire n9592;
wire n9593;
wire n9594;
wire n9595;
wire n9596;
wire n9597;
wire n9598;
wire n9599;
wire n9600;
wire n9601;
wire n9602;
wire n9603;
wire n9604;
wire n9605;
wire n9606;
wire n9607;
wire n9608;
wire n9609;
wire n9610;
wire n9611;
wire n9612;
wire n9613;
wire n9614;
wire n9615;
wire n9616;
wire n9617;
wire n9618;
wire n9619;
wire n9620;
wire n9621;
wire n9622;
wire n9623;
wire n9624;
wire n9625;
wire n9626;
wire n9627;
wire n9628;
wire n9629;
wire n9630;
wire n9631;
wire n9632;
wire n9633;
wire n9634;
wire n9635;
wire n9636;
wire n9637;
wire n9638;
wire n9639;
wire n9640;
wire n9641;
wire n9642;
wire n9643;
wire n9644;
wire n9645;
wire n9646;
wire n9647;
wire n9648;
wire n9649;
wire n9650;
wire n9651;
wire n9652;
wire n9653;
wire n9654;
wire n9655;
wire n9656;
wire n9657;
wire n9658;
wire n9659;
wire n9660;
wire n9661;
wire n9662;
wire n9663;
wire n9664;
wire n9665;
wire n9666;
wire n9667;
wire n9668;
wire n9669;
wire n9670;
wire n9671;
wire n9672;
wire n9673;
wire n9674;
wire n9675;
wire n9676;
wire n9677;
wire n9678;
wire n9679;
wire n9680;
wire n9681;
wire n9682;
wire n9683;
wire n9684;
wire n9685;
wire n9686;
wire n9687;
wire n9688;
wire n9689;
wire n9690;
wire n9691;
wire n9692;
wire n9693;
wire n9694;
wire n9695;
wire n9696;
wire n9697;
wire n9698;
wire n9699;
wire n9700;
wire n9701;
wire n9702;
wire n9703;
wire n9704;
wire n9705;
wire n9706;
wire n9707;
wire n9708;
wire n9709;
wire n9710;
wire n9711;
wire n9712;
wire n9713;
wire n9714;
wire n9715;
wire n9716;
wire n9717;
wire n9718;
wire n9719;
wire n9720;
wire n9721;
wire n9722;
wire n9723;
wire n9724;
wire n9725;
wire n9726;
wire n9727;
wire n9728;
wire n9729;
wire n9730;
wire n9731;
wire n9732;
wire n9733;
wire n9734;
wire n9735;
wire n9736;
wire n9737;
wire n9738;
wire n9739;
wire n9740;
wire n9741;
wire n9742;
wire n9743;
wire n9744;
wire n9745;
wire n9746;
wire n9747;
wire n9748;
wire n9749;
wire n9750;
wire n9751;
wire n9752;
wire n9753;
wire n9754;
wire n9755;
wire n9756;
wire n9757;
wire n9758;
wire n9759;
wire n9760;
wire n9761;
wire n9762;
wire n9763;
wire n9764;
wire n9765;
wire n9766;
wire n9767;
wire n9768;
wire n9769;
wire n9770;
wire n9771;
wire n9772;
wire n9773;
wire n9774;
wire n9775;
wire n9776;
wire n9777;
wire n9778;
wire n9779;
wire n9780;
wire n9781;
wire n9782;
wire n9783;
wire n9784;
wire n9785;
wire n9786;
wire n9787;
wire n9788;
wire n9789;
wire n9790;
wire n9791;
wire n9792;
wire n9793;
wire n9794;
wire n9795;
wire n9796;
wire n9797;
wire n9798;
wire n9799;
wire n9800;
wire n9801;
wire n9802;
wire n9803;
wire n9804;
wire n9805;
wire n9806;
wire n9807;
wire n9808;
wire n9809;
wire n9810;
wire n9811;
wire n9812;
wire n9813;
wire n9814;
wire n9815;
wire n9816;
wire n9817;
wire n9818;
wire n9819;
wire n9820;
wire n9821;
wire n9822;
wire n9823;
wire n9824;
wire n9825;
wire n9826;
wire n9827;
wire n9828;
wire n9829;
wire n9830;
wire n9831;
wire n9832;
wire n9833;
wire n9834;
wire n9835;
wire n9836;
wire n9837;
wire n9838;
wire n9839;
wire n9840;
wire n9841;
wire n9842;
wire n9843;
wire n9844;
wire n9845;
wire n9846;
wire n9847;
wire n9848;
wire n9849;
wire n9850;
wire n9851;
wire n9852;
wire n9853;
wire n9854;
wire n9855;
wire n9856;
wire n9857;
wire n9858;
wire n9859;
wire n9860;
wire n9861;
wire n9862;
wire n9863;
wire n9864;
wire n9865;
wire n9866;
wire n9867;
wire n9868;
wire n9869;
wire n9870;
wire n9871;
wire n9872;
wire n9873;
wire n9874;
wire n9875;
wire n9876;
wire n9877;
wire n9878;
wire n9879;
wire n9880;
wire n9881;
wire n9882;
wire n9883;
wire n9884;
wire n9885;
wire n9886;
wire n9887;
wire n9888;
wire n9889;
wire n9890;
wire n9891;
wire n9892;
wire n9893;
wire n9894;
wire n9895;
wire n9896;
wire n9897;
wire n9898;
wire n9899;
wire n9900;
wire n9901;
wire n9902;
wire n9903;
wire n9904;
wire n9905;
wire n9906;
wire n9907;
wire n9908;
wire n9909;
wire n9910;
wire n9911;
wire n9912;
wire n9913;
wire n9914;
wire n9915;
wire n9916;
wire n9917;
wire n9918;
wire n9919;
wire n9920;
wire n9921;
wire n9922;
wire n9923;
wire n9924;
wire n9925;
wire n9926;
wire n9927;
wire n9928;
wire n9929;
wire n9930;
wire n9931;
wire n9932;
wire n9933;
wire n9934;
wire n9935;
wire n9936;
wire n9937;
wire n9938;
wire n9939;
wire n9940;
wire n9942;
wire n9943;
wire n9945;
wire n9946;
wire n9947;
wire n9948;
wire n9949;
wire n9950;
wire n9951;
wire n9952;
wire n9953;
wire n9954;
wire n9955;
wire n9956;
wire n9957;
wire n9958;
wire n9959;
wire n9960;
wire n9961;
wire n9962;
wire n9963;
wire n9964;
wire n9965;
wire n9966;
wire n9967;
wire n9968;
wire n9969;
wire n9970;
wire n9971;
wire n9972;
wire n9973;
wire n9974;
wire n9975;
wire n9976;
wire n9977;
wire n9978;
wire n9979;
wire n9980;
wire n9981;
wire n9982;
wire n9983;
wire n9984;
wire n9985;
wire n9986;
wire n9987;
wire n9988;
wire n9989;
wire n9990;
wire n9991;
wire n9992;
wire n9993;
wire n9994;
wire n9995;
wire n9996;
wire n9997;
wire n9998;
wire n9999;
wire n10000;
wire n10001;
wire n10002;
wire n10003;
wire n10004;
wire n10005;
wire n10006;
wire n10007;
wire n10008;
wire n10009;
wire n10010;
wire n10011;
wire n10012;
wire n10013;
wire n10014;
wire n10015;
wire n10016;
wire n10017;
wire n10018;
wire n10019;
wire n10020;
wire n10021;
wire n10022;
wire n10023;
wire n10024;
wire n10025;
wire n10026;
wire n10027;
wire n10028;
wire n10029;
wire n10030;
wire n10031;
wire n10032;
wire n10033;
wire n10034;
wire n10035;
wire n10036;
wire n10037;
wire n10038;
wire n10039;
wire n10040;
wire n10041;
wire n10042;
wire n10043;
wire n10044;
wire n10045;
wire n10046;
wire n10047;
wire n10048;
wire n10049;
wire n10050;
wire n10051;
wire n10052;
wire n10053;
wire n10054;
wire n10055;
wire n10056;
wire n10057;
wire n10058;
wire n10059;
wire n10060;
wire n10061;
wire n10062;
wire n10063;
wire n10064;
wire n10065;
wire n10066;
wire n10067;
wire n10068;
wire n10069;
wire n10070;
wire n10071;
wire n10072;
wire n10073;
wire n10074;
wire n10075;
wire n10076;
wire n10077;
wire n10078;
wire n10079;
wire n10080;
wire n10081;
wire n10082;
wire n10083;
wire n10084;
wire n10085;
wire n10086;
wire n10087;
wire n10088;
wire n10089;
wire n10090;
wire n10091;
wire n10092;
wire n10093;
wire n10094;
wire n10095;
wire n10096;
wire n10097;
wire n10098;
wire n10099;
wire n10100;
wire n10101;
wire n10102;
wire n10103;
wire n10104;
wire n10105;
wire n10106;
wire n10107;
wire n10108;
wire n10109;
wire n10110;
wire n10111;
wire n10112;
wire n10113;
wire n10114;
wire n10115;
wire n10116;
wire n10117;
wire n10118;
wire n10119;
wire n10120;
wire n10121;
wire n10122;
wire n10123;
wire n10124;
wire n10125;
wire n10126;
wire n10127;
wire n10128;
wire n10129;
wire n10130;
wire n10131;
wire n10132;
wire n10133;
wire n10134;
wire n10135;
wire n10136;
wire n10137;
wire n10138;
wire n10139;
wire n10140;
wire n10141;
wire n10142;
wire n10143;
wire n10144;
wire n10145;
wire n10146;
wire n10147;
wire n10148;
wire n10149;
wire n10150;
wire n10151;
wire n10152;
wire n10153;
wire n10154;
wire n10155;
wire n10156;
wire n10157;
wire n10158;
wire n10159;
wire n10160;
wire n10161;
wire n10162;
wire n10163;
wire n10164;
wire n10165;
wire n10166;
wire n10167;
wire n10168;
wire n10169;
wire n10170;
wire n10171;
wire n10172;
wire n10173;
wire n10174;
wire n10175;
wire n10176;
wire n10177;
wire n10178;
wire n10179;
wire n10180;
wire n10181;
wire n10182;
wire n10183;
wire n10184;
wire n10185;
wire n10186;
wire n10187;
wire n10188;
wire n10189;
wire n10190;
wire n10191;
wire n10192;
wire n10193;
wire n10194;
wire n10195;
wire n10196;
wire n10197;
wire n10198;
wire n10199;
wire n10200;
wire n10201;
wire n10202;
wire n10203;
wire n10204;
wire n10205;
wire n10206;
wire n10207;
wire n10208;
wire n10209;
wire n10210;
wire n10211;
wire n10212;
wire n10213;
wire n10214;
wire n10215;
wire n10216;
wire n10217;
wire n10218;
wire n10219;
wire n10220;
wire n10221;
wire n10222;
wire n10223;
wire n10224;
wire n10225;
wire n10226;
wire n10227;
wire n10228;
wire n10229;
wire n10230;
wire n10231;
wire n10232;
wire n10233;
wire n10234;
wire n10235;
wire n10236;
wire n10237;
wire n10238;
wire n10239;
wire n10240;
wire n10241;
wire n10242;
wire n10243;
wire n10244;
wire n10245;
wire n10246;
wire n10247;
wire n10248;
wire n10249;
wire n10250;
wire n10251;
wire n10252;
wire n10253;
wire n10254;
wire n10255;
wire n10256;
wire n10257;
wire n10258;
wire n10259;
wire n10260;
wire n10261;
wire n10262;
wire n10263;
wire n10264;
wire n10265;
wire n10266;
wire n10267;
wire n10268;
wire n10269;
wire n10270;
wire n10271;
wire n10272;
wire n10273;
wire n10274;
wire n10275;
wire n10276;
wire n10277;
wire n10278;
wire n10279;
wire n10280;
wire n10281;
wire n10282;
wire n10283;
wire n10284;
wire n10285;
wire n10286;
wire n10287;
wire n10288;
wire n10289;
wire n10290;
wire n10291;
wire n10292;
wire n10293;
wire n10294;
wire n10295;
wire n10296;
wire n10297;
wire n10298;
wire n10299;
wire n10300;
wire n10301;
wire n10302;
wire n10303;
wire n10304;
wire n10305;
wire n10306;
wire n10307;
wire n10308;
wire n10309;
wire n10310;
wire n10311;
wire n10312;
wire n10313;
wire n10314;
wire n10315;
wire n10316;
wire n10317;
wire n10318;
wire n10319;
wire n10320;
wire n10321;
wire n10322;
wire n10323;
wire n10324;
wire n10325;
wire n10326;
wire n10327;
wire n10328;
wire n10329;
wire n10330;
wire n10331;
wire n10332;
wire n10333;
wire n10334;
wire n10335;
wire n10336;
wire n10337;
wire n10338;
wire n10339;
wire n10340;
wire n10341;
wire n10342;
wire n10343;
wire n10344;
wire n10345;
wire n10346;
wire n10347;
wire n10348;
wire n10349;
wire n10350;
wire n10351;
wire n10352;
wire n10353;
wire n10354;
wire n10355;
wire n10356;
wire n10357;
wire n10358;
wire n10359;
wire n10360;
wire n10361;
wire n10362;
wire n10363;
wire n10364;
wire n10365;
wire n10366;
wire n10367;
wire n10368;
wire n10369;
wire n10370;
wire n10371;
wire n10372;
wire n10373;
wire n10374;
wire n10375;
wire n10376;
wire n10377;
wire n10378;
wire n10379;
wire n10380;
wire n10381;
wire n10382;
wire n10383;
wire n10384;
wire n10385;
wire n10386;
wire n10387;
wire n10388;
wire n10389;
wire n10390;
wire n10391;
wire n10392;
wire n10393;
wire n10394;
wire n10395;
wire n10396;
wire n10397;
wire n10398;
wire n10399;
wire n10400;
wire n10401;
wire n10402;
wire n10403;
wire n10404;
wire n10405;
wire n10406;
wire n10407;
wire n10408;
wire n10409;
wire n10410;
wire n10411;
wire n10412;
wire n10413;
wire n10414;
wire n10415;
wire n10416;
wire n10417;
wire n10418;
wire n10419;
wire n10420;
wire n10421;
wire n10422;
wire n10423;
wire n10424;
wire n10425;
wire n10426;
wire n10427;
wire n10428;
wire n10429;
wire n10430;
wire n10431;
wire n10432;
wire n10433;
wire n10434;
wire n10435;
wire n10436;
wire n10437;
wire n10438;
wire n10439;
wire n10440;
wire n10441;
wire n10442;
wire n10443;
wire n10444;
wire n10445;
wire n10446;
wire n10447;
wire n10448;
wire n10449;
wire n10450;
wire n10451;
wire n10452;
wire n10453;
wire n10454;
wire n10455;
wire n10456;
wire n10457;
wire n10458;
wire n10459;
wire n10460;
wire n10461;
wire n10462;
wire n10463;
wire n10464;
wire n10465;
wire n10466;
wire n10467;
wire n10468;
wire n10469;
wire n10470;
wire n10471;
wire n10472;
wire n10473;
wire n10474;
wire n10475;
wire n10476;
wire n10477;
wire n10478;
wire n10479;
wire n10480;
wire n10481;
wire n10482;
wire n10483;
wire n10484;
wire n10485;
wire n10486;
wire n10487;
wire n10488;
wire n10489;
wire n10490;
wire n10491;
wire n10492;
wire n10493;
wire n10494;
wire n10495;
wire n10496;
wire n10497;
wire n10498;
wire n10499;
wire n10500;
wire n10501;
wire n10502;
wire n10503;
wire n10504;
wire n10505;
wire n10506;
wire n10507;
wire n10508;
wire n10509;
wire n10510;
wire n10511;
wire n10512;
wire n10513;
wire n10514;
wire n10515;
wire n10516;
wire n10517;
wire n10518;
wire n10519;
wire n10520;
wire n10521;
wire n10522;
wire n10523;
wire n10524;
wire n10525;
wire n10526;
wire n10527;
wire n10528;
wire n10529;
wire n10530;
wire n10531;
wire n10532;
wire n10533;
wire n10534;
wire n10535;
wire n10536;
wire n10537;
wire n10538;
wire n10539;
wire n10540;
wire n10541;
wire n10542;
wire n10543;
wire n10544;
wire n10545;
wire n10546;
wire n10547;
wire n10548;
wire n10549;
wire n10550;
wire n10551;
wire n10552;
wire n10555;
wire n10556;
wire n10557;
wire n10558;
wire n10559;
wire n10560;
wire n10561;
wire n10562;
wire n10563;
wire n10564;
wire n10565;
wire n10566;
wire n10567;
wire n10569;
wire n10570;
wire n10571;
wire n10572;
wire n10573;
wire n10576;
wire n10577;
wire n10578;
wire n10579;
wire n10580;
wire n10581;
wire n10582;
wire n10583;
wire n10584;
wire n10585;
wire n10586;
wire n10587;
wire n10588;
wire n10591;
wire n10592;
wire n10593;
wire n10594;
wire n10595;
wire n10596;
wire n10597;
wire n10598;
wire n10599;
wire n10600;
wire n10601;
wire n10602;
wire n10603;
wire n10604;
wire n10605;
wire n10606;
wire n10607;
wire n10608;
wire n10609;
wire n10610;
wire n10611;
wire n10612;
wire n10613;
wire n10614;
wire n10615;
wire n10616;
wire n10619;
wire n10620;
wire n10621;
wire n10622;
wire n10623;
wire n10624;
wire n10625;
wire n10626;
wire n10627;
wire n10628;
wire n10629;
wire n10630;
wire n10631;
wire n10633;
wire n10634;
wire n10635;
wire n10636;
wire n10637;
wire n10640;
wire n10641;
wire n10642;
wire n10643;
wire n10644;
wire n10645;
wire n10646;
wire n10647;
wire n10648;
wire n10649;
wire n10650;
wire n10651;
wire n10652;
wire n10655;
wire n10656;
wire n10657;
wire n10658;
wire n10659;
wire n10660;
wire n10661;
wire n10662;
wire n10663;
wire n10664;
wire n10665;
wire n10666;
wire n10667;
wire n10668;
wire n10669;
wire n10670;
wire n10671;
wire n10672;
wire n10673;
wire n10674;
wire n10675;
wire n10676;
wire n10677;
wire n10678;
wire n10679;
wire n10680;
wire n10683;
wire n10684;
wire n10685;
wire n10686;
wire n10687;
wire n10688;
wire n10689;
wire n10690;
wire n10691;
wire n10692;
wire n10693;
wire n10694;
wire n10695;
wire n10697;
wire n10698;
wire n10699;
wire n10700;
wire n10701;
wire n10704;
wire n10705;
wire n10706;
wire n10707;
wire n10708;
wire n10709;
wire n10710;
wire n10711;
wire n10712;
wire n10713;
wire n10714;
wire n10715;
wire n10716;
wire n10719;
wire n10720;
wire n10721;
wire n10722;
wire n10723;
wire n10724;
wire n10725;
wire n10726;
wire n10727;
wire n10728;
wire n10729;
wire n10730;
wire n10731;
wire n10732;
wire n10733;
wire n10734;
wire n10735;
wire n10736;
wire n10737;
wire n10738;
wire n10739;
wire n10740;
wire n10741;
wire n10742;
wire n10743;
wire n10744;
wire n10747;
wire n10748;
wire n10749;
wire n10750;
wire n10751;
wire n10752;
wire n10753;
wire n10754;
wire n10755;
wire n10756;
wire n10757;
wire n10758;
wire n10759;
wire n10761;
wire n10762;
wire n10763;
wire n10764;
wire n10765;
wire n10768;
wire n10769;
wire n10770;
wire n10771;
wire n10772;
wire n10773;
wire n10774;
wire n10775;
wire n10776;
wire n10777;
wire n10778;
wire n10779;
wire n10780;
wire n10783;
wire n10784;
wire n10785;
wire n10786;
wire n10787;
wire n10788;
wire n10789;
wire n10790;
wire n10791;
wire n10792;
wire n10793;
wire n10794;
wire n10795;
wire n10796;
wire n10797;
wire n10798;
wire n10799;
wire n10800;
wire n10801;
wire n10802;
wire n10803;
wire n10804;
wire n10805;
wire n10806;
wire n10807;
wire n10808;
wire n10809;
wire n10812;
wire n10813;
wire n10814;
wire n10815;
wire n10816;
wire n10817;
wire n10818;
wire n10819;
wire n10820;
wire n10821;
wire n10822;
wire n10823;
wire n10824;
wire n10826;
wire n10827;
wire n10828;
wire n10829;
wire n10830;
wire n10833;
wire n10834;
wire n10835;
wire n10836;
wire n10837;
wire n10838;
wire n10839;
wire n10840;
wire n10841;
wire n10842;
wire n10843;
wire n10844;
wire n10845;
wire n10846;
wire n10849;
wire n10850;
wire n10851;
wire n10852;
wire n10853;
wire n10854;
wire n10855;
wire n10856;
wire n10857;
wire n10858;
wire n10859;
wire n10860;
wire n10861;
wire n10862;
wire n10863;
wire n10864;
wire n10865;
wire n10866;
wire n10867;
wire n10868;
wire n10869;
wire n10870;
wire n10871;
wire n10872;
wire n10873;
wire n10874;
wire n10875;
wire n10876;
wire n10879;
wire n10880;
wire n10881;
wire n10882;
wire n10883;
wire n10884;
wire n10885;
wire n10886;
wire n10887;
wire n10888;
wire n10889;
wire n10890;
wire n10891;
wire n10892;
wire n10894;
wire n10895;
wire n10896;
wire n10897;
wire n10898;
wire n10901;
wire n10902;
wire n10903;
wire n10904;
wire n10905;
wire n10906;
wire n10907;
wire n10908;
wire n10909;
wire n10910;
wire n10911;
wire n10912;
wire n10913;
wire n10916;
wire n10917;
wire n10918;
wire n10919;
wire n10920;
wire n10921;
wire n10922;
wire n10923;
wire n10924;
wire n10925;
wire n10926;
wire n10927;
wire n10928;
wire n10929;
wire n10930;
wire n10931;
wire n10932;
wire n10933;
wire n10934;
wire n10935;
wire n10936;
wire n10937;
wire n10938;
wire n10939;
wire n10940;
wire n10941;
wire n10944;
wire n10945;
wire n10946;
wire n10947;
wire n10948;
wire n10949;
wire n10950;
wire n10951;
wire n10952;
wire n10953;
wire n10954;
wire n10955;
wire n10956;
wire n10958;
wire n10959;
wire n10960;
wire n10961;
wire n10962;
wire n10965;
wire n10966;
wire n10967;
wire n10968;
wire n10969;
wire n10970;
wire n10971;
wire n10972;
wire n10973;
wire n10974;
wire n10975;
wire n10976;
wire n10977;
wire n10980;
wire n10981;
wire n10982;
wire n10983;
wire n10984;
wire n10985;
wire n10986;
wire n10987;
wire n10988;
wire n10989;
wire n10990;
wire n10991;
wire n10992;
wire n10993;
wire n10994;
wire n10995;
wire n10996;
wire n10997;
wire n10998;
wire n10999;
wire n11000;
wire n11001;
wire n11002;
wire n11003;
wire n11004;
wire n11005;
wire n11008;
wire n11009;
wire n11010;
wire n11011;
wire n11012;
wire n11013;
wire n11014;
wire n11015;
wire n11016;
wire n11017;
wire n11018;
wire n11019;
wire n11020;
wire n11021;
wire n11023;
wire n11024;
wire n11025;
wire n11026;
wire n11027;
wire n11030;
wire n11031;
wire n11032;
wire n11033;
wire n11034;
wire n11035;
wire n11036;
wire n11037;
wire n11038;
wire n11039;
wire n11040;
wire n11041;
wire n11042;
wire n11043;
wire n11046;
wire n11047;
wire n11048;
wire n11049;
wire n11050;
wire n11051;
wire n11052;
wire n11053;
wire n11054;
wire n11055;
wire n11056;
wire n11057;
wire n11058;
wire n11059;
wire n11060;
wire n11061;
wire n11062;
wire n11063;
wire n11064;
wire n11065;
wire n11066;
wire n11067;
wire n11068;
wire n11069;
wire n11070;
wire n11071;
wire n11072;
wire n11073;
wire n11074;
wire n11075;
wire n11076;
wire n11077;
wire n11078;
wire n11079;
wire n11080;
wire n11081;
wire n11082;
wire n11083;
wire n11084;
wire n11085;
wire n11086;
wire n11087;
wire n11088;
wire n11089;
wire n11090;
wire n11091;
wire n11092;
wire n11093;
wire n11094;
wire n11095;
wire n11096;
wire n11097;
wire n11098;
wire n11099;
wire n11100;
wire n11101;
wire n11102;
wire n11103;
wire n11104;
wire n11105;
wire n11106;
wire n11107;
wire n11108;
wire n11109;
wire n11110;
wire n11111;
wire n11112;
wire n11113;
wire n11114;
wire n11115;
wire n11116;
wire n11117;
wire n11118;
wire n11119;
wire n11120;
wire n11121;
wire n11122;
wire n11123;
wire n11124;
wire n11125;
wire n11126;
wire n11127;
wire n11128;
wire n11129;
wire n11130;
wire n11131;
wire n11132;
wire n11133;
wire n11134;
wire n11135;
wire n11136;
wire n11137;
wire n11138;
wire n11139;
wire n11140;
wire n11141;
wire n11142;
wire n11143;
wire n11144;
wire n11145;
wire n11146;
wire n11147;
wire n11148;
wire n11149;
wire n11150;
wire n11151;
wire n11152;
wire n11153;
wire n11154;
wire n11155;
wire n11156;
wire n11157;
wire n11158;
wire n11159;
wire n11160;
wire n11161;
wire n11162;
wire n11165;
wire n11166;
wire n11167;
wire n11168;
wire n11169;
wire n11170;
wire n11171;
wire n11172;
wire n11173;
wire n11175;
wire n11176;
wire n11177;
wire n11178;
wire n11179;
wire n11182;
wire n11183;
wire n11184;
wire n11185;
wire n11186;
wire n11187;
wire n11188;
wire n11189;
wire n11190;
wire n11193;
wire n11194;
wire n11195;
wire n11196;
wire n11197;
wire n11198;
wire n11199;
wire n11200;
wire n11201;
wire n11202;
wire n11203;
wire n11204;
wire n11205;
wire n11206;
wire n11207;
wire n11208;
wire n11209;
wire n11212;
wire n11213;
wire n11214;
wire n11215;
wire n11216;
wire n11217;
wire n11218;
wire n11219;
wire n11220;
wire n11222;
wire n11223;
wire n11224;
wire n11225;
wire n11226;
wire n11229;
wire n11230;
wire n11231;
wire n11232;
wire n11233;
wire n11234;
wire n11235;
wire n11236;
wire n11237;
wire n11240;
wire n11241;
wire n11242;
wire n11243;
wire n11244;
wire n11245;
wire n11246;
wire n11247;
wire n11248;
wire n11249;
wire n11250;
wire n11251;
wire n11252;
wire n11253;
wire n11254;
wire n11255;
wire n11256;
wire n11259;
wire n11260;
wire n11261;
wire n11262;
wire n11263;
wire n11264;
wire n11265;
wire n11266;
wire n11267;
wire n11269;
wire n11270;
wire n11271;
wire n11272;
wire n11273;
wire n11276;
wire n11277;
wire n11278;
wire n11279;
wire n11280;
wire n11281;
wire n11282;
wire n11283;
wire n11284;
wire n11287;
wire n11288;
wire n11289;
wire n11290;
wire n11291;
wire n11292;
wire n11293;
wire n11294;
wire n11295;
wire n11296;
wire n11297;
wire n11298;
wire n11299;
wire n11300;
wire n11301;
wire n11302;
wire n11303;
wire n11306;
wire n11307;
wire n11308;
wire n11309;
wire n11310;
wire n11311;
wire n11312;
wire n11313;
wire n11314;
wire n11316;
wire n11317;
wire n11318;
wire n11319;
wire n11320;
wire n11323;
wire n11324;
wire n11325;
wire n11326;
wire n11327;
wire n11328;
wire n11329;
wire n11330;
wire n11331;
wire n11334;
wire n11335;
wire n11336;
wire n11337;
wire n11338;
wire n11339;
wire n11340;
wire n11341;
wire n11342;
wire n11343;
wire n11344;
wire n11345;
wire n11346;
wire n11347;
wire n11348;
wire n11349;
wire n11350;
wire n11353;
wire n11354;
wire n11355;
wire n11356;
wire n11357;
wire n11358;
wire n11359;
wire n11360;
wire n11361;
wire n11363;
wire n11364;
wire n11365;
wire n11366;
wire n11367;
wire n11370;
wire n11371;
wire n11372;
wire n11373;
wire n11374;
wire n11375;
wire n11376;
wire n11377;
wire n11380;
wire n11381;
wire n11382;
wire n11383;
wire n11384;
wire n11385;
wire n11386;
wire n11387;
wire n11388;
wire n11389;
wire n11390;
wire n11391;
wire n11392;
wire n11393;
wire n11394;
wire n11395;
wire n11398;
wire n11399;
wire n11400;
wire n11401;
wire n11402;
wire n11403;
wire n11404;
wire n11405;
wire n11406;
wire n11408;
wire n11409;
wire n11410;
wire n11411;
wire n11412;
wire n11415;
wire n11416;
wire n11417;
wire n11418;
wire n11419;
wire n11420;
wire n11421;
wire n11422;
wire n11423;
wire n11426;
wire n11427;
wire n11428;
wire n11429;
wire n11430;
wire n11431;
wire n11432;
wire n11433;
wire n11434;
wire n11435;
wire n11436;
wire n11437;
wire n11438;
wire n11439;
wire n11440;
wire n11441;
wire n11442;
wire n11445;
wire n11446;
wire n11447;
wire n11448;
wire n11449;
wire n11450;
wire n11451;
wire n11452;
wire n11453;
wire n11455;
wire n11456;
wire n11457;
wire n11458;
wire n11459;
wire n11462;
wire n11463;
wire n11464;
wire n11465;
wire n11466;
wire n11467;
wire n11468;
wire n11469;
wire n11470;
wire n11473;
wire n11474;
wire n11475;
wire n11476;
wire n11477;
wire n11478;
wire n11479;
wire n11480;
wire n11481;
wire n11482;
wire n11483;
wire n11484;
wire n11485;
wire n11486;
wire n11487;
wire n11488;
wire n11491;
wire n11492;
wire n11493;
wire n11494;
wire n11495;
wire n11496;
wire n11497;
wire n11498;
wire n11499;
wire n11501;
wire n11502;
wire n11503;
wire n11504;
wire n11505;
wire n11508;
wire n11509;
wire n11510;
wire n11511;
wire n11512;
wire n11513;
wire n11514;
wire n11515;
wire n11516;
wire n11519;
wire n11520;
wire n11521;
wire n11522;
wire n11523;
wire n11524;
wire n11525;
wire n11526;
wire n11527;
wire n11528;
wire n11529;
wire n11530;
wire n11531;
wire n11532;
wire n11533;
wire n11534;
wire n11535;
wire n11536;
wire n11537;
wire n11538;
wire n11539;
wire n11540;
wire n11541;
wire n11542;
wire n11543;
wire n11544;
wire n11545;
wire n11546;
wire n11547;
wire n11548;
wire n11549;
wire n11550;
wire n11551;
wire n11552;
wire n11553;
wire n11554;
wire n11555;
wire n11556;
wire n11557;
wire n11558;
wire n11559;
wire n11560;
wire n11561;
wire n11562;
wire n11563;
wire n11564;
wire n11565;
wire n11566;
wire n11567;
wire n11568;
wire n11569;
wire n11570;
wire n11571;
wire n11572;
wire n11573;
wire n11574;
wire n11575;
wire n11576;
wire n11577;
wire n11578;
wire n11579;
wire n11580;
wire n11581;
wire n11582;
wire n11583;
wire n11584;
wire n11585;
wire n11586;
wire n11587;
wire n11588;
wire n11589;
wire n11590;
wire n11591;
wire n11592;
wire n11593;
wire n11594;
wire n11595;
wire n11596;
wire n11597;
wire n11598;
wire n11599;
wire n11600;
wire n11601;
wire n11602;
wire n11603;
wire n11604;
wire n11605;
wire n11606;
wire n11607;
wire n11608;
wire n11609;
wire n11610;
wire n11611;
wire n11612;
wire n11613;
wire n11614;
wire n11615;
wire n11616;
wire n11617;
wire n11618;
wire n11619;
wire n11620;
wire n11621;
wire n11622;
wire n11623;
wire n11624;
wire n11625;
wire n11626;
wire n11627;
wire n11628;
wire n11629;
wire n11630;
wire n11631;
wire n11632;
wire n11633;
wire n11634;
wire n11635;
wire n11636;
wire n11637;
wire n11638;
wire n11639;
wire n11640;
wire n11641;
wire n11642;
wire n11643;
wire n11644;
wire n11645;
wire n11646;
wire n11647;
wire n11648;
wire n11649;
wire n11650;
wire n11651;
wire n11652;
wire n11653;
wire n11654;
wire n11655;
wire n11656;
wire n11657;
wire n11658;
wire n11659;
wire n11660;
wire n11661;
wire n11662;
wire n11663;
wire n11664;
wire n11665;
wire n11666;
wire n11667;
wire n11668;
wire n11669;
wire n11670;
wire n11671;
wire n11672;
wire n11673;
wire n11674;
wire n11675;
wire n11676;
wire n11677;
wire n11678;
wire n11679;
wire n11680;
wire n11681;
wire n11682;
wire n11683;
wire n11684;
wire n11685;
wire n11686;
wire n11687;
wire n11688;
wire n11689;
wire n11690;
wire n11691;
wire n11692;
wire n11693;
wire n11694;
wire n11695;
wire n11696;
wire n11697;
wire n11698;
wire n11699;
wire n11700;
wire n11701;
wire n11702;
wire n11703;
wire n11704;
wire n11705;
wire n11706;
wire n11707;
wire n11708;
wire n11709;
wire n11710;
wire n11711;
wire n11712;
wire n11713;
wire n11714;
wire n11715;
wire n11716;
wire n11717;
wire n11718;
wire n11719;
wire n11720;
wire n11721;
wire n11722;
wire n11723;
wire n11724;
wire n11725;
wire n11726;
wire n11727;
wire n11728;
wire n11729;
wire n11730;
wire n11731;
wire n11732;
wire n11733;
wire n11734;
wire n11735;
wire n11736;
wire n11737;
wire n11738;
wire n11739;
wire n11740;
wire n11741;
wire n11742;
wire n11743;
wire n11744;
wire n11745;
wire n11746;
wire n11748;
wire n11749;
wire n11750;
wire n11752;
wire n11753;
wire n11754;
wire n11755;
wire n11757;
wire n11758;
wire n11759;
wire n11760;
wire n11762;
wire n11763;
wire n11764;
wire n11765;
wire n11767;
wire n11768;
wire n11769;
wire n11770;
wire n11771;
wire n11772;
wire n11773;
wire n11774;
wire n11775;
wire n11778;
wire n11779;
wire n11781;
wire n11782;
wire n11784;
wire n11785;
wire n11787;
wire n11788;
wire n11789;
wire n11790;
wire n11792;
wire n11793;
wire n11795;
wire n11796;
wire n11798;
wire n11799;
wire n11801;
wire n11802;
wire n11804;
wire n11805;
wire n11806;
wire n11807;
wire n11808;
wire n11809;
wire n11810;
wire n11811;
wire n11812;
wire n11815;
wire n11816;
wire n11818;
wire n11819;
wire n11821;
wire n11822;
wire n11824;
wire n11825;
wire n11826;
wire n11827;
wire n11829;
wire n11830;
wire n11832;
wire n11833;
wire n11835;
wire n11836;
wire n11838;
wire n11839;
wire n11841;
wire n11842;
wire n11843;
wire n11844;
wire n11845;
wire n11846;
wire n11847;
wire n11848;
wire n11849;
wire n11852;
wire n11853;
wire n11855;
wire n11856;
wire n11858;
wire n11859;
wire n11861;
wire n11862;
wire n11863;
wire n11864;
wire n11866;
wire n11867;
wire n11869;
wire n11870;
wire n11872;
wire n11873;
wire n11875;
wire n11876;
wire n11878;
wire n11879;
wire n11880;
wire n11881;
wire n11882;
wire n11883;
wire n11884;
wire n11885;
wire n11886;
wire n11889;
wire n11890;
wire n11892;
wire n11893;
wire n11895;
wire n11896;
wire n11898;
wire n11899;
wire n11900;
wire n11901;
wire n11903;
wire n11904;
wire n11906;
wire n11907;
wire n11909;
wire n11910;
wire n11912;
wire n11913;
wire n11915;
wire n11916;
wire n11917;
wire n11918;
wire n11919;
wire n11920;
wire n11921;
wire n11922;
wire n11923;
wire n11926;
wire n11927;
wire n11929;
wire n11930;
wire n11932;
wire n11933;
wire n11935;
wire n11936;
wire n11937;
wire n11938;
wire n11940;
wire n11941;
wire n11943;
wire n11944;
wire n11946;
wire n11947;
wire n11949;
wire n11950;
wire n11952;
wire n11953;
wire n11954;
wire n11955;
wire n11956;
wire n11957;
wire n11958;
wire n11959;
wire n11960;
wire n11963;
wire n11964;
wire n11966;
wire n11967;
wire n11969;
wire n11970;
wire n11972;
wire n11973;
wire n11974;
wire n11975;
wire n11977;
wire n11978;
wire n11980;
wire n11981;
wire n11983;
wire n11984;
wire n11986;
wire n11987;
wire n11989;
wire n11990;
wire n11991;
wire n11992;
wire n11993;
wire n11994;
wire n11995;
wire n11996;
wire n11997;
wire n12000;
wire n12001;
wire n12003;
wire n12004;
wire n12006;
wire n12007;
wire n12009;
wire n12010;
wire n12011;
wire n12012;
wire n12014;
wire n12015;
wire n12017;
wire n12018;
wire n12020;
wire n12021;
wire n12023;
wire n12024;
wire n12026;
wire n12027;
wire n12028;
wire n12029;
wire n12030;
wire n12031;
wire n12032;
wire n12033;
wire n12036;
wire n12037;
wire n12039;
wire n12040;
wire n12042;
wire n12043;
wire n12045;
wire n12046;
wire n12047;
wire n12048;
wire n12050;
wire n12051;
wire n12053;
wire n12054;
wire n12056;
wire n12057;
wire n12059;
wire n12060;
wire n12062;
wire n12063;
wire n12064;
wire n12065;
wire n12066;
wire n12067;
wire n12068;
wire n12069;
wire n12070;
wire n12071;
wire n12072;
wire n12073;
wire n12074;
wire n12075;
wire n12076;
wire n12077;
wire n12078;
wire n12079;
wire n12080;
wire n12081;
wire n12082;
wire n12083;
wire n12084;
wire n12085;
wire n12086;
wire n12087;
wire n12088;
wire n12089;
wire n12090;
wire n12091;
wire n12092;
wire n12093;
wire n12094;
wire n12095;
wire n12096;
wire n12097;
wire n12098;
wire n12099;
wire n12100;
wire n12101;
wire n12102;
wire n12103;
wire n12104;
wire n12105;
wire n12106;
wire n12107;
wire n12108;
wire n12109;
wire n12110;
wire n12111;
wire n12112;
wire n12113;
wire n12114;
wire n12115;
wire n12116;
wire n12117;
wire n12118;
wire n12119;
wire n12120;
wire n12121;
wire n12122;
wire n12123;
wire n12125;
wire n12126;
wire n12128;
wire n12129;
wire n12130;
wire n12132;
wire n12133;
wire n12135;
wire n12136;
wire n12137;
wire n12138;
wire n12139;
wire n12140;
wire n12141;
wire n12142;
wire n12143;
wire n12146;
wire n12147;
wire n12149;
wire n12150;
wire n12152;
wire n12153;
wire n12155;
wire n12156;
wire n12157;
wire n12158;
wire n12160;
wire n12161;
wire n12163;
wire n12164;
wire n12166;
wire n12167;
wire n12169;
wire n12170;
wire n12172;
wire n12173;
wire n12174;
wire n12175;
wire n12176;
wire n12177;
wire n12178;
wire n12179;
wire n12180;
wire n12183;
wire n12184;
wire n12186;
wire n12187;
wire n12189;
wire n12190;
wire n12192;
wire n12193;
wire n12194;
wire n12195;
wire n12197;
wire n12198;
wire n12200;
wire n12201;
wire n12203;
wire n12204;
wire n12206;
wire n12207;
wire n12209;
wire n12210;
wire n12211;
wire n12212;
wire n12213;
wire n12214;
wire n12215;
wire n12216;
wire n12217;
wire n12220;
wire n12221;
wire n12223;
wire n12224;
wire n12226;
wire n12227;
wire n12229;
wire n12230;
wire n12231;
wire n12232;
wire n12234;
wire n12235;
wire n12237;
wire n12238;
wire n12240;
wire n12241;
wire n12243;
wire n12244;
wire n12246;
wire n12247;
wire n12248;
wire n12249;
wire n12250;
wire n12251;
wire n12252;
wire n12253;
wire n12254;
wire n12257;
wire n12258;
wire n12260;
wire n12261;
wire n12263;
wire n12264;
wire n12266;
wire n12267;
wire n12268;
wire n12269;
wire n12271;
wire n12272;
wire n12274;
wire n12275;
wire n12277;
wire n12278;
wire n12280;
wire n12281;
wire n12283;
wire n12284;
wire n12285;
wire n12286;
wire n12287;
wire n12288;
wire n12289;
wire n12290;
wire n12291;
wire n12294;
wire n12295;
wire n12297;
wire n12298;
wire n12300;
wire n12301;
wire n12303;
wire n12304;
wire n12305;
wire n12306;
wire n12308;
wire n12309;
wire n12311;
wire n12312;
wire n12314;
wire n12315;
wire n12317;
wire n12318;
wire n12320;
wire n12321;
wire n12322;
wire n12323;
wire n12324;
wire n12325;
wire n12326;
wire n12327;
wire n12328;
wire n12331;
wire n12332;
wire n12334;
wire n12335;
wire n12337;
wire n12338;
wire n12340;
wire n12341;
wire n12342;
wire n12343;
wire n12345;
wire n12346;
wire n12348;
wire n12349;
wire n12351;
wire n12352;
wire n12354;
wire n12355;
wire n12357;
wire n12358;
wire n12359;
wire n12360;
wire n12361;
wire n12362;
wire n12363;
wire n12364;
wire n12365;
wire n12368;
wire n12369;
wire n12371;
wire n12372;
wire n12374;
wire n12375;
wire n12377;
wire n12378;
wire n12379;
wire n12380;
wire n12382;
wire n12383;
wire n12385;
wire n12386;
wire n12388;
wire n12389;
wire n12391;
wire n12392;
wire n12394;
wire n12395;
wire n12396;
wire n12397;
wire n12398;
wire n12399;
wire n12400;
wire n12401;
wire n12404;
wire n12405;
wire n12407;
wire n12408;
wire n12410;
wire n12411;
wire n12413;
wire n12414;
wire n12415;
wire n12416;
wire n12418;
wire n12419;
wire n12421;
wire n12422;
wire n12424;
wire n12425;
wire n12427;
wire n12428;
wire n12430;
wire n12431;
wire n12432;
wire n12433;
wire n12434;
wire n12435;
wire n12436;
wire n12437;
wire n12438;
wire n12439;
wire n12440;
wire n12441;
wire n12442;
wire n12443;
wire n12444;
wire n12445;
wire n12446;
wire n12447;
wire n12448;
wire n12449;
wire n12450;
wire n12451;
wire n12452;
wire n12453;
wire n12454;
wire n12456;
wire n12457;
wire n12458;
wire n12459;
wire n12460;
wire n12461;
wire n12462;
wire n12463;
wire n12464;
wire n12465;
wire n12466;
wire n12467;
wire n12468;
wire n12469;
wire n12470;
wire n12471;
wire n12472;
wire n12473;
wire n12474;
wire n12475;
wire n12476;
wire n12477;
wire n12478;
wire n12479;
wire n12480;
wire n12481;
wire n12482;
wire n12483;
wire n12484;
wire n12485;
wire n12486;
wire n12487;
wire n12488;
wire n12489;
wire n12490;
wire n12491;
wire n12492;
wire n12493;
wire n12494;
wire n12495;
wire n12496;
wire n12497;
wire n12498;
wire n12499;
wire n12500;
wire n12501;
wire n12502;
wire n12503;
wire n12504;
wire n12505;
wire n12506;
wire n12507;
wire n12508;
wire n12509;
wire n12510;
wire n12511;
wire n12512;
wire n12513;
wire n12514;
wire n12515;
wire n12516;
wire n12517;
wire n12518;
wire n12519;
wire n12520;
wire n12521;
wire n12522;
wire n12523;
wire n12524;
wire n12525;
wire n12526;
wire n12527;
wire n12528;
wire n12529;
wire n12530;
wire n12531;
wire n12532;
wire n12533;
wire n12534;
wire n12535;
wire n12536;
wire n12537;
wire n12538;
wire n12539;
wire n12540;
wire n12541;
wire n12542;
wire n12543;
wire n12544;
wire n12545;
wire n12546;
wire n12547;
wire n12548;
wire n12549;
wire n12550;
wire n12551;
wire n12552;
wire n12553;
wire n12554;
wire n12555;
wire n12556;
wire n12557;
wire n12558;
wire n12559;
wire n12560;
wire n12561;
wire n12562;
wire n12563;
wire n12564;
wire n12565;
wire n12566;
wire n12567;
wire n12568;
wire n12569;
wire n12570;
wire n12571;
wire n12572;
wire n12573;
wire n12574;
wire n12575;
wire n12576;
wire n12577;
wire n12578;
wire n12579;
wire n12580;
wire n12581;
wire n12582;
wire n12583;
wire n12584;
wire n12585;
wire n12586;
wire n12587;
wire n12588;
wire n12589;
wire n12590;
wire n12591;
wire n12592;
wire n12593;
wire n12594;
wire n12595;
wire n12596;
wire n12597;
wire n12598;
wire n12599;
wire n12600;
wire n12601;
wire n12602;
wire n12603;
wire n12604;
wire n12605;
wire n12606;
wire n12607;
wire n12608;
wire n12609;
wire n12610;
wire n12611;
wire n12612;
wire n12613;
wire n12614;
wire n12615;
wire n12616;
wire n12617;
wire n12618;
wire n12619;
wire n12620;
wire n12621;
wire n12622;
wire n12623;
wire n12624;
wire n12625;
wire n12626;
wire n12627;
wire n12628;
wire n12629;
wire n12630;
wire n12631;
wire n12632;
wire n12633;
wire n12634;
wire n12635;
wire n12636;
wire n12637;
wire n12638;
wire n12639;
wire n12640;
wire n12641;
wire n12642;
wire n12643;
wire n12644;
wire n12645;
wire n12646;
wire n12647;
wire n12648;
wire n12649;
wire n12650;
wire n12651;
wire n12652;
wire n12653;
wire n12654;
wire n12655;
wire n12656;
wire n12657;
wire n12658;
wire n12659;
wire n12660;
wire n12661;
wire n12662;
wire n12663;
wire n12664;
wire n12665;
wire n12666;
wire n12667;
wire n12668;
wire n12669;
wire n12670;
wire n12671;
wire n12672;
wire n12673;
wire n12674;
wire n12675;
wire n12676;
wire n12677;
wire n12678;
wire n12679;
wire n12680;
wire n12681;
wire n12682;
wire n12683;
wire n12684;
wire n12685;
wire n12686;
wire n12687;
wire n12688;
wire n12689;
wire n12690;
wire n12691;
wire n12692;
wire n12693;
wire n12694;
wire n12695;
wire n12696;
wire n12697;
wire n12698;
wire n12699;
wire n12700;
wire n12701;
wire n12702;
wire n12703;
wire n12704;
wire n12705;
wire n12706;
wire n12707;
wire n12708;
wire n12709;
wire n12710;
wire n12711;
wire n12712;
wire n12713;
wire n12714;
wire n12715;
wire n12716;
wire n12717;
wire n12718;
wire n12719;
wire n12720;
wire n12721;
wire n12722;
wire n12723;
wire n12724;
wire n12725;
wire n12726;
wire n12727;
wire n12728;
wire n12729;
wire n12730;
wire n12731;
wire n12732;
wire n12733;
wire n12734;
wire n12735;
wire n12736;
wire n12737;
wire n12738;
wire n12739;
wire n12740;
wire n12741;
wire n12742;
wire n12743;
wire n12744;
wire n12745;
wire n12746;
wire n12747;
wire n12748;
wire n12749;
wire n12750;
wire n12751;
wire n12752;
wire n12753;
wire n12754;
wire n12755;
wire n12756;
wire n12757;
wire n12758;
wire n12759;
wire n12760;
wire n12761;
wire n12762;
wire n12763;
wire n12764;
wire n12765;
wire n12766;
wire n12767;
wire n12768;
wire n12769;
wire n12770;
wire n12771;
wire n12772;
wire n12773;
wire n12774;
wire n12775;
wire n12776;
wire n12777;
wire n12778;
wire n12779;
wire n12780;
wire n12781;
wire n12782;
wire n12783;
wire n12784;
wire n12785;
wire n12786;
wire n12787;
wire n12788;
wire n12789;
wire n12790;
wire n12791;
wire n12792;
wire n12793;
wire n12794;
wire n12795;
wire n12796;
wire n12797;
wire n12798;
wire n12799;
wire n12800;
wire n12801;
wire n12802;
wire n12803;
wire n12804;
wire n12805;
wire n12806;
wire n12807;
wire n12808;
wire n12809;
wire n12810;
wire n12811;
wire n12812;
wire n12813;
wire n12814;
wire n12815;
wire n12816;
wire n12817;
wire n12818;
wire n12819;
wire n12820;
wire n12821;
wire n12822;
wire n12823;
wire n12825;
wire n12826;
wire n12827;
wire n12828;
wire n12829;
wire n12830;
wire n12832;
wire n12833;
wire n12834;
wire n12835;
wire n12836;
wire n12837;
wire n12838;
wire n12839;
wire n12840;
wire n12841;
wire n12842;
wire n12843;
wire n12844;
wire n12845;
wire n12846;
wire n12847;
wire n12848;
wire n12849;
wire n12850;
wire n12851;
wire n12852;
wire n12853;
wire n12854;
wire n12855;
wire n12856;
wire n12857;
wire n12858;
wire n12859;
wire n12860;
wire n12861;
wire n12862;
wire n12863;
wire n12864;
wire n12865;
wire n12866;
wire n12867;
wire n12868;
wire n12869;
wire n12870;
wire n12871;
wire n12872;
wire n12873;
wire n12875;
wire n12876;
wire n12878;
wire n12879;
wire n12880;
wire n12881;
wire n12882;
wire n12883;
wire n12884;
wire n12885;
wire n12886;
wire n12887;
wire n12888;
wire n12889;
wire n12890;
wire n12891;
wire n12892;
wire n12893;
wire n12894;
wire n12895;
wire n12896;
wire n12897;
wire n12898;
wire n12899;
wire n12900;
wire n12901;
wire n12902;
wire n12903;
wire n12904;
wire n12905;
wire n12906;
wire n12907;
wire n12908;
wire n12909;
wire n12910;
wire n12911;
wire n12912;
wire n12913;
wire n12914;
wire n12915;
wire n12916;
wire n12917;
wire n12918;
wire n12919;
wire n12920;
wire n12921;
wire n12922;
wire n12923;
wire n12924;
wire n12925;
wire n12926;
wire n12927;
wire n12928;
wire n12929;
wire n12930;
wire n12931;
wire n12932;
wire n12933;
wire n12934;
wire n12935;
wire n12936;
wire n12937;
wire n12938;
wire n12939;
wire n12940;
wire n12941;
wire n12942;
wire n12943;
wire n12944;
wire n12945;
wire n12946;
wire n12947;
wire n12948;
wire n12949;
wire n12950;
wire n12951;
wire n12952;
wire n12953;
wire n12954;
wire n12955;
wire n12956;
wire n12957;
wire n12958;
wire n12959;
wire n12960;
wire n12961;
wire n12962;
wire n12963;
wire n12964;
wire n12965;
wire n12966;
wire n12967;
wire n12968;
wire n12969;
wire n12970;
wire n12971;
wire n12972;
wire n12973;
wire n12974;
wire n12975;
wire n12976;
wire n12977;
wire n12978;
wire n12979;
wire n12980;
wire n12981;
wire n12982;
wire n12983;
wire n12984;
wire n12985;
wire n12986;
wire n12987;
wire n12988;
wire n12989;
wire n12990;
wire n12991;
wire n12992;
wire n12993;
wire n12994;
wire n12995;
wire n12996;
wire n12997;
wire n12998;
wire n12999;
wire n13000;
wire n13001;
wire n13002;
wire n13003;
wire n13004;
wire n13005;
wire n13006;
wire n13007;
wire n13008;
wire n13009;
wire n13010;
wire n13011;
wire n13012;
wire n13013;
wire n13014;
wire n13015;
wire n13016;
wire n13017;
wire n13018;
wire n13019;
wire n13020;
wire n13021;
wire n13022;
wire n13023;
wire n13024;
wire n13025;
wire n13026;
wire n13027;
wire n13028;
wire n13029;
wire n13030;
wire n13031;
wire n13032;
wire n13033;
wire n13034;
wire n13035;
wire n13036;
wire n13037;
wire n13038;
wire n13039;
wire n13040;
wire n13041;
wire n13042;
wire n13043;
wire n13044;
wire n13045;
wire n13046;
wire n13047;
wire n13048;
wire n13049;
wire n13050;
wire n13051;
wire n13052;
wire n13053;
wire n13054;
wire n13055;
wire n13056;
wire n13057;
wire n13058;
wire n13059;
wire n13060;
wire n13061;
wire n13062;
wire n13063;
wire n13064;
wire n13065;
wire n13066;
wire n13068;
wire n13069;
wire n13071;
wire n13072;
wire n13073;
wire n13074;
wire n13075;
wire n13076;
wire n13077;
wire n13078;
wire n13079;
wire n13080;
wire n13081;
wire n13082;
wire n13083;
wire n13084;
wire n13085;
wire n13086;
wire n13087;
wire n13088;
wire n13089;
wire n13090;
wire n13091;
wire n13092;
wire n13093;
wire n13094;
wire n13095;
wire n13096;
wire n13097;
wire n13098;
wire n13099;
wire n13100;
wire n13101;
wire n13102;
wire n13103;
wire n13104;
wire n13105;
wire n13106;
wire n13107;
wire n13108;
wire n13109;
wire n13110;
wire n13111;
wire n13112;
wire n13113;
wire n13114;
wire n13115;
wire n13116;
wire n13117;
wire n13118;
wire n13119;
wire n13120;
wire n13121;
wire n13122;
wire n13123;
wire n13124;
wire n13125;
wire n13126;
wire n13127;
wire n13128;
wire n13129;
wire n13130;
wire n13131;
wire n13132;
wire n13133;
wire n13134;
wire n13135;
wire n13136;
wire n13137;
wire n13138;
wire n13139;
wire n13140;
wire n13141;
wire n13142;
wire n13143;
wire n13144;
wire n13145;
wire n13146;
wire n13147;
wire n13148;
wire n13149;
wire n13150;
wire n13151;
wire n13152;
wire n13153;
wire n13154;
wire n13155;
wire n13156;
wire n13157;
wire n13158;
wire n13159;
wire n13160;
wire n13161;
wire n13162;
wire n13163;
wire n13164;
wire n13165;
wire n13166;
wire n13167;
wire n13168;
wire n13169;
wire n13170;
wire n13171;
wire n13172;
wire n13173;
wire n13174;
wire n13175;
wire n13176;
wire n13177;
wire n13178;
wire n13180;
wire n13181;
wire n13183;
wire n13184;
wire n13185;
wire n13186;
wire n13187;
wire n13188;
wire n13189;
wire n13190;
wire n13191;
wire n13192;
wire n13193;
wire n13194;
wire n13195;
wire n13196;
wire n13197;
wire n13198;
wire n13199;
wire n13200;
wire n13201;
wire n13202;
wire n13203;
wire n13204;
wire n13205;
wire n13206;
wire n13207;
wire n13208;
wire n13209;
wire n13210;
wire n13211;
wire n13212;
wire n13213;
wire n13214;
wire n13215;
wire n13216;
wire n13217;
wire n13218;
wire n13219;
wire n13220;
wire n13221;
wire n13222;
wire n13223;
wire n13224;
wire n13225;
wire n13226;
wire n13227;
wire n13228;
wire n13229;
wire n13230;
wire n13231;
wire n13232;
wire n13233;
wire n13234;
wire n13235;
wire n13236;
wire n13237;
wire n13238;
wire n13239;
wire n13240;
wire n13241;
wire n13242;
wire n13243;
wire n13244;
wire n13245;
wire n13246;
wire n13247;
wire n13248;
wire n13249;
wire n13250;
wire n13251;
wire n13252;
wire n13253;
wire n13254;
wire n13255;
wire n13256;
wire n13257;
wire n13258;
wire n13259;
wire n13260;
wire n13261;
wire n13262;
wire n13263;
wire n13264;
wire n13265;
wire n13266;
wire n13267;
wire n13268;
wire n13269;
wire n13270;
wire n13271;
wire n13272;
wire n13273;
wire n13274;
wire n13275;
wire n13276;
wire n13277;
wire n13278;
wire n13279;
wire n13280;
wire n13281;
wire n13282;
wire n13283;
wire n13284;
wire n13285;
wire n13286;
wire n13287;
wire n13288;
wire n13289;
wire n13290;
wire n13292;
wire n13293;
wire n13295;
wire n13296;
wire n13297;
wire n13298;
wire n13299;
wire n13300;
wire n13301;
wire n13302;
wire n13303;
wire n13304;
wire n13305;
wire n13306;
wire n13307;
wire n13308;
wire n13309;
wire n13310;
wire n13311;
wire n13312;
wire n13313;
wire n13314;
wire n13315;
wire n13316;
wire n13317;
wire n13318;
wire n13319;
wire n13320;
wire n13321;
wire n13322;
wire n13323;
wire n13324;
wire n13325;
wire n13326;
wire n13327;
wire n13328;
wire n13329;
wire n13330;
wire n13331;
wire n13332;
wire n13333;
wire n13334;
wire n13335;
wire n13336;
wire n13337;
wire n13338;
wire n13339;
wire n13340;
wire n13341;
wire n13342;
wire n13343;
wire n13344;
wire n13345;
wire n13346;
wire n13347;
wire n13348;
wire n13349;
wire n13350;
wire n13351;
wire n13352;
wire n13353;
wire n13354;
wire n13355;
wire n13356;
wire n13357;
wire n13358;
wire n13359;
wire n13360;
wire n13361;
wire n13362;
wire n13363;
wire n13364;
wire n13365;
wire n13366;
wire n13367;
wire n13368;
wire n13369;
wire n13370;
wire n13371;
wire n13372;
wire n13373;
wire n13374;
wire n13375;
wire n13376;
wire n13377;
wire n13378;
wire n13379;
wire n13380;
wire n13381;
wire n13382;
wire n13383;
wire n13384;
wire n13385;
wire n13386;
wire n13387;
wire n13388;
wire n13389;
wire n13390;
wire n13391;
wire n13392;
wire n13393;
wire n13394;
wire n13395;
wire n13396;
wire n13397;
wire n13398;
wire n13399;
wire n13400;
wire n13401;
wire n13402;
wire n13404;
wire n13405;
wire n13407;
wire n13408;
wire n13409;
wire n13410;
wire n13411;
wire n13412;
wire n13413;
wire n13414;
wire n13415;
wire n13416;
wire n13417;
wire n13418;
wire n13419;
wire n13420;
wire n13421;
wire n13422;
wire n13423;
wire n13424;
wire n13425;
wire n13426;
wire n13427;
wire n13428;
wire n13429;
wire n13430;
wire n13431;
wire n13432;
wire n13433;
wire n13434;
wire n13435;
wire n13436;
wire n13437;
wire n13438;
wire n13439;
wire n13440;
wire n13441;
wire n13442;
wire n13443;
wire n13444;
wire n13445;
wire n13446;
wire n13447;
wire n13448;
wire n13449;
wire n13450;
wire n13451;
wire n13452;
wire n13453;
wire n13454;
wire n13455;
wire n13456;
wire n13457;
wire n13458;
wire n13459;
wire n13460;
wire n13461;
wire n13462;
wire n13463;
wire n13464;
wire n13465;
wire n13466;
wire n13467;
wire n13468;
wire n13469;
wire n13470;
wire n13471;
wire n13472;
wire n13473;
wire n13474;
wire n13475;
wire n13476;
wire n13477;
wire n13478;
wire n13479;
wire n13480;
wire n13481;
wire n13482;
wire n13483;
wire n13484;
wire n13485;
wire n13486;
wire n13487;
wire n13488;
wire n13489;
wire n13490;
wire n13491;
wire n13492;
wire n13493;
wire n13494;
wire n13495;
wire n13496;
wire n13497;
wire n13498;
wire n13499;
wire n13500;
wire n13501;
wire n13502;
wire n13503;
wire n13504;
wire n13505;
wire n13506;
wire n13507;
wire n13508;
wire n13509;
wire n13510;
wire n13512;
wire n13513;
wire n13515;
wire n13516;
wire n13517;
wire n13518;
wire n13519;
wire n13520;
wire n13521;
wire n13522;
wire n13523;
wire n13524;
wire n13525;
wire n13526;
wire n13527;
wire n13528;
wire n13529;
wire n13530;
wire n13531;
wire n13532;
wire n13533;
wire n13534;
wire n13535;
wire n13536;
wire n13537;
wire n13538;
wire n13539;
wire n13540;
wire n13541;
wire n13542;
wire n13543;
wire n13544;
wire n13545;
wire n13546;
wire n13547;
wire n13548;
wire n13549;
wire n13550;
wire n13551;
wire n13552;
wire n13553;
wire n13554;
wire n13555;
wire n13556;
wire n13557;
wire n13558;
wire n13559;
wire n13560;
wire n13561;
wire n13562;
wire n13563;
wire n13564;
wire n13565;
wire n13566;
wire n13567;
wire n13568;
wire n13569;
wire n13570;
wire n13571;
wire n13572;
wire n13573;
wire n13574;
wire n13575;
wire n13576;
wire n13577;
wire n13578;
wire n13579;
wire n13580;
wire n13581;
wire n13582;
wire n13583;
wire n13584;
wire n13585;
wire n13586;
wire n13587;
wire n13588;
wire n13589;
wire n13590;
wire n13591;
wire n13592;
wire n13593;
wire n13594;
wire n13595;
wire n13596;
wire n13597;
wire n13598;
wire n13599;
wire n13600;
wire n13601;
wire n13602;
wire n13603;
wire n13604;
wire n13605;
wire n13606;
wire n13607;
wire n13608;
wire n13609;
wire n13610;
wire n13611;
wire n13612;
wire n13613;
wire n13614;
wire n13615;
wire n13616;
wire n13617;
wire n13618;
wire n13620;
wire n13621;
wire n13623;
wire n13624;
wire n13625;
wire n13626;
wire n13627;
wire n13628;
wire n13629;
wire n13630;
wire n13631;
wire n13632;
wire n13633;
wire n13634;
wire n13635;
wire n13636;
wire n13637;
wire n13638;
wire n13639;
wire n13640;
wire n13641;
wire n13642;
wire n13643;
wire n13644;
wire n13645;
wire n13646;
wire n13647;
wire n13648;
wire n13649;
wire n13650;
wire n13651;
wire n13652;
wire n13653;
wire n13654;
wire n13655;
wire n13656;
wire n13657;
wire n13658;
wire n13659;
wire n13660;
wire n13661;
wire n13662;
wire n13663;
wire n13664;
wire n13665;
wire n13666;
wire n13667;
wire n13668;
wire n13669;
wire n13670;
wire n13671;
wire n13672;
wire n13673;
wire n13674;
wire n13675;
wire n13676;
wire n13677;
wire n13678;
wire n13679;
wire n13680;
wire n13681;
wire n13682;
wire n13683;
wire n13684;
wire n13685;
wire n13686;
wire n13687;
wire n13688;
wire n13689;
wire n13690;
wire n13691;
wire n13692;
wire n13693;
wire n13694;
wire n13695;
wire n13696;
wire n13697;
wire n13698;
wire n13699;
wire n13700;
wire n13701;
wire n13702;
wire n13703;
wire n13704;
wire n13705;
wire n13706;
wire n13707;
wire n13708;
wire n13709;
wire n13710;
wire n13711;
wire n13712;
wire n13713;
wire n13714;
wire n13715;
wire n13716;
wire n13717;
wire n13718;
wire n13719;
wire n13720;
wire n13721;
wire n13722;
wire n13723;
wire n13724;
wire n13725;
wire n13727;
wire n13728;
wire n13730;
wire n13731;
wire n13732;
wire n13733;
wire n13734;
wire n13735;
wire n13736;
wire n13737;
wire n13738;
wire n13739;
wire n13740;
wire n13741;
wire n13742;
wire n13743;
wire n13744;
wire n13745;
wire n13746;
wire n13747;
wire n13748;
wire n13749;
wire n13750;
wire n13751;
wire n13752;
wire n13753;
wire n13754;
wire n13755;
wire n13756;
wire n13757;
wire n13758;
wire n13759;
wire n13760;
wire n13761;
wire n13762;
wire n13763;
wire n13764;
wire n13765;
wire n13766;
wire n13767;
wire n13768;
wire n13769;
wire n13770;
wire n13771;
wire n13772;
wire n13773;
wire n13774;
wire n13775;
wire n13776;
wire n13777;
wire n13778;
wire n13779;
wire n13780;
wire n13781;
wire n13782;
wire n13783;
wire n13784;
wire n13785;
wire n13786;
wire n13787;
wire n13788;
wire n13789;
wire n13790;
wire n13791;
wire n13792;
wire n13793;
wire n13794;
wire n13795;
wire n13796;
wire n13797;
wire n13798;
wire n13799;
wire n13800;
wire n13801;
wire n13802;
wire n13803;
wire n13804;
wire n13805;
wire n13806;
wire n13807;
wire n13808;
wire n13809;
wire n13810;
wire n13811;
wire n13812;
wire n13813;
wire n13814;
wire n13815;
wire n13816;
wire n13817;
wire n13818;
wire n13819;
wire n13820;
wire n13821;
wire n13822;
wire n13823;
wire n13824;
wire n13825;
wire n13826;
wire n13827;
wire n13828;
wire n13829;
wire n13830;
wire n13831;
wire n13832;
wire n13833;
wire n13834;
wire n13835;
wire n13836;
wire n13837;
wire n13838;
wire n13839;
wire n13840;
wire n13841;
wire n13842;
wire n13843;
wire n13844;
wire n13845;
wire n13846;
wire n13847;
wire n13848;
wire n13849;
wire n13850;
wire n13851;
wire n13852;
wire n13853;
wire n13854;
wire n13855;
wire n13856;
wire n13857;
wire n13858;
wire n13859;
wire n13860;
wire n13861;
wire n13862;
wire n13863;
wire n13864;
wire n13865;
wire n13866;
wire n13867;
wire n13868;
wire n13869;
wire n13870;
wire n13871;
wire n13872;
wire n13873;
wire n13874;
wire n13875;
wire n13876;
wire n13877;
wire n13878;
wire n13879;
wire n13880;
wire n13881;
wire n13882;
wire n13883;
wire n13884;
wire n13885;
wire n13886;
wire n13887;
wire n13889;
wire n13891;
wire n13893;
wire n13895;
wire n13897;
wire n13898;
wire n13900;
wire n13901;
wire n13902;
wire n13903;
wire n13904;
wire n13905;
wire n13907;
wire n13910;
wire n13911;
wire n13913;
wire n13914;
wire n13915;
wire n13916;
wire n13917;
wire n13918;
wire n13920;
wire n13921;
wire n13923;
wire n13924;
wire n13925;
wire n13926;
wire n13928;
wire n13929;
wire n13930;
wire n13931;
wire n13932;
wire n13933;
wire n13935;
wire n13936;
wire n13937;
wire n13938;
wire n13939;
wire n13940;
wire n13941;
wire n13942;
wire n13943;
wire n13944;
wire n13945;
wire n13946;
wire n13947;
wire n13948;
wire n13949;
wire n13950;
wire n13951;
wire n13952;
wire n13953;
wire n13955;
wire n13957;
wire n13959;
wire n13961;
wire n13963;
wire n13965;
wire n13967;
wire n13969;
wire n13971;
wire n13973;
wire n13975;
wire n13977;
wire n13979;
wire n13981;
wire n13983;
wire n13985;
wire n13986;
wire n13987;
wire n13988;
wire n13990;
wire n13991;
wire n13992;
wire n13993;
wire n13994;
wire n13995;
wire n13996;
wire n13998;
wire n13999;
wire n14000;
wire n14001;
wire n14003;
wire n14004;
wire n14005;
wire n14006;
wire n14007;
wire n14009;
wire n14011;
wire n14013;
wire n14015;
wire n14017;
wire n14019;
wire n14021;
wire n14023;
wire n14025;
wire n14027;
wire n14029;
wire n14031;
wire n14033;
wire n14035;
wire n14037;
wire n14039;
wire n14040;
wire n14041;
wire n14042;
wire n14044;
wire n14046;
wire n14048;
wire n14050;
wire n14052;
wire n14054;
wire n14056;
wire n14058;
wire n14060;
wire n14062;
wire n14064;
wire n14066;
wire n14068;
wire n14070;
wire n14072;
wire n14074;
wire n14075;
wire n14076;
wire n14078;
wire n14080;
wire n14082;
wire n14084;
wire n14086;
wire n14088;
wire n14090;
wire n14092;
wire n14094;
wire n14096;
wire n14098;
wire n14100;
wire n14102;
wire n14104;
wire n14106;
wire n14108;
wire n14109;
wire n14110;
wire n14111;
wire n14112;
wire n14113;
wire n14116;
wire n14117;
wire n14118;
wire n14119;
wire n14120;
wire n14123;
wire n14124;
wire n14125;
wire n14126;
wire n14131;
wire n14132;
wire n14133;
wire n14134;
wire n14135;
wire n14136;
wire n14137;
wire n14138;
wire n14139;
wire n14140;
wire n14141;
wire n14142;
wire n14143;
wire n14144;
wire n14145;
wire n14147;
wire n14148;
wire n14149;
wire n14150;
wire n14151;
wire n14152;
wire n14153;
wire n14154;
wire n14156;
wire n14157;
wire n14158;
wire n14159;
wire n14160;
wire n14161;
wire n14162;
wire n14163;
wire n14164;
wire n14165;
wire n14166;
wire n14167;
wire n14168;
wire n14169;
wire n14171;
wire n14172;
wire n14173;
wire n14174;
wire n14176;
wire n14177;
wire n14178;
wire n14179;
wire n14180;
wire n14181;
wire n14182;
wire n14183;
wire n14184;
wire n14185;
wire n14186;
wire n14187;
wire n14188;
wire n14189;
wire n14190;
wire n14191;
wire n14192;
wire n14193;
wire n14194;
wire n14195;
wire n14196;
wire n14197;
wire n14199;
wire n14200;
wire n14201;
wire n14203;
wire n14205;
wire n14206;
wire n14207;
wire n14208;
wire n14210;
wire n14211;
wire n14212;
wire n14217;
wire n14218;
wire n14221;
wire n14224;
wire n14225;
wire n14226;
wire n14227;
wire n14228;
wire n14229;
wire n14230;
wire n14231;
wire n14232;
wire n14233;
wire n14234;
wire n14235;
wire n14236;
wire n14237;
wire n14238;
wire n14239;
wire n14241;
wire n14242;
wire n14243;
wire n14244;
wire n14245;
wire n14246;
wire n14247;
wire n14248;
wire n14249;
wire n14250;
wire n14251;
wire n14252;
wire n14254;
wire n14255;
wire n14256;
wire n14257;
wire n14258;
wire n14259;
wire n14260;
wire n14261;
wire n14262;
wire n14263;
wire n14264;
wire n14265;
wire n14266;
wire n14267;
wire n14268;
wire n14269;
wire n14270;
wire n14271;
wire n14272;
wire n14273;
wire n14274;
wire n14275;
wire n14276;
wire n14277;
wire n14278;
wire n14279;
wire n14280;
wire n14281;
wire n14282;
wire n14283;
wire n14284;
wire n14286;
wire n14288;
wire n14289;
wire n14291;
wire n14293;
wire n14294;
wire n14295;
wire n14296;
wire n14297;
wire n14298;
wire n14299;
wire n14300;
wire n14301;
wire n14303;
wire n14305;
wire n14306;
wire n14308;
wire n14310;
wire n14311;
wire n14312;
wire n14313;
wire n14315;
wire n14316;
wire n14317;
wire n14318;
wire n14319;
wire n14321;
wire n14322;
wire n14324;
wire n14325;
wire n14326;
wire n14327;
wire n14328;
wire n14329;
wire n14330;
wire n14331;
wire n14332;
wire n14333;
wire n14334;
wire n14335;
wire n14336;
wire n14337;
wire n14338;
wire n14339;
wire n14340;
wire n14342;
wire n14343;
wire n14344;
wire n14345;
wire n14346;
wire n14347;
wire n14348;
wire n14349;
wire n14350;
wire n14352;
wire n14353;
wire n14355;
wire n14356;
wire n14358;
wire n14359;
wire n14361;
wire n14362;
wire n14363;
wire n14364;
wire n14365;
wire n14366;
wire n14367;
wire n14368;
wire n14369;
wire n14370;
wire n14371;
wire n14372;
wire n14374;
wire n14375;
wire n14376;
wire n14377;
wire n14378;
wire n14379;
wire n14380;
wire n14381;
wire n14382;
wire n14383;
wire n14384;
wire n14385;
wire n14386;
wire n14387;
wire n14388;
wire n14389;
wire n14390;
wire n14391;
wire n14393;
wire n14394;
wire n14395;
wire n14396;
wire n14397;
wire n14398;
wire n14399;
wire n14400;
wire n14401;
wire n14402;
wire n14403;
wire n14404;
wire n14405;
wire n14406;
wire n14407;
wire n14408;
wire n14409;
wire n14410;
wire n14412;
wire n14413;
wire n14414;
wire n14415;
wire n14416;
wire n14417;
wire n14418;
wire n14419;
wire n14421;
wire n14422;
wire n14423;
wire n14424;
wire n14425;
wire n14426;
wire n14427;
wire n14429;
wire n14430;
wire n14431;
wire n14432;
wire n14433;
wire n14434;
wire n14435;
wire n14437;
wire n14438;
wire n14439;
wire n14440;
wire n14442;
wire n14443;
wire n14444;
wire n14445;
wire n14446;
wire n14447;
wire n14448;
wire n14449;
wire n14450;
wire n14451;
wire n14452;
wire n14453;
wire n14454;
wire n14455;
wire n14456;
wire n14457;
wire n14458;
wire n14459;
wire n14460;
wire n14462;
wire n14464;
wire n14466;
wire n14468;
wire n14469;
wire n14470;
wire n14472;
wire n14473;
wire n14475;
wire n14476;
wire n14477;
wire n14478;
wire n14479;
wire n14481;
wire n14482;
wire n14483;
wire n14484;
wire n14485;
wire n14487;
wire n14488;
wire n14489;
wire n14490;
wire n14491;
wire n14492;
wire n14493;
wire n14494;
wire n14495;
wire n14496;
wire n14497;
wire n14498;
wire n14499;
wire n14500;
wire n14501;
wire n14502;
wire n14503;
wire n14504;
wire n14505;
wire n14506;
wire n14508;
wire n14509;
wire n14511;
wire n14512;
wire n14513;
wire n14514;
wire n14515;
wire n14516;
wire n14517;
wire n14518;
wire n14519;
wire n14520;
wire n14521;
wire n14522;
wire n14523;
wire n14525;
wire n14527;
wire n14529;
wire n14531;
wire n14532;
wire n14533;
wire n14535;
wire n14536;
wire n14537;
wire n14538;
wire n14539;
wire n14540;
wire n14542;
wire n14543;
wire n14544;
wire n14545;
wire n14546;
wire n14548;
wire n14549;
wire n14550;
wire n14551;
wire n14552;
wire n14553;
wire n14554;
wire n14555;
wire n14558;
wire n14559;
wire n14560;
wire n14561;
wire n14563;
wire n14564;
wire n14565;
wire n14566;
wire n14567;
wire n14568;
wire n14569;
wire n14570;
wire n14571;
wire n14572;
wire n14573;
wire n14574;
wire n14575;
wire n14576;
wire n14577;
wire n14578;
wire n14579;
wire n14580;
wire n14581;
wire n14583;
wire n14585;
wire n14587;
wire n14589;
wire n14590;
wire n14591;
wire n14593;
wire n14594;
wire n14596;
wire n14597;
wire n14598;
wire n14599;
wire n14600;
wire n14602;
wire n14603;
wire n14604;
wire n14605;
wire n14606;
wire n14608;
wire n14609;
wire n14610;
wire n14611;
wire n14612;
wire n14613;
wire n14614;
wire n14615;
wire n14616;
wire n14617;
wire n14619;
wire n14620;
wire n14621;
wire n14622;
wire n14623;
wire n14624;
wire n14625;
wire n14626;
wire n14627;
wire n14628;
wire n14629;
wire n14630;
wire n14631;
wire n14632;
wire n14633;
wire n14634;
wire n14635;
wire n14636;
wire n14637;
wire n14638;
wire n14639;
wire n14640;
wire n14641;
wire n14643;
wire n14644;
wire n14646;
wire n14647;
wire n14649;
wire n14651;
wire n14652;
wire n14653;
wire n14654;
wire n14655;
wire n14656;
wire n14657;
wire n14658;
wire n14659;
wire n14661;
wire n14663;
wire n14664;
wire n14666;
wire n14668;
wire n14669;
wire n14670;
wire n14671;
wire n14672;
wire n14673;
wire n14674;
wire n14675;
wire n14677;
wire n14679;
wire n14680;
wire n14682;
wire n14684;
wire n14685;
wire n14686;
wire n14687;
wire n14688;
wire n14689;
wire n14690;
wire n14691;
wire n14693;
wire n14695;
wire n14696;
wire n14698;
wire n14700;
wire n14701;
wire n14702;
wire n14703;
wire n14704;
wire n14705;
wire n14706;
wire n14707;
wire n14709;
wire n14711;
wire n14712;
wire n14714;
wire n14716;
wire n14717;
wire n14718;
wire n14719;
wire n14720;
wire n14721;
wire n14722;
wire n14723;
wire n14724;
wire n14726;
wire n14728;
wire n14730;
wire n14732;
wire n14733;
wire n14734;
wire n14736;
wire n14737;
wire n14739;
wire n14740;
wire n14741;
wire n14742;
wire n14743;
wire n14745;
wire n14746;
wire n14747;
wire n14748;
wire n14749;
wire n14751;
wire n14752;
wire n14753;
wire n14754;
wire n14755;
wire n14756;
wire n14757;
wire n14758;
wire n14759;
wire n14761;
wire n14762;
wire n14763;
wire n14764;
wire n14765;
wire n14766;
wire n14768;
wire n14769;
wire n14770;
wire n14771;
wire n14772;
wire n14773;
wire n14774;
wire n14775;
wire n14776;
wire n14777;
wire n14778;
wire n14779;
wire n14781;
wire n14782;
wire n14783;
wire n14784;
wire n14785;
wire n14786;
wire n14788;
wire n14790;
wire n14791;
wire n14792;
wire n14793;
wire n14794;
wire n14795;
wire n14797;
wire n14799;
wire n14801;
wire n14803;
wire n14804;
wire n14805;
wire n14807;
wire n14808;
wire n14809;
wire n14810;
wire n14811;
wire n14812;
wire n14814;
wire n14815;
wire n14816;
wire n14817;
wire n14818;
wire n14820;
wire n14821;
wire n14822;
wire n14823;
wire n14824;
wire n14825;
wire n14827;
wire n14829;
wire n14831;
wire n14833;
wire n14834;
wire n14835;
wire n14837;
wire n14838;
wire n14840;
wire n14841;
wire n14842;
wire n14843;
wire n14844;
wire n14846;
wire n14847;
wire n14848;
wire n14849;
wire n14850;
wire n14852;
wire n14853;
wire n14854;
wire n14856;
wire n14858;
wire n14860;
wire n14861;
wire n14862;
wire n14863;
wire n14864;
wire n14866;
wire n14867;
wire n14869;
wire n14871;
wire n14873;
wire n14875;
wire n14877;
wire n14878;
wire n14879;
wire n14882;
wire n14883;
wire n14884;
wire n14885;
wire n14886;
wire n14887;
wire n14888;
wire n14889;
wire n14890;
wire n14892;
wire n14894;
wire n14895;
wire n14896;
wire n14897;
wire n14898;
wire n14899;
wire n14900;
wire n14901;
wire n14902;
wire n14903;
wire n14905;
wire n14906;
wire n14907;
wire n14908;
wire n14910;
wire n14911;
wire n14912;
wire n14913;
wire n14914;
wire n14915;
wire n14916;
wire n14917;
wire n14918;
wire n14919;
wire n14920;
wire n14921;
wire n14922;
wire n14923;
wire n14924;
wire n14926;
wire n14928;
wire n14930;
wire n14932;
wire n14933;
wire n14934;
wire n14936;
wire n14937;
wire n14939;
wire n14940;
wire n14941;
wire n14942;
wire n14943;
wire n14945;
wire n14946;
wire n14947;
wire n14948;
wire n14949;
wire n14951;
wire n14952;
wire n14953;
wire n14954;
wire n14955;
wire n14956;
wire n14957;
wire n14958;
wire n14959;
wire n14960;
wire n14962;
wire n14963;
wire n14964;
wire n14965;
wire n14966;
wire n14967;
wire n14968;
wire n14969;
wire n14970;
wire n14971;
wire n14972;
wire n14973;
wire n14974;
wire n14975;
wire n14976;
wire n14977;
wire n14979;
wire n14981;
wire n14983;
wire n14984;
wire n14985;
wire n14986;
wire n14987;
wire n14989;
wire n14990;
wire n14992;
wire n14994;
wire n14996;
wire n14998;
wire n15000;
wire n15001;
wire n15002;
wire n15005;
wire n15006;
wire n15007;
wire n15008;
wire n15009;
wire n15010;
wire n15011;
wire n15012;
wire n15013;
wire n15014;
wire n15015;
wire n15016;
wire n15018;
wire n15020;
wire n15021;
wire n15023;
wire n15025;
wire n15026;
wire n15027;
wire n15028;
wire n15029;
wire n15030;
wire n15032;
wire n15033;
wire n15035;
wire n15037;
wire n15038;
wire n15039;
wire n15040;
wire n15041;
wire n15042;
wire n15043;
wire n15045;
wire n15047;
wire n15048;
wire n15050;
wire n15052;
wire n15053;
wire n15054;
wire n15055;
wire n15056;
wire n15057;
wire n15058;
wire n15059;
wire n15060;
wire n15062;
wire n15064;
wire n15065;
wire n15067;
wire n15069;
wire n15070;
wire n15071;
wire n15072;
wire n15073;
wire n15074;
wire n15075;
wire n15076;
wire n15078;
wire n15080;
wire n15081;
wire n15083;
wire n15085;
wire n15086;
wire n15087;
wire n15088;
wire n15089;
wire n15090;
wire n15091;
wire n15092;
wire n15093;
wire n15094;
wire n15095;
wire n15096;
wire n15098;
wire n15099;
wire n15101;
wire n15102;
wire n15103;
wire n15104;
wire n15105;
wire n15106;
wire n15108;
wire n15109;
wire n15110;
wire n15112;
wire n15114;
wire n15115;
wire n15116;
wire n15118;
wire n15119;
wire n15120;
wire n15121;
wire n15122;
wire n15123;
wire n15125;
wire n15127;
wire n15129;
wire n15131;
wire n15132;
wire n15133;
wire n15135;
wire n15136;
wire n15138;
wire n15139;
wire n15140;
wire n15141;
wire n15142;
wire n15144;
wire n15145;
wire n15146;
wire n15147;
wire n15148;
wire n15150;
wire n15151;
wire n15152;
wire n15153;
wire n15154;
wire n15155;
wire n15157;
wire n15159;
wire n15161;
wire n15163;
wire n15164;
wire n15165;
wire n15167;
wire n15168;
wire n15170;
wire n15171;
wire n15172;
wire n15173;
wire n15174;
wire n15176;
wire n15177;
wire n15178;
wire n15179;
wire n15180;
wire n15182;
wire n15183;
wire n15184;
wire n15186;
wire n15187;
wire n15189;
wire n15190;
wire n15191;
wire n15192;
wire n15193;
wire n15194;
wire n15195;
wire n15197;
wire n15199;
wire n15201;
wire n15203;
wire n15204;
wire n15205;
wire n15207;
wire n15208;
wire n15209;
wire n15210;
wire n15211;
wire n15212;
wire n15214;
wire n15215;
wire n15216;
wire n15217;
wire n15218;
wire n15220;
wire n15221;
wire n15222;
wire n15223;
wire n15224;
wire n15225;
wire n15226;
wire n15227;
wire n15229;
wire n15230;
wire n15231;
wire n15232;
wire n15234;
wire n15235;
wire n15236;
wire n15237;
wire n15238;
wire n15239;
wire n15240;
wire n15241;
wire n15242;
wire n15243;
wire n15244;
wire n15245;
wire n15246;
wire n15247;
wire n15248;
wire n15250;
wire n15252;
wire n15254;
wire n15256;
wire n15257;
wire n15258;
wire n15260;
wire n15261;
wire n15263;
wire n15264;
wire n15265;
wire n15266;
wire n15267;
wire n15269;
wire n15270;
wire n15271;
wire n15272;
wire n15273;
wire n15275;
wire n15276;
wire n15277;
wire n15278;
wire n15279;
wire n15280;
wire n15281;
wire n15282;
wire n15283;
wire n15284;
wire n15286;
wire n15287;
wire n15288;
wire n15289;
wire n15290;
wire n15291;
wire n15292;
wire n15293;
wire n15294;
wire n15295;
wire n15296;
wire n15297;
wire n15298;
wire n15299;
wire n15300;
wire n15301;
wire n15302;
wire n15303;
wire n15304;
wire n15305;
wire n15307;
wire n15308;
wire n15310;
wire n15311;
wire n15313;
wire n15315;
wire n15316;
wire n15317;
wire n15318;
wire n15319;
wire n15320;
wire n15321;
wire n15322;
wire n15323;
wire n15325;
wire n15327;
wire n15328;
wire n15330;
wire n15332;
wire n15333;
wire n15334;
wire n15335;
wire n15336;
wire n15337;
wire n15338;
wire n15339;
wire n15341;
wire n15343;
wire n15344;
wire n15346;
wire n15348;
wire n15349;
wire n15350;
wire n15351;
wire n15352;
wire n15353;
wire n15354;
wire n15355;
wire n15357;
wire n15359;
wire n15360;
wire n15362;
wire n15364;
wire n15365;
wire n15366;
wire n15367;
wire n15368;
wire n15369;
wire n15370;
wire n15371;
wire n15373;
wire n15375;
wire n15376;
wire n15378;
wire n15380;
wire n15381;
wire n15382;
wire n15383;
wire n15384;
wire n15385;
wire n15386;
wire n15387;
wire n15389;
wire n15391;
wire n15393;
wire n15395;
wire n15396;
wire n15397;
wire n15399;
wire n15400;
wire n15402;
wire n15403;
wire n15404;
wire n15405;
wire n15406;
wire n15408;
wire n15409;
wire n15410;
wire n15411;
wire n15412;
wire n15414;
wire n15415;
wire n15416;
wire n15417;
wire n15418;
wire n15419;
wire n15420;
wire n15421;
wire n15422;
wire n15424;
wire n15425;
wire n15426;
wire n15427;
wire n15428;
wire n15429;
wire n15431;
wire n15432;
wire n15433;
wire n15434;
wire n15435;
wire n15436;
wire n15437;
wire n15438;
wire n15439;
wire n15440;
wire n15441;
wire n15442;
wire n15444;
wire n15445;
wire n15446;
wire n15447;
wire n15448;
wire n15449;
wire n15451;
wire n15453;
wire n15454;
wire n15455;
wire n15456;
wire n15457;
wire n15458;
wire n15460;
wire n15462;
wire n15464;
wire n15466;
wire n15467;
wire n15468;
wire n15470;
wire n15471;
wire n15472;
wire n15473;
wire n15474;
wire n15475;
wire n15477;
wire n15478;
wire n15479;
wire n15480;
wire n15481;
wire n15483;
wire n15484;
wire n15485;
wire n15486;
wire n15487;
wire n15488;
wire n15490;
wire n15492;
wire n15494;
wire n15496;
wire n15497;
wire n15498;
wire n15500;
wire n15501;
wire n15503;
wire n15504;
wire n15505;
wire n15506;
wire n15507;
wire n15509;
wire n15510;
wire n15511;
wire n15512;
wire n15513;
wire n15515;
wire n15516;
wire n15517;
wire n15518;
wire n15520;
wire n15522;
wire n15524;
wire n15525;
wire n15526;
wire n15527;
wire n15528;
wire n15530;
wire n15531;
wire n15533;
wire n15535;
wire n15537;
wire n15539;
wire n15541;
wire n15542;
wire n15543;
wire n15546;
wire n15547;
wire n15548;
wire n15549;
wire n15550;
wire n15551;
wire n15552;
wire n15553;
wire n15554;
wire n15556;
wire n15558;
wire n15559;
wire n15560;
wire n15561;
wire n15562;
wire n15563;
wire n15564;
wire n15565;
wire n15566;
wire n15567;
wire n15569;
wire n15570;
wire n15571;
wire n15572;
wire n15574;
wire n15575;
wire n15576;
wire n15577;
wire n15578;
wire n15579;
wire n15580;
wire n15581;
wire n15582;
wire n15583;
wire n15584;
wire n15585;
wire n15586;
wire n15587;
wire n15588;
wire n15590;
wire n15592;
wire n15594;
wire n15596;
wire n15597;
wire n15598;
wire n15600;
wire n15601;
wire n15603;
wire n15604;
wire n15605;
wire n15606;
wire n15607;
wire n15609;
wire n15610;
wire n15611;
wire n15612;
wire n15613;
wire n15615;
wire n15616;
wire n15617;
wire n15618;
wire n15619;
wire n15620;
wire n15621;
wire n15622;
wire n15623;
wire n15624;
wire n15626;
wire n15627;
wire n15628;
wire n15629;
wire n15630;
wire n15631;
wire n15632;
wire n15633;
wire n15634;
wire n15635;
wire n15636;
wire n15637;
wire n15638;
wire n15639;
wire n15640;
wire n15641;
wire n15642;
wire n15643;
wire n15644;
wire n15646;
wire n15647;
wire n15649;
wire n15650;
wire n15652;
wire n15654;
wire n15655;
wire n15656;
wire n15657;
wire n15658;
wire n15659;
wire n15660;
wire n15661;
wire n15662;
wire n15664;
wire n15666;
wire n15667;
wire n15669;
wire n15671;
wire n15672;
wire n15673;
wire n15674;
wire n15675;
wire n15676;
wire n15677;
wire n15678;
wire n15680;
wire n15682;
wire n15683;
wire n15685;
wire n15687;
wire n15688;
wire n15689;
wire n15690;
wire n15691;
wire n15692;
wire n15693;
wire n15694;
wire n15696;
wire n15698;
wire n15699;
wire n15701;
wire n15703;
wire n15704;
wire n15705;
wire n15706;
wire n15707;
wire n15708;
wire n15709;
wire n15710;
wire n15712;
wire n15714;
wire n15715;
wire n15717;
wire n15719;
wire n15720;
wire n15721;
wire n15722;
wire n15723;
wire n15724;
wire n15725;
wire n15726;
wire n15728;
wire n15730;
wire n15732;
wire n15734;
wire n15735;
wire n15736;
wire n15738;
wire n15739;
wire n15741;
wire n15742;
wire n15743;
wire n15744;
wire n15745;
wire n15747;
wire n15748;
wire n15749;
wire n15750;
wire n15751;
wire n15753;
wire n15754;
wire n15755;
wire n15756;
wire n15757;
wire n15758;
wire n15759;
wire n15760;
wire n15761;
wire n15763;
wire n15764;
wire n15765;
wire n15766;
wire n15767;
wire n15768;
wire n15770;
wire n15771;
wire n15772;
wire n15773;
wire n15774;
wire n15775;
wire n15776;
wire n15777;
wire n15778;
wire n15779;
wire n15780;
wire n15781;
wire n15783;
wire n15784;
wire n15785;
wire n15786;
wire n15787;
wire n15788;
wire n15790;
wire n15792;
wire n15793;
wire n15794;
wire n15795;
wire n15796;
wire n15797;
wire n15799;
wire n15801;
wire n15803;
wire n15805;
wire n15806;
wire n15807;
wire n15809;
wire n15810;
wire n15811;
wire n15812;
wire n15813;
wire n15814;
wire n15816;
wire n15817;
wire n15818;
wire n15819;
wire n15820;
wire n15822;
wire n15823;
wire n15824;
wire n15825;
wire n15826;
wire n15827;
wire n15829;
wire n15831;
wire n15833;
wire n15835;
wire n15836;
wire n15837;
wire n15839;
wire n15840;
wire n15842;
wire n15843;
wire n15844;
wire n15845;
wire n15846;
wire n15848;
wire n15849;
wire n15850;
wire n15851;
wire n15852;
wire n15854;
wire n15855;
wire n15856;
wire n15857;
wire n15859;
wire n15861;
wire n15863;
wire n15864;
wire n15865;
wire n15866;
wire n15867;
wire n15869;
wire n15870;
wire n15872;
wire n15874;
wire n15876;
wire n15878;
wire n15880;
wire n15881;
wire n15882;
wire n15885;
wire n15886;
wire n15887;
wire n15888;
wire n15889;
wire n15890;
wire n15891;
wire n15892;
wire n15893;
wire n15895;
wire n15897;
wire n15898;
wire n15899;
wire n15900;
wire n15901;
wire n15902;
wire n15903;
wire n15904;
wire n15905;
wire n15906;
wire n15908;
wire n15909;
wire n15910;
wire n15911;
wire n15913;
wire n15914;
wire n15915;
wire n15916;
wire n15917;
wire n15918;
wire n15919;
wire n15920;
wire n15921;
wire n15922;
wire n15923;
wire n15924;
wire n15925;
wire n15926;
wire n15927;
wire n15929;
wire n15931;
wire n15933;
wire n15935;
wire n15936;
wire n15937;
wire n15939;
wire n15940;
wire n15942;
wire n15943;
wire n15944;
wire n15945;
wire n15946;
wire n15948;
wire n15949;
wire n15950;
wire n15951;
wire n15952;
wire n15954;
wire n15955;
wire n15956;
wire n15957;
wire n15958;
wire n15959;
wire n15960;
wire n15961;
wire n15962;
wire n15963;
wire n15965;
wire n15966;
wire n15967;
wire n15968;
wire n15969;
wire n15970;
wire n15971;
wire n15972;
wire n15973;
wire n15974;
wire n15975;
wire n15976;
wire n15977;
wire n15978;
wire n15979;
wire n15980;
wire n15981;
wire n15982;
wire n15983;
wire n15984;
wire n15986;
wire n15987;
wire n15989;
wire n15990;
wire n15992;
wire n15994;
wire n15995;
wire n15996;
wire n15997;
wire n15998;
wire n15999;
wire n16000;
wire n16001;
wire n16002;
wire n16004;
wire n16006;
wire n16007;
wire n16009;
wire n16011;
wire n16012;
wire n16013;
wire n16014;
wire n16015;
wire n16016;
wire n16017;
wire n16018;
wire n16020;
wire n16022;
wire n16023;
wire n16025;
wire n16027;
wire n16028;
wire n16029;
wire n16030;
wire n16031;
wire n16032;
wire n16033;
wire n16034;
wire n16036;
wire n16038;
wire n16039;
wire n16041;
wire n16043;
wire n16044;
wire n16045;
wire n16046;
wire n16047;
wire n16048;
wire n16049;
wire n16050;
wire n16052;
wire n16054;
wire n16055;
wire n16057;
wire n16059;
wire n16060;
wire n16061;
wire n16062;
wire n16063;
wire n16064;
wire n16065;
wire n16066;
wire n16068;
wire n16070;
wire n16072;
wire n16074;
wire n16075;
wire n16076;
wire n16078;
wire n16079;
wire n16081;
wire n16082;
wire n16083;
wire n16084;
wire n16085;
wire n16087;
wire n16088;
wire n16089;
wire n16090;
wire n16091;
wire n16093;
wire n16094;
wire n16095;
wire n16096;
wire n16097;
wire n16098;
wire n16099;
wire n16100;
wire n16101;
wire n16103;
wire n16104;
wire n16105;
wire n16106;
wire n16107;
wire n16108;
wire n16110;
wire n16111;
wire n16112;
wire n16113;
wire n16114;
wire n16115;
wire n16116;
wire n16117;
wire n16118;
wire n16119;
wire n16120;
wire n16121;
wire n16123;
wire n16124;
wire n16125;
wire n16126;
wire n16127;
wire n16128;
wire n16130;
wire n16132;
wire n16133;
wire n16134;
wire n16135;
wire n16136;
wire n16137;
wire n16139;
wire n16141;
wire n16143;
wire n16145;
wire n16146;
wire n16147;
wire n16149;
wire n16150;
wire n16151;
wire n16152;
wire n16153;
wire n16154;
wire n16156;
wire n16157;
wire n16158;
wire n16159;
wire n16160;
wire n16162;
wire n16163;
wire n16164;
wire n16165;
wire n16166;
wire n16167;
wire n16169;
wire n16171;
wire n16173;
wire n16175;
wire n16176;
wire n16177;
wire n16179;
wire n16180;
wire n16182;
wire n16183;
wire n16184;
wire n16185;
wire n16186;
wire n16188;
wire n16189;
wire n16190;
wire n16191;
wire n16192;
wire n16194;
wire n16195;
wire n16196;
wire n16197;
wire n16199;
wire n16201;
wire n16203;
wire n16204;
wire n16205;
wire n16206;
wire n16207;
wire n16209;
wire n16210;
wire n16212;
wire n16214;
wire n16216;
wire n16218;
wire n16220;
wire n16221;
wire n16222;
wire n16225;
wire n16226;
wire n16227;
wire n16228;
wire n16229;
wire n16230;
wire n16231;
wire n16232;
wire n16233;
wire n16235;
wire n16237;
wire n16238;
wire n16239;
wire n16240;
wire n16241;
wire n16242;
wire n16243;
wire n16244;
wire n16245;
wire n16246;
wire n16248;
wire n16249;
wire n16250;
wire n16251;
wire n16253;
wire n16254;
wire n16255;
wire n16256;
wire n16257;
wire n16258;
wire n16259;
wire n16260;
wire n16261;
wire n16262;
wire n16263;
wire n16264;
wire n16265;
wire n16266;
wire n16267;
wire n16269;
wire n16271;
wire n16273;
wire n16275;
wire n16276;
wire n16277;
wire n16279;
wire n16280;
wire n16282;
wire n16283;
wire n16284;
wire n16285;
wire n16286;
wire n16288;
wire n16289;
wire n16290;
wire n16291;
wire n16292;
wire n16294;
wire n16295;
wire n16296;
wire n16297;
wire n16298;
wire n16299;
wire n16300;
wire n16301;
wire n16302;
wire n16303;
wire n16305;
wire n16306;
wire n16307;
wire n16308;
wire n16309;
wire n16310;
wire n16311;
wire n16312;
wire n16313;
wire n16314;
wire n16315;
wire n16316;
wire n16317;
wire n16318;
wire n16319;
wire n16320;
wire n16321;
wire n16322;
wire n16323;
wire n16324;
wire n16326;
wire n16327;
wire n16329;
wire n16330;
wire n16332;
wire n16334;
wire n16335;
wire n16336;
wire n16337;
wire n16338;
wire n16339;
wire n16340;
wire n16341;
wire n16342;
wire n16344;
wire n16346;
wire n16347;
wire n16349;
wire n16351;
wire n16352;
wire n16353;
wire n16354;
wire n16355;
wire n16356;
wire n16357;
wire n16358;
wire n16360;
wire n16362;
wire n16363;
wire n16365;
wire n16367;
wire n16368;
wire n16369;
wire n16370;
wire n16371;
wire n16372;
wire n16373;
wire n16374;
wire n16376;
wire n16378;
wire n16379;
wire n16381;
wire n16383;
wire n16384;
wire n16385;
wire n16386;
wire n16387;
wire n16388;
wire n16389;
wire n16390;
wire n16392;
wire n16394;
wire n16395;
wire n16397;
wire n16399;
wire n16400;
wire n16401;
wire n16402;
wire n16403;
wire n16404;
wire n16405;
wire n16406;
wire n16408;
wire n16410;
wire n16412;
wire n16414;
wire n16415;
wire n16416;
wire n16418;
wire n16419;
wire n16421;
wire n16422;
wire n16423;
wire n16424;
wire n16425;
wire n16427;
wire n16428;
wire n16429;
wire n16430;
wire n16431;
wire n16433;
wire n16434;
wire n16435;
wire n16436;
wire n16437;
wire n16438;
wire n16439;
wire n16440;
wire n16441;
wire n16443;
wire n16444;
wire n16445;
wire n16446;
wire n16447;
wire n16448;
wire n16450;
wire n16451;
wire n16452;
wire n16453;
wire n16454;
wire n16455;
wire n16456;
wire n16457;
wire n16458;
wire n16459;
wire n16460;
wire n16461;
wire n16463;
wire n16464;
wire n16465;
wire n16466;
wire n16467;
wire n16468;
wire n16470;
wire n16472;
wire n16473;
wire n16474;
wire n16475;
wire n16476;
wire n16477;
wire n16479;
wire n16481;
wire n16483;
wire n16485;
wire n16486;
wire n16487;
wire n16489;
wire n16490;
wire n16491;
wire n16492;
wire n16493;
wire n16494;
wire n16496;
wire n16497;
wire n16498;
wire n16499;
wire n16500;
wire n16502;
wire n16503;
wire n16504;
wire n16505;
wire n16506;
wire n16507;
wire n16509;
wire n16511;
wire n16513;
wire n16515;
wire n16516;
wire n16517;
wire n16519;
wire n16520;
wire n16522;
wire n16523;
wire n16524;
wire n16525;
wire n16526;
wire n16528;
wire n16529;
wire n16530;
wire n16531;
wire n16532;
wire n16534;
wire n16535;
wire n16536;
wire n16537;
wire n16539;
wire n16541;
wire n16543;
wire n16544;
wire n16545;
wire n16546;
wire n16547;
wire n16549;
wire n16550;
wire n16552;
wire n16554;
wire n16556;
wire n16558;
wire n16560;
wire n16561;
wire n16562;
wire n16565;
wire n16566;
wire n16567;
wire n16568;
wire n16569;
wire n16570;
wire n16571;
wire n16572;
wire n16573;
wire n16575;
wire n16577;
wire n16578;
wire n16579;
wire n16580;
wire n16581;
wire n16582;
wire n16583;
wire n16584;
wire n16585;
wire n16586;
wire n16588;
wire n16589;
wire n16590;
wire n16591;
wire n16593;
wire n16594;
wire n16595;
wire n16596;
wire n16597;
wire n16598;
wire n16599;
wire n16600;
wire n16601;
wire n16602;
wire n16603;
wire n16604;
wire n16605;
wire n16606;
wire n16607;
wire n16608;
wire n16609;
wire n16613;
wire n16614;
wire n16615;
wire n16616;
wire n16617;
wire n16618;
wire n16619;
wire n16620;
wire n16621;
wire n16625;
wire n16626;
wire n16627;
wire n16628;
wire n16629;
wire n16630;
wire n16632;
wire n16633;
wire n16634;
wire n16635;
wire n16637;
wire n16638;
wire n16639;
wire n16640;
wire n16641;
wire n16642;
wire n16643;
wire n16644;
wire n16645;
wire n16646;
wire n16647;
wire n16648;
wire n16649;
wire n16650;
wire n16651;
wire n16652;
wire n16653;
wire n16654;
wire n16655;
wire n16656;
wire n16657;
wire n16658;
wire n16659;
wire n16660;
wire n16661;
wire n16662;
wire n16663;
wire n16664;
wire n16665;
wire n16666;
wire n16667;
wire n16668;
wire n16669;
wire n16670;
wire n16671;
wire n16672;
wire n16673;
wire n16674;
wire n16676;
wire n16677;
wire n16678;
wire n16679;
wire n16680;
wire n16681;
wire n16682;
wire n16683;
wire n16684;
wire n16685;
wire n16686;
wire n16687;
wire n16688;
wire n16689;
wire n16690;
wire n16691;
wire n16692;
wire n16694;
wire n16695;
wire n16697;
wire n16698;
wire n16700;
wire n16702;
wire n16703;
wire n16704;
wire n16705;
wire n16706;
wire n16707;
wire n16708;
wire n16709;
wire n16710;
wire n16712;
wire n16714;
wire n16715;
wire n16717;
wire n16719;
wire n16720;
wire n16721;
wire n16722;
wire n16723;
wire n16724;
wire n16725;
wire n16726;
wire n16728;
wire n16730;
wire n16731;
wire n16733;
wire n16735;
wire n16736;
wire n16737;
wire n16738;
wire n16739;
wire n16740;
wire n16741;
wire n16742;
wire n16744;
wire n16746;
wire n16747;
wire n16749;
wire n16751;
wire n16752;
wire n16753;
wire n16754;
wire n16755;
wire n16756;
wire n16757;
wire n16758;
wire n16760;
wire n16762;
wire n16763;
wire n16765;
wire n16767;
wire n16768;
wire n16769;
wire n16770;
wire n16771;
wire n16772;
wire n16773;
wire n16774;
wire n16776;
wire n16778;
wire n16780;
wire n16782;
wire n16783;
wire n16784;
wire n16786;
wire n16787;
wire n16789;
wire n16790;
wire n16791;
wire n16792;
wire n16793;
wire n16795;
wire n16796;
wire n16797;
wire n16798;
wire n16799;
wire n16801;
wire n16802;
wire n16803;
wire n16804;
wire n16805;
wire n16806;
wire n16807;
wire n16808;
wire n16809;
wire n16811;
wire n16812;
wire n16813;
wire n16814;
wire n16815;
wire n16816;
wire n16818;
wire n16819;
wire n16820;
wire n16821;
wire n16822;
wire n16823;
wire n16824;
wire n16825;
wire n16826;
wire n16827;
wire n16828;
wire n16829;
wire n16831;
wire n16832;
wire n16833;
wire n16834;
wire n16835;
wire n16836;
wire n16838;
wire n16840;
wire n16841;
wire n16842;
wire n16843;
wire n16844;
wire n16845;
wire n16847;
wire n16849;
wire n16851;
wire n16853;
wire n16854;
wire n16855;
wire n16857;
wire n16858;
wire n16859;
wire n16860;
wire n16861;
wire n16862;
wire n16864;
wire n16865;
wire n16866;
wire n16867;
wire n16868;
wire n16870;
wire n16871;
wire n16872;
wire n16873;
wire n16874;
wire n16875;
wire n16877;
wire n16879;
wire n16881;
wire n16883;
wire n16884;
wire n16885;
wire n16887;
wire n16888;
wire n16890;
wire n16891;
wire n16892;
wire n16893;
wire n16894;
wire n16896;
wire n16897;
wire n16898;
wire n16899;
wire n16900;
wire n16902;
wire n16903;
wire n16904;
wire n16905;
wire n16907;
wire n16909;
wire n16911;
wire n16912;
wire n16913;
wire n16914;
wire n16915;
wire n16917;
wire n16918;
wire n16920;
wire n16922;
wire n16924;
wire n16926;
wire n16928;
wire n16929;
wire n16930;
wire n16933;
wire n16934;
wire n16935;
wire n16936;
wire n16937;
wire n16938;
wire n16939;
wire n16940;
wire n16941;
wire n16943;
wire n16945;
wire n16946;
wire n16947;
wire n16948;
wire n16949;
wire n16950;
wire n16951;
wire n16952;
wire n16953;
wire n16954;
wire n16956;
wire n16957;
wire n16958;
wire n16959;
wire n16960;
wire n16961;
wire n16962;
wire n16963;
wire n16964;
wire n16965;
wire n16966;
wire n16967;
wire n16968;
wire n16969;
wire n16970;
wire n16971;
wire n16972;
wire n16973;
wire n16974;
wire n16976;
wire n16978;
wire n16980;
wire n16982;
wire n16983;
wire n16984;
wire n16986;
wire n16987;
wire n16989;
wire n16990;
wire n16991;
wire n16992;
wire n16993;
wire n16995;
wire n16996;
wire n16997;
wire n16998;
wire n16999;
wire n17001;
wire n17002;
wire n17003;
wire n17004;
wire n17005;
wire n17006;
wire n17007;
wire n17008;
wire n17009;
wire n17010;
wire n17012;
wire n17013;
wire n17014;
wire n17015;
wire n17016;
wire n17017;
wire n17018;
wire n17019;
wire n17020;
wire n17021;
wire n17022;
wire n17023;
wire n17024;
wire n17025;
wire n17026;
wire n17027;
wire n17028;
wire n17029;
wire n17030;
wire n17031;
wire n17032;
wire n17033;
wire n17034;
wire n17035;
wire n17036;
wire n17037;
wire n17038;
wire n17039;
wire n17040;
wire n17041;
wire n17042;
wire n17043;
wire n17044;
wire n17045;
wire n17046;
wire n17047;
wire n17048;
wire n17049;
wire n17050;
wire n17051;
wire n17052;
wire n17053;
wire n17054;
wire n17055;
wire n17056;
wire n17057;
wire n17058;
wire n17059;
wire n17060;
wire n17061;
wire n17062;
wire n17063;
wire n17064;
wire n17065;
wire n17066;
wire n17067;
wire n17068;
wire n17069;
wire n17070;
wire n17071;
wire n17072;
wire n17073;
wire n17074;
wire n17075;
wire n17076;
wire n17077;
wire n17078;
wire n17079;
wire n17080;
wire n17081;
wire n17082;
wire n17083;
wire n17084;
wire n17085;
wire n17086;
wire n17087;
wire n17088;
wire n17089;
wire n17090;
wire n17091;
wire n17092;
wire n17093;
wire n17094;
wire n17095;
wire n17096;
wire n17097;
wire n17098;
wire n17099;
wire n17100;
wire n17101;
wire n17102;
wire n17103;
wire n17104;
wire n17105;
wire n17106;
wire n17107;
wire n17108;
wire n17109;
wire n17110;
wire n17111;
wire n17112;
wire n17113;
wire n17114;
wire n17115;
wire n17116;
wire n17117;
wire n17118;
wire n17119;
wire n17120;
wire n17121;
wire n17122;
wire n17123;
wire n17124;
wire n17125;
wire n17126;
wire n17127;
wire n17128;
wire n17129;
wire n17130;
wire n17131;
wire n17132;
wire n17133;
wire n17134;
wire n17135;
wire n17136;
wire n17137;
wire n17138;
wire n17139;
wire n17140;
wire n17141;
wire n17142;
wire n17143;
wire n17144;
wire n17145;
wire n17146;
wire n17147;
wire n17148;
wire n17149;
wire n17150;
wire n17151;
wire n17152;
wire n17153;
wire n17154;
wire n17155;
wire n17156;
wire n17157;
wire n17158;
wire n17159;
wire n17160;
wire n17161;
wire n17162;
wire n17163;
wire n17164;
wire n17165;
wire n17166;
wire n17167;
wire n17168;
wire n17169;
wire n17170;
wire n17171;
wire n17172;
wire n17173;
wire n17174;
wire n17175;
wire n17176;
wire n17177;
wire n17178;
wire n17179;
wire n17180;
wire n17181;
wire n17182;
wire n17183;
wire n17184;
wire n17185;
wire n17186;
wire n17187;
wire n17188;
wire n17189;
wire n17190;
wire n17191;
wire n17192;
wire n17193;
wire n17194;
wire n17195;
wire n17196;
wire n17197;
wire n17198;
wire n17199;
wire n17200;
wire n17201;
wire n17202;
wire n17203;
wire n17204;
wire n17205;
wire n17206;
wire n17207;
wire n17208;
wire n17209;
wire n17210;
wire n17211;
wire n17212;
wire n17213;
wire n17214;
wire n17215;
wire n17216;
wire n17217;
wire n17218;
wire n17219;
wire n17220;
wire n17221;
wire n17222;
wire n17223;
wire n17224;
wire n17225;
wire n17226;
wire n17227;
wire n17228;
wire n17229;
wire n17230;
wire n17231;
wire n17232;
wire n17233;
wire n17234;
wire n17235;
wire n17236;
wire n17237;
wire n17238;
wire n17239;
wire n17240;
wire n17241;
wire n17242;
wire n17243;
wire n17244;
wire n17245;
wire n17246;
wire n17247;
wire n17248;
wire n17249;
wire n17250;
wire n17251;
wire n17252;
wire n17253;
wire n17254;
wire n17255;
wire n17256;
wire n17257;
wire n17258;
wire n17259;
wire n17260;
wire n17261;
wire n17262;
wire n17263;
wire n17264;
wire n17265;
wire n17266;
wire n17267;
wire n17268;
wire n17269;
wire n17270;
wire n17271;
wire n17272;
wire n17273;
wire n17274;
wire n17275;
wire n17276;
wire n17277;
wire n17278;
wire n17279;
wire n17280;
wire n17281;
wire n17282;
wire n17283;
wire n17284;
wire n17285;
wire n17286;
wire n17287;
wire n17288;
wire n17289;
wire n17290;
wire n17291;
wire n17292;
wire n17293;
wire n17294;
wire n17295;
wire n17296;
wire n17297;
wire n17298;
wire n17299;
wire n17300;
wire n17301;
wire n17302;
wire n17303;
wire n17304;
wire n17305;
wire n17306;
wire n17307;
wire n17308;
wire n17309;
wire n17310;
wire n17311;
wire n17312;
wire n17313;
wire n17314;
wire n17315;
wire n17316;
wire n17317;
wire n17318;
wire n17319;
wire n17320;
wire n17321;
wire n17322;
wire n17323;
wire n17324;
wire n17325;
wire n17326;
wire n17327;
wire n17328;
wire n17329;
wire n17330;
wire n17331;
wire n17332;
wire n17333;
wire n17334;
wire n17335;
wire n17336;
wire n17337;
wire n17338;
wire n17339;
wire n17340;
wire n17341;
wire n17342;
wire n17343;
wire n17344;
wire n17345;
wire n17346;
wire n17347;
wire n17348;
wire n17349;
wire n17350;
wire n17351;
wire n17352;
wire n17353;
wire n17354;
wire n17355;
wire n17356;
wire n17357;
wire n17358;
wire n17359;
wire n17360;
wire n17361;
wire n17362;
wire n17363;
wire n17364;
wire n17365;
wire n17366;
wire n17367;
wire n17368;
wire n17369;
wire n17370;
wire n17371;
wire n17372;
wire n17373;
wire n17374;
wire n17375;
wire n17376;
wire n17377;
wire n17378;
wire n17379;
wire n17380;
wire n17381;
wire n17382;
wire n17383;
wire n17384;
wire n17385;
wire n17386;
wire n17387;
wire n17388;
wire n17389;
wire n17390;
wire n17391;
wire n17392;
wire n17393;
wire n17394;
wire n17395;
wire n17396;
wire n17397;
wire n17398;
wire n17399;
wire n17401;
wire n17402;
wire n17403;
wire n17405;
wire n17406;
wire n17408;
wire n17410;
wire n17411;
wire n17412;
wire n17413;
wire n17414;
wire n17415;
wire n17418;
wire n17419;
wire n17420;
wire n17421;
wire n17422;
wire n17423;
wire n17424;
wire n17425;
wire n17426;
wire n17427;
wire n17428;
wire n17429;
wire n17430;
wire n17431;
wire n17432;
wire n17433;
wire n17434;
wire n17435;
wire n17436;
wire n17437;
wire n17438;
wire n17439;
wire n17440;
wire n17441;
wire n17442;
wire n17443;
wire n17444;
wire n17445;
wire n17446;
wire n17447;
wire n17448;
wire n17449;
wire n17450;
wire n17451;
wire n17452;
wire n17454;
wire n17455;
wire n17456;
wire n17458;
wire n17459;
wire n17461;
wire n17463;
wire n17464;
wire n17465;
wire n17466;
wire n17467;
wire n17468;
wire n17471;
wire n17472;
wire n17473;
wire n17474;
wire n17475;
wire n17476;
wire n17477;
wire n17478;
wire n17479;
wire n17480;
wire n17481;
wire n17482;
wire n17483;
wire n17484;
wire n17485;
wire n17486;
wire n17487;
wire n17488;
wire n17489;
wire n17490;
wire n17491;
wire n17492;
wire n17493;
wire n17494;
wire n17495;
wire n17496;
wire n17497;
wire n17498;
wire n17500;
wire n17501;
wire n17502;
wire n17504;
wire n17505;
wire n17507;
wire n17509;
wire n17510;
wire n17511;
wire n17512;
wire n17513;
wire n17514;
wire n17517;
wire n17518;
wire n17519;
wire n17520;
wire n17521;
wire n17522;
wire n17523;
wire n17524;
wire n17525;
wire n17526;
wire n17527;
wire n17528;
wire n17529;
wire n17530;
wire n17531;
wire n17532;
wire n17533;
wire n17534;
wire n17535;
wire n17536;
wire n17537;
wire n17538;
wire n17539;
wire n17540;
wire n17541;
wire n17542;
wire n17543;
wire n17544;
wire n17545;
wire n17547;
wire n17548;
wire n17549;
wire n17551;
wire n17552;
wire n17554;
wire n17556;
wire n17557;
wire n17558;
wire n17559;
wire n17560;
wire n17561;
wire n17564;
wire n17565;
wire n17566;
wire n17567;
wire n17568;
wire n17569;
wire n17570;
wire n17571;
wire n17572;
wire n17573;
wire n17574;
wire n17575;
wire n17576;
wire n17577;
wire n17578;
wire n17579;
wire n17580;
wire n17581;
wire n17582;
wire n17583;
wire n17584;
wire n17585;
wire n17586;
wire n17587;
wire n17588;
wire n17589;
wire n17590;
wire n17591;
wire n17593;
wire n17594;
wire n17595;
wire n17597;
wire n17598;
wire n17600;
wire n17602;
wire n17603;
wire n17604;
wire n17605;
wire n17606;
wire n17607;
wire n17608;
wire n17609;
wire n17610;
wire n17611;
wire n17612;
wire n17613;
wire n17614;
wire n17615;
wire n17616;
wire n17617;
wire n17618;
wire n17619;
wire n17620;
wire n17621;
wire n17622;
wire n17623;
wire n17624;
wire n17625;
wire n17626;
wire n17627;
wire n17628;
wire n17629;
wire n17630;
wire n17631;
wire n17632;
wire n17633;
wire n17635;
wire n17636;
wire n17637;
wire n17639;
wire n17640;
wire n17642;
wire n17644;
wire n17645;
wire n17646;
wire n17647;
wire n17648;
wire n17649;
wire n17650;
wire n17651;
wire n17652;
wire n17653;
wire n17654;
wire n17655;
wire n17656;
wire n17657;
wire n17658;
wire n17659;
wire n17660;
wire n17661;
wire n17662;
wire n17663;
wire n17664;
wire n17666;
wire n17667;
wire n17668;
wire n17670;
wire n17671;
wire n17673;
wire n17675;
wire n17676;
wire n17677;
wire n17678;
wire n17679;
wire n17680;
wire n17681;
wire n17682;
wire n17683;
wire n17684;
wire n17685;
wire n17686;
wire n17687;
wire n17688;
wire n17689;
wire n17690;
wire n17691;
wire n17692;
wire n17693;
wire n17694;
wire n17696;
wire n17697;
wire n17698;
wire n17700;
wire n17701;
wire n17703;
wire n17705;
wire n17706;
wire n17707;
wire n17708;
wire n17709;
wire n17710;
wire n17711;
wire n17712;
wire n17713;
wire n17714;
wire n17715;
wire n17716;
wire n17717;
wire n17718;
wire n17719;
wire n17720;
wire n17721;
wire n17722;
wire n17723;
wire n17724;
wire n17725;
wire n17726;
wire n17727;
wire n17728;
wire n17729;
wire n17730;
wire n17731;
wire n17732;
wire n17733;
wire n17734;
wire n17735;
wire n17736;
wire n17737;
wire n17738;
wire n17739;
wire n17740;
wire n17741;
wire n17742;
wire n17744;
wire n17745;
wire n17746;
wire n17747;
wire n17748;
wire n17749;
wire n17750;
wire n17751;
wire n17752;
wire n17753;
wire n17754;
wire n17755;
wire n17756;
wire n17757;
wire n17758;
wire n17759;
wire n17760;
wire n17762;
wire n17763;
wire n17764;
wire n17765;
wire n17766;
wire n17767;
wire n17768;
wire n17769;
wire n17770;
wire n17771;
wire n17772;
wire n17773;
wire n17774;
wire n17775;
wire n17776;
wire n17777;
wire n17778;
wire n17779;
wire n17780;
wire n17781;
wire n17782;
wire n17783;
wire n17784;
wire n17785;
wire n17786;
wire n17787;
wire n17788;
wire n17790;
wire n17792;
wire n17793;
wire n17794;
wire n17795;
wire n17796;
wire n17797;
wire n17798;
wire n17799;
wire n17800;
wire n17801;
wire n17802;
wire n17803;
wire n17804;
wire n17805;
wire n17806;
wire n17807;
wire n17808;
wire n17809;
wire n17810;
wire n17811;
wire n17812;
wire n17813;
wire n17814;
wire n17815;
wire n17816;
wire n17817;
wire n17818;
wire n17819;
wire n17820;
wire n17821;
wire n17822;
wire n17823;
wire n17824;
wire n17825;
wire n17826;
wire n17827;
wire n17828;
wire n17829;
wire n17830;
wire n17831;
wire n17832;
wire n17833;
wire n17834;
wire n17835;
wire n17836;
wire n17837;
wire n17838;
wire n17839;
wire n17840;
wire n17841;
wire n17842;
wire n17843;
wire n17844;
wire n17845;
wire n17846;
wire n17847;
wire n17848;
wire n17849;
wire n17850;
wire n17851;
wire n17852;
wire n17853;
wire n17854;
wire n17855;
wire n17856;
wire n17857;
wire n17858;
wire n17859;
wire n17860;
wire n17861;
wire n17862;
wire n17863;
wire n17864;
wire n17865;
wire n17866;
wire n17867;
wire n17868;
wire n17869;
wire n17870;
wire n17871;
wire n17872;
wire n17873;
wire n17874;
wire n17875;
wire n17876;
wire n17877;
wire n17878;
wire n17879;
wire n17880;
wire n17881;
wire n17882;
wire n17883;
wire n17884;
wire n17885;
wire n17886;
wire n17887;
wire n17889;
wire n17890;
wire n17891;
wire n17892;
wire n17893;
wire n17894;
wire n17895;
wire n17896;
wire n17897;
wire n17899;
wire n17900;
wire n17901;
wire n17902;
wire n17903;
wire n17904;
wire n17905;
wire n17906;
wire n17907;
wire n17908;
wire n17909;
wire n17910;
wire n17911;
wire n17912;
wire n17913;
wire n17914;
wire n17915;
wire n17916;
wire n17917;
wire n17918;
wire n17920;
wire n17922;
wire n17924;
wire n17925;
wire n17926;
wire n17927;
wire n17928;
wire n17929;
wire n17930;
wire n17931;
wire n17932;
wire n17933;
wire n17934;
wire n17935;
wire n17936;
wire n17937;
wire n17938;
wire n17939;
wire n17940;
wire n17941;
wire n17942;
wire n17943;
wire n17944;
wire n17945;
wire n17946;
wire n17947;
wire n17948;
wire n17949;
wire n17950;
wire n17951;
wire n17952;
wire n17953;
wire n17954;
wire n17955;
wire n17956;
wire n17957;
wire n17958;
wire n17959;
wire n17960;
wire n17961;
wire n17962;
wire n17963;
wire n17964;
wire n17965;
wire n17966;
wire n17967;
wire n17968;
wire n17969;
wire n17970;
wire n17971;
wire n17972;
wire n17973;
wire n17974;
wire n17975;
wire n17976;
wire n17977;
wire n17978;
wire n17979;
wire n17980;
wire n17981;
wire n17982;
wire n17983;
wire n17984;
wire n17985;
wire n17986;
wire n17987;
wire n17988;
wire n17989;
wire n17990;
wire n17991;
wire n17992;
wire n17993;
wire n17994;
wire n17995;
wire n17996;
wire n17997;
wire n17998;
wire n17999;
wire n18000;
wire n18001;
wire n18003;
wire n18004;
wire n18005;
wire n18006;
wire n18007;
wire n18008;
wire n18009;
wire n18010;
wire n18011;
wire n18012;
wire n18013;
wire n18014;
wire n18015;
wire n18016;
wire n18017;
wire n18019;
wire n18020;
wire n18021;
wire n18022;
wire n18023;
wire n18024;
wire n18025;
wire n18026;
wire n18027;
wire n18028;
wire n18029;
wire n18030;
wire n18031;
wire n18032;
wire n18033;
wire n18034;
wire n18035;
wire n18036;
wire n18037;
wire n18038;
wire n18039;
wire n18040;
wire n18041;
wire n18043;
wire n18045;
wire n18047;
wire n18048;
wire n18049;
wire n18050;
wire n18051;
wire n18052;
wire n18053;
wire n18054;
wire n18055;
wire n18056;
wire n18057;
wire n18058;
wire n18059;
wire n18060;
wire n18061;
wire n18062;
wire n18063;
wire n18064;
wire n18065;
wire n18066;
wire n18067;
wire n18068;
wire n18069;
wire n18070;
wire n18071;
wire n18072;
wire n18073;
wire n18074;
wire n18075;
wire n18076;
wire n18077;
wire n18078;
wire n18079;
wire n18080;
wire n18081;
wire n18082;
wire n18083;
wire n18084;
wire n18085;
wire n18086;
wire n18087;
wire n18088;
wire n18089;
wire n18090;
wire n18091;
wire n18092;
wire n18093;
wire n18094;
wire n18095;
wire n18096;
wire n18097;
wire n18098;
wire n18099;
wire n18100;
wire n18101;
wire n18102;
wire n18103;
wire n18104;
wire n18105;
wire n18106;
wire n18107;
wire n18108;
wire n18109;
wire n18110;
wire n18111;
wire n18112;
wire n18113;
wire n18114;
wire n18115;
wire n18116;
wire n18117;
wire n18118;
wire n18119;
wire n18120;
wire n18121;
wire n18122;
wire n18123;
wire n18124;
wire n18126;
wire n18127;
wire n18128;
wire n18129;
wire n18130;
wire n18131;
wire n18132;
wire n18133;
wire n18134;
wire n18136;
wire n18137;
wire n18138;
wire n18139;
wire n18140;
wire n18141;
wire n18142;
wire n18143;
wire n18144;
wire n18145;
wire n18146;
wire n18147;
wire n18148;
wire n18149;
wire n18150;
wire n18151;
wire n18152;
wire n18153;
wire n18154;
wire n18155;
wire n18157;
wire n18159;
wire n18161;
wire n18162;
wire n18163;
wire n18164;
wire n18165;
wire n18166;
wire n18167;
wire n18168;
wire n18169;
wire n18170;
wire n18171;
wire n18172;
wire n18173;
wire n18174;
wire n18175;
wire n18176;
wire n18177;
wire n18178;
wire n18179;
wire n18180;
wire n18181;
wire n18182;
wire n18183;
wire n18184;
wire n18185;
wire n18186;
wire n18187;
wire n18188;
wire n18189;
wire n18190;
wire n18191;
wire n18192;
wire n18193;
wire n18194;
wire n18195;
wire n18196;
wire n18197;
wire n18198;
wire n18199;
wire n18200;
wire n18201;
wire n18202;
wire n18203;
wire n18204;
wire n18205;
wire n18206;
wire n18207;
wire n18208;
wire n18209;
wire n18210;
wire n18211;
wire n18212;
wire n18213;
wire n18214;
wire n18215;
wire n18216;
wire n18217;
wire n18218;
wire n18219;
wire n18220;
wire n18221;
wire n18222;
wire n18223;
wire n18224;
wire n18225;
wire n18226;
wire n18227;
wire n18228;
wire n18229;
wire n18230;
wire n18231;
wire n18232;
wire n18233;
wire n18234;
wire n18235;
wire n18236;
wire n18237;
wire n18238;
wire n18240;
wire n18241;
wire n18242;
wire n18243;
wire n18244;
wire n18245;
wire n18246;
wire n18247;
wire n18248;
wire n18250;
wire n18251;
wire n18252;
wire n18253;
wire n18254;
wire n18255;
wire n18256;
wire n18257;
wire n18258;
wire n18259;
wire n18260;
wire n18261;
wire n18262;
wire n18263;
wire n18264;
wire n18265;
wire n18266;
wire n18267;
wire n18268;
wire n18269;
wire n18271;
wire n18273;
wire n18275;
wire n18276;
wire n18277;
wire n18278;
wire n18279;
wire n18280;
wire n18281;
wire n18282;
wire n18283;
wire n18284;
wire n18285;
wire n18286;
wire n18287;
wire n18288;
wire n18289;
wire n18290;
wire n18291;
wire n18292;
wire n18293;
wire n18294;
wire n18295;
wire n18296;
wire n18297;
wire n18298;
wire n18299;
wire n18300;
wire n18301;
wire n18302;
wire n18303;
wire n18304;
wire n18305;
wire n18306;
wire n18307;
wire n18308;
wire n18309;
wire n18310;
wire n18311;
wire n18312;
wire n18313;
wire n18314;
wire n18315;
wire n18316;
wire n18317;
wire n18318;
wire n18319;
wire n18320;
wire n18321;
wire n18322;
wire n18323;
wire n18324;
wire n18325;
wire n18326;
wire n18327;
wire n18328;
wire n18329;
wire n18330;
wire n18331;
wire n18332;
wire n18333;
wire n18334;
wire n18335;
wire n18336;
wire n18337;
wire n18338;
wire n18339;
wire n18340;
wire n18341;
wire n18342;
wire n18343;
wire n18344;
wire n18345;
wire n18346;
wire n18347;
wire n18348;
wire n18349;
wire n18350;
wire n18351;
wire n18352;
wire n18354;
wire n18355;
wire n18356;
wire n18357;
wire n18358;
wire n18359;
wire n18360;
wire n18361;
wire n18362;
wire n18364;
wire n18365;
wire n18366;
wire n18367;
wire n18368;
wire n18369;
wire n18370;
wire n18371;
wire n18372;
wire n18373;
wire n18374;
wire n18375;
wire n18376;
wire n18377;
wire n18378;
wire n18379;
wire n18380;
wire n18381;
wire n18382;
wire n18383;
wire n18385;
wire n18387;
wire n18389;
wire n18390;
wire n18391;
wire n18392;
wire n18393;
wire n18394;
wire n18395;
wire n18396;
wire n18397;
wire n18398;
wire n18399;
wire n18400;
wire n18401;
wire n18402;
wire n18403;
wire n18404;
wire n18405;
wire n18406;
wire n18407;
wire n18408;
wire n18409;
wire n18410;
wire n18411;
wire n18412;
wire n18413;
wire n18414;
wire n18415;
wire n18416;
wire n18417;
wire n18418;
wire n18419;
wire n18420;
wire n18421;
wire n18422;
wire n18423;
wire n18424;
wire n18425;
wire n18426;
wire n18427;
wire n18428;
wire n18429;
wire n18430;
wire n18431;
wire n18432;
wire n18433;
wire n18434;
wire n18435;
wire n18436;
wire n18437;
wire n18438;
wire n18439;
wire n18440;
wire n18441;
wire n18442;
wire n18443;
wire n18444;
wire n18445;
wire n18446;
wire n18447;
wire n18448;
wire n18449;
wire n18450;
wire n18451;
wire n18452;
wire n18453;
wire n18454;
wire n18455;
wire n18456;
wire n18457;
wire n18458;
wire n18459;
wire n18460;
wire n18461;
wire n18462;
wire n18463;
wire n18464;
wire n18465;
wire n18466;
wire n18468;
wire n18469;
wire n18470;
wire n18471;
wire n18472;
wire n18473;
wire n18474;
wire n18475;
wire n18476;
wire n18478;
wire n18479;
wire n18480;
wire n18481;
wire n18482;
wire n18483;
wire n18484;
wire n18485;
wire n18486;
wire n18487;
wire n18488;
wire n18489;
wire n18490;
wire n18491;
wire n18492;
wire n18493;
wire n18494;
wire n18495;
wire n18496;
wire n18497;
wire n18499;
wire n18501;
wire n18503;
wire n18504;
wire n18505;
wire n18506;
wire n18507;
wire n18508;
wire n18509;
wire n18510;
wire n18511;
wire n18512;
wire n18513;
wire n18514;
wire n18515;
wire n18516;
wire n18517;
wire n18518;
wire n18519;
wire n18520;
wire n18521;
wire n18522;
wire n18523;
wire n18524;
wire n18525;
wire n18526;
wire n18527;
wire n18528;
wire n18529;
wire n18530;
wire n18531;
wire n18532;
wire n18533;
wire n18534;
wire n18535;
wire n18536;
wire n18537;
wire n18538;
wire n18539;
wire n18540;
wire n18541;
wire n18542;
wire n18543;
wire n18544;
wire n18545;
wire n18546;
wire n18547;
wire n18548;
wire n18549;
wire n18550;
wire n18551;
wire n18552;
wire n18553;
wire n18554;
wire n18555;
wire n18556;
wire n18557;
wire n18558;
wire n18559;
wire n18560;
wire n18561;
wire n18562;
wire n18563;
wire n18564;
wire n18565;
wire n18566;
wire n18567;
wire n18568;
wire n18569;
wire n18570;
wire n18571;
wire n18572;
wire n18573;
wire n18574;
wire n18575;
wire n18576;
wire n18577;
wire n18578;
wire n18579;
wire n18581;
wire n18582;
wire n18583;
wire n18584;
wire n18585;
wire n18586;
wire n18587;
wire n18588;
wire n18589;
wire n18591;
wire n18592;
wire n18593;
wire n18594;
wire n18595;
wire n18596;
wire n18597;
wire n18598;
wire n18599;
wire n18600;
wire n18601;
wire n18602;
wire n18603;
wire n18604;
wire n18605;
wire n18606;
wire n18607;
wire n18608;
wire n18609;
wire n18610;
wire n18612;
wire n18614;
wire n18616;
wire n18617;
wire n18618;
wire n18619;
wire n18620;
wire n18621;
wire n18622;
wire n18623;
wire n18624;
wire n18625;
wire n18626;
wire n18627;
wire n18628;
wire n18629;
wire n18630;
wire n18631;
wire n18632;
wire n18633;
wire n18634;
wire n18635;
wire n18636;
wire n18637;
wire n18638;
wire n18639;
wire n18640;
wire n18641;
wire n18642;
wire n18643;
wire n18644;
wire n18645;
wire n18646;
wire n18647;
wire n18648;
wire n18649;
wire n18650;
wire n18651;
wire n18652;
wire n18653;
wire n18654;
wire n18655;
wire n18656;
wire n18657;
wire n18658;
wire n18659;
wire n18660;
wire n18661;
wire n18662;
wire n18663;
wire n18664;
wire n18665;
wire n18666;
wire n18667;
wire n18668;
wire n18669;
wire n18670;
wire n18671;
wire n18672;
wire n18673;
wire n18674;
wire n18675;
wire n18676;
wire n18677;
wire n18678;
wire n18679;
wire n18680;
wire n18681;
wire n18682;
wire n18683;
wire n18684;
wire n18685;
wire n18686;
wire n18687;
wire n18688;
wire n18689;
wire n18690;
wire n18691;
wire n18692;
wire n18693;
wire n18694;
wire n18695;
wire n18696;
wire n18697;
wire n18698;
wire n18699;
wire n18700;
wire n18701;
wire n18702;
wire n18703;
wire n18704;
wire n18705;
wire n18706;
wire n18707;
wire n18708;
wire n18709;
wire n18710;
wire n18711;
wire n18712;
wire n18713;
wire n18714;
wire n18715;
wire n18716;
wire n18717;
wire n18718;
wire n18719;
wire n18720;
wire n18721;
wire n18722;
wire n18723;
wire n18724;
wire n18725;
wire n18726;
wire n18727;
wire n18728;
wire n18729;
wire n18730;
wire n18731;
wire n18732;
wire n18733;
wire n18734;
wire n18735;
wire n18736;
wire n18737;
wire n18738;
wire n18739;
wire n18740;
wire n18741;
wire n18742;
wire n18743;
wire n18744;
wire n18745;
wire n18747;
wire n18748;
wire n18749;
wire n18750;
wire n18751;
wire n18752;
wire n18753;
wire n18754;
wire n18755;
wire n18756;
wire n18757;
wire n18758;
wire n18759;
wire n18760;
wire n18761;
wire n18762;
wire n18763;
wire n18764;
wire n18765;
wire n18766;
wire n18767;
wire n18768;
wire n18769;
wire n18770;
wire n18771;
wire n18772;
wire n18773;
wire n18774;
wire n18775;
wire n18776;
wire n18777;
wire n18778;
wire n18779;
wire n18780;
wire n18781;
wire n18782;
wire n18783;
wire n18784;
wire n18785;
wire n18786;
wire n18787;
wire n18789;
wire n18790;
wire n18791;
wire n18792;
wire n18793;
wire n18794;
wire n18795;
wire n18796;
wire n18797;
wire n18798;
wire n18799;
wire n18800;
wire n18801;
wire n18802;
wire n18803;
wire n18804;
wire n18805;
wire n18806;
wire n18807;
wire n18808;
wire n18809;
wire n18810;
wire n18811;
wire n18812;
wire n18813;
wire n18814;
wire n18815;
wire n18816;
wire n18817;
wire n18818;
wire n18819;
wire n18820;
wire n18821;
wire n18822;
wire n18823;
wire n18824;
wire n18825;
wire n18826;
wire n18827;
wire n18828;
wire n18829;
wire n18830;
wire n18832;
wire n18833;
wire n18834;
wire n18835;
wire n18836;
wire n18837;
wire n18838;
wire n18839;
wire n18840;
wire n18841;
wire n18842;
wire n18843;
wire n18844;
wire n18845;
wire n18846;
wire n18847;
wire n18848;
wire n18849;
wire n18850;
wire n18851;
wire n18852;
wire n18853;
wire n18854;
wire n18855;
wire n18856;
wire n18857;
wire n18858;
wire n18859;
wire n18860;
wire n18861;
wire n18862;
wire n18863;
wire n18864;
wire n18865;
wire n18866;
wire n18867;
wire n18868;
wire n18869;
wire n18870;
wire n18871;
wire n18872;
wire n18873;
wire n18875;
wire n18876;
wire n18877;
wire n18878;
wire n18879;
wire n18880;
wire n18881;
wire n18882;
wire n18883;
wire n18884;
wire n18885;
wire n18886;
wire n18887;
wire n18888;
wire n18889;
wire n18890;
wire n18891;
wire n18892;
wire n18893;
wire n18894;
wire n18895;
wire n18896;
wire n18897;
wire n18898;
wire n18899;
wire n18900;
wire n18901;
wire n18902;
wire n18903;
wire n18904;
wire n18905;
wire n18906;
wire n18907;
wire n18908;
wire n18909;
wire n18910;
wire n18911;
wire n18912;
wire n18913;
wire n18914;
wire n18915;
wire n18916;
wire n18918;
wire n18919;
wire n18920;
wire n18921;
wire n18922;
wire n18923;
wire n18924;
wire n18925;
wire n18926;
wire n18927;
wire n18928;
wire n18929;
wire n18930;
wire n18931;
wire n18932;
wire n18933;
wire n18934;
wire n18935;
wire n18936;
wire n18937;
wire n18938;
wire n18939;
wire n18940;
wire n18941;
wire n18942;
wire n18943;
wire n18944;
wire n18945;
wire n18946;
wire n18947;
wire n18948;
wire n18949;
wire n18950;
wire n18951;
wire n18952;
wire n18953;
wire n18954;
wire n18955;
wire n18956;
wire n18957;
wire n18958;
wire n18959;
wire n18961;
wire n18962;
wire n18963;
wire n18964;
wire n18965;
wire n18966;
wire n18967;
wire n18968;
wire n18969;
wire n18970;
wire n18971;
wire n18972;
wire n18973;
wire n18974;
wire n18975;
wire n18976;
wire n18977;
wire n18978;
wire n18979;
wire n18980;
wire n18981;
wire n18982;
wire n18983;
wire n18984;
wire n18985;
wire n18986;
wire n18987;
wire n18988;
wire n18989;
wire n18990;
wire n18991;
wire n18992;
wire n18993;
wire n18994;
wire n18995;
wire n18996;
wire n18997;
wire n18998;
wire n18999;
wire n19000;
wire n19001;
wire n19002;
wire n19004;
wire n19005;
wire n19006;
wire n19007;
wire n19008;
wire n19009;
wire n19010;
wire n19011;
wire n19012;
wire n19013;
wire n19014;
wire n19015;
wire n19016;
wire n19017;
wire n19018;
wire n19019;
wire n19020;
wire n19021;
wire n19022;
wire n19023;
wire n19024;
wire n19025;
wire n19026;
wire n19027;
wire n19028;
wire n19029;
wire n19030;
wire n19031;
wire n19032;
wire n19033;
wire n19034;
wire n19035;
wire n19036;
wire n19037;
wire n19038;
wire n19039;
wire n19040;
wire n19041;
wire n19042;
wire n19043;
wire n19044;
wire n19046;
wire n19047;
wire n19048;
wire n19049;
wire n19050;
wire n19051;
wire n19052;
wire n19053;
wire n19054;
wire n19055;
wire n19056;
wire n19057;
wire n19058;
wire n19059;
wire n19060;
wire n19061;
wire n19062;
wire n19063;
wire n19064;
wire n19065;
wire n19066;
wire n19067;
wire n19068;
wire n19069;
wire n19070;
wire n19071;
wire n19072;
wire n19073;
wire n19074;
wire n19075;
wire n19076;
wire n19077;
wire n19078;
wire n19079;
wire n19080;
wire n19081;
wire n19082;
wire n19083;
wire n19084;
wire n19085;
wire n19086;
wire n19087;
wire n19088;
wire n19089;
wire n19090;
wire n19091;
wire n19092;
wire n19093;
wire n19094;
wire n19095;
wire n19096;
wire n19097;
wire n19098;
wire n19099;
wire n19100;
wire n19101;
wire n19102;
wire n19103;
wire n19104;
wire n19105;
wire n19106;
wire n19107;
wire n19108;
wire n19109;
wire n19110;
wire n19111;
wire n19112;
wire n19113;
wire n19114;
wire n19115;
wire n19116;
wire n19117;
wire n19118;
wire n19119;
wire n19120;
wire n19121;
wire n19122;
wire n19123;
wire n19124;
wire n19125;
wire n19126;
wire n19127;
wire n19128;
wire n19129;
wire n19130;
wire n19131;
wire n19132;
wire n19133;
wire n19134;
wire n19135;
wire n19136;
wire n19137;
wire n19138;
wire n19139;
wire n19140;
wire n19141;
wire n19142;
wire n19143;
wire n19144;
wire n19145;
wire n19146;
wire n19147;
wire n19148;
wire n19149;
wire n19150;
wire n19151;
wire n19152;
wire n19153;
wire n19154;
wire n19155;
wire n19156;
wire n19157;
wire n19158;
wire n19159;
wire n19160;
wire n19161;
wire n19162;
wire n19163;
wire n19164;
wire n19165;
wire n19166;
wire n19167;
wire n19168;
wire n19169;
wire n19170;
wire n19171;
wire n19172;
wire n19173;
wire n19174;
wire n19175;
wire n19176;
wire n19177;
wire n19178;
wire n19179;
wire n19180;
wire n19181;
wire n19182;
wire n19183;
wire n19184;
wire n19185;
wire n19186;
wire n19187;
wire n19188;
wire n19189;
wire n19190;
wire n19191;
wire n19192;
wire n19193;
wire n19194;
wire n19195;
wire n19196;
wire n19197;
wire n19198;
wire n19199;
wire n19200;
wire n19201;
wire n19202;
wire n19203;
wire n19204;
wire n19205;
wire n19206;
wire n19207;
wire n19209;
wire n19210;
wire n19211;
wire n19212;
wire n19213;
wire n19214;
wire n19216;
wire n19217;
wire n19218;
wire n19219;
wire n19220;
wire n19221;
wire n19222;
wire n19223;
wire n19224;
wire n19225;
wire n19226;
wire n19227;
wire n19228;
wire n19229;
wire n19230;
wire n19231;
wire n19232;
wire n19233;
wire n19234;
wire n19235;
wire n19236;
wire n19237;
wire n19238;
wire n19239;
wire n19240;
wire n19241;
wire n19242;
wire n19243;
wire n19244;
wire n19245;
wire n19246;
wire n19247;
wire n19248;
wire n19249;
wire n19250;
wire n19251;
wire n19252;
wire n19253;
wire n19254;
wire n19255;
wire n19256;
wire n19257;
wire n19258;
wire n19260;
wire n19261;
wire n19262;
wire n19263;
wire n19264;
wire n19265;
wire n19266;
wire n19267;
wire n19268;
wire n19269;
wire n19270;
wire n19271;
wire n19272;
wire n19273;
wire n19274;
wire n19275;
wire n19276;
wire n19277;
wire n19278;
wire n19279;
wire n19280;
wire n19281;
wire n19282;
wire n19283;
wire n19284;
wire n19285;
wire n19286;
wire n19287;
wire n19289;
wire n19290;
wire n19291;
wire n19292;
wire n19293;
wire n19294;
wire n19296;
wire n19297;
wire n19298;
wire n19299;
wire n19300;
wire n19301;
wire n19302;
wire n19303;
wire n19304;
wire n19305;
wire n19306;
wire n19307;
wire n19308;
wire n19309;
wire n19310;
wire n19311;
wire n19312;
wire n19313;
wire n19314;
wire n19315;
wire n19316;
wire n19317;
wire n19318;
wire n19319;
wire n19320;
wire n19321;
wire n19322;
wire n19323;
wire n19324;
wire n19325;
wire n19326;
wire n19327;
wire n19328;
wire n19329;
wire n19330;
wire n19331;
wire n19332;
wire n19333;
wire n19334;
wire n19335;
wire n19336;
wire n19337;
wire n19339;
wire n19340;
wire n19341;
wire n19342;
wire n19343;
wire n19344;
wire n19345;
wire n19346;
wire n19347;
wire n19348;
wire n19349;
wire n19350;
wire n19351;
wire n19352;
wire n19353;
wire n19354;
wire n19355;
wire n19356;
wire n19357;
wire n19358;
wire n19359;
wire n19360;
wire n19362;
wire n19363;
wire n19364;
wire n19365;
wire n19366;
wire n19367;
wire n19369;
wire n19370;
wire n19371;
wire n19372;
wire n19373;
wire n19374;
wire n19375;
wire n19376;
wire n19377;
wire n19378;
wire n19379;
wire n19380;
wire n19381;
wire n19382;
wire n19383;
wire n19384;
wire n19385;
wire n19386;
wire n19387;
wire n19388;
wire n19389;
wire n19390;
wire n19391;
wire n19392;
wire n19393;
wire n19394;
wire n19395;
wire n19396;
wire n19397;
wire n19398;
wire n19399;
wire n19400;
wire n19401;
wire n19402;
wire n19403;
wire n19404;
wire n19405;
wire n19406;
wire n19407;
wire n19408;
wire n19409;
wire n19410;
wire n19412;
wire n19413;
wire n19414;
wire n19415;
wire n19416;
wire n19417;
wire n19418;
wire n19419;
wire n19420;
wire n19421;
wire n19422;
wire n19423;
wire n19424;
wire n19425;
wire n19426;
wire n19427;
wire n19428;
wire n19429;
wire n19430;
wire n19431;
wire n19432;
wire n19433;
wire n19434;
wire n19435;
wire n19436;
wire n19437;
wire n19438;
wire n19439;
wire n19440;
wire n19441;
wire n19442;
wire n19443;
wire n19444;
wire n19446;
wire n19447;
wire n19448;
wire n19449;
wire n19450;
wire n19451;
wire n19453;
wire n19454;
wire n19455;
wire n19456;
wire n19457;
wire n19458;
wire n19459;
wire n19460;
wire n19461;
wire n19462;
wire n19463;
wire n19464;
wire n19465;
wire n19466;
wire n19467;
wire n19468;
wire n19469;
wire n19470;
wire n19471;
wire n19472;
wire n19473;
wire n19474;
wire n19475;
wire n19476;
wire n19477;
wire n19478;
wire n19479;
wire n19480;
wire n19481;
wire n19482;
wire n19483;
wire n19484;
wire n19485;
wire n19486;
wire n19487;
wire n19488;
wire n19489;
wire n19490;
wire n19491;
wire n19493;
wire n19494;
wire n19495;
wire n19496;
wire n19497;
wire n19498;
wire n19499;
wire n19500;
wire n19501;
wire n19502;
wire n19503;
wire n19504;
wire n19505;
wire n19506;
wire n19507;
wire n19508;
wire n19509;
wire n19510;
wire n19511;
wire n19512;
wire n19513;
wire n19514;
wire n19516;
wire n19517;
wire n19518;
wire n19519;
wire n19520;
wire n19521;
wire n19523;
wire n19524;
wire n19525;
wire n19526;
wire n19527;
wire n19528;
wire n19529;
wire n19530;
wire n19531;
wire n19532;
wire n19533;
wire n19534;
wire n19535;
wire n19536;
wire n19537;
wire n19538;
wire n19539;
wire n19540;
wire n19541;
wire n19542;
wire n19543;
wire n19544;
wire n19545;
wire n19546;
wire n19547;
wire n19548;
wire n19549;
wire n19550;
wire n19551;
wire n19552;
wire n19553;
wire n19554;
wire n19555;
wire n19556;
wire n19557;
wire n19558;
wire n19559;
wire n19560;
wire n19561;
wire n19563;
wire n19564;
wire n19565;
wire n19566;
wire n19567;
wire n19568;
wire n19569;
wire n19570;
wire n19571;
wire n19572;
wire n19573;
wire n19574;
wire n19575;
wire n19576;
wire n19577;
wire n19578;
wire n19579;
wire n19580;
wire n19581;
wire n19582;
wire n19583;
wire n19584;
wire n19585;
wire n19587;
wire n19588;
wire n19589;
wire n19590;
wire n19591;
wire n19592;
wire n19594;
wire n19595;
wire n19596;
wire n19597;
wire n19598;
wire n19599;
wire n19600;
wire n19601;
wire n19602;
wire n19603;
wire n19604;
wire n19605;
wire n19606;
wire n19607;
wire n19608;
wire n19609;
wire n19610;
wire n19611;
wire n19612;
wire n19613;
wire n19614;
wire n19615;
wire n19616;
wire n19617;
wire n19618;
wire n19619;
wire n19620;
wire n19621;
wire n19622;
wire n19623;
wire n19624;
wire n19625;
wire n19626;
wire n19627;
wire n19628;
wire n19629;
wire n19630;
wire n19631;
wire n19632;
wire n19634;
wire n19635;
wire n19636;
wire n19637;
wire n19638;
wire n19639;
wire n19640;
wire n19641;
wire n19642;
wire n19643;
wire n19644;
wire n19645;
wire n19646;
wire n19647;
wire n19648;
wire n19649;
wire n19650;
wire n19651;
wire n19652;
wire n19653;
wire n19654;
wire n19655;
wire n19657;
wire n19658;
wire n19659;
wire n19660;
wire n19661;
wire n19662;
wire n19664;
wire n19665;
wire n19666;
wire n19667;
wire n19668;
wire n19669;
wire n19670;
wire n19671;
wire n19672;
wire n19673;
wire n19674;
wire n19675;
wire n19676;
wire n19677;
wire n19678;
wire n19679;
wire n19680;
wire n19681;
wire n19682;
wire n19683;
wire n19684;
wire n19685;
wire n19686;
wire n19687;
wire n19688;
wire n19689;
wire n19690;
wire n19691;
wire n19692;
wire n19693;
wire n19694;
wire n19695;
wire n19696;
wire n19697;
wire n19698;
wire n19699;
wire n19700;
wire n19701;
wire n19702;
wire n19704;
wire n19705;
wire n19706;
wire n19707;
wire n19708;
wire n19709;
wire n19710;
wire n19711;
wire n19712;
wire n19713;
wire n19714;
wire n19715;
wire n19716;
wire n19717;
wire n19718;
wire n19719;
wire n19720;
wire n19721;
wire n19722;
wire n19723;
wire n19724;
wire n19725;
wire n19726;
wire n19727;
wire n19728;
wire n19729;
wire n19730;
wire n19731;
wire n19732;
wire n19733;
wire n19734;
wire n19735;
wire n19736;
wire n19737;
wire n19738;
wire n19739;
wire n19741;
wire n19742;
wire n19743;
wire n19744;
wire n19745;
wire n19746;
wire n19748;
wire n19749;
wire n19750;
wire n19751;
wire n19752;
wire n19753;
wire n19754;
wire n19755;
wire n19756;
wire n19757;
wire n19758;
wire n19759;
wire n19760;
wire n19761;
wire n19762;
wire n19763;
wire n19764;
wire n19765;
wire n19766;
wire n19767;
wire n19768;
wire n19769;
wire n19770;
wire n19771;
wire n19772;
wire n19773;
wire n19774;
wire n19775;
wire n19776;
wire n19777;
wire n19778;
wire n19779;
wire n19780;
wire n19781;
wire n19782;
wire n19783;
wire n19784;
wire n19785;
wire n19786;
wire n19788;
wire n19789;
wire n19790;
wire n19791;
wire n19792;
wire n19793;
wire n19794;
wire n19795;
wire n19796;
wire n19797;
wire n19798;
wire n19799;
wire n19800;
wire n19801;
wire n19802;
wire n19803;
wire n19804;
wire n19805;
wire n19806;
wire n19807;
wire n19808;
wire n19809;
wire n19810;
wire n19811;
wire n19812;
wire n19813;
wire n19814;
wire n19815;
wire n19816;
wire n19817;
wire n19818;
wire n19819;
wire n19820;
wire n19821;
wire n19822;
wire n19823;
wire n19824;
wire n19825;
wire n19826;
wire n19827;
wire n19828;
wire n19829;
wire n19830;
wire n19831;
wire n19832;
wire n19833;
wire n19834;
wire n19835;
wire n19836;
wire n19837;
wire n19838;
wire n19839;
wire n19840;
wire n19841;
wire n19842;
wire n19843;
wire n19844;
wire n19845;
wire n19846;
wire n19847;
wire n19848;
wire n19849;
wire n19850;
wire n19851;
wire n19852;
wire n19853;
wire n19854;
wire n19855;
wire n19856;
wire n19857;
wire n19858;
wire n19859;
wire n19860;
wire n19861;
wire n19862;
wire n19863;
wire n19864;
wire n19865;
wire n19866;
wire n19867;
wire n19868;
wire n19869;
wire n19870;
wire n19871;
wire n19872;
wire n19873;
wire n19874;
wire n19875;
wire n19876;
wire n19877;
wire n19878;
wire n19879;
wire n19880;
wire n19881;
wire n19882;
wire n19883;
wire n19884;
wire n19885;
wire n19886;
wire n19887;
wire n19888;
wire n19889;
wire n19890;
wire n19891;
wire n19892;
wire n19893;
wire n19894;
wire n19895;
wire n19896;
wire n19897;
wire n19898;
wire n19899;
wire n19900;
wire n19901;
wire n19902;
wire n19903;
wire n19904;
wire n19905;
wire n19906;
wire n19907;
wire n19908;
wire n19909;
wire n19910;
wire n19911;
wire n19912;
wire n19913;
wire n19914;
wire n19915;
wire n19916;
wire n19917;
wire n19918;
wire n19919;
wire n19920;
wire n19921;
wire n19922;
wire n19923;
wire n19924;
wire n19925;
wire n19926;
wire n19927;
wire n19928;
wire n19929;
wire n19930;
wire n19931;
wire n19932;
wire n19933;
wire n19934;
wire n19935;
wire n19936;
wire n19937;
wire n19938;
wire n19939;
wire n19940;
wire n19941;
wire n19942;
wire n19943;
wire n19944;
wire n19945;
wire n19946;
wire n19947;
wire n19948;
wire n19949;
wire n19950;
wire n19951;
wire n19952;
wire n19953;
wire n19954;
wire n19955;
wire n19956;
wire n19957;
wire n19958;
wire n19959;
wire n19960;
wire n19961;
wire n19962;
wire n19963;
wire n19964;
wire n19965;
wire n19966;
wire n19967;
wire n19968;
wire n19969;
wire n19970;
wire n19971;
wire n19972;
wire n19973;
wire n19974;
wire n19975;
wire n19976;
wire n19977;
wire n19978;
wire n19979;
wire n19980;
wire n19981;
wire n19982;
wire n19983;
wire n19984;
wire n19985;
wire n19986;
wire n19987;
wire n19988;
wire n19989;
wire n19990;
wire n19991;
wire n19992;
wire n19993;
wire n19994;
wire n19995;
wire n19996;
wire n19997;
wire n19998;
wire n19999;
wire n20000;
wire n20001;
wire n20002;
wire n20003;
wire n20004;
wire n20005;
wire n20006;
wire n20007;
wire n20008;
wire n20009;
wire n20010;
wire n20011;
wire n20012;
wire n20013;
wire n20014;
wire n20015;
wire n20016;
wire n20017;
wire n20018;
wire n20019;
wire n20020;
wire n20021;
wire n20022;
wire n20023;
wire n20024;
wire n20025;
wire n20026;
wire n20027;
wire n20028;
wire n20029;
wire n20030;
wire n20031;
wire n20032;
wire n20033;
wire n20034;
wire n20035;
wire n20036;
wire n20037;
wire n20038;
wire n20039;
wire n20040;
wire n20041;
wire n20042;
wire n20043;
wire n20044;
wire n20045;
wire n20046;
wire n20047;
wire n20048;
wire n20049;
wire n20050;
wire n20051;
wire n20052;
wire n20053;
wire n20054;
wire n20055;
wire n20056;
wire n20057;
wire n20058;
wire n20059;
wire n20060;
wire n20061;
wire n20062;
wire n20063;
wire n20064;
wire n20065;
wire n20066;
wire n20067;
wire n20068;
wire n20069;
wire n20070;
wire n20071;
wire n20072;
wire n20073;
wire n20074;
wire n20075;
wire n20076;
wire n20077;
wire n20078;
wire n20079;
wire n20080;
wire n20081;
wire n20082;
wire n20083;
wire n20084;
wire n20085;
wire n20086;
wire n20087;
wire n20088;
wire n20089;
wire n20090;
wire n20091;
wire n20092;
wire n20093;
wire n20094;
wire n20095;
wire n20096;
wire n20097;
wire n20098;
wire n20099;
wire n20100;
wire n20101;
wire n20102;
wire n20103;
wire n20104;
wire n20105;
wire n20106;
wire n20107;
wire n20108;
wire n20109;
wire n20110;
wire n20111;
wire n20112;
wire n20113;
wire n20114;
wire n20115;
wire n20116;
wire n20117;
wire n20118;
wire n20119;
wire n20120;
wire n20121;
wire n20122;
wire n20123;
wire n20124;
wire n20125;
wire n20126;
wire n20127;
wire n20128;
wire n20129;
wire n20130;
wire n20131;
wire n20132;
wire n20133;
wire n20134;
wire n20135;
wire n20136;
wire n20137;
wire n20138;
wire n20139;
wire n20140;
wire n20141;
wire n20142;
wire n20143;
wire n20144;
wire n20145;
wire n20146;
wire n20147;
wire n20148;
wire n20149;
wire n20150;
wire n20151;
wire n20152;
wire n20153;
wire n20154;
wire n20155;
wire n20156;
wire n20157;
wire n20158;
wire n20159;
wire n20160;
wire n20161;
wire n20162;
wire n20163;
wire n20164;
wire n20165;
wire n20166;
wire n20167;
wire n20168;
wire n20169;
wire n20170;
wire n20171;
wire n20172;
wire n20173;
wire n20174;
wire n20175;
wire n20176;
wire n20177;
wire n20178;
wire n20179;
wire n20180;
wire n20181;
wire n20182;
wire n20183;
wire n20184;
wire n20185;
wire n20186;
wire n20187;
wire n20188;
wire n20189;
wire n20190;
wire n20191;
wire n20192;
wire n20193;
wire n20194;
wire n20195;
wire n20196;
wire n20197;
wire n20198;
wire n20199;
wire n20200;
wire n20201;
wire n20202;
wire n20203;
wire n20204;
wire n20205;
wire n20206;
wire n20207;
wire n20208;
wire n20209;
wire n20210;
wire n20211;
wire n20212;
wire n20213;
wire n20214;
wire n20215;
wire n20216;
wire n20217;
wire n20218;
wire n20219;
wire n20220;
wire n20221;
wire n20222;
wire n20223;
wire n20224;
wire n20225;
wire n20226;
wire n20227;
wire n20228;
wire n20229;
wire n20230;
wire n20231;
wire n20232;
wire n20233;
wire n20234;
wire n20235;
wire n20236;
wire n20237;
wire n20238;
wire n20239;
wire n20240;
wire n20241;
wire n20242;
wire n20243;
wire n20244;
wire n20245;
wire n20246;
wire n20247;
wire n20248;
wire n20249;
wire n20250;
wire n20251;
wire n20252;
wire n20253;
wire n20254;
wire n20255;
wire n20256;
wire n20257;
wire n20258;
wire n20259;
wire n20260;
wire n20261;
wire n20262;
wire n20263;
wire n20264;
wire n20265;
wire n20266;
wire n20267;
wire n20268;
wire n20269;
wire n20270;
wire n20271;
wire n20272;
wire n20273;
wire n20274;
wire n20275;
wire n20276;
wire n20277;
wire n20278;
wire n20279;
wire n20280;
wire n20281;
wire n20282;
wire n20283;
wire n20284;
wire n20285;
wire n20286;
wire n20287;
wire n20288;
wire n20289;
wire n20290;
wire n20291;
wire n20292;
wire n20293;
wire n20294;
wire n20295;
wire n20296;
wire n20297;
wire n20298;
wire n20299;
wire n20300;
wire n20301;
wire n20302;
wire n20303;
wire n20304;
wire n20305;
wire n20306;
wire n20307;
wire n20308;
wire n20309;
wire n20310;
wire n20311;
wire n20312;
wire n20313;
wire n20314;
wire n20315;
wire n20316;
wire n20317;
wire n20318;
wire n20319;
wire n20320;
wire n20321;
wire n20322;
wire n20323;
wire n20324;
wire n20325;
wire n20326;
wire n20327;
wire n20328;
wire n20329;
wire n20330;
wire n20331;
wire n20332;
wire n20333;
wire n20334;
wire n20335;
wire n20336;
wire n20337;
wire n20338;
wire n20339;
wire n20340;
wire n20341;
wire n20342;
wire n20343;
wire n20344;
wire n20345;
wire n20346;
wire n20347;
wire n20348;
wire n20349;
wire n20350;
wire n20351;
wire n20352;
wire n20353;
wire n20354;
wire n20355;
wire n20356;
wire n20357;
wire n20358;
wire n20359;
wire n20360;
wire n20361;
wire n20362;
wire n20363;
wire n20364;
wire n20365;
wire n20366;
wire n20367;
wire n20368;
wire n20369;
wire n20370;
wire n20371;
wire n20372;
wire n20373;
wire n20374;
wire n20375;
wire n20376;
wire n20377;
wire n20378;
wire n20379;
wire n20380;
wire n20381;
wire n20382;
wire n20383;
wire n20384;
wire n20385;
wire n20386;
wire n20387;
wire n20388;
wire n20389;
wire n20390;
wire n20391;
wire n20392;
wire n20393;
wire n20394;
wire n20395;
wire n20396;
wire n20397;
wire n20398;
wire n20399;
wire n20400;
wire n20401;
wire n20402;
wire n20403;
wire n20404;
wire n20405;
wire n20406;
wire n20407;
wire n20408;
wire n20409;
wire n20410;
wire n20411;
wire n20412;
wire n20413;
wire n20414;
wire n20415;
wire n20416;
wire n20417;
wire n20418;
wire n20419;
wire n20420;
wire n20421;
wire n20422;
wire n20423;
wire n20424;
wire n20425;
wire n20426;
wire n20427;
wire n20428;
wire n20429;
wire n20430;
wire n20431;
wire n20432;
wire n20433;
wire n20434;
wire n20435;
wire n20436;
wire n20437;
wire n20438;
wire n20439;
wire n20440;
wire n20441;
wire n20442;
wire n20443;
wire n20444;
wire n20445;
wire n20446;
wire n20447;
wire n20448;
wire n20449;
wire n20450;
wire n20451;
wire n20452;
wire n20453;
wire n20454;
wire n20455;
wire n20456;
wire n20457;
wire n20458;
wire n20459;
wire n20460;
wire n20461;
wire n20462;
wire n20463;
wire n20464;
wire n20465;
wire n20466;
wire n20467;
wire n20468;
wire n20469;
wire n20470;
wire n20471;
wire n20472;
wire n20473;
wire n20474;
wire n20475;
wire n20476;
wire n20477;
wire n20478;
wire n20479;
wire n20480;
wire n20481;
wire n20482;
wire n20483;
wire n20484;
wire n20485;
wire n20486;
wire n20487;
wire n20488;
wire n20489;
wire n20490;
wire n20491;
wire n20492;
wire n20493;
wire n20494;
wire n20495;
wire n20496;
wire n20497;
wire n20498;
wire n20499;
wire n20500;
wire n20501;
wire n20502;
wire n20503;
wire n20504;
wire n20505;
wire n20506;
wire n20507;
wire n20508;
wire n20509;
wire n20510;
wire n20511;
wire n20512;
wire n20513;
wire n20514;
wire n20515;
wire n20516;
wire n20517;
wire n20518;
wire n20519;
wire n20520;
wire n20521;
wire n20522;
wire n20523;
wire n20524;
wire n20525;
wire n20526;
wire n20527;
wire n20528;
wire n20529;
wire n20530;
wire n20531;
wire n20532;
wire n20533;
wire n20534;
wire n20535;
wire n20536;
wire n20537;
wire n20538;
wire n20539;
wire n20540;
wire n20541;
wire n20542;
wire n20543;
wire n20544;
wire n20545;
wire n20546;
wire n20547;
wire n20548;
wire n20549;
wire n20550;
wire n20551;
wire n20552;
wire n20553;
wire n20554;
wire n20555;
wire n20556;
wire n20557;
wire n20558;
wire n20559;
wire n20560;
wire n20561;
wire n20562;
wire n20563;
wire n20564;
wire n20565;
wire n20566;
wire n20567;
wire n20568;
wire n20569;
wire n20570;
wire n20571;
wire n20572;
wire n20573;
wire n20574;
wire n20575;
wire n20576;
wire n20577;
wire n20578;
wire n20579;
wire n20580;
wire n20581;
wire n20582;
wire n20583;
wire n20584;
wire n20585;
wire n20586;
wire n20587;
wire n20588;
wire n20589;
wire n20590;
wire n20591;
wire n20592;
wire n20593;
wire n20594;
wire n20595;
wire n20596;
wire n20597;
wire n20598;
wire n20599;
wire n20600;
wire n20601;
wire n20602;
wire n20603;
wire n20604;
wire n20605;
wire n20606;
wire n20607;
wire n20608;
wire n20609;
wire n20610;
wire n20611;
wire n20612;
wire n20613;
wire n20614;
wire n20615;
wire n20616;
wire n20617;
wire n20618;
wire n20619;
wire n20620;
wire n20621;
wire n20622;
wire n20623;
wire n20624;
wire n20625;
wire n20626;
wire n20627;
wire n20628;
wire n20629;
wire n20630;
wire n20631;
wire n20632;
wire n20633;
wire n20634;
wire n20635;
wire n20636;
wire n20637;
wire n20638;
wire n20639;
wire n20640;
wire n20641;
wire n20642;
wire n20643;
wire n20644;
wire n20645;
wire n20646;
wire n20647;
wire n20648;
wire n20649;
wire n20650;
wire n20651;
wire n20652;
wire n20653;
wire n20654;
wire n20655;
wire n20656;
wire n20657;
wire n20658;
wire n20659;
wire n20660;
wire n20661;
wire n20662;
wire n20663;
wire n20664;
wire n20665;
wire n20666;
wire n20667;
wire n20668;
wire n20669;
wire n20670;
wire n20671;
wire n20672;
wire n20673;
wire n20674;
wire n20675;
wire n20676;
wire n20677;
wire n20678;
wire n20679;
wire n20680;
wire n20681;
wire n20682;
wire n20683;
wire n20684;
wire n20685;
wire n20686;
wire n20687;
wire n20688;
wire n20689;
wire n20690;
wire n20691;
wire n20692;
wire n20693;
wire n20694;
wire n20695;
wire n20696;
wire n20697;
wire n20698;
wire n20699;
wire n20700;
wire n20701;
wire n20702;
wire n20703;
wire n20704;
wire n20705;
wire n20706;
wire n20707;
wire n20708;
wire n20709;
wire n20710;
wire n20711;
wire n20712;
wire n20713;
wire n20714;
wire n20715;
wire n20716;
wire n20717;
wire n20718;
wire n20719;
wire n20720;
wire n20721;
wire n20722;
wire n20723;
wire n20724;
wire n20725;
wire n20726;
wire n20727;
wire n20728;
wire n20729;
wire n20730;
wire n20731;
wire n20732;
wire n20733;
wire n20734;
wire n20735;
wire n20736;
wire n20737;
wire n20738;
wire n20739;
wire n20740;
wire n20741;
wire n20742;
wire n20743;
wire n20744;
wire n20745;
wire n20746;
wire n20747;
wire n20748;
wire n20749;
wire n20750;
wire n20751;
wire n20752;
wire n20753;
wire n20754;
wire n20755;
wire n20756;
wire n20757;
wire n20758;
wire n20759;
wire n20760;
wire n20761;
wire n20762;
wire n20763;
wire n20764;
wire n20765;
wire n20766;
wire n20767;
wire n20768;
wire n20769;
wire n20770;
wire n20771;
wire n20772;
wire n20773;
wire n20774;
wire n20775;
wire n20776;
wire n20777;
wire n20778;
wire n20779;
wire n20780;
wire n20781;
wire n20782;
wire n20783;
wire n20784;
wire n20785;
wire n20786;
wire n20787;
wire n20788;
wire n20789;
wire n20790;
wire n20791;
wire n20792;
wire n20793;
wire n20794;
wire n20795;
wire n20796;
wire n20797;
wire n20798;
wire n20799;
wire n20800;
wire n20801;
wire n20802;
wire n20803;
wire n20804;
wire n20805;
wire n20806;
wire n20807;
wire n20808;
wire n20809;
wire n20810;
wire n20811;
wire n20812;
wire n20813;
wire n20814;
wire n20815;
wire n20816;
wire n20817;
wire n20818;
wire n20819;
wire n20820;
wire n20821;
wire n20822;
wire n20823;
wire n20824;
wire n20825;
wire n20826;
wire n20827;
wire n20828;
wire n20829;
wire n20830;
wire n20831;
wire n20832;
wire n20833;
wire n20834;
wire n20835;
wire n20836;
wire n20837;
wire n20838;
wire n20839;
wire n20840;
wire n20841;
wire n20842;
wire n20843;
wire n20844;
wire n20845;
wire n20846;
wire n20847;
wire n20848;
wire n20849;
wire n20850;
wire n20851;
wire n20852;
wire n20853;
wire n20854;
wire n20855;
wire n20856;
wire n20857;
wire n20858;
wire n20859;
wire n20860;
wire n20861;
wire n20862;
wire n20863;
wire n20864;
wire n20865;
wire n20866;
wire n20867;
wire n20868;
wire n20869;
wire n20870;
wire n20871;
wire n20872;
wire n20873;
wire n20874;
wire n20875;
wire n20876;
wire n20877;
wire n20878;
wire n20879;
wire n20880;
wire n20881;
wire n20882;
wire n20883;
wire n20884;
wire n20885;
wire n20886;
wire n20887;
wire n20888;
wire n20889;
wire n20890;
wire n20891;
wire n20892;
wire n20893;
wire n20894;
wire n20895;
wire n20896;
wire n20897;
wire n20898;
wire n20899;
wire n20900;
wire n20901;
wire n20902;
wire n20903;
wire n20904;
wire n20905;
wire n20906;
wire n20907;
wire n20908;
wire n20909;
wire n20910;
wire n20911;
wire n20912;
wire n20913;
wire n20914;
wire n20915;
wire n20916;
wire n20917;
wire n20918;
wire n20919;
wire n20920;
wire n20921;
wire n20922;
wire n20923;
wire n20924;
wire n20925;
wire n20926;
wire n20927;
wire n20928;
wire n20929;
wire n20930;
wire n20931;
wire n20932;
wire n20933;
wire n20934;
wire n20935;
wire n20936;
wire n20937;
wire n20938;
wire n20939;
wire n20940;
wire n20941;
wire n20942;
wire n20943;
wire n20944;
wire n20945;
wire n20946;
wire n20947;
wire n20948;
wire n20949;
wire n20950;
wire n20951;
wire n20952;
wire n20953;
wire n20954;
wire n20955;
wire n20956;
wire n20957;
wire n20958;
wire n20959;
wire n20960;
wire n20961;
wire n20962;
wire n20963;
wire n20964;
wire n20965;
wire n20966;
wire n20967;
wire n20968;
wire n20969;
wire n20970;
wire n20971;
wire n20972;
wire n20973;
wire n20974;
wire n20975;
wire n20976;
wire n20977;
wire n20978;
wire n20979;
wire n20980;
wire n20981;
wire n20982;
wire n20983;
wire n20984;
wire n20985;
wire n20986;
wire n20987;
wire n20988;
wire n20989;
wire n20990;
wire n20991;
wire n20992;
wire n20993;
wire n20994;
wire n20995;
wire n20996;
wire n20997;
wire n20998;
wire n20999;
wire n21000;
wire n21001;
wire n21002;
wire n21003;
wire n21004;
wire n21005;
wire n21006;
wire n21007;
wire n21008;
wire n21009;
wire n21010;
wire n21011;
wire n21012;
wire n21013;
wire n21014;
wire n21015;
wire n21016;
wire n21017;
wire n21018;
wire n21019;
wire n21020;
wire n21021;
wire n21022;
wire n21023;
wire n21024;
wire n21025;
wire n21026;
wire n21027;
wire n21028;
wire n21029;
wire n21030;
wire n21031;
wire n21032;
wire n21033;
wire n21034;
wire n21035;
wire n21036;
wire n21037;
wire n21038;
wire n21039;
wire n21040;
wire n21041;
wire n21042;
wire n21043;
wire n21044;
wire n21045;
wire n21046;
wire n21047;
wire n21048;
wire n21049;
wire n21050;
wire n21051;
wire n21052;
wire n21053;
wire n21054;
wire n21055;
wire n21056;
wire n21057;
wire n21058;
wire n21059;
wire n21060;
wire n21061;
wire n21062;
wire n21063;
wire n21064;
wire n21065;
wire n21066;
wire n21067;
wire n21068;
wire n21069;
wire n21070;
wire n21071;
wire n21072;
wire n21073;
wire n21074;
wire n21075;
wire n21076;
wire n21077;
wire n21078;
wire n21079;
wire n21080;
wire n21081;
wire n21082;
wire n21083;
wire n21084;
wire n21085;
wire n21086;
wire n21087;
wire n21088;
wire n21089;
wire n21090;
wire n21091;
wire n21092;
wire n21093;
wire n21094;
wire n21095;
wire n21096;
wire n21097;
wire n21098;
wire n21099;
wire n21100;
wire n21101;
wire n21102;
wire n21103;
wire n21104;
wire n21105;
wire n21106;
wire n21107;
wire n21108;
wire n21109;
wire n21110;
wire n21111;
wire n21112;
wire n21113;
wire n21114;
wire n21115;
wire n21116;
wire n21117;
wire n21118;
wire n21119;
wire n21120;
wire n21121;
wire n21122;
wire n21123;
wire n21124;
wire n21125;
wire n21126;
wire n21127;
wire n21128;
wire n21129;
wire n21130;
wire n21131;
wire n21132;
wire n21133;
wire n21134;
wire n21135;
wire n21136;
wire n21137;
wire n21138;
wire n21139;
wire n21140;
wire n21141;
wire n21142;
wire n21143;
wire n21144;
wire n21145;
wire n21146;
wire n21147;
wire n21148;
wire n21149;
wire n21150;
wire n21151;
wire n21152;
wire n21153;
wire n21154;
wire n21155;
wire n21156;
wire n21157;
wire n21158;
wire n21159;
wire n21160;
wire n21161;
wire n21162;
wire n21163;
wire n21164;
wire n21165;
wire n21166;
wire n21167;
wire n21168;
wire n21169;
wire n21170;
wire n21171;
wire n21172;
wire n21173;
wire n21174;
wire n21175;
wire n21176;
wire n21177;
wire n21178;
wire n21179;
wire n21180;
wire n21181;
wire n21182;
wire n21183;
wire n21184;
wire n21185;
wire n21186;
wire n21187;
wire n21188;
wire n21189;
wire n21190;
wire n21191;
wire n21192;
wire n21193;
wire n21194;
wire n21195;
wire n21196;
wire n21197;
wire n21198;
wire n21199;
wire n21200;
wire n21201;
wire n21202;
wire n21203;
wire n21204;
wire n21205;
wire n21206;
wire n21207;
wire n21208;
wire n21209;
wire n21210;
wire n21211;
wire n21212;
wire n21213;
wire n21214;
wire n21215;
wire n21216;
wire n21217;
wire n21218;
wire n21219;
wire n21220;
wire n21221;
wire n21222;
wire n21223;
wire n21224;
wire n21225;
wire n21226;
wire n21227;
wire n21228;
wire n21229;
wire n21230;
wire n21231;
wire n21232;
wire n21233;
wire n21234;
wire n21235;
wire n21236;
wire n21237;
wire n21238;
wire n21239;
wire n21240;
wire n21241;
wire n21242;
wire n21243;
wire n21244;
wire n21245;
wire n21246;
wire n21247;
wire n21248;
wire n21249;
wire n21250;
wire n21251;
wire n21252;
wire n21253;
wire n21254;
wire n21255;
wire n21256;
wire n21257;
wire n21258;
wire n21259;
wire n21260;
wire n21261;
wire n21262;
wire n21263;
wire n21264;
wire n21265;
wire n21266;
wire n21267;
wire n21268;
wire n21269;
wire n21270;
wire n21271;
wire n21272;
wire n21273;
wire n21274;
wire n21275;
wire n21276;
wire n21277;
wire n21278;
wire n21279;
wire n21280;
wire n21281;
wire n21282;
wire n21283;
wire n21284;
wire n21285;
wire n21286;
wire n21287;
wire n21288;
wire n21289;
wire n21290;
wire n21291;
wire n21292;
wire n21293;
wire n21294;
wire n21295;
wire n21296;
wire n21297;
wire n21298;
wire n21299;
wire n21300;
wire n21301;
wire n21302;
wire n21303;
wire n21304;
wire n21305;
wire n21306;
wire n21307;
wire n21308;
wire n21309;
wire n21310;
wire n21311;
wire n21312;
wire n21313;
wire n21314;
wire n21315;
wire n21316;
wire n21317;
wire n21318;
wire n21319;
wire n21320;
wire n21321;
wire n21322;
wire n21323;
wire n21324;
wire n21325;
wire n21326;
wire n21327;
wire n21328;
wire n21329;
wire n21330;
wire n21331;
wire n21332;
wire n21333;
wire n21334;
wire n21335;
wire n21336;
wire n21337;
wire n21338;
wire n21339;
wire n21340;
wire n21341;
wire n21342;
wire n21343;
wire n21344;
wire n21345;
wire n21346;
wire n21347;
wire n21348;
wire n21349;
wire n21350;
wire n21351;
wire n21352;
wire n21353;
wire n21354;
wire n21355;
wire n21356;
wire n21357;
wire n21358;
wire n21359;
wire n21360;
wire n21361;
wire n21362;
wire n21363;
wire n21364;
wire n21365;
wire n21366;
wire n21367;
wire n21368;
wire n21369;
wire n21370;
wire n21371;
wire n21372;
wire n21373;
wire n21374;
wire n21375;
wire n21376;
wire n21377;
wire n21378;
wire n21379;
wire n21380;
wire n21381;
wire n21382;
wire n21383;
wire n21384;
wire n21385;
wire n21386;
wire n21387;
wire n21388;
wire n21389;
wire n21390;
wire n21391;
wire n21392;
wire n21393;
wire n21394;
wire n21395;
wire n21396;
wire n21397;
wire n21398;
wire n21399;
wire n21400;
wire n21401;
wire n21402;
wire n21403;
wire n21404;
wire n21405;
wire n21406;
wire n21407;
wire n21408;
wire n21409;
wire n21410;
wire n21411;
wire n21412;
wire n21413;
wire n21414;
wire n21415;
wire n21416;
wire n21417;
wire n21418;
wire n21419;
wire n21420;
wire n21421;
wire n21422;
wire n21423;
wire n21424;
wire n21425;
wire n21426;
wire n21427;
wire n21428;
wire n21429;
wire n21430;
wire n21431;
wire n21432;
wire n21433;
wire n21434;
wire n21435;
wire n21436;
wire n21437;
wire n21438;
wire n21439;
wire n21440;
wire n21441;
wire n21442;
wire n21443;
wire n21444;
wire n21445;
wire n21446;
wire n21447;
wire n21448;
wire n21449;
wire n21450;
wire n21451;
wire n21452;
wire n21453;
wire n21454;
wire n21455;
wire n21456;
wire n21457;
wire n21458;
wire n21459;
wire n21460;
wire n21461;
wire n21462;
wire n21463;
wire n21464;
wire n21465;
wire n21466;
wire n21467;
wire n21468;
wire n21469;
wire n21470;
wire n21471;
wire n21472;
wire n21473;
wire n21474;
wire n21475;
wire n21476;
wire n21477;
wire n21478;
wire n21479;
wire n21480;
wire n21481;
wire n21482;
wire n21483;
wire n21484;
wire n21485;
wire n21486;
wire n21487;
wire n21488;
wire n21489;
wire n21490;
wire n21491;
wire n21492;
wire n21493;
wire n21494;
wire n21495;
wire n21496;
wire n21497;
wire n21498;
wire n21499;
wire n21500;
xor (out,n0,n19817);
wire s0n0,s1n0,notn0;
or (n0,s0n0,s1n0);
not(notn0,n14125);
and (s0n0,notn0,n1);
and (s1n0,n14125,n13868);
wire s0n1,s1n1,notn1;
or (n1,s0n1,s1n1);
not(notn1,n8689);
and (s0n1,notn1,n2);
and (s1n1,n8689,n8697);
wire s0n2,s1n2,notn2;
or (n2,s0n2,s1n2);
not(notn2,n8696);
and (s0n2,notn2,n3);
and (s1n2,n8696,n4);
wire s0n4,s1n4,notn4;
or (n4,s0n4,s1n4);
not(notn4,n577);
and (s0n4,notn4,n5);
and (s1n4,n577,n8692);
or (n5,n6,n8690);
and (n6,n7,n567);
wire s0n7,s1n7,notn7;
or (n7,s0n7,s1n7);
not(notn7,n8689);
and (s0n7,notn7,n8);
and (s1n7,n8689,n2878);
wire s0n8,s1n8,notn8;
or (n8,s0n8,s1n8);
not(notn8,n2705);
and (s0n8,notn8,n9);
and (s1n8,n2705,n2700);
xor (n9,n10,n2677);
xor (n10,n11,n2578);
xor (n11,n12,n1680);
xor (n12,n13,n1585);
xor (n13,n14,n1241);
xor (n14,n15,n1074);
wire s0n15,s1n15,notn15;
or (n15,s0n15,s1n15);
not(notn15,n928);
and (s0n15,notn15,1'b0);
and (s1n15,n928,n17);
xor (n17,n18,n746);
wire s0n18,s1n18,notn18;
or (n18,s0n18,s1n18);
not(notn18,n592);
and (s0n18,notn18,1'b0);
and (s1n18,n592,n19);
wire s0n19,s1n19,notn19;
or (n19,s0n19,s1n19);
not(notn19,n575);
and (s0n19,notn19,n20);
and (s1n19,n575,n562);
wire s0n20,s1n20,notn20;
or (n20,s0n20,s1n20);
not(notn20,n22);
and (s0n20,notn20,1'b0);
and (s1n20,n22,n21);
and (n22,n23,n556);
and (n23,n24,n40);
or (n24,n25,n30,n34,n37);
and (n25,n26,n27);
and (n27,n28,n29);
and (n30,n31,n32);
and (n32,n33,n29);
not (n33,n28);
and (n34,n35,n36);
nor (n36,n33,n29);
and (n37,n38,n39);
nor (n39,n28,n29);
and (n40,n41,n555);
not (n41,n42);
wire s0n42,s1n42,notn42;
or (n42,s0n42,s1n42);
not(notn42,n554);
and (s0n42,notn42,n43);
and (s1n42,n554,1'b0);
wire s0n43,s1n43,notn43;
or (n43,s0n43,s1n43);
not(notn43,n184);
and (s0n43,notn43,n44);
and (s1n43,n184,n45);
wire s0n45,s1n45,notn45;
or (n45,s0n45,s1n45);
not(notn45,n547);
and (s0n45,notn45,n46);
and (s1n45,n547,n521);
or (n46,n47,n489,n520,1'b0,1'b0,1'b0,1'b0,1'b0);
or (n47,n48,n488);
or (n48,n49,n487);
or (n49,n50,n486);
or (n50,n51,n484);
or (n51,n52,n483);
or (n52,n53,n481);
or (n53,n54,n479);
nor (n54,n55,n404,n413,n425,n437,n448,n459,n470);
or (n55,1'b0,n56,n398,n402);
and (n56,n57,n397);
wire s0n57,s1n57,notn57;
or (n57,s0n57,s1n57);
not(notn57,n388);
and (s0n57,notn57,n58);
and (s1n57,n388,n296);
wire s0n58,s1n58,notn58;
or (n58,s0n58,s1n58);
not(notn58,n255);
and (s0n58,notn58,1'b0);
and (s1n58,n255,n59);
or (n59,n60,n236,n240,n244,n247,n250,n252,1'b0);
and (n60,n61,n63);
not (n61,n62);
and (n63,n64,n209,n220,n230);
wire s0n64,s1n64,notn64;
or (n64,s0n64,s1n64);
not(notn64,n98);
and (s0n64,notn64,n65);
and (s1n64,n98,1'b0);
wire s0n65,s1n65,notn65;
or (n65,s0n65,s1n65);
not(notn65,n96);
and (s0n65,notn65,n66);
and (s1n65,n96,n94);
wire s0n66,s1n66,notn66;
or (n66,s0n66,s1n66);
not(notn66,n90);
and (s0n66,notn66,n67);
and (s1n66,n90,n84);
wire s0n67,s1n67,notn67;
or (n67,s0n67,s1n67);
not(notn67,n83);
and (s0n67,notn67,n68);
and (s1n67,n83,1'b0);
wire s0n68,s1n68,notn68;
or (n68,s0n68,s1n68);
not(notn68,n82);
and (s0n68,notn68,n69);
and (s1n68,n82,1'b1);
wire s0n69,s1n69,notn69;
or (n69,s0n69,s1n69);
not(notn69,n81);
and (s0n69,notn69,n70);
and (s1n69,n81,1'b0);
wire s0n70,s1n70,notn70;
or (n70,s0n70,s1n70);
not(notn70,n80);
and (s0n70,notn70,n71);
and (s1n70,n80,1'b1);
wire s0n71,s1n71,notn71;
or (n71,s0n71,s1n71);
not(notn71,n79);
and (s0n71,notn71,n72);
and (s1n71,n79,1'b0);
wire s0n72,s1n72,notn72;
or (n72,s0n72,s1n72);
not(notn72,n78);
and (s0n72,notn72,n73);
and (s1n72,n78,1'b1);
wire s0n73,s1n73,notn73;
or (n73,s0n73,s1n73);
not(notn73,n77);
and (s0n73,notn73,n74);
and (s1n73,n77,1'b0);
wire s0n74,s1n74,notn74;
or (n74,s0n74,s1n74);
not(notn74,n76);
and (s0n74,notn74,n61);
and (s1n74,n76,1'b1);
wire s0n84,s1n84,notn84;
or (n84,s0n84,s1n84);
not(notn84,n89);
and (s0n84,notn84,n85);
and (s1n84,n89,1'b0);
wire s0n85,s1n85,notn85;
or (n85,s0n85,s1n85);
not(notn85,n88);
and (s0n85,notn85,n86);
and (s1n85,n88,1'b1);
not (n86,n87);
or (n90,n91,n93);
or (n91,n92,n87);
or (n92,n89,n88);
not (n94,n95);
or (n96,n95,n97);
not (n98,n99);
or (n99,n100,n207);
or (n100,n101,n205);
or (n101,n102,n199);
or (n102,n103,n198);
or (n103,n104,n194);
or (n104,n105,n193);
or (n105,n106,n188);
or (n106,n107,n187);
or (n107,n108,n186);
or (n108,n109,n184);
or (n109,n110,n178);
or (n110,n111,n177);
or (n111,n112,n176);
or (n112,n113,n175);
or (n113,n114,n174);
or (n114,n115,n173);
or (n115,n116,n172);
or (n116,n117,n171);
or (n117,n118,n168);
or (n118,n119,n162);
or (n119,n120,n161);
or (n120,n121,n160);
or (n121,n122,n159);
or (n122,n123,n158);
or (n123,n124,n157);
or (n124,n125,n155);
or (n125,n126,n153);
or (n126,n127,n147);
or (n127,n128,n146);
or (n128,n129,n145);
or (n129,n130,n144);
or (n130,n131,n143);
or (n131,n132,n141);
or (n132,n133,n139);
nor (n133,n134,n135,n137,n138);
not (n135,n136);
nor (n139,n134,n135,n140,n138);
not (n140,n137);
and (n141,n134,n136,n137,n142);
not (n142,n138);
and (n143,n134,n135,n137,n142);
nor (n144,n134,n136,n140,n138);
and (n145,n134,n135,n137,n138);
and (n146,n134,n136,n137,n138);
nor (n147,n148,n150,n151,n152);
not (n148,n149);
nor (n153,n148,n154,n151,n152);
not (n154,n150);
and (n155,n148,n150,n151,n156);
not (n156,n152);
and (n157,n149,n150,n151,n156);
and (n158,n149,n154,n151,n156);
and (n159,n148,n154,n151,n152);
and (n160,n149,n154,n151,n152);
and (n161,n149,n150,n151,n152);
nor (n162,n163,n165,n166,n167);
not (n163,n164);
and (n168,n164,n165,n169,n170);
not (n169,n166);
not (n170,n167);
and (n171,n163,n165,n169,n170);
and (n172,n164,n165,n166,n170);
nor (n173,n164,n165,n169,n170);
and (n174,n163,n165,n166,n167);
and (n175,n163,n165,n169,n167);
and (n176,n164,n165,n169,n167);
nor (n177,n163,n165,n166,n170);
nor (n178,n179,n181,n182,n183);
not (n179,n180);
nor (n184,n180,n185,n182,n183);
not (n185,n181);
and (n186,n179,n185,n182,n183);
and (n187,n180,n185,n182,n183);
nor (n188,n189,n190,n192);
not (n190,n191);
and (n193,n189,n191,n192);
and (n194,n195,n196);
not (n196,n197);
nor (n198,n195,n196);
nor (n199,n200,n201,n203,n204);
not (n201,n202);
and (n205,n200,n202,n203,n206);
not (n206,n204);
and (n207,n208,n201,n203,n206);
not (n208,n200);
wire s0n209,s1n209,notn209;
or (n209,s0n209,s1n209);
not(notn209,n98);
and (s0n209,notn209,n210);
and (s1n209,n98,1'b0);
wire s0n210,s1n210,notn210;
or (n210,s0n210,s1n210);
not(notn210,n96);
and (s0n210,notn210,n211);
and (s1n210,n96,1'b0);
wire s0n211,s1n211,notn211;
or (n211,s0n211,s1n211);
not(notn211,n90);
and (s0n211,notn211,n212);
and (s1n211,n90,n92);
wire s0n212,s1n212,notn212;
or (n212,s0n212,s1n212);
not(notn212,n83);
and (s0n212,notn212,n213);
and (s1n212,n83,1'b1);
wire s0n213,s1n213,notn213;
or (n213,s0n213,s1n213);
not(notn213,n82);
and (s0n213,notn213,n214);
and (s1n213,n82,1'b1);
wire s0n214,s1n214,notn214;
or (n214,s0n214,s1n214);
not(notn214,n81);
and (s0n214,notn214,n215);
and (s1n214,n81,1'b0);
wire s0n215,s1n215,notn215;
or (n215,s0n215,s1n215);
not(notn215,n80);
and (s0n215,notn215,n216);
and (s1n215,n80,1'b0);
wire s0n216,s1n216,notn216;
or (n216,s0n216,s1n216);
not(notn216,n79);
and (s0n216,notn216,n217);
and (s1n216,n79,1'b1);
wire s0n217,s1n217,notn217;
or (n217,s0n217,s1n217);
not(notn217,n78);
and (s0n217,notn217,n218);
and (s1n217,n78,1'b1);
wire s0n218,s1n218,notn218;
or (n218,s0n218,s1n218);
not(notn218,n77);
and (s0n218,notn218,n219);
and (s1n218,n77,1'b0);
not (n219,n76);
wire s0n220,s1n220,notn220;
or (n220,s0n220,s1n220);
not(notn220,n98);
and (s0n220,notn220,n221);
and (s1n220,n98,1'b0);
wire s0n221,s1n221,notn221;
or (n221,s0n221,s1n221);
not(notn221,n96);
and (s0n221,notn221,n222);
and (s1n221,n96,1'b0);
wire s0n222,s1n222,notn222;
or (n222,s0n222,s1n222);
not(notn222,n90);
and (s0n222,notn222,n223);
and (s1n222,n90,n229);
wire s0n223,s1n223,notn223;
or (n223,s0n223,s1n223);
not(notn223,n83);
and (s0n223,notn223,n224);
and (s1n223,n83,1'b1);
wire s0n224,s1n224,notn224;
or (n224,s0n224,s1n224);
not(notn224,n82);
and (s0n224,notn224,n225);
and (s1n224,n82,1'b1);
wire s0n225,s1n225,notn225;
or (n225,s0n225,s1n225);
not(notn225,n81);
and (s0n225,notn225,n226);
and (s1n225,n81,1'b0);
wire s0n226,s1n226,notn226;
or (n226,s0n226,s1n226);
not(notn226,n80);
and (s0n226,notn226,n227);
and (s1n226,n80,1'b0);
wire s0n227,s1n227,notn227;
or (n227,s0n227,s1n227);
not(notn227,n79);
and (s0n227,notn227,n228);
and (s1n227,n79,1'b0);
not (n228,n78);
not (n229,n92);
not (n230,n231);
wire s0n231,s1n231,notn231;
or (n231,s0n231,s1n231);
not(notn231,n98);
and (s0n231,notn231,n232);
and (s1n231,n98,1'b0);
wire s0n232,s1n232,notn232;
or (n232,s0n232,s1n232);
not(notn232,n96);
and (s0n232,notn232,n233);
and (s1n232,n96,1'b0);
wire s0n233,s1n233,notn233;
or (n233,s0n233,s1n233);
not(notn233,n90);
and (s0n233,notn233,n234);
and (s1n233,n90,1'b0);
wire s0n234,s1n234,notn234;
or (n234,s0n234,s1n234);
not(notn234,n83);
and (s0n234,notn234,n235);
and (s1n234,n83,1'b0);
not (n235,n82);
and (n236,n237,n238);
not (n237,n77);
and (n238,n239,n209,n220,n230);
not (n239,n64);
and (n240,n241,n242);
not (n241,n79);
and (n242,n64,n243,n220,n230);
not (n243,n209);
and (n244,n245,n246);
not (n245,n81);
and (n246,n239,n243,n220,n230);
and (n247,n248,n249);
not (n248,n83);
nor (n249,n239,n243,n220,n231);
and (n250,n86,n251);
nor (n251,n64,n243,n220,n231);
and (n252,n253,n254);
not (n253,n89);
nor (n254,n239,n209,n220,n231);
or (n255,n256,n285);
wire s0n256,s1n256,notn256;
or (n256,s0n256,s1n256);
not(notn256,n283);
and (s0n256,notn256,n257);
and (s1n256,n283,1'b0);
wire s0n257,s1n257,notn257;
or (n257,s0n257,s1n257);
not(notn257,n282);
and (s0n257,notn257,n258);
and (s1n257,n282,n277);
wire s0n258,s1n258,notn258;
or (n258,s0n258,s1n258);
not(notn258,n276);
and (s0n258,notn258,n259);
and (s1n258,n276,n265);
wire s0n259,s1n259,notn259;
or (n259,s0n259,s1n259);
not(notn259,n264);
and (s0n259,notn259,n260);
and (s1n259,n264,n127);
or (n260,n261,n158);
or (n261,n262,n157);
or (n262,n263,n155);
or (n263,n147,n153);
or (n264,n134,n136,n137,n138);
or (n265,1'b0,1'b0,n266,n272,n274);
and (n266,n267,n270);
or (n267,1'b0,1'b0,n268,n188);
and (n268,n269,n191,n192);
not (n269,n189);
and (n270,n179,n185,n182,n271);
not (n271,n183);
and (n272,n195,n273);
and (n273,n180,n185,n182,n271);
or (n274,n275,n186);
or (n275,n178,n184);
or (n276,n180,n181,n182,n183);
or (n277,n278,n177);
or (n278,n279,n175);
or (n279,n280,n172);
or (n280,n281,n171);
or (n281,n162,n168);
or (n282,n164,n165,n166,n167);
not (n283,n284);
wire s0n285,s1n285,notn285;
or (n285,s0n285,s1n285);
not(notn285,n283);
and (s0n285,notn285,n286);
and (s1n285,n283,1'b0);
wire s0n286,s1n286,notn286;
or (n286,s0n286,s1n286);
not(notn286,n282);
and (s0n286,notn286,n287);
and (s1n286,n282,n295);
wire s0n287,s1n287,notn287;
or (n287,s0n287,s1n287);
not(notn287,n276);
and (s0n287,notn287,n288);
and (s1n287,n276,n291);
wire s0n288,s1n288,notn288;
or (n288,s0n288,s1n288);
not(notn288,n264);
and (s0n288,notn288,n289);
and (s1n288,n264,1'b0);
or (n289,n290,n161);
or (n290,n159,n160);
or (n291,1'b0,n187,n292,n294,1'b0);
and (n292,n293,n270);
or (n293,1'b0,n193,n268,1'b0);
and (n294,n197,n273);
or (n295,n174,n176);
not (n296,n297);
nor (n297,n58,n298,n314,n334,n351,n365,n376,n384);
wire s0n298,s1n298,notn298;
or (n298,s0n298,s1n298);
not(notn298,n255);
and (s0n298,notn298,1'b0);
and (s1n298,n255,n299);
or (n299,n300,n302,n304,n306,n308,n310,n312,1'b0);
and (n300,n301,n63);
xnor (n301,n76,n62);
and (n302,n303,n238);
xnor (n303,n78,n77);
and (n304,n305,n242);
xnor (n305,n80,n79);
and (n306,n307,n246);
xnor (n307,n82,n81);
and (n308,n309,n249);
xnor (n309,n93,n83);
and (n310,n311,n251);
xnor (n311,n88,n87);
and (n312,n313,n254);
xnor (n313,n97,n89);
wire s0n314,s1n314,notn314;
or (n314,s0n314,s1n314);
not(notn314,n255);
and (s0n314,notn314,1'b0);
and (s1n314,n255,n315);
or (n315,n316,n319,n322,n325,n328,n331,1'b0,1'b0);
and (n316,n317,n63);
xnor (n317,n77,n318);
or (n318,n76,n62);
and (n319,n320,n238);
xnor (n320,n79,n321);
or (n321,n78,n77);
and (n322,n323,n242);
xnor (n323,n81,n324);
or (n324,n80,n79);
and (n325,n326,n246);
xnor (n326,n83,n327);
or (n327,n82,n81);
and (n328,n329,n249);
xnor (n329,n87,n330);
or (n330,n93,n83);
and (n331,n332,n251);
xnor (n332,n89,n333);
or (n333,n88,n87);
wire s0n334,s1n334,notn334;
or (n334,s0n334,s1n334);
not(notn334,n255);
and (s0n334,notn334,1'b0);
and (s1n334,n255,n335);
or (n335,n336,n339,n342,n345,n348,1'b0,1'b0,1'b0);
and (n336,n337,n63);
xnor (n337,n78,n338);
or (n338,n77,n318);
and (n339,n340,n238);
xnor (n340,n80,n341);
or (n341,n79,n321);
and (n342,n343,n242);
xnor (n343,n82,n344);
or (n344,n81,n324);
and (n345,n346,n246);
xnor (n346,n93,n347);
or (n347,n83,n327);
and (n348,n349,n249);
xnor (n349,n88,n350);
or (n350,n87,n330);
wire s0n351,s1n351,notn351;
or (n351,s0n351,s1n351);
not(notn351,n255);
and (s0n351,notn351,1'b0);
and (s1n351,n255,n352);
or (n352,n353,n356,n359,n362,1'b0,1'b0,1'b0,1'b0);
and (n353,n354,n63);
xnor (n354,n79,n355);
or (n355,n78,n338);
and (n356,n357,n238);
xnor (n357,n81,n358);
or (n358,n80,n341);
and (n359,n360,n242);
xnor (n360,n83,n361);
or (n361,n82,n344);
and (n362,n363,n246);
xnor (n363,n87,n364);
or (n364,n93,n347);
wire s0n365,s1n365,notn365;
or (n365,s0n365,s1n365);
not(notn365,n255);
and (s0n365,notn365,1'b0);
and (s1n365,n255,n366);
or (n366,n367,n370,n373,1'b0,1'b0,1'b0,1'b0,1'b0);
and (n367,n368,n63);
xnor (n368,n80,n369);
or (n369,n79,n355);
and (n370,n371,n238);
xnor (n371,n82,n372);
or (n372,n81,n358);
and (n373,n374,n242);
xnor (n374,n93,n375);
or (n375,n83,n361);
wire s0n376,s1n376,notn376;
or (n376,s0n376,s1n376);
not(notn376,n255);
and (s0n376,notn376,1'b0);
and (s1n376,n255,n377);
or (n377,n378,n381,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0);
and (n378,n379,n63);
xnor (n379,n81,n380);
or (n380,n80,n369);
and (n381,n382,n238);
xnor (n382,n83,n383);
or (n383,n82,n372);
wire s0n384,s1n384,notn384;
or (n384,s0n384,s1n384);
not(notn384,n255);
and (s0n384,notn384,1'b0);
and (s1n384,n255,n385);
and (n385,n386,n63);
xnor (n386,n82,n387);
or (n387,n81,n380);
nor (n388,n389,n391,n394);
not (n389,n390);
not (n391,n392);
xor (n392,n393,n390);
xor (n394,n395,n396);
and (n396,n393,n390);
and (n397,n256,n285);
and (n398,n399,n400);
xor (n399,n298,n58);
nor (n400,n256,n401);
not (n401,n285);
and (n402,n58,n403);
and (n403,n256,n401);
not (n404,n405);
or (n405,1'b0,n406,n408,n412);
and (n406,n407,n397);
wire s0n407,s1n407,notn407;
or (n407,s0n407,s1n407);
not(notn407,n388);
and (s0n407,notn407,n298);
and (s1n407,n388,1'b0);
and (n408,n409,n400);
xor (n409,n410,n411);
not (n410,n314);
not (n411,n298);
and (n412,n298,n403);
or (n413,1'b0,n414,n416,n424);
and (n414,n415,n397);
wire s0n415,s1n415,notn415;
or (n415,s0n415,s1n415);
not(notn415,n388);
and (s0n415,notn415,n314);
and (s1n415,n388,1'b0);
and (n416,n417,n400);
wire s0n417,s1n417,notn417;
or (n417,s0n417,s1n417);
not(notn417,n58);
and (s0n417,notn417,n418);
and (s1n417,n58,n421);
xor (n418,n419,n420);
not (n419,n334);
and (n420,n410,n411);
xor (n421,n334,n422);
and (n422,n314,n423);
and (n423,n298,n58);
and (n424,n314,n403);
not (n425,n426);
or (n426,1'b0,n427,n429,n436);
and (n427,n428,n397);
wire s0n428,s1n428,notn428;
or (n428,s0n428,s1n428);
not(notn428,n388);
and (s0n428,notn428,n334);
and (s1n428,n388,1'b0);
and (n429,n430,n400);
wire s0n430,s1n430,notn430;
or (n430,s0n430,s1n430);
not(notn430,n58);
and (s0n430,notn430,n431);
and (s1n430,n58,n434);
xor (n431,n432,n433);
not (n432,n351);
and (n433,n419,n420);
xor (n434,n351,n435);
and (n435,n334,n422);
and (n436,n334,n403);
or (n437,1'b0,n438,n440,n447);
and (n438,n439,n397);
wire s0n439,s1n439,notn439;
or (n439,s0n439,s1n439);
not(notn439,n388);
and (s0n439,notn439,n351);
and (s1n439,n388,1'b0);
and (n440,n441,n400);
wire s0n441,s1n441,notn441;
or (n441,s0n441,s1n441);
not(notn441,n58);
and (s0n441,notn441,n442);
and (s1n441,n58,n445);
xor (n442,n443,n444);
not (n443,n365);
and (n444,n432,n433);
xor (n445,n365,n446);
and (n446,n351,n435);
and (n447,n351,n403);
or (n448,1'b0,n449,n451,n458);
and (n449,n450,n397);
wire s0n450,s1n450,notn450;
or (n450,s0n450,s1n450);
not(notn450,n388);
and (s0n450,notn450,n365);
and (s1n450,n388,1'b0);
and (n451,n452,n400);
wire s0n452,s1n452,notn452;
or (n452,s0n452,s1n452);
not(notn452,n58);
and (s0n452,notn452,n453);
and (s1n452,n58,n456);
xor (n453,n454,n455);
not (n454,n376);
and (n455,n443,n444);
xor (n456,n376,n457);
and (n457,n365,n446);
and (n458,n365,n403);
or (n459,1'b0,n460,n462,n469);
and (n460,n461,n397);
wire s0n461,s1n461,notn461;
or (n461,s0n461,s1n461);
not(notn461,n388);
and (s0n461,notn461,n376);
and (s1n461,n388,1'b0);
and (n462,n463,n400);
wire s0n463,s1n463,notn463;
or (n463,s0n463,s1n463);
not(notn463,n58);
and (s0n463,notn463,n464);
and (s1n463,n58,n467);
xor (n464,n465,n466);
not (n465,n384);
and (n466,n454,n455);
xor (n467,n384,n468);
and (n468,n376,n457);
and (n469,n376,n403);
or (n470,1'b0,n471,n473,n478);
and (n471,n472,n397);
wire s0n472,s1n472,notn472;
or (n472,s0n472,s1n472);
not(notn472,n388);
and (s0n472,notn472,n384);
and (s1n472,n388,1'b0);
and (n473,n474,n400);
wire s0n474,s1n474,notn474;
or (n474,s0n474,s1n474);
not(notn474,n58);
and (s0n474,notn474,n475);
and (s1n474,n58,n477);
not (n475,n476);
and (n476,n465,n466);
and (n477,n384,n468);
and (n478,n384,n403);
nor (n479,n480,n404,n413,n425,n437,n448,n459,n470);
not (n480,n55);
nor (n481,n55,n405,n482,n425,n437,n448,n459,n470);
not (n482,n413);
nor (n483,n480,n405,n482,n425,n437,n448,n459,n470);
nor (n484,n55,n404,n482,n426,n485,n448,n459,n470);
not (n485,n437);
nor (n486,n480,n404,n482,n426,n485,n448,n459,n470);
nor (n487,n55,n405,n413,n425,n485,n448,n459,n470);
nor (n488,n480,n405,n413,n425,n485,n448,n459,n470);
or (n489,n490,n505);
or (n490,n491,n504);
or (n491,n492,n503);
or (n492,n493,n502);
or (n493,n494,n501);
or (n494,n495,n500);
or (n495,n496,n499);
or (n496,n497,n498);
nor (n497,n55,n404,n482,n426,n437,n448,n459,n470);
nor (n498,n480,n404,n482,n426,n437,n448,n459,n470);
nor (n499,n55,n405,n413,n425,n437,n448,n459,n470);
nor (n500,n480,n405,n413,n425,n437,n448,n459,n470);
nor (n501,n55,n404,n413,n426,n485,n448,n459,n470);
nor (n502,n480,n404,n413,n426,n485,n448,n459,n470);
nor (n503,n55,n405,n482,n426,n485,n448,n459,n470);
nor (n504,n480,n405,n482,n426,n485,n448,n459,n470);
or (n505,n506,n519);
or (n506,n507,n518);
or (n507,n508,n517);
or (n508,n509,n516);
or (n509,n510,n515);
or (n510,n511,n514);
or (n511,n512,n513);
nor (n512,n55,n404,n482,n425,n437,n448,n459,n470);
nor (n513,n480,n404,n482,n425,n437,n448,n459,n470);
nor (n514,n55,n405,n413,n426,n485,n448,n459,n470);
nor (n515,n480,n405,n413,n426,n485,n448,n459,n470);
nor (n516,n55,n404,n413,n425,n485,n448,n459,n470);
nor (n517,n480,n404,n413,n425,n485,n448,n459,n470);
nor (n518,n55,n405,n482,n425,n485,n448,n459,n470);
nor (n519,n480,n405,n482,n425,n485,n448,n459,n470);
nor (n520,n480,n405,n482,n426,n437,n448,n459,n470);
or (n521,1'b0,n522,n529,n536,n297);
or (n522,n523,n487);
or (n523,n524,n486);
or (n524,n525,n484);
or (n525,n526,n504);
or (n526,n527,n481);
or (n527,n528,n479);
or (n528,n500,n54);
or (n529,n530,n503);
or (n530,n531,n502);
or (n531,n532,n501);
or (n532,n533,n515);
or (n533,n534,n499);
or (n534,n535,n498);
or (n535,n520,n497);
or (n536,n537,n514);
or (n537,n538,n513);
or (n538,n539,n512);
or (n539,n540,n483);
or (n540,n541,n546);
or (n541,n542,n545);
or (n542,n543,n544);
nor (n543,n480,n405,n413,n426,n437,n448,n459,n470);
nor (n544,n55,n404,n413,n426,n437,n448,n459,n470);
nor (n545,n480,n404,n413,n426,n437,n448,n459,n470);
nor (n546,n55,n405,n482,n426,n437,n448,n459,n470);
or (n547,n548,n553);
nor (n548,n549,n550,n552);
not (n550,n551);
and (n553,n549,n551,n552);
nor (n554,n179,n185,n182,n183);
nor (n556,n557,n559,n560,n561);
not (n557,n558);
or (n562,1'b0,n563,n565,n569,n572);
and (n563,n564,n556);
and (n565,n566,n567);
nor (n567,n558,n568,n560,n561);
not (n568,n559);
and (n569,n570,n571);
nor (n571,n557,n568,n560,n561);
and (n572,n21,n573);
and (n573,n557,n568,n560,n574);
not (n574,n561);
and (n575,n40,n576);
not (n576,n577);
wire s0n577,s1n577,notn577;
or (n577,s0n577,s1n577);
not(notn577,n590);
and (s0n577,notn577,n23);
and (s1n577,n590,n578);
or (n578,n579,n583,n586,n588);
and (n579,n26,n580);
and (n580,n581,n582);
and (n583,n31,n584);
and (n584,n585,n582);
not (n585,n581);
and (n586,n35,n587);
nor (n587,n585,n582);
and (n588,n38,n589);
nor (n589,n581,n582);
and (n590,n41,n591);
not (n591,n555);
and (n592,n593,n649);
not (n593,n594);
wire s0n594,s1n594,notn594;
or (n594,s0n594,s1n594);
not(notn594,n40);
and (s0n594,notn594,1'b0);
and (s1n594,n40,n595);
wire s0n595,s1n595,notn595;
or (n595,s0n595,s1n595);
not(notn595,n648);
and (s0n595,notn595,n596);
and (s1n595,n648,n639);
or (n596,n597,n615,n626,n637);
and (n597,n598,n27);
wire s0n598,s1n598,notn598;
or (n598,s0n598,s1n598);
not(notn598,n577);
and (s0n598,notn598,n599);
and (s1n598,n577,n600);
or (n600,n601,n606,n610,n613);
and (n601,n602,n603);
nor (n603,n604,n605);
and (n606,n607,n608);
nor (n608,n609,n605);
not (n609,n604);
and (n610,n611,n612);
and (n612,n609,n605);
and (n613,n599,n614);
and (n614,n604,n605);
and (n615,n616,n32);
wire s0n616,s1n616,notn616;
or (n616,s0n616,s1n616);
not(notn616,n577);
and (s0n616,notn616,n617);
and (s1n616,n577,n618);
or (n618,n619,n621,n623,n625);
and (n619,n620,n603);
and (n621,n622,n608);
and (n623,n624,n612);
and (n625,n617,n614);
and (n626,n627,n36);
wire s0n627,s1n627,notn627;
or (n627,s0n627,s1n627);
not(notn627,n577);
and (s0n627,notn627,n628);
and (s1n627,n577,n629);
or (n629,n630,n632,n634,n636);
and (n630,n631,n603);
and (n632,n633,n608);
and (n634,n635,n612);
and (n636,n628,n614);
and (n637,n638,n39);
wire s0n638,s1n638,notn638;
or (n638,s0n638,s1n638);
not(notn638,n577);
and (s0n638,notn638,n639);
and (s1n638,n577,n640);
or (n640,n641,n643,n645,n647);
and (n641,n642,n603);
and (n643,n644,n608);
and (n645,n646,n612);
and (n647,n639,n614);
and (n649,n650,n698);
not (n650,n651);
wire s0n651,s1n651,notn651;
or (n651,s0n651,s1n651);
not(notn651,n40);
and (s0n651,notn651,1'b0);
and (s1n651,n40,n652);
wire s0n652,s1n652,notn652;
or (n652,s0n652,s1n652);
not(notn652,n648);
and (s0n652,notn652,n653);
and (s1n652,n648,n689);
or (n653,n654,n665,n676,n687);
and (n654,n655,n27);
wire s0n655,s1n655,notn655;
or (n655,s0n655,s1n655);
not(notn655,n577);
and (s0n655,notn655,n656);
and (s1n655,n577,n657);
or (n657,n658,n660,n662,n664);
and (n658,n659,n603);
and (n660,n661,n608);
and (n662,n663,n612);
and (n664,n656,n614);
and (n665,n666,n32);
wire s0n666,s1n666,notn666;
or (n666,s0n666,s1n666);
not(notn666,n577);
and (s0n666,notn666,n667);
and (s1n666,n577,n668);
or (n668,n669,n671,n673,n675);
and (n669,n670,n603);
and (n671,n672,n608);
and (n673,n674,n612);
and (n675,n667,n614);
and (n676,n677,n36);
wire s0n677,s1n677,notn677;
or (n677,s0n677,s1n677);
not(notn677,n577);
and (s0n677,notn677,n678);
and (s1n677,n577,n679);
or (n679,n680,n682,n684,n686);
and (n680,n681,n603);
and (n682,n683,n608);
and (n684,n685,n612);
and (n686,n678,n614);
and (n687,n688,n39);
wire s0n688,s1n688,notn688;
or (n688,s0n688,s1n688);
not(notn688,n577);
and (s0n688,notn688,n689);
and (s1n688,n577,n690);
or (n690,n691,n693,n695,n697);
and (n691,n692,n603);
and (n693,n694,n608);
and (n695,n696,n612);
and (n697,n689,n614);
not (n698,n699);
wire s0n699,s1n699,notn699;
or (n699,s0n699,s1n699);
not(notn699,n40);
and (s0n699,notn699,1'b0);
and (s1n699,n40,n700);
wire s0n700,s1n700,notn700;
or (n700,s0n700,s1n700);
not(notn700,n648);
and (s0n700,notn700,n701);
and (s1n700,n648,n737);
or (n701,n702,n713,n724,n735);
and (n702,n703,n27);
wire s0n703,s1n703,notn703;
or (n703,s0n703,s1n703);
not(notn703,n577);
and (s0n703,notn703,n704);
and (s1n703,n577,n705);
or (n705,n706,n708,n710,n712);
and (n706,n707,n603);
and (n708,n709,n608);
and (n710,n711,n612);
and (n712,n704,n614);
and (n713,n714,n32);
wire s0n714,s1n714,notn714;
or (n714,s0n714,s1n714);
not(notn714,n577);
and (s0n714,notn714,n715);
and (s1n714,n577,n716);
or (n716,n717,n719,n721,n723);
and (n717,n718,n603);
and (n719,n720,n608);
and (n721,n722,n612);
and (n723,n715,n614);
and (n724,n725,n36);
wire s0n725,s1n725,notn725;
or (n725,s0n725,s1n725);
not(notn725,n577);
and (s0n725,notn725,n726);
and (s1n725,n577,n727);
or (n727,n728,n730,n732,n734);
and (n728,n729,n603);
and (n730,n731,n608);
and (n732,n733,n612);
and (n734,n726,n614);
and (n735,n736,n39);
wire s0n736,s1n736,notn736;
or (n736,s0n736,s1n736);
not(notn736,n577);
and (s0n736,notn736,n737);
and (s1n736,n577,n738);
or (n738,n739,n741,n743,n745);
and (n739,n740,n603);
and (n741,n742,n608);
and (n743,n744,n612);
and (n745,n737,n614);
or (n746,n747,n869,n927);
and (n747,n748,n763);
xor (n748,n749,n761);
wire s0n749,s1n749,notn749;
or (n749,s0n749,s1n749);
not(notn749,n592);
and (s0n749,notn749,1'b0);
and (s1n749,n592,n750);
wire s0n750,s1n750,notn750;
or (n750,s0n750,s1n750);
not(notn750,n575);
and (s0n750,notn750,n751);
and (s1n750,n575,n753);
wire s0n751,s1n751,notn751;
or (n751,s0n751,s1n751);
not(notn751,n22);
and (s0n751,notn751,1'b0);
and (s1n751,n22,n752);
or (n753,1'b0,n754,n756,n758,n760);
and (n754,n755,n556);
and (n756,n757,n567);
and (n758,n759,n571);
and (n760,n752,n573);
wire s0n761,s1n761,notn761;
or (n761,s0n761,s1n761);
not(notn761,n762);
and (s0n761,notn761,1'b0);
and (s1n761,n762,n19);
xor (n762,n593,n649);
and (n763,n764,n766);
wire s0n764,s1n764,notn764;
or (n764,s0n764,s1n764);
not(notn764,n765);
and (s0n764,notn764,1'b0);
and (s1n764,n765,n19);
xor (n765,n650,n698);
or (n766,n767,n770,n868);
and (n767,n768,n769);
wire s0n768,s1n768,notn768;
or (n768,s0n768,s1n768);
not(notn768,n765);
and (s0n768,notn768,1'b0);
and (s1n768,n765,n750);
wire s0n769,s1n769,notn769;
or (n769,s0n769,s1n769);
not(notn769,n699);
and (s0n769,notn769,1'b0);
and (s1n769,n699,n19);
and (n770,n769,n771);
or (n771,n772,n786,n867);
and (n772,n773,n785);
wire s0n773,s1n773,notn773;
or (n773,s0n773,s1n773);
not(notn773,n765);
and (s0n773,notn773,1'b0);
and (s1n773,n765,n774);
wire s0n774,s1n774,notn774;
or (n774,s0n774,s1n774);
not(notn774,n575);
and (s0n774,notn774,n775);
and (s1n774,n575,n777);
wire s0n775,s1n775,notn775;
or (n775,s0n775,s1n775);
not(notn775,n22);
and (s0n775,notn775,1'b0);
and (s1n775,n22,n776);
or (n777,1'b0,n778,n780,n782,n784);
and (n778,n779,n556);
and (n780,n781,n567);
and (n782,n783,n571);
and (n784,n776,n573);
wire s0n785,s1n785,notn785;
or (n785,s0n785,s1n785);
not(notn785,n699);
and (s0n785,notn785,1'b0);
and (s1n785,n699,n750);
and (n786,n785,n787);
or (n787,n788,n802,n866);
and (n788,n789,n801);
wire s0n789,s1n789,notn789;
or (n789,s0n789,s1n789);
not(notn789,n765);
and (s0n789,notn789,1'b0);
and (s1n789,n765,n790);
wire s0n790,s1n790,notn790;
or (n790,s0n790,s1n790);
not(notn790,n575);
and (s0n790,notn790,n791);
and (s1n790,n575,n793);
wire s0n791,s1n791,notn791;
or (n791,s0n791,s1n791);
not(notn791,n22);
and (s0n791,notn791,1'b0);
and (s1n791,n22,n792);
or (n793,1'b0,n794,n796,n798,n800);
and (n794,n795,n556);
and (n796,n797,n567);
and (n798,n799,n571);
and (n800,n792,n573);
wire s0n801,s1n801,notn801;
or (n801,s0n801,s1n801);
not(notn801,n699);
and (s0n801,notn801,1'b0);
and (s1n801,n699,n774);
and (n802,n801,n803);
or (n803,n804,n818,n865);
and (n804,n805,n817);
wire s0n805,s1n805,notn805;
or (n805,s0n805,s1n805);
not(notn805,n765);
and (s0n805,notn805,1'b0);
and (s1n805,n765,n806);
wire s0n806,s1n806,notn806;
or (n806,s0n806,s1n806);
not(notn806,n575);
and (s0n806,notn806,n807);
and (s1n806,n575,n809);
wire s0n807,s1n807,notn807;
or (n807,s0n807,s1n807);
not(notn807,n22);
and (s0n807,notn807,1'b0);
and (s1n807,n22,n808);
or (n809,1'b0,n810,n812,n814,n816);
and (n810,n811,n556);
and (n812,n813,n567);
and (n814,n815,n571);
and (n816,n808,n573);
wire s0n817,s1n817,notn817;
or (n817,s0n817,s1n817);
not(notn817,n699);
and (s0n817,notn817,1'b0);
and (s1n817,n699,n790);
and (n818,n817,n819);
or (n819,n820,n834,n836);
and (n820,n821,n833);
wire s0n821,s1n821,notn821;
or (n821,s0n821,s1n821);
not(notn821,n765);
and (s0n821,notn821,1'b0);
and (s1n821,n765,n822);
wire s0n822,s1n822,notn822;
or (n822,s0n822,s1n822);
not(notn822,n575);
and (s0n822,notn822,n823);
and (s1n822,n575,n825);
wire s0n823,s1n823,notn823;
or (n823,s0n823,s1n823);
not(notn823,n22);
and (s0n823,notn823,1'b0);
and (s1n823,n22,n824);
or (n825,1'b0,n826,n828,n830,n832);
and (n826,n827,n556);
and (n828,n829,n567);
and (n830,n831,n571);
and (n832,n824,n573);
wire s0n833,s1n833,notn833;
or (n833,s0n833,s1n833);
not(notn833,n699);
and (s0n833,notn833,1'b0);
and (s1n833,n699,n806);
and (n834,n833,n835);
or (n835,n836,n850,n851);
and (n836,n837,n849);
wire s0n837,s1n837,notn837;
or (n837,s0n837,s1n837);
not(notn837,n765);
and (s0n837,notn837,1'b0);
and (s1n837,n765,n838);
wire s0n838,s1n838,notn838;
or (n838,s0n838,s1n838);
not(notn838,n575);
and (s0n838,notn838,n839);
and (s1n838,n575,n841);
wire s0n839,s1n839,notn839;
or (n839,s0n839,s1n839);
not(notn839,n22);
and (s0n839,notn839,1'b0);
and (s1n839,n22,n840);
or (n841,1'b0,n842,n844,n846,n848);
and (n842,n843,n556);
and (n844,n845,n567);
and (n846,n847,n571);
and (n848,n840,n573);
wire s0n849,s1n849,notn849;
or (n849,s0n849,s1n849);
not(notn849,n699);
and (s0n849,notn849,1'b0);
and (s1n849,n699,n822);
and (n850,n849,n851);
and (n851,n852,n864);
wire s0n852,s1n852,notn852;
or (n852,s0n852,s1n852);
not(notn852,n765);
and (s0n852,notn852,1'b0);
and (s1n852,n765,n853);
wire s0n853,s1n853,notn853;
or (n853,s0n853,s1n853);
not(notn853,n575);
and (s0n853,notn853,n854);
and (s1n853,n575,n856);
wire s0n854,s1n854,notn854;
or (n854,s0n854,s1n854);
not(notn854,n22);
and (s0n854,notn854,1'b0);
and (s1n854,n22,n855);
or (n856,1'b0,n857,n859,n861,n863);
and (n857,n858,n556);
and (n859,n860,n567);
and (n861,n862,n571);
and (n863,n855,n573);
wire s0n864,s1n864,notn864;
or (n864,s0n864,s1n864);
not(notn864,n699);
and (s0n864,notn864,1'b0);
and (s1n864,n699,n838);
and (n865,n805,n819);
and (n866,n789,n803);
and (n867,n773,n787);
and (n868,n768,n771);
and (n869,n763,n870);
or (n870,n871,n876,n926);
and (n871,n872,n875);
xor (n872,n873,n874);
wire s0n873,s1n873,notn873;
or (n873,s0n873,s1n873);
not(notn873,n592);
and (s0n873,notn873,1'b0);
and (s1n873,n592,n774);
wire s0n874,s1n874,notn874;
or (n874,s0n874,s1n874);
not(notn874,n762);
and (s0n874,notn874,1'b0);
and (s1n874,n762,n750);
xor (n875,n764,n766);
and (n876,n875,n877);
or (n877,n878,n884,n925);
and (n878,n879,n882);
xor (n879,n880,n881);
wire s0n880,s1n880,notn880;
or (n880,s0n880,s1n880);
not(notn880,n592);
and (s0n880,notn880,1'b0);
and (s1n880,n592,n790);
wire s0n881,s1n881,notn881;
or (n881,s0n881,s1n881);
not(notn881,n762);
and (s0n881,notn881,1'b0);
and (s1n881,n762,n774);
xor (n882,n883,n771);
xor (n883,n768,n769);
and (n884,n882,n885);
or (n885,n886,n892,n924);
and (n886,n887,n890);
xor (n887,n888,n889);
wire s0n888,s1n888,notn888;
or (n888,s0n888,s1n888);
not(notn888,n592);
and (s0n888,notn888,1'b0);
and (s1n888,n592,n806);
wire s0n889,s1n889,notn889;
or (n889,s0n889,s1n889);
not(notn889,n762);
and (s0n889,notn889,1'b0);
and (s1n889,n762,n790);
xor (n890,n891,n787);
xor (n891,n773,n785);
and (n892,n890,n893);
or (n893,n894,n900,n923);
and (n894,n895,n898);
xor (n895,n896,n897);
wire s0n896,s1n896,notn896;
or (n896,s0n896,s1n896);
not(notn896,n592);
and (s0n896,notn896,1'b0);
and (s1n896,n592,n822);
wire s0n897,s1n897,notn897;
or (n897,s0n897,s1n897);
not(notn897,n762);
and (s0n897,notn897,1'b0);
and (s1n897,n762,n806);
xor (n898,n899,n803);
xor (n899,n789,n801);
and (n900,n898,n901);
or (n901,n902,n908,n922);
and (n902,n903,n906);
xor (n903,n904,n905);
wire s0n904,s1n904,notn904;
or (n904,s0n904,s1n904);
not(notn904,n592);
and (s0n904,notn904,1'b0);
and (s1n904,n592,n838);
wire s0n905,s1n905,notn905;
or (n905,s0n905,s1n905);
not(notn905,n762);
and (s0n905,notn905,1'b0);
and (s1n905,n762,n822);
xor (n906,n907,n819);
xor (n907,n805,n817);
and (n908,n906,n909);
or (n909,n910,n916,n921);
and (n910,n911,n914);
xor (n911,n912,n913);
wire s0n912,s1n912,notn912;
or (n912,s0n912,s1n912);
not(notn912,n592);
and (s0n912,notn912,1'b0);
and (s1n912,n592,n853);
wire s0n913,s1n913,notn913;
or (n913,s0n913,s1n913);
not(notn913,n762);
and (s0n913,notn913,1'b0);
and (s1n913,n762,n838);
xor (n914,n915,n835);
xor (n915,n821,n833);
and (n916,n914,n917);
and (n917,n918,n919);
wire s0n918,s1n918,notn918;
or (n918,s0n918,s1n918);
not(notn918,n762);
and (s0n918,notn918,1'b0);
and (s1n918,n762,n853);
xor (n919,n920,n851);
xor (n920,n837,n849);
and (n921,n911,n917);
and (n922,n903,n909);
and (n923,n895,n901);
and (n924,n887,n893);
and (n925,n879,n885);
and (n926,n872,n877);
and (n927,n748,n870);
and (n928,n929,n977);
not (n929,n930);
wire s0n930,s1n930,notn930;
or (n930,s0n930,s1n930);
not(notn930,n40);
and (s0n930,notn930,1'b0);
and (s1n930,n40,n931);
wire s0n931,s1n931,notn931;
or (n931,s0n931,s1n931);
not(notn931,n648);
and (s0n931,notn931,n932);
and (s1n931,n648,n968);
or (n932,n933,n944,n955,n966);
and (n933,n934,n27);
wire s0n934,s1n934,notn934;
or (n934,s0n934,s1n934);
not(notn934,n577);
and (s0n934,notn934,n935);
and (s1n934,n577,n936);
or (n936,n937,n939,n941,n943);
and (n937,n938,n603);
and (n939,n940,n608);
and (n941,n942,n612);
and (n943,n935,n614);
and (n944,n945,n32);
wire s0n945,s1n945,notn945;
or (n945,s0n945,s1n945);
not(notn945,n577);
and (s0n945,notn945,n946);
and (s1n945,n577,n947);
or (n947,n948,n950,n952,n954);
and (n948,n949,n603);
and (n950,n951,n608);
and (n952,n953,n612);
and (n954,n946,n614);
and (n955,n956,n36);
wire s0n956,s1n956,notn956;
or (n956,s0n956,s1n956);
not(notn956,n577);
and (s0n956,notn956,n957);
and (s1n956,n577,n958);
or (n958,n959,n961,n963,n965);
and (n959,n960,n603);
and (n961,n962,n608);
and (n963,n964,n612);
and (n965,n957,n614);
and (n966,n967,n39);
wire s0n967,s1n967,notn967;
or (n967,s0n967,s1n967);
not(notn967,n577);
and (s0n967,notn967,n968);
and (s1n967,n577,n969);
or (n969,n970,n972,n974,n976);
and (n970,n971,n603);
and (n972,n973,n608);
and (n974,n975,n612);
and (n976,n968,n614);
and (n977,n978,n1026);
not (n978,n979);
wire s0n979,s1n979,notn979;
or (n979,s0n979,s1n979);
not(notn979,n40);
and (s0n979,notn979,1'b0);
and (s1n979,n40,n980);
wire s0n980,s1n980,notn980;
or (n980,s0n980,s1n980);
not(notn980,n648);
and (s0n980,notn980,n981);
and (s1n980,n648,n1017);
or (n981,n982,n993,n1004,n1015);
and (n982,n983,n27);
wire s0n983,s1n983,notn983;
or (n983,s0n983,s1n983);
not(notn983,n577);
and (s0n983,notn983,n984);
and (s1n983,n577,n985);
or (n985,n986,n988,n990,n992);
and (n986,n987,n603);
and (n988,n989,n608);
and (n990,n991,n612);
and (n992,n984,n614);
and (n993,n994,n32);
wire s0n994,s1n994,notn994;
or (n994,s0n994,s1n994);
not(notn994,n577);
and (s0n994,notn994,n995);
and (s1n994,n577,n996);
or (n996,n997,n999,n1001,n1003);
and (n997,n998,n603);
and (n999,n1000,n608);
and (n1001,n1002,n612);
and (n1003,n995,n614);
and (n1004,n1005,n36);
wire s0n1005,s1n1005,notn1005;
or (n1005,s0n1005,s1n1005);
not(notn1005,n577);
and (s0n1005,notn1005,n1006);
and (s1n1005,n577,n1007);
or (n1007,n1008,n1010,n1012,n1014);
and (n1008,n1009,n603);
and (n1010,n1011,n608);
and (n1012,n1013,n612);
and (n1014,n1006,n614);
and (n1015,n1016,n39);
wire s0n1016,s1n1016,notn1016;
or (n1016,s0n1016,s1n1016);
not(notn1016,n577);
and (s0n1016,notn1016,n1017);
and (s1n1016,n577,n1018);
or (n1018,n1019,n1021,n1023,n1025);
and (n1019,n1020,n603);
and (n1021,n1022,n608);
and (n1023,n1024,n612);
and (n1025,n1017,n614);
not (n1026,n1027);
wire s0n1027,s1n1027,notn1027;
or (n1027,s0n1027,s1n1027);
not(notn1027,n40);
and (s0n1027,notn1027,1'b0);
and (s1n1027,n40,n1028);
wire s0n1028,s1n1028,notn1028;
or (n1028,s0n1028,s1n1028);
not(notn1028,n648);
and (s0n1028,notn1028,n1029);
and (s1n1028,n648,n1065);
or (n1029,n1030,n1041,n1052,n1063);
and (n1030,n1031,n27);
wire s0n1031,s1n1031,notn1031;
or (n1031,s0n1031,s1n1031);
not(notn1031,n577);
and (s0n1031,notn1031,n1032);
and (s1n1031,n577,n1033);
or (n1033,n1034,n1036,n1038,n1040);
and (n1034,n1035,n603);
and (n1036,n1037,n608);
and (n1038,n1039,n612);
and (n1040,n1032,n614);
and (n1041,n1042,n32);
wire s0n1042,s1n1042,notn1042;
or (n1042,s0n1042,s1n1042);
not(notn1042,n577);
and (s0n1042,notn1042,n1043);
and (s1n1042,n577,n1044);
or (n1044,n1045,n1047,n1049,n1051);
and (n1045,n1046,n603);
and (n1047,n1048,n608);
and (n1049,n1050,n612);
and (n1051,n1043,n614);
and (n1052,n1053,n36);
wire s0n1053,s1n1053,notn1053;
or (n1053,s0n1053,s1n1053);
not(notn1053,n577);
and (s0n1053,notn1053,n1054);
and (s1n1053,n577,n1055);
or (n1055,n1056,n1058,n1060,n1062);
and (n1056,n1057,n603);
and (n1058,n1059,n608);
and (n1060,n1061,n612);
and (n1062,n1054,n614);
and (n1063,n1064,n39);
wire s0n1064,s1n1064,notn1064;
or (n1064,s0n1064,s1n1064);
not(notn1064,n577);
and (s0n1064,notn1064,n1065);
and (s1n1064,n577,n1066);
or (n1066,n1067,n1069,n1071,n1073);
and (n1067,n1068,n603);
and (n1069,n1070,n608);
and (n1071,n1072,n612);
and (n1073,n1065,n614);
or (n1074,n1075,n1155,n1240);
and (n1075,n1076,n1082);
xor (n1076,n1077,n1080);
wire s0n1077,s1n1077,notn1077;
or (n1077,s0n1077,s1n1077);
not(notn1077,n928);
and (s0n1077,notn1077,1'b0);
and (s1n1077,n928,n1078);
xor (n1078,n1079,n870);
xor (n1079,n748,n763);
wire s0n1080,s1n1080,notn1080;
or (n1080,s0n1080,s1n1080);
not(notn1080,n1081);
and (s0n1080,notn1080,1'b0);
and (s1n1080,n1081,n17);
xor (n1081,n929,n977);
and (n1082,n1083,n1085);
wire s0n1083,s1n1083,notn1083;
or (n1083,s0n1083,s1n1083);
not(notn1083,n1084);
and (s0n1083,notn1083,1'b0);
and (s1n1083,n1084,n17);
xor (n1084,n978,n1026);
or (n1085,n1086,n1089,n1154);
and (n1086,n1087,n1088);
wire s0n1087,s1n1087,notn1087;
or (n1087,s0n1087,s1n1087);
not(notn1087,n1084);
and (s0n1087,notn1087,1'b0);
and (s1n1087,n1084,n1078);
wire s0n1088,s1n1088,notn1088;
or (n1088,s0n1088,s1n1088);
not(notn1088,n1027);
and (s0n1088,notn1088,1'b0);
and (s1n1088,n1027,n17);
and (n1089,n1088,n1090);
or (n1090,n1091,n1096,n1153);
and (n1091,n1092,n1095);
wire s0n1092,s1n1092,notn1092;
or (n1092,s0n1092,s1n1092);
not(notn1092,n1084);
and (s0n1092,notn1092,1'b0);
and (s1n1092,n1084,n1093);
xor (n1093,n1094,n877);
xor (n1094,n872,n875);
wire s0n1095,s1n1095,notn1095;
or (n1095,s0n1095,s1n1095);
not(notn1095,n1027);
and (s0n1095,notn1095,1'b0);
and (s1n1095,n1027,n1078);
and (n1096,n1095,n1097);
or (n1097,n1098,n1103,n1152);
and (n1098,n1099,n1102);
wire s0n1099,s1n1099,notn1099;
or (n1099,s0n1099,s1n1099);
not(notn1099,n1084);
and (s0n1099,notn1099,1'b0);
and (s1n1099,n1084,n1100);
xor (n1100,n1101,n885);
xor (n1101,n879,n882);
wire s0n1102,s1n1102,notn1102;
or (n1102,s0n1102,s1n1102);
not(notn1102,n1027);
and (s0n1102,notn1102,1'b0);
and (s1n1102,n1027,n1093);
and (n1103,n1102,n1104);
or (n1104,n1105,n1110,n1151);
and (n1105,n1106,n1109);
wire s0n1106,s1n1106,notn1106;
or (n1106,s0n1106,s1n1106);
not(notn1106,n1084);
and (s0n1106,notn1106,1'b0);
and (s1n1106,n1084,n1107);
xor (n1107,n1108,n893);
xor (n1108,n887,n890);
wire s0n1109,s1n1109,notn1109;
or (n1109,s0n1109,s1n1109);
not(notn1109,n1027);
and (s0n1109,notn1109,1'b0);
and (s1n1109,n1027,n1100);
and (n1110,n1109,n1111);
or (n1111,n1112,n1117,n1150);
and (n1112,n1113,n1116);
wire s0n1113,s1n1113,notn1113;
or (n1113,s0n1113,s1n1113);
not(notn1113,n1084);
and (s0n1113,notn1113,1'b0);
and (s1n1113,n1084,n1114);
xor (n1114,n1115,n901);
xor (n1115,n895,n898);
wire s0n1116,s1n1116,notn1116;
or (n1116,s0n1116,s1n1116);
not(notn1116,n1027);
and (s0n1116,notn1116,1'b0);
and (s1n1116,n1027,n1107);
and (n1117,n1116,n1118);
or (n1118,n1119,n1124,n1149);
and (n1119,n1120,n1123);
wire s0n1120,s1n1120,notn1120;
or (n1120,s0n1120,s1n1120);
not(notn1120,n1084);
and (s0n1120,notn1120,1'b0);
and (s1n1120,n1084,n1121);
xor (n1121,n1122,n909);
xor (n1122,n903,n906);
wire s0n1123,s1n1123,notn1123;
or (n1123,s0n1123,s1n1123);
not(notn1123,n1027);
and (s0n1123,notn1123,1'b0);
and (s1n1123,n1027,n1114);
and (n1124,n1123,n1125);
or (n1125,n1126,n1131,n1148);
and (n1126,n1127,n1130);
wire s0n1127,s1n1127,notn1127;
or (n1127,s0n1127,s1n1127);
not(notn1127,n1084);
and (s0n1127,notn1127,1'b0);
and (s1n1127,n1084,n1128);
xor (n1128,n1129,n917);
xor (n1129,n911,n914);
wire s0n1130,s1n1130,notn1130;
or (n1130,s0n1130,s1n1130);
not(notn1130,n1027);
and (s0n1130,notn1130,1'b0);
and (s1n1130,n1027,n1121);
and (n1131,n1130,n1132);
or (n1132,n1133,n1137,n1139);
and (n1133,n1134,n1136);
wire s0n1134,s1n1134,notn1134;
or (n1134,s0n1134,s1n1134);
not(notn1134,n1084);
and (s0n1134,notn1134,1'b0);
and (s1n1134,n1084,n1135);
xor (n1135,n918,n919);
wire s0n1136,s1n1136,notn1136;
or (n1136,s0n1136,s1n1136);
not(notn1136,n1027);
and (s0n1136,notn1136,1'b0);
and (s1n1136,n1027,n1128);
and (n1137,n1136,n1138);
or (n1138,n1139,n1143,n1144);
and (n1139,n1140,n1142);
wire s0n1140,s1n1140,notn1140;
or (n1140,s0n1140,s1n1140);
not(notn1140,n1084);
and (s0n1140,notn1140,1'b0);
and (s1n1140,n1084,n1141);
xor (n1141,n852,n864);
wire s0n1142,s1n1142,notn1142;
or (n1142,s0n1142,s1n1142);
not(notn1142,n1027);
and (s0n1142,notn1142,1'b0);
and (s1n1142,n1027,n1135);
and (n1143,n1142,n1144);
and (n1144,n1145,n1147);
wire s0n1145,s1n1145,notn1145;
or (n1145,s0n1145,s1n1145);
not(notn1145,n1084);
and (s0n1145,notn1145,1'b0);
and (s1n1145,n1084,n1146);
wire s0n1146,s1n1146,notn1146;
or (n1146,s0n1146,s1n1146);
not(notn1146,n699);
and (s0n1146,notn1146,1'b0);
and (s1n1146,n699,n853);
wire s0n1147,s1n1147,notn1147;
or (n1147,s0n1147,s1n1147);
not(notn1147,n1027);
and (s0n1147,notn1147,1'b0);
and (s1n1147,n1027,n1141);
and (n1148,n1127,n1132);
and (n1149,n1120,n1125);
and (n1150,n1113,n1118);
and (n1151,n1106,n1111);
and (n1152,n1099,n1104);
and (n1153,n1092,n1097);
and (n1154,n1087,n1090);
and (n1155,n1082,n1156);
or (n1156,n1157,n1162,n1239);
and (n1157,n1158,n1161);
xor (n1158,n1159,n1160);
wire s0n1159,s1n1159,notn1159;
or (n1159,s0n1159,s1n1159);
not(notn1159,n928);
and (s0n1159,notn1159,1'b0);
and (s1n1159,n928,n1093);
wire s0n1160,s1n1160,notn1160;
or (n1160,s0n1160,s1n1160);
not(notn1160,n1081);
and (s0n1160,notn1160,1'b0);
and (s1n1160,n1081,n1078);
xor (n1161,n1083,n1085);
and (n1162,n1161,n1163);
or (n1163,n1164,n1170,n1238);
and (n1164,n1165,n1168);
xor (n1165,n1166,n1167);
wire s0n1166,s1n1166,notn1166;
or (n1166,s0n1166,s1n1166);
not(notn1166,n928);
and (s0n1166,notn1166,1'b0);
and (s1n1166,n928,n1100);
wire s0n1167,s1n1167,notn1167;
or (n1167,s0n1167,s1n1167);
not(notn1167,n1081);
and (s0n1167,notn1167,1'b0);
and (s1n1167,n1081,n1093);
xor (n1168,n1169,n1090);
xor (n1169,n1087,n1088);
and (n1170,n1168,n1171);
or (n1171,n1172,n1178,n1237);
and (n1172,n1173,n1176);
xor (n1173,n1174,n1175);
wire s0n1174,s1n1174,notn1174;
or (n1174,s0n1174,s1n1174);
not(notn1174,n928);
and (s0n1174,notn1174,1'b0);
and (s1n1174,n928,n1107);
wire s0n1175,s1n1175,notn1175;
or (n1175,s0n1175,s1n1175);
not(notn1175,n1081);
and (s0n1175,notn1175,1'b0);
and (s1n1175,n1081,n1100);
xor (n1176,n1177,n1097);
xor (n1177,n1092,n1095);
and (n1178,n1176,n1179);
or (n1179,n1180,n1186,n1236);
and (n1180,n1181,n1184);
xor (n1181,n1182,n1183);
wire s0n1182,s1n1182,notn1182;
or (n1182,s0n1182,s1n1182);
not(notn1182,n928);
and (s0n1182,notn1182,1'b0);
and (s1n1182,n928,n1114);
wire s0n1183,s1n1183,notn1183;
or (n1183,s0n1183,s1n1183);
not(notn1183,n1081);
and (s0n1183,notn1183,1'b0);
and (s1n1183,n1081,n1107);
xor (n1184,n1185,n1104);
xor (n1185,n1099,n1102);
and (n1186,n1184,n1187);
or (n1187,n1188,n1194,n1235);
and (n1188,n1189,n1192);
xor (n1189,n1190,n1191);
wire s0n1190,s1n1190,notn1190;
or (n1190,s0n1190,s1n1190);
not(notn1190,n928);
and (s0n1190,notn1190,1'b0);
and (s1n1190,n928,n1121);
wire s0n1191,s1n1191,notn1191;
or (n1191,s0n1191,s1n1191);
not(notn1191,n1081);
and (s0n1191,notn1191,1'b0);
and (s1n1191,n1081,n1114);
xor (n1192,n1193,n1111);
xor (n1193,n1106,n1109);
and (n1194,n1192,n1195);
or (n1195,n1196,n1202,n1234);
and (n1196,n1197,n1200);
xor (n1197,n1198,n1199);
wire s0n1198,s1n1198,notn1198;
or (n1198,s0n1198,s1n1198);
not(notn1198,n928);
and (s0n1198,notn1198,1'b0);
and (s1n1198,n928,n1128);
wire s0n1199,s1n1199,notn1199;
or (n1199,s0n1199,s1n1199);
not(notn1199,n1081);
and (s0n1199,notn1199,1'b0);
and (s1n1199,n1081,n1121);
xor (n1200,n1201,n1118);
xor (n1201,n1113,n1116);
and (n1202,n1200,n1203);
or (n1203,n1204,n1210,n1233);
and (n1204,n1205,n1208);
xor (n1205,n1206,n1207);
wire s0n1206,s1n1206,notn1206;
or (n1206,s0n1206,s1n1206);
not(notn1206,n928);
and (s0n1206,notn1206,1'b0);
and (s1n1206,n928,n1135);
wire s0n1207,s1n1207,notn1207;
or (n1207,s0n1207,s1n1207);
not(notn1207,n1081);
and (s0n1207,notn1207,1'b0);
and (s1n1207,n1081,n1128);
xor (n1208,n1209,n1125);
xor (n1209,n1120,n1123);
and (n1210,n1208,n1211);
or (n1211,n1212,n1218,n1232);
and (n1212,n1213,n1216);
xor (n1213,n1214,n1215);
wire s0n1214,s1n1214,notn1214;
or (n1214,s0n1214,s1n1214);
not(notn1214,n928);
and (s0n1214,notn1214,1'b0);
and (s1n1214,n928,n1141);
wire s0n1215,s1n1215,notn1215;
or (n1215,s0n1215,s1n1215);
not(notn1215,n1081);
and (s0n1215,notn1215,1'b0);
and (s1n1215,n1081,n1135);
xor (n1216,n1217,n1132);
xor (n1217,n1127,n1130);
and (n1218,n1216,n1219);
or (n1219,n1220,n1226,n1231);
and (n1220,n1221,n1224);
xor (n1221,n1222,n1223);
wire s0n1222,s1n1222,notn1222;
or (n1222,s0n1222,s1n1222);
not(notn1222,n928);
and (s0n1222,notn1222,1'b0);
and (s1n1222,n928,n1146);
wire s0n1223,s1n1223,notn1223;
or (n1223,s0n1223,s1n1223);
not(notn1223,n1081);
and (s0n1223,notn1223,1'b0);
and (s1n1223,n1081,n1141);
xor (n1224,n1225,n1138);
xor (n1225,n1134,n1136);
and (n1226,n1224,n1227);
and (n1227,n1228,n1229);
wire s0n1228,s1n1228,notn1228;
or (n1228,s0n1228,s1n1228);
not(notn1228,n1081);
and (s0n1228,notn1228,1'b0);
and (s1n1228,n1081,n1146);
xor (n1229,n1230,n1144);
xor (n1230,n1140,n1142);
and (n1231,n1221,n1227);
and (n1232,n1213,n1219);
and (n1233,n1205,n1211);
and (n1234,n1197,n1203);
and (n1235,n1189,n1195);
and (n1236,n1181,n1187);
and (n1237,n1173,n1179);
and (n1238,n1165,n1171);
and (n1239,n1158,n1163);
and (n1240,n1076,n1156);
xor (n1241,n1242,n1420);
wire s0n1242,s1n1242,notn1242;
or (n1242,s0n1242,s1n1242);
not(notn1242,n928);
and (s0n1242,notn1242,1'b0);
and (s1n1242,n928,n1243);
or (n1243,n1244,n1373,n1419);
and (n1244,n1245,n1257);
wire s0n1245,s1n1245,notn1245;
or (n1245,s0n1245,s1n1245);
not(notn1245,n594);
and (s0n1245,notn1245,1'b0);
and (s1n1245,n594,n1246);
wire s0n1246,s1n1246,notn1246;
or (n1246,s0n1246,s1n1246);
not(notn1246,n575);
and (s0n1246,notn1246,n1247);
and (s1n1246,n575,n1249);
wire s0n1247,s1n1247,notn1247;
or (n1247,s0n1247,s1n1247);
not(notn1247,n22);
and (s0n1247,notn1247,1'b0);
and (s1n1247,n22,n1248);
or (n1249,1'b0,n1250,n1252,n1254,n1256);
and (n1250,n1251,n556);
and (n1252,n1253,n567);
and (n1254,n1255,n571);
and (n1256,n1248,n573);
and (n1257,n1258,n1259);
wire s0n1258,s1n1258,notn1258;
or (n1258,s0n1258,s1n1258);
not(notn1258,n651);
and (s0n1258,notn1258,1'b0);
and (s1n1258,n651,n1246);
or (n1259,n1260,n1274,n1372);
and (n1260,n1261,n1273);
wire s0n1261,s1n1261,notn1261;
or (n1261,s0n1261,s1n1261);
not(notn1261,n651);
and (s0n1261,notn1261,1'b0);
and (s1n1261,n651,n1262);
wire s0n1262,s1n1262,notn1262;
or (n1262,s0n1262,s1n1262);
not(notn1262,n575);
and (s0n1262,notn1262,n1263);
and (s1n1262,n575,n1265);
wire s0n1263,s1n1263,notn1263;
or (n1263,s0n1263,s1n1263);
not(notn1263,n22);
and (s0n1263,notn1263,1'b0);
and (s1n1263,n22,n1264);
or (n1265,1'b0,n1266,n1268,n1270,n1272);
and (n1266,n1267,n556);
and (n1268,n1269,n567);
and (n1270,n1271,n571);
and (n1272,n1264,n573);
wire s0n1273,s1n1273,notn1273;
or (n1273,s0n1273,s1n1273);
not(notn1273,n699);
and (s0n1273,notn1273,1'b0);
and (s1n1273,n699,n1246);
and (n1274,n1273,n1275);
or (n1275,n1276,n1290,n1371);
and (n1276,n1277,n1289);
wire s0n1277,s1n1277,notn1277;
or (n1277,s0n1277,s1n1277);
not(notn1277,n651);
and (s0n1277,notn1277,1'b0);
and (s1n1277,n651,n1278);
wire s0n1278,s1n1278,notn1278;
or (n1278,s0n1278,s1n1278);
not(notn1278,n575);
and (s0n1278,notn1278,n1279);
and (s1n1278,n575,n1281);
wire s0n1279,s1n1279,notn1279;
or (n1279,s0n1279,s1n1279);
not(notn1279,n22);
and (s0n1279,notn1279,1'b0);
and (s1n1279,n22,n1280);
or (n1281,1'b0,n1282,n1284,n1286,n1288);
and (n1282,n1283,n556);
and (n1284,n1285,n567);
and (n1286,n1287,n571);
and (n1288,n1280,n573);
wire s0n1289,s1n1289,notn1289;
or (n1289,s0n1289,s1n1289);
not(notn1289,n699);
and (s0n1289,notn1289,1'b0);
and (s1n1289,n699,n1262);
and (n1290,n1289,n1291);
or (n1291,n1292,n1306,n1370);
and (n1292,n1293,n1305);
wire s0n1293,s1n1293,notn1293;
or (n1293,s0n1293,s1n1293);
not(notn1293,n651);
and (s0n1293,notn1293,1'b0);
and (s1n1293,n651,n1294);
wire s0n1294,s1n1294,notn1294;
or (n1294,s0n1294,s1n1294);
not(notn1294,n575);
and (s0n1294,notn1294,n1295);
and (s1n1294,n575,n1297);
wire s0n1295,s1n1295,notn1295;
or (n1295,s0n1295,s1n1295);
not(notn1295,n22);
and (s0n1295,notn1295,1'b0);
and (s1n1295,n22,n1296);
or (n1297,1'b0,n1298,n1300,n1302,n1304);
and (n1298,n1299,n556);
and (n1300,n1301,n567);
and (n1302,n1303,n571);
and (n1304,n1296,n573);
wire s0n1305,s1n1305,notn1305;
or (n1305,s0n1305,s1n1305);
not(notn1305,n699);
and (s0n1305,notn1305,1'b0);
and (s1n1305,n699,n1278);
and (n1306,n1305,n1307);
or (n1307,n1308,n1322,n1369);
and (n1308,n1309,n1321);
wire s0n1309,s1n1309,notn1309;
or (n1309,s0n1309,s1n1309);
not(notn1309,n651);
and (s0n1309,notn1309,1'b0);
and (s1n1309,n651,n1310);
wire s0n1310,s1n1310,notn1310;
or (n1310,s0n1310,s1n1310);
not(notn1310,n575);
and (s0n1310,notn1310,n1311);
and (s1n1310,n575,n1313);
wire s0n1311,s1n1311,notn1311;
or (n1311,s0n1311,s1n1311);
not(notn1311,n22);
and (s0n1311,notn1311,1'b0);
and (s1n1311,n22,n1312);
or (n1313,1'b0,n1314,n1316,n1318,n1320);
and (n1314,n1315,n556);
and (n1316,n1317,n567);
and (n1318,n1319,n571);
and (n1320,n1312,n573);
wire s0n1321,s1n1321,notn1321;
or (n1321,s0n1321,s1n1321);
not(notn1321,n699);
and (s0n1321,notn1321,1'b0);
and (s1n1321,n699,n1294);
and (n1322,n1321,n1323);
or (n1323,n1324,n1338,n1340);
and (n1324,n1325,n1337);
wire s0n1325,s1n1325,notn1325;
or (n1325,s0n1325,s1n1325);
not(notn1325,n651);
and (s0n1325,notn1325,1'b0);
and (s1n1325,n651,n1326);
wire s0n1326,s1n1326,notn1326;
or (n1326,s0n1326,s1n1326);
not(notn1326,n575);
and (s0n1326,notn1326,n1327);
and (s1n1326,n575,n1329);
wire s0n1327,s1n1327,notn1327;
or (n1327,s0n1327,s1n1327);
not(notn1327,n22);
and (s0n1327,notn1327,1'b0);
and (s1n1327,n22,n1328);
or (n1329,1'b0,n1330,n1332,n1334,n1336);
and (n1330,n1331,n556);
and (n1332,n1333,n567);
and (n1334,n1335,n571);
and (n1336,n1328,n573);
wire s0n1337,s1n1337,notn1337;
or (n1337,s0n1337,s1n1337);
not(notn1337,n699);
and (s0n1337,notn1337,1'b0);
and (s1n1337,n699,n1310);
and (n1338,n1337,n1339);
or (n1339,n1340,n1354,n1355);
and (n1340,n1341,n1353);
wire s0n1341,s1n1341,notn1341;
or (n1341,s0n1341,s1n1341);
not(notn1341,n651);
and (s0n1341,notn1341,1'b0);
and (s1n1341,n651,n1342);
wire s0n1342,s1n1342,notn1342;
or (n1342,s0n1342,s1n1342);
not(notn1342,n575);
and (s0n1342,notn1342,n1343);
and (s1n1342,n575,n1345);
wire s0n1343,s1n1343,notn1343;
or (n1343,s0n1343,s1n1343);
not(notn1343,n22);
and (s0n1343,notn1343,1'b0);
and (s1n1343,n22,n1344);
or (n1345,1'b0,n1346,n1348,n1350,n1352);
and (n1346,n1347,n556);
and (n1348,n1349,n567);
and (n1350,n1351,n571);
and (n1352,n1344,n573);
wire s0n1353,s1n1353,notn1353;
or (n1353,s0n1353,s1n1353);
not(notn1353,n699);
and (s0n1353,notn1353,1'b0);
and (s1n1353,n699,n1326);
and (n1354,n1353,n1355);
and (n1355,n1356,n1368);
wire s0n1356,s1n1356,notn1356;
or (n1356,s0n1356,s1n1356);
not(notn1356,n651);
and (s0n1356,notn1356,1'b0);
and (s1n1356,n651,n1357);
wire s0n1357,s1n1357,notn1357;
or (n1357,s0n1357,s1n1357);
not(notn1357,n575);
and (s0n1357,notn1357,n1358);
and (s1n1357,n575,n1360);
wire s0n1358,s1n1358,notn1358;
or (n1358,s0n1358,s1n1358);
not(notn1358,n22);
and (s0n1358,notn1358,1'b0);
and (s1n1358,n22,n1359);
or (n1360,1'b0,n1361,n1363,n1365,n1367);
and (n1361,n1362,n556);
and (n1363,n1364,n567);
and (n1365,n1366,n571);
and (n1367,n1359,n573);
wire s0n1368,s1n1368,notn1368;
or (n1368,s0n1368,s1n1368);
not(notn1368,n699);
and (s0n1368,notn1368,1'b0);
and (s1n1368,n699,n1342);
and (n1369,n1309,n1323);
and (n1370,n1293,n1307);
and (n1371,n1277,n1291);
and (n1372,n1261,n1275);
and (n1373,n1257,n1374);
or (n1374,n1375,n1378,n1418);
and (n1375,n1376,n1377);
wire s0n1376,s1n1376,notn1376;
or (n1376,s0n1376,s1n1376);
not(notn1376,n594);
and (s0n1376,notn1376,1'b0);
and (s1n1376,n594,n1262);
xor (n1377,n1258,n1259);
and (n1378,n1377,n1379);
or (n1379,n1380,n1384,n1417);
and (n1380,n1381,n1382);
wire s0n1381,s1n1381,notn1381;
or (n1381,s0n1381,s1n1381);
not(notn1381,n594);
and (s0n1381,notn1381,1'b0);
and (s1n1381,n594,n1278);
xor (n1382,n1383,n1275);
xor (n1383,n1261,n1273);
and (n1384,n1382,n1385);
or (n1385,n1386,n1390,n1416);
and (n1386,n1387,n1388);
wire s0n1387,s1n1387,notn1387;
or (n1387,s0n1387,s1n1387);
not(notn1387,n594);
and (s0n1387,notn1387,1'b0);
and (s1n1387,n594,n1294);
xor (n1388,n1389,n1291);
xor (n1389,n1277,n1289);
and (n1390,n1388,n1391);
or (n1391,n1392,n1396,n1415);
and (n1392,n1393,n1394);
wire s0n1393,s1n1393,notn1393;
or (n1393,s0n1393,s1n1393);
not(notn1393,n594);
and (s0n1393,notn1393,1'b0);
and (s1n1393,n594,n1310);
xor (n1394,n1395,n1307);
xor (n1395,n1293,n1305);
and (n1396,n1394,n1397);
or (n1397,n1398,n1402,n1414);
and (n1398,n1399,n1400);
wire s0n1399,s1n1399,notn1399;
or (n1399,s0n1399,s1n1399);
not(notn1399,n594);
and (s0n1399,notn1399,1'b0);
and (s1n1399,n594,n1326);
xor (n1400,n1401,n1323);
xor (n1401,n1309,n1321);
and (n1402,n1400,n1403);
or (n1403,n1404,n1408,n1413);
and (n1404,n1405,n1406);
wire s0n1405,s1n1405,notn1405;
or (n1405,s0n1405,s1n1405);
not(notn1405,n594);
and (s0n1405,notn1405,1'b0);
and (s1n1405,n594,n1342);
xor (n1406,n1407,n1339);
xor (n1407,n1325,n1337);
and (n1408,n1406,n1409);
and (n1409,n1410,n1411);
wire s0n1410,s1n1410,notn1410;
or (n1410,s0n1410,s1n1410);
not(notn1410,n594);
and (s0n1410,notn1410,1'b0);
and (s1n1410,n594,n1357);
xor (n1411,n1412,n1355);
xor (n1412,n1341,n1353);
and (n1413,n1405,n1409);
and (n1414,n1399,n1403);
and (n1415,n1393,n1397);
and (n1416,n1387,n1391);
and (n1417,n1381,n1385);
and (n1418,n1376,n1379);
and (n1419,n1245,n1374);
or (n1420,n1421,n1499,n1584);
and (n1421,n1422,n1427);
xor (n1422,n1423,n1426);
wire s0n1423,s1n1423,notn1423;
or (n1423,s0n1423,s1n1423);
not(notn1423,n928);
and (s0n1423,notn1423,1'b0);
and (s1n1423,n928,n1424);
xor (n1424,n1425,n1374);
xor (n1425,n1245,n1257);
wire s0n1426,s1n1426,notn1426;
or (n1426,s0n1426,s1n1426);
not(notn1426,n1081);
and (s0n1426,notn1426,1'b0);
and (s1n1426,n1081,n1243);
and (n1427,n1428,n1429);
wire s0n1428,s1n1428,notn1428;
or (n1428,s0n1428,s1n1428);
not(notn1428,n1084);
and (s0n1428,notn1428,1'b0);
and (s1n1428,n1084,n1243);
or (n1429,n1430,n1433,n1498);
and (n1430,n1431,n1432);
wire s0n1431,s1n1431,notn1431;
or (n1431,s0n1431,s1n1431);
not(notn1431,n1084);
and (s0n1431,notn1431,1'b0);
and (s1n1431,n1084,n1424);
wire s0n1432,s1n1432,notn1432;
or (n1432,s0n1432,s1n1432);
not(notn1432,n1027);
and (s0n1432,notn1432,1'b0);
and (s1n1432,n1027,n1243);
and (n1433,n1432,n1434);
or (n1434,n1435,n1440,n1497);
and (n1435,n1436,n1439);
wire s0n1436,s1n1436,notn1436;
or (n1436,s0n1436,s1n1436);
not(notn1436,n1084);
and (s0n1436,notn1436,1'b0);
and (s1n1436,n1084,n1437);
xor (n1437,n1438,n1379);
xor (n1438,n1376,n1377);
wire s0n1439,s1n1439,notn1439;
or (n1439,s0n1439,s1n1439);
not(notn1439,n1027);
and (s0n1439,notn1439,1'b0);
and (s1n1439,n1027,n1424);
and (n1440,n1439,n1441);
or (n1441,n1442,n1447,n1496);
and (n1442,n1443,n1446);
wire s0n1443,s1n1443,notn1443;
or (n1443,s0n1443,s1n1443);
not(notn1443,n1084);
and (s0n1443,notn1443,1'b0);
and (s1n1443,n1084,n1444);
xor (n1444,n1445,n1385);
xor (n1445,n1381,n1382);
wire s0n1446,s1n1446,notn1446;
or (n1446,s0n1446,s1n1446);
not(notn1446,n1027);
and (s0n1446,notn1446,1'b0);
and (s1n1446,n1027,n1437);
and (n1447,n1446,n1448);
or (n1448,n1449,n1454,n1495);
and (n1449,n1450,n1453);
wire s0n1450,s1n1450,notn1450;
or (n1450,s0n1450,s1n1450);
not(notn1450,n1084);
and (s0n1450,notn1450,1'b0);
and (s1n1450,n1084,n1451);
xor (n1451,n1452,n1391);
xor (n1452,n1387,n1388);
wire s0n1453,s1n1453,notn1453;
or (n1453,s0n1453,s1n1453);
not(notn1453,n1027);
and (s0n1453,notn1453,1'b0);
and (s1n1453,n1027,n1444);
and (n1454,n1453,n1455);
or (n1455,n1456,n1461,n1494);
and (n1456,n1457,n1460);
wire s0n1457,s1n1457,notn1457;
or (n1457,s0n1457,s1n1457);
not(notn1457,n1084);
and (s0n1457,notn1457,1'b0);
and (s1n1457,n1084,n1458);
xor (n1458,n1459,n1397);
xor (n1459,n1393,n1394);
wire s0n1460,s1n1460,notn1460;
or (n1460,s0n1460,s1n1460);
not(notn1460,n1027);
and (s0n1460,notn1460,1'b0);
and (s1n1460,n1027,n1451);
and (n1461,n1460,n1462);
or (n1462,n1463,n1468,n1493);
and (n1463,n1464,n1467);
wire s0n1464,s1n1464,notn1464;
or (n1464,s0n1464,s1n1464);
not(notn1464,n1084);
and (s0n1464,notn1464,1'b0);
and (s1n1464,n1084,n1465);
xor (n1465,n1466,n1403);
xor (n1466,n1399,n1400);
wire s0n1467,s1n1467,notn1467;
or (n1467,s0n1467,s1n1467);
not(notn1467,n1027);
and (s0n1467,notn1467,1'b0);
and (s1n1467,n1027,n1458);
and (n1468,n1467,n1469);
or (n1469,n1470,n1475,n1492);
and (n1470,n1471,n1474);
wire s0n1471,s1n1471,notn1471;
or (n1471,s0n1471,s1n1471);
not(notn1471,n1084);
and (s0n1471,notn1471,1'b0);
and (s1n1471,n1084,n1472);
xor (n1472,n1473,n1409);
xor (n1473,n1405,n1406);
wire s0n1474,s1n1474,notn1474;
or (n1474,s0n1474,s1n1474);
not(notn1474,n1027);
and (s0n1474,notn1474,1'b0);
and (s1n1474,n1027,n1465);
and (n1475,n1474,n1476);
or (n1476,n1477,n1481,n1483);
and (n1477,n1478,n1480);
wire s0n1478,s1n1478,notn1478;
or (n1478,s0n1478,s1n1478);
not(notn1478,n1084);
and (s0n1478,notn1478,1'b0);
and (s1n1478,n1084,n1479);
xor (n1479,n1410,n1411);
wire s0n1480,s1n1480,notn1480;
or (n1480,s0n1480,s1n1480);
not(notn1480,n1027);
and (s0n1480,notn1480,1'b0);
and (s1n1480,n1027,n1472);
and (n1481,n1480,n1482);
or (n1482,n1483,n1487,n1488);
and (n1483,n1484,n1486);
wire s0n1484,s1n1484,notn1484;
or (n1484,s0n1484,s1n1484);
not(notn1484,n1084);
and (s0n1484,notn1484,1'b0);
and (s1n1484,n1084,n1485);
xor (n1485,n1356,n1368);
wire s0n1486,s1n1486,notn1486;
or (n1486,s0n1486,s1n1486);
not(notn1486,n1027);
and (s0n1486,notn1486,1'b0);
and (s1n1486,n1027,n1479);
and (n1487,n1486,n1488);
and (n1488,n1489,n1491);
wire s0n1489,s1n1489,notn1489;
or (n1489,s0n1489,s1n1489);
not(notn1489,n1084);
and (s0n1489,notn1489,1'b0);
and (s1n1489,n1084,n1490);
wire s0n1490,s1n1490,notn1490;
or (n1490,s0n1490,s1n1490);
not(notn1490,n699);
and (s0n1490,notn1490,1'b0);
and (s1n1490,n699,n1357);
wire s0n1491,s1n1491,notn1491;
or (n1491,s0n1491,s1n1491);
not(notn1491,n1027);
and (s0n1491,notn1491,1'b0);
and (s1n1491,n1027,n1485);
and (n1492,n1471,n1476);
and (n1493,n1464,n1469);
and (n1494,n1457,n1462);
and (n1495,n1450,n1455);
and (n1496,n1443,n1448);
and (n1497,n1436,n1441);
and (n1498,n1431,n1434);
and (n1499,n1427,n1500);
or (n1500,n1501,n1506,n1583);
and (n1501,n1502,n1505);
xor (n1502,n1503,n1504);
wire s0n1503,s1n1503,notn1503;
or (n1503,s0n1503,s1n1503);
not(notn1503,n928);
and (s0n1503,notn1503,1'b0);
and (s1n1503,n928,n1437);
wire s0n1504,s1n1504,notn1504;
or (n1504,s0n1504,s1n1504);
not(notn1504,n1081);
and (s0n1504,notn1504,1'b0);
and (s1n1504,n1081,n1424);
xor (n1505,n1428,n1429);
and (n1506,n1505,n1507);
or (n1507,n1508,n1514,n1582);
and (n1508,n1509,n1512);
xor (n1509,n1510,n1511);
wire s0n1510,s1n1510,notn1510;
or (n1510,s0n1510,s1n1510);
not(notn1510,n928);
and (s0n1510,notn1510,1'b0);
and (s1n1510,n928,n1444);
wire s0n1511,s1n1511,notn1511;
or (n1511,s0n1511,s1n1511);
not(notn1511,n1081);
and (s0n1511,notn1511,1'b0);
and (s1n1511,n1081,n1437);
xor (n1512,n1513,n1434);
xor (n1513,n1431,n1432);
and (n1514,n1512,n1515);
or (n1515,n1516,n1522,n1581);
and (n1516,n1517,n1520);
xor (n1517,n1518,n1519);
wire s0n1518,s1n1518,notn1518;
or (n1518,s0n1518,s1n1518);
not(notn1518,n928);
and (s0n1518,notn1518,1'b0);
and (s1n1518,n928,n1451);
wire s0n1519,s1n1519,notn1519;
or (n1519,s0n1519,s1n1519);
not(notn1519,n1081);
and (s0n1519,notn1519,1'b0);
and (s1n1519,n1081,n1444);
xor (n1520,n1521,n1441);
xor (n1521,n1436,n1439);
and (n1522,n1520,n1523);
or (n1523,n1524,n1530,n1580);
and (n1524,n1525,n1528);
xor (n1525,n1526,n1527);
wire s0n1526,s1n1526,notn1526;
or (n1526,s0n1526,s1n1526);
not(notn1526,n928);
and (s0n1526,notn1526,1'b0);
and (s1n1526,n928,n1458);
wire s0n1527,s1n1527,notn1527;
or (n1527,s0n1527,s1n1527);
not(notn1527,n1081);
and (s0n1527,notn1527,1'b0);
and (s1n1527,n1081,n1451);
xor (n1528,n1529,n1448);
xor (n1529,n1443,n1446);
and (n1530,n1528,n1531);
or (n1531,n1532,n1538,n1579);
and (n1532,n1533,n1536);
xor (n1533,n1534,n1535);
wire s0n1534,s1n1534,notn1534;
or (n1534,s0n1534,s1n1534);
not(notn1534,n928);
and (s0n1534,notn1534,1'b0);
and (s1n1534,n928,n1465);
wire s0n1535,s1n1535,notn1535;
or (n1535,s0n1535,s1n1535);
not(notn1535,n1081);
and (s0n1535,notn1535,1'b0);
and (s1n1535,n1081,n1458);
xor (n1536,n1537,n1455);
xor (n1537,n1450,n1453);
and (n1538,n1536,n1539);
or (n1539,n1540,n1546,n1578);
and (n1540,n1541,n1544);
xor (n1541,n1542,n1543);
wire s0n1542,s1n1542,notn1542;
or (n1542,s0n1542,s1n1542);
not(notn1542,n928);
and (s0n1542,notn1542,1'b0);
and (s1n1542,n928,n1472);
wire s0n1543,s1n1543,notn1543;
or (n1543,s0n1543,s1n1543);
not(notn1543,n1081);
and (s0n1543,notn1543,1'b0);
and (s1n1543,n1081,n1465);
xor (n1544,n1545,n1462);
xor (n1545,n1457,n1460);
and (n1546,n1544,n1547);
or (n1547,n1548,n1554,n1577);
and (n1548,n1549,n1552);
xor (n1549,n1550,n1551);
wire s0n1550,s1n1550,notn1550;
or (n1550,s0n1550,s1n1550);
not(notn1550,n928);
and (s0n1550,notn1550,1'b0);
and (s1n1550,n928,n1479);
wire s0n1551,s1n1551,notn1551;
or (n1551,s0n1551,s1n1551);
not(notn1551,n1081);
and (s0n1551,notn1551,1'b0);
and (s1n1551,n1081,n1472);
xor (n1552,n1553,n1469);
xor (n1553,n1464,n1467);
and (n1554,n1552,n1555);
or (n1555,n1556,n1562,n1576);
and (n1556,n1557,n1560);
xor (n1557,n1558,n1559);
wire s0n1558,s1n1558,notn1558;
or (n1558,s0n1558,s1n1558);
not(notn1558,n928);
and (s0n1558,notn1558,1'b0);
and (s1n1558,n928,n1485);
wire s0n1559,s1n1559,notn1559;
or (n1559,s0n1559,s1n1559);
not(notn1559,n1081);
and (s0n1559,notn1559,1'b0);
and (s1n1559,n1081,n1479);
xor (n1560,n1561,n1476);
xor (n1561,n1471,n1474);
and (n1562,n1560,n1563);
or (n1563,n1564,n1570,n1575);
and (n1564,n1565,n1568);
xor (n1565,n1566,n1567);
wire s0n1566,s1n1566,notn1566;
or (n1566,s0n1566,s1n1566);
not(notn1566,n928);
and (s0n1566,notn1566,1'b0);
and (s1n1566,n928,n1490);
wire s0n1567,s1n1567,notn1567;
or (n1567,s0n1567,s1n1567);
not(notn1567,n1081);
and (s0n1567,notn1567,1'b0);
and (s1n1567,n1081,n1485);
xor (n1568,n1569,n1482);
xor (n1569,n1478,n1480);
and (n1570,n1568,n1571);
and (n1571,n1572,n1573);
wire s0n1572,s1n1572,notn1572;
or (n1572,s0n1572,s1n1572);
not(notn1572,n1081);
and (s0n1572,notn1572,1'b0);
and (s1n1572,n1081,n1490);
xor (n1573,n1574,n1488);
xor (n1574,n1484,n1486);
and (n1575,n1565,n1571);
and (n1576,n1557,n1563);
and (n1577,n1549,n1555);
and (n1578,n1541,n1547);
and (n1579,n1533,n1539);
and (n1580,n1525,n1531);
and (n1581,n1517,n1523);
and (n1582,n1509,n1515);
and (n1583,n1502,n1507);
and (n1584,n1422,n1500);
or (n1585,n1586,n1591,n1679);
and (n1586,n1587,n1589);
xor (n1587,n1588,n1156);
xor (n1588,n1076,n1082);
xor (n1589,n1590,n1500);
xor (n1590,n1422,n1427);
and (n1591,n1589,n1592);
or (n1592,n1593,n1598,n1678);
and (n1593,n1594,n1596);
xor (n1594,n1595,n1163);
xor (n1595,n1158,n1161);
xor (n1596,n1597,n1507);
xor (n1597,n1502,n1505);
and (n1598,n1596,n1599);
or (n1599,n1600,n1605,n1677);
and (n1600,n1601,n1603);
xor (n1601,n1602,n1171);
xor (n1602,n1165,n1168);
xor (n1603,n1604,n1515);
xor (n1604,n1509,n1512);
and (n1605,n1603,n1606);
or (n1606,n1607,n1612,n1676);
and (n1607,n1608,n1610);
xor (n1608,n1609,n1179);
xor (n1609,n1173,n1176);
xor (n1610,n1611,n1523);
xor (n1611,n1517,n1520);
and (n1612,n1610,n1613);
or (n1613,n1614,n1619,n1675);
and (n1614,n1615,n1617);
xor (n1615,n1616,n1187);
xor (n1616,n1181,n1184);
xor (n1617,n1618,n1531);
xor (n1618,n1525,n1528);
and (n1619,n1617,n1620);
or (n1620,n1621,n1626,n1674);
and (n1621,n1622,n1624);
xor (n1622,n1623,n1195);
xor (n1623,n1189,n1192);
xor (n1624,n1625,n1539);
xor (n1625,n1533,n1536);
and (n1626,n1624,n1627);
or (n1627,n1628,n1633,n1673);
and (n1628,n1629,n1631);
xor (n1629,n1630,n1203);
xor (n1630,n1197,n1200);
xor (n1631,n1632,n1547);
xor (n1632,n1541,n1544);
and (n1633,n1631,n1634);
or (n1634,n1635,n1640,n1672);
and (n1635,n1636,n1638);
xor (n1636,n1637,n1211);
xor (n1637,n1205,n1208);
xor (n1638,n1639,n1555);
xor (n1639,n1549,n1552);
and (n1640,n1638,n1641);
or (n1641,n1642,n1647,n1671);
and (n1642,n1643,n1645);
xor (n1643,n1644,n1219);
xor (n1644,n1213,n1216);
xor (n1645,n1646,n1563);
xor (n1646,n1557,n1560);
and (n1647,n1645,n1648);
or (n1648,n1649,n1654,n1670);
and (n1649,n1650,n1652);
xor (n1650,n1651,n1227);
xor (n1651,n1221,n1224);
xor (n1652,n1653,n1571);
xor (n1653,n1565,n1568);
and (n1654,n1652,n1655);
or (n1655,n1656,n1659,n1669);
and (n1656,n1657,n1658);
xor (n1657,n1228,n1229);
xor (n1658,n1572,n1573);
and (n1659,n1658,n1660);
or (n1660,n1661,n1664,n1668);
and (n1661,n1662,n1663);
xor (n1662,n1145,n1147);
xor (n1663,n1489,n1491);
and (n1664,n1663,n1665);
and (n1665,n1666,n1667);
wire s0n1666,s1n1666,notn1666;
or (n1666,s0n1666,s1n1666);
not(notn1666,n1027);
and (s0n1666,notn1666,1'b0);
and (s1n1666,n1027,n1146);
wire s0n1667,s1n1667,notn1667;
or (n1667,s0n1667,s1n1667);
not(notn1667,n1027);
and (s0n1667,notn1667,1'b0);
and (s1n1667,n1027,n1490);
and (n1668,n1662,n1665);
and (n1669,n1657,n1660);
and (n1670,n1650,n1655);
and (n1671,n1643,n1648);
and (n1672,n1636,n1641);
and (n1673,n1629,n1634);
and (n1674,n1622,n1627);
and (n1675,n1615,n1620);
and (n1676,n1608,n1613);
and (n1677,n1601,n1606);
and (n1678,n1594,n1599);
and (n1679,n1587,n1592);
xor (n1680,n1681,n2483);
xor (n1681,n1682,n2076);
or (n1682,n1683,n2008,n2075);
and (n1683,n1684,n1885);
wire s0n1684,s1n1684,notn1684;
or (n1684,s0n1684,s1n1684);
not(notn1684,n930);
and (s0n1684,notn1684,1'b0);
and (s1n1684,n930,n1685);
xor (n1685,n1686,n1698);
wire s0n1686,s1n1686,notn1686;
or (n1686,s0n1686,s1n1686);
not(notn1686,n592);
and (s0n1686,notn1686,1'b0);
and (s1n1686,n592,n1687);
wire s0n1687,s1n1687,notn1687;
or (n1687,s0n1687,s1n1687);
not(notn1687,n575);
and (s0n1687,notn1687,n1688);
and (s1n1687,n575,n1690);
wire s0n1688,s1n1688,notn1688;
or (n1688,s0n1688,s1n1688);
not(notn1688,n22);
and (s0n1688,notn1688,1'b0);
and (s1n1688,n22,n1689);
or (n1690,1'b0,n1691,n1693,n1695,n1697);
and (n1691,n1692,n556);
and (n1693,n1694,n567);
and (n1695,n1696,n571);
and (n1697,n1689,n573);
or (n1698,n1699,n1736);
and (n1699,n1700,n1737);
xor (n1700,n1701,n1715);
xor (n1701,n1702,n1714);
wire s0n1702,s1n1702,notn1702;
or (n1702,s0n1702,s1n1702);
not(notn1702,n592);
and (s0n1702,notn1702,1'b0);
and (s1n1702,n592,n1703);
wire s0n1703,s1n1703,notn1703;
or (n1703,s0n1703,s1n1703);
not(notn1703,n575);
and (s0n1703,notn1703,n1704);
and (s1n1703,n575,n1706);
wire s0n1704,s1n1704,notn1704;
or (n1704,s0n1704,s1n1704);
not(notn1704,n22);
and (s0n1704,notn1704,1'b0);
and (s1n1704,n22,n1705);
or (n1706,1'b0,n1707,n1709,n1711,n1713);
and (n1707,n1708,n556);
and (n1709,n1710,n567);
and (n1711,n1712,n571);
and (n1713,n1705,n573);
wire s0n1714,s1n1714,notn1714;
or (n1714,s0n1714,s1n1714);
not(notn1714,n762);
and (s0n1714,notn1714,1'b0);
and (s1n1714,n762,n1687);
or (n1715,n1716,n1736);
and (n1716,n1717,n1733);
xor (n1717,n1718,n1719);
wire s0n1718,s1n1718,notn1718;
or (n1718,s0n1718,s1n1718);
not(notn1718,n762);
and (s0n1718,notn1718,1'b0);
and (s1n1718,n762,n1703);
xor (n1719,n1720,n1721);
wire s0n1720,s1n1720,notn1720;
or (n1720,s0n1720,s1n1720);
not(notn1720,n765);
and (s0n1720,notn1720,1'b0);
and (s1n1720,n765,n1687);
wire s0n1721,s1n1721,notn1721;
or (n1721,s0n1721,s1n1721);
not(notn1721,n592);
and (s0n1721,notn1721,1'b0);
and (s1n1721,n592,n1722);
wire s0n1722,s1n1722,notn1722;
or (n1722,s0n1722,s1n1722);
not(notn1722,n575);
and (s0n1722,notn1722,n1723);
and (s1n1722,n575,n1725);
wire s0n1723,s1n1723,notn1723;
or (n1723,s0n1723,s1n1723);
not(notn1723,n22);
and (s0n1723,notn1723,1'b0);
and (s1n1723,n22,n1724);
or (n1725,1'b0,n1726,n1728,n1730,n1732);
and (n1726,n1727,n556);
and (n1728,n1729,n567);
and (n1730,n1731,n571);
and (n1732,n1724,n573);
and (n1733,n1734,n1735);
wire s0n1734,s1n1734,notn1734;
or (n1734,s0n1734,s1n1734);
not(notn1734,n765);
and (s0n1734,notn1734,1'b0);
and (s1n1734,n765,n1703);
wire s0n1735,s1n1735,notn1735;
or (n1735,s0n1735,s1n1735);
not(notn1735,n699);
and (s0n1735,notn1735,1'b0);
and (s1n1735,n699,n1687);
and (n1736,n1718,n1719);
nand (n1737,n1738,n1884);
or (n1738,n1739,n1879);
nor (n1739,n1740,n1878);
and (n1740,n1741,n1867);
nand (n1741,n1742,n1866);
or (n1742,n1743,n1800);
not (n1743,n1744);
or (n1744,n1745,n1778);
xor (n1745,n1746,n1775);
xor (n1746,n1747,n1759);
wire s0n1747,s1n1747,notn1747;
or (n1747,s0n1747,s1n1747);
not(notn1747,n762);
and (s0n1747,notn1747,1'b0);
and (s1n1747,n762,n1748);
wire s0n1748,s1n1748,notn1748;
or (n1748,s0n1748,s1n1748);
not(notn1748,n575);
and (s0n1748,notn1748,n1749);
and (s1n1748,n575,n1751);
wire s0n1749,s1n1749,notn1749;
or (n1749,s0n1749,s1n1749);
not(notn1749,n22);
and (s0n1749,notn1749,1'b0);
and (s1n1749,n22,n1750);
or (n1751,1'b0,n1752,n1754,n1756,n1758);
and (n1752,n1753,n556);
and (n1754,n1755,n567);
and (n1756,n1757,n571);
and (n1758,n1750,n573);
xor (n1759,n1760,n1763);
xor (n1760,n1761,n1762);
wire s0n1761,s1n1761,notn1761;
or (n1761,s0n1761,s1n1761);
not(notn1761,n765);
and (s0n1761,notn1761,1'b0);
and (s1n1761,n765,n1722);
wire s0n1762,s1n1762,notn1762;
or (n1762,s0n1762,s1n1762);
not(notn1762,n699);
and (s0n1762,notn1762,1'b0);
and (s1n1762,n699,n1703);
wire s0n1763,s1n1763,notn1763;
or (n1763,s0n1763,s1n1763);
not(notn1763,n592);
and (s0n1763,notn1763,1'b0);
and (s1n1763,n592,n1764);
wire s0n1764,s1n1764,notn1764;
or (n1764,s0n1764,s1n1764);
not(notn1764,n575);
and (s0n1764,notn1764,n1765);
and (s1n1764,n575,n1767);
wire s0n1765,s1n1765,notn1765;
or (n1765,s0n1765,s1n1765);
not(notn1765,n22);
and (s0n1765,notn1765,1'b0);
and (s1n1765,n22,n1766);
or (n1767,1'b0,n1768,n1770,n1772,n1774);
and (n1768,n1769,n556);
and (n1770,n1771,n567);
and (n1772,n1773,n571);
and (n1774,n1766,n573);
and (n1775,n1776,n1777);
wire s0n1776,s1n1776,notn1776;
or (n1776,s0n1776,s1n1776);
not(notn1776,n765);
and (s0n1776,notn1776,1'b0);
and (s1n1776,n765,n1748);
wire s0n1777,s1n1777,notn1777;
or (n1777,s0n1777,s1n1777);
not(notn1777,n699);
and (s0n1777,notn1777,1'b0);
and (s1n1777,n699,n1722);
or (n1778,n1779,n1799);
and (n1779,n1780,n1796);
xor (n1780,n1781,n1782);
wire s0n1781,s1n1781,notn1781;
or (n1781,s0n1781,s1n1781);
not(notn1781,n762);
and (s0n1781,notn1781,1'b0);
and (s1n1781,n762,n1764);
xor (n1782,n1783,n1784);
xor (n1783,n1776,n1777);
wire s0n1784,s1n1784,notn1784;
or (n1784,s0n1784,s1n1784);
not(notn1784,n592);
and (s0n1784,notn1784,1'b0);
and (s1n1784,n592,n1785);
wire s0n1785,s1n1785,notn1785;
or (n1785,s0n1785,s1n1785);
not(notn1785,n575);
and (s0n1785,notn1785,n1786);
and (s1n1785,n575,n1788);
wire s0n1786,s1n1786,notn1786;
or (n1786,s0n1786,s1n1786);
not(notn1786,n22);
and (s0n1786,notn1786,1'b0);
and (s1n1786,n22,n1787);
or (n1788,1'b0,n1789,n1791,n1793,n1795);
and (n1789,n1790,n556);
and (n1791,n1792,n567);
and (n1793,n1794,n571);
and (n1795,n1787,n573);
and (n1796,n1797,n1798);
wire s0n1797,s1n1797,notn1797;
or (n1797,s0n1797,s1n1797);
not(notn1797,n765);
and (s0n1797,notn1797,1'b0);
and (s1n1797,n765,n1764);
wire s0n1798,s1n1798,notn1798;
or (n1798,s0n1798,s1n1798);
not(notn1798,n699);
and (s0n1798,notn1798,1'b0);
and (s1n1798,n699,n1748);
and (n1799,n1781,n1782);
not (n1800,n1801);
nand (n1801,n1802,n1862,n1865);
nand (n1802,n1803,n1827,n1859);
or (n1803,n1804,n1805);
xor (n1804,n1780,n1796);
or (n1805,n1806,n1826);
and (n1806,n1807,n1812);
xor (n1807,n1808,n1809);
wire s0n1808,s1n1808,notn1808;
or (n1808,s0n1808,s1n1808);
not(notn1808,n762);
and (s0n1808,notn1808,1'b0);
and (s1n1808,n762,n1785);
and (n1809,n1810,n1811);
wire s0n1810,s1n1810,notn1810;
or (n1810,s0n1810,s1n1810);
not(notn1810,n765);
and (s0n1810,notn1810,1'b0);
and (s1n1810,n765,n1785);
wire s0n1811,s1n1811,notn1811;
or (n1811,s0n1811,s1n1811);
not(notn1811,n699);
and (s0n1811,notn1811,1'b0);
and (s1n1811,n699,n1764);
xor (n1812,n1813,n1814);
xor (n1813,n1797,n1798);
wire s0n1814,s1n1814,notn1814;
or (n1814,s0n1814,s1n1814);
not(notn1814,n592);
and (s0n1814,notn1814,1'b0);
and (s1n1814,n592,n1815);
wire s0n1815,s1n1815,notn1815;
or (n1815,s0n1815,s1n1815);
not(notn1815,n575);
and (s0n1815,notn1815,n1816);
and (s1n1815,n575,n1818);
wire s0n1816,s1n1816,notn1816;
or (n1816,s0n1816,s1n1816);
not(notn1816,n22);
and (s0n1816,notn1816,1'b0);
and (s1n1816,n22,n1817);
or (n1818,1'b0,n1819,n1821,n1823,n1825);
and (n1819,n1820,n556);
and (n1821,n1822,n567);
and (n1823,n1824,n571);
and (n1825,n1817,n573);
and (n1826,n1808,n1809);
or (n1827,n1828,n1858);
and (n1828,n1829,n1853);
xor (n1829,n1830,n1833);
and (n1830,n1831,n1832);
wire s0n1831,s1n1831,notn1831;
or (n1831,s0n1831,s1n1831);
not(notn1831,n765);
and (s0n1831,notn1831,1'b0);
and (s1n1831,n765,n1815);
wire s0n1832,s1n1832,notn1832;
or (n1832,s0n1832,s1n1832);
not(notn1832,n699);
and (s0n1832,notn1832,1'b0);
and (s1n1832,n699,n1785);
or (n1833,n1834,n1852);
and (n1834,n1835,n1851);
xor (n1835,n1836,n1850);
and (n1836,n1837,n1849);
wire s0n1837,s1n1837,notn1837;
or (n1837,s0n1837,s1n1837);
not(notn1837,n765);
and (s0n1837,notn1837,1'b0);
and (s1n1837,n765,n1838);
wire s0n1838,s1n1838,notn1838;
or (n1838,s0n1838,s1n1838);
not(notn1838,n575);
and (s0n1838,notn1838,n1839);
and (s1n1838,n575,n1841);
wire s0n1839,s1n1839,notn1839;
or (n1839,s0n1839,s1n1839);
not(notn1839,n22);
and (s0n1839,notn1839,1'b0);
and (s1n1839,n22,n1840);
or (n1841,1'b0,n1842,n1844,n1846,n1848);
and (n1842,n1843,n556);
and (n1844,n1845,n567);
and (n1846,n1847,n571);
and (n1848,n1840,n573);
wire s0n1849,s1n1849,notn1849;
or (n1849,s0n1849,s1n1849);
not(notn1849,n699);
and (s0n1849,notn1849,1'b0);
and (s1n1849,n699,n1815);
wire s0n1850,s1n1850,notn1850;
or (n1850,s0n1850,s1n1850);
not(notn1850,n762);
and (s0n1850,notn1850,1'b0);
and (s1n1850,n762,n1838);
xor (n1851,n1831,n1832);
and (n1852,n1836,n1850);
xor (n1853,n1854,n1857);
xor (n1854,n1855,n1856);
wire s0n1855,s1n1855,notn1855;
or (n1855,s0n1855,s1n1855);
not(notn1855,n592);
and (s0n1855,notn1855,1'b0);
and (s1n1855,n592,n1838);
xor (n1856,n1810,n1811);
wire s0n1857,s1n1857,notn1857;
or (n1857,s0n1857,s1n1857);
not(notn1857,n762);
and (s0n1857,notn1857,1'b0);
and (s1n1857,n762,n1815);
and (n1858,n1830,n1833);
or (n1859,n1860,n1861);
xor (n1860,n1807,n1812);
and (n1861,n1854,n1857);
nand (n1862,n1863,n1803);
not (n1863,n1864);
nand (n1864,n1860,n1861);
nand (n1865,n1804,n1805);
nand (n1866,n1745,n1778);
or (n1867,n1868,n1875);
xor (n1868,n1869,n1874);
xor (n1869,n1870,n1871);
wire s0n1870,s1n1870,notn1870;
or (n1870,s0n1870,s1n1870);
not(notn1870,n762);
and (s0n1870,notn1870,1'b0);
and (s1n1870,n762,n1722);
xor (n1871,n1872,n1873);
xor (n1872,n1734,n1735);
wire s0n1873,s1n1873,notn1873;
or (n1873,s0n1873,s1n1873);
not(notn1873,n592);
and (s0n1873,notn1873,1'b0);
and (s1n1873,n592,n1748);
and (n1874,n1761,n1762);
or (n1875,n1876,n1877);
and (n1876,n1746,n1775);
and (n1877,n1747,n1759);
and (n1878,n1868,n1875);
nor (n1879,n1880,n1883);
or (n1880,n1881,n1882);
and (n1881,n1869,n1874);
and (n1882,n1870,n1871);
xor (n1883,n1717,n1733);
nand (n1884,n1880,n1883);
and (n1885,n1886,n1887);
wire s0n1886,s1n1886,notn1886;
or (n1886,s0n1886,s1n1886);
not(notn1886,n979);
and (s0n1886,notn1886,1'b0);
and (s1n1886,n979,n1685);
or (n1887,n1888,n1892,n2007);
and (n1888,n1889,n1891);
wire s0n1889,s1n1889,notn1889;
or (n1889,s0n1889,s1n1889);
not(notn1889,n979);
and (s0n1889,notn1889,1'b0);
and (s1n1889,n979,n1890);
xor (n1890,n1700,n1737);
wire s0n1891,s1n1891,notn1891;
or (n1891,s0n1891,s1n1891);
not(notn1891,n1027);
and (s0n1891,notn1891,1'b0);
and (s1n1891,n1027,n1685);
and (n1892,n1891,n1893);
or (n1893,n1894,n1949,n2006);
and (n1894,n1895,n1948);
wire s0n1895,s1n1895,notn1895;
or (n1895,s0n1895,s1n1895);
not(notn1895,n979);
and (s0n1895,notn1895,1'b0);
and (s1n1895,n979,n1896);
xor (n1896,n1897,n1916);
xor (n1897,n1898,n1899);
xor (n1898,n1721,n1718);
xor (n1899,n1720,n1900);
or (n1900,n1733,n1901,n1915);
and (n1901,n1735,n1902);
or (n1902,n1874,n1903,n1914);
and (n1903,n1762,n1904);
or (n1904,n1775,n1905,n1913);
and (n1905,n1777,n1906);
or (n1906,n1796,n1907,n1912);
and (n1907,n1798,n1908);
or (n1908,n1809,n1909,n1830);
and (n1909,n1811,n1910);
or (n1910,n1830,n1911,n1836);
and (n1911,n1832,n1836);
and (n1912,n1797,n1908);
and (n1913,n1776,n1906);
and (n1914,n1761,n1904);
and (n1915,n1734,n1902);
or (n1916,n1917,n1920,n1947);
and (n1917,n1918,n1919);
xor (n1918,n1873,n1870);
xor (n1919,n1872,n1902);
and (n1920,n1919,n1921);
or (n1921,n1922,n1925,n1946);
and (n1922,n1923,n1924);
xor (n1923,n1763,n1747);
xor (n1924,n1760,n1904);
and (n1925,n1924,n1926);
or (n1926,n1927,n1930,n1945);
and (n1927,n1928,n1929);
xor (n1928,n1784,n1781);
xor (n1929,n1783,n1906);
and (n1930,n1929,n1931);
or (n1931,n1932,n1935,n1944);
and (n1932,n1933,n1934);
xor (n1933,n1814,n1808);
xor (n1934,n1813,n1908);
and (n1935,n1934,n1936);
or (n1936,n1937,n1940,n1943);
and (n1937,n1938,n1939);
xor (n1938,n1855,n1857);
xor (n1939,n1856,n1910);
and (n1940,n1939,n1941);
and (n1941,n1850,n1942);
xor (n1942,n1851,n1836);
and (n1943,n1938,n1941);
and (n1944,n1933,n1936);
and (n1945,n1928,n1931);
and (n1946,n1923,n1926);
and (n1947,n1918,n1921);
and (n1948,n1890,n1027);
and (n1949,n1948,n1950);
or (n1950,n1951,n1957,n2005);
and (n1951,n1952,n1956);
wire s0n1952,s1n1952,notn1952;
or (n1952,s0n1952,s1n1952);
not(notn1952,n979);
and (s0n1952,notn1952,1'b0);
and (s1n1952,n979,n1953);
xor (n1953,n1954,n1741);
nor (n1954,n1955,n1878);
not (n1955,n1867);
wire s0n1956,s1n1956,notn1956;
or (n1956,s0n1956,s1n1956);
not(notn1956,n1027);
and (s0n1956,notn1956,1'b0);
and (s1n1956,n1027,n1896);
and (n1957,n1956,n1958);
or (n1958,n1959,n1964,n2004);
and (n1959,n1960,n1963);
wire s0n1960,s1n1960,notn1960;
or (n1960,s0n1960,s1n1960);
not(notn1960,n979);
and (s0n1960,notn1960,1'b0);
and (s1n1960,n979,n1961);
xnor (n1961,n1801,n1962);
nand (n1962,n1744,n1866);
and (n1963,n1953,n1027);
and (n1964,n1963,n1965);
or (n1965,n1966,n1971,n2003);
and (n1966,n1967,n1970);
wire s0n1967,s1n1967,notn1967;
or (n1967,s0n1967,s1n1967);
not(notn1967,n979);
and (s0n1967,notn1967,1'b0);
and (s1n1967,n979,n1968);
xor (n1968,n1969,n1931);
xor (n1969,n1928,n1929);
and (n1970,n1961,n1027);
and (n1971,n1970,n1972);
or (n1972,n1973,n1978,n2002);
and (n1973,n1974,n1977);
wire s0n1974,s1n1974,notn1974;
or (n1974,s0n1974,s1n1974);
not(notn1974,n979);
and (s0n1974,notn1974,1'b0);
and (s1n1974,n979,n1975);
xor (n1975,n1976,n1936);
xor (n1976,n1933,n1934);
wire s0n1977,s1n1977,notn1977;
or (n1977,s0n1977,s1n1977);
not(notn1977,n1027);
and (s0n1977,notn1977,1'b0);
and (s1n1977,n1027,n1968);
and (n1978,n1977,n1979);
or (n1979,n1980,n1984,n2001);
and (n1980,n1981,n1983);
wire s0n1981,s1n1981,notn1981;
or (n1981,s0n1981,s1n1981);
not(notn1981,n979);
and (s0n1981,notn1981,1'b0);
and (s1n1981,n979,n1982);
xor (n1982,n1829,n1853);
wire s0n1983,s1n1983,notn1983;
or (n1983,s0n1983,s1n1983);
not(notn1983,n1027);
and (s0n1983,notn1983,1'b0);
and (s1n1983,n1027,n1975);
and (n1984,n1983,n1985);
or (n1985,n1986,n1990,n1992);
and (n1986,n1987,n1989);
wire s0n1987,s1n1987,notn1987;
or (n1987,s0n1987,s1n1987);
not(notn1987,n979);
and (s0n1987,notn1987,1'b0);
and (s1n1987,n979,n1988);
xor (n1988,n1835,n1851);
and (n1989,n1982,n1027);
and (n1990,n1989,n1991);
or (n1991,n1992,n1996,n1997);
and (n1992,n1993,n1995);
wire s0n1993,s1n1993,notn1993;
or (n1993,s0n1993,s1n1993);
not(notn1993,n979);
and (s0n1993,notn1993,1'b0);
and (s1n1993,n979,n1994);
xor (n1994,n1837,n1849);
and (n1995,n1988,n1027);
and (n1996,n1995,n1997);
and (n1997,n1998,n2000);
wire s0n1998,s1n1998,notn1998;
or (n1998,s0n1998,s1n1998);
not(notn1998,n979);
and (s0n1998,notn1998,1'b0);
and (s1n1998,n979,n1999);
wire s0n1999,s1n1999,notn1999;
or (n1999,s0n1999,s1n1999);
not(notn1999,n699);
and (s0n1999,notn1999,1'b0);
and (s1n1999,n699,n1838);
wire s0n2000,s1n2000,notn2000;
or (n2000,s0n2000,s1n2000);
not(notn2000,n1027);
and (s0n2000,notn2000,1'b0);
and (s1n2000,n1027,n1994);
and (n2001,n1981,n1985);
and (n2002,n1974,n1979);
and (n2003,n1967,n1972);
and (n2004,n1960,n1965);
and (n2005,n1952,n1958);
and (n2006,n1895,n1950);
and (n2007,n1889,n1893);
and (n2008,n1885,n2009);
or (n2009,n2010,n2013,n2074);
and (n2010,n2011,n2012);
wire s0n2011,s1n2011,notn2011;
or (n2011,s0n2011,s1n2011);
not(notn2011,n930);
and (s0n2011,notn2011,1'b0);
and (s1n2011,n930,n1890);
xor (n2012,n1886,n1887);
and (n2013,n2012,n2014);
or (n2014,n2015,n2019,n2073);
and (n2015,n2016,n2017);
wire s0n2016,s1n2016,notn2016;
or (n2016,s0n2016,s1n2016);
not(notn2016,n930);
and (s0n2016,notn2016,1'b0);
and (s1n2016,n930,n1896);
xor (n2017,n2018,n1893);
xor (n2018,n1889,n1891);
and (n2019,n2017,n2020);
or (n2020,n2021,n2025,n2072);
and (n2021,n2022,n2023);
wire s0n2022,s1n2022,notn2022;
or (n2022,s0n2022,s1n2022);
not(notn2022,n930);
and (s0n2022,notn2022,1'b0);
and (s1n2022,n930,n1953);
xor (n2023,n2024,n1950);
xor (n2024,n1895,n1948);
and (n2025,n2023,n2026);
or (n2026,n2027,n2031,n2071);
and (n2027,n2028,n2029);
wire s0n2028,s1n2028,notn2028;
or (n2028,s0n2028,s1n2028);
not(notn2028,n930);
and (s0n2028,notn2028,1'b0);
and (s1n2028,n930,n1961);
xor (n2029,n2030,n1958);
xor (n2030,n1952,n1956);
and (n2031,n2029,n2032);
or (n2032,n2033,n2037,n2070);
and (n2033,n2034,n2035);
wire s0n2034,s1n2034,notn2034;
or (n2034,s0n2034,s1n2034);
not(notn2034,n930);
and (s0n2034,notn2034,1'b0);
and (s1n2034,n930,n1968);
xor (n2035,n2036,n1965);
xor (n2036,n1960,n1963);
and (n2037,n2035,n2038);
or (n2038,n2039,n2043,n2069);
and (n2039,n2040,n2041);
wire s0n2040,s1n2040,notn2040;
or (n2040,s0n2040,s1n2040);
not(notn2040,n930);
and (s0n2040,notn2040,1'b0);
and (s1n2040,n930,n1975);
xor (n2041,n2042,n1972);
xor (n2042,n1967,n1970);
and (n2043,n2041,n2044);
or (n2044,n2045,n2049,n2068);
and (n2045,n2046,n2047);
wire s0n2046,s1n2046,notn2046;
or (n2046,s0n2046,s1n2046);
not(notn2046,n930);
and (s0n2046,notn2046,1'b0);
and (s1n2046,n930,n1982);
xor (n2047,n2048,n1979);
xor (n2048,n1974,n1977);
and (n2049,n2047,n2050);
or (n2050,n2051,n2055,n2067);
and (n2051,n2052,n2053);
wire s0n2052,s1n2052,notn2052;
or (n2052,s0n2052,s1n2052);
not(notn2052,n930);
and (s0n2052,notn2052,1'b0);
and (s1n2052,n930,n1988);
xor (n2053,n2054,n1985);
xor (n2054,n1981,n1983);
and (n2055,n2053,n2056);
or (n2056,n2057,n2061,n2066);
and (n2057,n2058,n2059);
wire s0n2058,s1n2058,notn2058;
or (n2058,s0n2058,s1n2058);
not(notn2058,n930);
and (s0n2058,notn2058,1'b0);
and (s1n2058,n930,n1994);
xor (n2059,n2060,n1991);
xor (n2060,n1987,n1989);
and (n2061,n2059,n2062);
and (n2062,n2063,n2064);
wire s0n2063,s1n2063,notn2063;
or (n2063,s0n2063,s1n2063);
not(notn2063,n930);
and (s0n2063,notn2063,1'b0);
and (s1n2063,n930,n1999);
xor (n2064,n2065,n1997);
xor (n2065,n1993,n1995);
and (n2066,n2058,n2062);
and (n2067,n2052,n2056);
and (n2068,n2046,n2050);
and (n2069,n2040,n2044);
and (n2070,n2034,n2038);
and (n2071,n2028,n2032);
and (n2072,n2022,n2026);
and (n2073,n2016,n2020);
and (n2074,n2011,n2014);
and (n2075,n1684,n2009);
or (n2076,n2077,n2415,n2482);
and (n2077,n2078,n2264);
wire s0n2078,s1n2078,notn2078;
or (n2078,s0n2078,s1n2078);
not(notn2078,n930);
and (s0n2078,notn2078,1'b0);
and (s1n2078,n930,n2079);
or (n2079,n2080,n2210,n2263);
and (n2080,n2081,n2093);
and (n2081,n594,n2082);
wire s0n2082,s1n2082,notn2082;
or (n2082,s0n2082,s1n2082);
not(notn2082,n575);
and (s0n2082,notn2082,n2083);
and (s1n2082,n575,n2085);
wire s0n2083,s1n2083,notn2083;
or (n2083,s0n2083,s1n2083);
not(notn2083,n22);
and (s0n2083,notn2083,1'b0);
and (s1n2083,n22,n2084);
or (n2085,1'b0,n2086,n2088,n2090,n2092);
and (n2086,n2087,n556);
and (n2088,n2089,n567);
and (n2090,n2091,n571);
and (n2092,n2084,n573);
and (n2093,n2094,n2095);
wire s0n2094,s1n2094,notn2094;
or (n2094,s0n2094,s1n2094);
not(notn2094,n651);
and (s0n2094,notn2094,1'b0);
and (s1n2094,n651,n2082);
or (n2095,n2096,n2110,n2209);
and (n2096,n2097,n2109);
wire s0n2097,s1n2097,notn2097;
or (n2097,s0n2097,s1n2097);
not(notn2097,n651);
and (s0n2097,notn2097,1'b0);
and (s1n2097,n651,n2098);
wire s0n2098,s1n2098,notn2098;
or (n2098,s0n2098,s1n2098);
not(notn2098,n575);
and (s0n2098,notn2098,n2099);
and (s1n2098,n575,n2101);
wire s0n2099,s1n2099,notn2099;
or (n2099,s0n2099,s1n2099);
not(notn2099,n22);
and (s0n2099,notn2099,1'b0);
and (s1n2099,n22,n2100);
or (n2101,1'b0,n2102,n2104,n2106,n2108);
and (n2102,n2103,n556);
and (n2104,n2105,n567);
and (n2106,n2107,n571);
and (n2108,n2100,n573);
wire s0n2109,s1n2109,notn2109;
or (n2109,s0n2109,s1n2109);
not(notn2109,n699);
and (s0n2109,notn2109,1'b0);
and (s1n2109,n699,n2082);
and (n2110,n2109,n2111);
or (n2111,n2112,n2126,n2208);
and (n2112,n2113,n2125);
wire s0n2113,s1n2113,notn2113;
or (n2113,s0n2113,s1n2113);
not(notn2113,n651);
and (s0n2113,notn2113,1'b0);
and (s1n2113,n651,n2114);
wire s0n2114,s1n2114,notn2114;
or (n2114,s0n2114,s1n2114);
not(notn2114,n575);
and (s0n2114,notn2114,n2115);
and (s1n2114,n575,n2117);
wire s0n2115,s1n2115,notn2115;
or (n2115,s0n2115,s1n2115);
not(notn2115,n22);
and (s0n2115,notn2115,1'b0);
and (s1n2115,n22,n2116);
or (n2117,1'b0,n2118,n2120,n2122,n2124);
and (n2118,n2119,n556);
and (n2120,n2121,n567);
and (n2122,n2123,n571);
and (n2124,n2116,n573);
wire s0n2125,s1n2125,notn2125;
or (n2125,s0n2125,s1n2125);
not(notn2125,n699);
and (s0n2125,notn2125,1'b0);
and (s1n2125,n699,n2098);
and (n2126,n2125,n2127);
or (n2127,n2128,n2142,n2207);
and (n2128,n2129,n2141);
wire s0n2129,s1n2129,notn2129;
or (n2129,s0n2129,s1n2129);
not(notn2129,n651);
and (s0n2129,notn2129,1'b0);
and (s1n2129,n651,n2130);
wire s0n2130,s1n2130,notn2130;
or (n2130,s0n2130,s1n2130);
not(notn2130,n575);
and (s0n2130,notn2130,n2131);
and (s1n2130,n575,n2133);
wire s0n2131,s1n2131,notn2131;
or (n2131,s0n2131,s1n2131);
not(notn2131,n22);
and (s0n2131,notn2131,1'b0);
and (s1n2131,n22,n2132);
or (n2133,1'b0,n2134,n2136,n2138,n2140);
and (n2134,n2135,n556);
and (n2136,n2137,n567);
and (n2138,n2139,n571);
and (n2140,n2132,n573);
wire s0n2141,s1n2141,notn2141;
or (n2141,s0n2141,s1n2141);
not(notn2141,n699);
and (s0n2141,notn2141,1'b0);
and (s1n2141,n699,n2114);
and (n2142,n2141,n2143);
or (n2143,n2144,n2158,n2206);
and (n2144,n2145,n2157);
wire s0n2145,s1n2145,notn2145;
or (n2145,s0n2145,s1n2145);
not(notn2145,n651);
and (s0n2145,notn2145,1'b0);
and (s1n2145,n651,n2146);
wire s0n2146,s1n2146,notn2146;
or (n2146,s0n2146,s1n2146);
not(notn2146,n575);
and (s0n2146,notn2146,n2147);
and (s1n2146,n575,n2149);
wire s0n2147,s1n2147,notn2147;
or (n2147,s0n2147,s1n2147);
not(notn2147,n22);
and (s0n2147,notn2147,1'b0);
and (s1n2147,n22,n2148);
or (n2149,1'b0,n2150,n2152,n2154,n2156);
and (n2150,n2151,n556);
and (n2152,n2153,n567);
and (n2154,n2155,n571);
and (n2156,n2148,n573);
wire s0n2157,s1n2157,notn2157;
or (n2157,s0n2157,s1n2157);
not(notn2157,n699);
and (s0n2157,notn2157,1'b0);
and (s1n2157,n699,n2130);
and (n2158,n2157,n2159);
or (n2159,n2160,n2174,n2176);
and (n2160,n2161,n2173);
wire s0n2161,s1n2161,notn2161;
or (n2161,s0n2161,s1n2161);
not(notn2161,n651);
and (s0n2161,notn2161,1'b0);
and (s1n2161,n651,n2162);
wire s0n2162,s1n2162,notn2162;
or (n2162,s0n2162,s1n2162);
not(notn2162,n575);
and (s0n2162,notn2162,n2163);
and (s1n2162,n575,n2165);
wire s0n2163,s1n2163,notn2163;
or (n2163,s0n2163,s1n2163);
not(notn2163,n22);
and (s0n2163,notn2163,1'b0);
and (s1n2163,n22,n2164);
or (n2165,1'b0,n2166,n2168,n2170,n2172);
and (n2166,n2167,n556);
and (n2168,n2169,n567);
and (n2170,n2171,n571);
and (n2172,n2164,n573);
wire s0n2173,s1n2173,notn2173;
or (n2173,s0n2173,s1n2173);
not(notn2173,n699);
and (s0n2173,notn2173,1'b0);
and (s1n2173,n699,n2146);
and (n2174,n2173,n2175);
or (n2175,n2176,n2191,n2192);
and (n2176,n2177,n2190);
not (n2177,n2178);
nand (n2178,n651,n2179);
wire s0n2179,s1n2179,notn2179;
or (n2179,s0n2179,s1n2179);
not(notn2179,n575);
and (s0n2179,notn2179,n2180);
and (s1n2179,n575,n2182);
wire s0n2180,s1n2180,notn2180;
or (n2180,s0n2180,s1n2180);
not(notn2180,n22);
and (s0n2180,notn2180,1'b0);
and (s1n2180,n22,n2181);
or (n2182,1'b0,n2183,n2185,n2187,n2189);
and (n2183,n2184,n556);
and (n2185,n2186,n567);
and (n2187,n2188,n571);
and (n2189,n2181,n573);
wire s0n2190,s1n2190,notn2190;
or (n2190,s0n2190,s1n2190);
not(notn2190,n699);
and (s0n2190,notn2190,1'b0);
and (s1n2190,n699,n2162);
and (n2191,n2190,n2192);
and (n2192,n2193,n2205);
wire s0n2193,s1n2193,notn2193;
or (n2193,s0n2193,s1n2193);
not(notn2193,n651);
and (s0n2193,notn2193,1'b0);
and (s1n2193,n651,n2194);
wire s0n2194,s1n2194,notn2194;
or (n2194,s0n2194,s1n2194);
not(notn2194,n575);
and (s0n2194,notn2194,n2195);
and (s1n2194,n575,n2197);
wire s0n2195,s1n2195,notn2195;
or (n2195,s0n2195,s1n2195);
not(notn2195,n22);
and (s0n2195,notn2195,1'b0);
and (s1n2195,n22,n2196);
or (n2197,1'b0,n2198,n2200,n2202,n2204);
and (n2198,n2199,n556);
and (n2200,n2201,n567);
and (n2202,n2203,n571);
and (n2204,n2196,n573);
wire s0n2205,s1n2205,notn2205;
or (n2205,s0n2205,s1n2205);
not(notn2205,n699);
and (s0n2205,notn2205,1'b0);
and (s1n2205,n699,n2179);
and (n2206,n2145,n2159);
and (n2207,n2129,n2143);
and (n2208,n2113,n2127);
and (n2209,n2097,n2111);
and (n2210,n2093,n2211);
or (n2211,n2212,n2216,n2262);
and (n2212,n2213,n2215);
not (n2213,n2214);
nand (n2214,n594,n2098);
xor (n2215,n2094,n2095);
and (n2216,n2215,n2217);
or (n2217,n2218,n2223,n2261);
and (n2218,n2219,n2221);
not (n2219,n2220);
nand (n2220,n594,n2114);
xor (n2221,n2222,n2111);
xor (n2222,n2097,n2109);
and (n2223,n2221,n2224);
or (n2224,n2225,n2230,n2260);
and (n2225,n2226,n2228);
not (n2226,n2227);
nand (n2227,n594,n2130);
xor (n2228,n2229,n2127);
xor (n2229,n2113,n2125);
and (n2230,n2228,n2231);
or (n2231,n2232,n2237,n2259);
and (n2232,n2233,n2235);
not (n2233,n2234);
nand (n2234,n594,n2146);
xor (n2235,n2236,n2143);
xor (n2236,n2129,n2141);
and (n2237,n2235,n2238);
or (n2238,n2239,n2244,n2258);
and (n2239,n2240,n2242);
not (n2240,n2241);
nand (n2241,n594,n2162);
xor (n2242,n2243,n2159);
xor (n2243,n2145,n2157);
and (n2244,n2242,n2245);
or (n2245,n2246,n2251,n2257);
and (n2246,n2247,n2249);
not (n2247,n2248);
nand (n2248,n594,n2179);
xor (n2249,n2250,n2175);
xor (n2250,n2161,n2173);
and (n2251,n2249,n2252);
and (n2252,n2253,n2255);
not (n2253,n2254);
nand (n2254,n594,n2194);
xor (n2255,n2256,n2192);
xor (n2256,n2177,n2190);
and (n2257,n2247,n2252);
and (n2258,n2240,n2245);
and (n2259,n2233,n2238);
and (n2260,n2226,n2231);
and (n2261,n2219,n2224);
and (n2262,n2213,n2217);
and (n2263,n2081,n2211);
and (n2264,n2265,n2266);
wire s0n2265,s1n2265,notn2265;
or (n2265,s0n2265,s1n2265);
not(notn2265,n979);
and (s0n2265,notn2265,1'b0);
and (s1n2265,n979,n2079);
or (n2266,n2267,n2272,n2414);
and (n2267,n2268,n2271);
wire s0n2268,s1n2268,notn2268;
or (n2268,s0n2268,s1n2268);
not(notn2268,n979);
and (s0n2268,notn2268,1'b0);
and (s1n2268,n979,n2269);
xor (n2269,n2270,n2211);
xor (n2270,n2081,n2093);
wire s0n2271,s1n2271,notn2271;
or (n2271,s0n2271,s1n2271);
not(notn2271,n1027);
and (s0n2271,notn2271,1'b0);
and (s1n2271,n1027,n2079);
and (n2272,n2271,n2273);
or (n2273,n2274,n2360,n2413);
and (n2274,n2275,n2359);
wire s0n2275,s1n2275,notn2275;
or (n2275,s0n2275,s1n2275);
not(notn2275,n979);
and (s0n2275,notn2275,1'b0);
and (s1n2275,n979,n2276);
xor (n2276,n2277,n2290);
xor (n2277,n2278,n2286);
nand (n2278,n2279,n2283);
or (n2279,n2280,n2282);
and (n2280,n2281,n2220);
not (n2281,n2109);
not (n2282,n2097);
or (n2283,n2284,n2285);
not (n2284,n2141);
not (n2285,n2081);
not (n2286,n2287);
xnor (n2287,n2288,n2289);
not (n2288,n2213);
not (n2289,n2094);
or (n2290,n2291,n2358);
and (n2291,n2292,n2304);
xor (n2292,n2293,n2298);
nor (n2293,n2294,n2296);
and (n2294,n2295,n2097);
xor (n2295,n2281,n2220);
and (n2296,n2297,n2282);
not (n2297,n2295);
nand (n2298,n2299,n2301,n2303);
or (n2299,n2220,n2300);
not (n2300,n2129);
or (n2301,n2227,n2302);
not (n2302,n2125);
not (n2303,n2112);
nand (n2304,n2305,n2357);
or (n2305,n2306,n2318);
not (n2306,n2307);
nand (n2307,n2308,n2310);
xor (n2308,n2229,n2309);
not (n2309,n2226);
not (n2310,n2311);
nand (n2311,n2312,n2315,n2317);
or (n2312,n2313,n2314);
not (n2313,n2173);
not (n2314,n2219);
or (n2315,n2309,n2316);
not (n2316,n2145);
not (n2317,n2128);
not (n2318,n2319);
or (n2319,n2320,n2356);
and (n2320,n2321,n2331);
xor (n2321,n2322,n2328);
nand (n2322,n2323,n2325,n2327);
or (n2323,n2227,n2324);
not (n2324,n2190);
or (n2325,n2234,n2326);
not (n2326,n2161);
not (n2327,n2144);
nand (n2328,n2329,n2330);
or (n2329,n2234,n2236);
nand (n2330,n2236,n2234);
or (n2331,n2332,n2355);
and (n2332,n2333,n2342);
xor (n2333,n2334,n2340);
nand (n2334,n2335,n2337,n2339);
not (n2335,n2336);
and (n2336,n2240,n2177);
or (n2337,n2234,n2338);
not (n2338,n2205);
not (n2339,n2160);
xnor (n2340,n2341,n2243);
not (n2341,n2240);
or (n2342,n2343,n2354);
and (n2343,n2344,n2350);
xor (n2344,n2345,n2346);
nor (n2345,n2254,n2324);
xnor (n2346,n2347,n2326);
nand (n2347,n2348,n2349);
or (n2348,n2247,n2313);
nand (n2349,n2247,n2313);
nand (n2350,n2351,n2353);
or (n2351,n2352,n2178);
xnor (n2352,n2324,n2254);
not (n2353,n2192);
and (n2354,n2345,n2346);
and (n2355,n2334,n2340);
and (n2356,n2322,n2328);
or (n2357,n2308,n2310);
and (n2358,n2293,n2298);
wire s0n2359,s1n2359,notn2359;
or (n2359,s0n2359,s1n2359);
not(notn2359,n1027);
and (s0n2359,notn2359,1'b0);
and (s1n2359,n1027,n2269);
and (n2360,n2359,n2361);
or (n2361,n2362,n2366,n2412);
and (n2362,n2363,n2365);
wire s0n2363,s1n2363,notn2363;
or (n2363,s0n2363,s1n2363);
not(notn2363,n979);
and (s0n2363,notn2363,1'b0);
and (s1n2363,n979,n2364);
xor (n2364,n2292,n2304);
wire s0n2365,s1n2365,notn2365;
or (n2365,s0n2365,s1n2365);
not(notn2365,n1027);
and (s0n2365,notn2365,1'b0);
and (s1n2365,n1027,n2276);
and (n2366,n2365,n2367);
or (n2367,n2368,n2373,n2411);
and (n2368,n2369,n2372);
wire s0n2369,s1n2369,notn2369;
or (n2369,s0n2369,s1n2369);
not(notn2369,n979);
and (s0n2369,notn2369,1'b0);
and (s1n2369,n979,n2370);
xor (n2370,n2371,n2231);
xor (n2371,n2226,n2228);
wire s0n2372,s1n2372,notn2372;
or (n2372,s0n2372,s1n2372);
not(notn2372,n1027);
and (s0n2372,notn2372,1'b0);
and (s1n2372,n1027,n2364);
and (n2373,n2372,n2374);
or (n2374,n2375,n2379,n2410);
and (n2375,n2376,n2378);
wire s0n2376,s1n2376,notn2376;
or (n2376,s0n2376,s1n2376);
not(notn2376,n979);
and (s0n2376,notn2376,1'b0);
and (s1n2376,n979,n2377);
xor (n2377,n2321,n2331);
wire s0n2378,s1n2378,notn2378;
or (n2378,s0n2378,s1n2378);
not(notn2378,n1027);
and (s0n2378,notn2378,1'b0);
and (s1n2378,n1027,n2370);
and (n2379,n2378,n2380);
or (n2380,n2381,n2385,n2409);
and (n2381,n2382,n2384);
wire s0n2382,s1n2382,notn2382;
or (n2382,s0n2382,s1n2382);
not(notn2382,n979);
and (s0n2382,notn2382,1'b0);
and (s1n2382,n979,n2383);
xor (n2383,n2333,n2342);
wire s0n2384,s1n2384,notn2384;
or (n2384,s0n2384,s1n2384);
not(notn2384,n1027);
and (s0n2384,notn2384,1'b0);
and (s1n2384,n1027,n2377);
and (n2385,n2384,n2386);
or (n2386,n2387,n2391,n2408);
and (n2387,n2388,n2390);
wire s0n2388,s1n2388,notn2388;
or (n2388,s0n2388,s1n2388);
not(notn2388,n979);
and (s0n2388,notn2388,1'b0);
and (s1n2388,n979,n2389);
xor (n2389,n2344,n2350);
wire s0n2390,s1n2390,notn2390;
or (n2390,s0n2390,s1n2390);
not(notn2390,n1027);
and (s0n2390,notn2390,1'b0);
and (s1n2390,n1027,n2383);
and (n2391,n2390,n2392);
or (n2392,n2393,n2397,n2399);
and (n2393,n2394,n2396);
wire s0n2394,s1n2394,notn2394;
or (n2394,s0n2394,s1n2394);
not(notn2394,n979);
and (s0n2394,notn2394,1'b0);
and (s1n2394,n979,n2395);
xor (n2395,n2253,n2255);
wire s0n2396,s1n2396,notn2396;
or (n2396,s0n2396,s1n2396);
not(notn2396,n1027);
and (s0n2396,notn2396,1'b0);
and (s1n2396,n1027,n2389);
and (n2397,n2396,n2398);
or (n2398,n2399,n2403,n2404);
and (n2399,n2400,n2402);
wire s0n2400,s1n2400,notn2400;
or (n2400,s0n2400,s1n2400);
not(notn2400,n979);
and (s0n2400,notn2400,1'b0);
and (s1n2400,n979,n2401);
xor (n2401,n2193,n2205);
wire s0n2402,s1n2402,notn2402;
or (n2402,s0n2402,s1n2402);
not(notn2402,n1027);
and (s0n2402,notn2402,1'b0);
and (s1n2402,n1027,n2395);
and (n2403,n2402,n2404);
and (n2404,n2405,n2407);
wire s0n2405,s1n2405,notn2405;
or (n2405,s0n2405,s1n2405);
not(notn2405,n979);
and (s0n2405,notn2405,1'b0);
and (s1n2405,n979,n2406);
wire s0n2406,s1n2406,notn2406;
or (n2406,s0n2406,s1n2406);
not(notn2406,n699);
and (s0n2406,notn2406,1'b0);
and (s1n2406,n699,n2194);
wire s0n2407,s1n2407,notn2407;
or (n2407,s0n2407,s1n2407);
not(notn2407,n1027);
and (s0n2407,notn2407,1'b0);
and (s1n2407,n1027,n2401);
and (n2408,n2388,n2392);
and (n2409,n2382,n2386);
and (n2410,n2376,n2380);
and (n2411,n2369,n2374);
and (n2412,n2363,n2367);
and (n2413,n2275,n2361);
and (n2414,n2268,n2273);
and (n2415,n2264,n2416);
or (n2416,n2417,n2420,n2481);
and (n2417,n2418,n2419);
wire s0n2418,s1n2418,notn2418;
or (n2418,s0n2418,s1n2418);
not(notn2418,n930);
and (s0n2418,notn2418,1'b0);
and (s1n2418,n930,n2269);
xor (n2419,n2265,n2266);
and (n2420,n2419,n2421);
or (n2421,n2422,n2426,n2480);
and (n2422,n2423,n2424);
wire s0n2423,s1n2423,notn2423;
or (n2423,s0n2423,s1n2423);
not(notn2423,n930);
and (s0n2423,notn2423,1'b0);
and (s1n2423,n930,n2276);
xor (n2424,n2425,n2273);
xor (n2425,n2268,n2271);
and (n2426,n2424,n2427);
or (n2427,n2428,n2432,n2479);
and (n2428,n2429,n2430);
wire s0n2429,s1n2429,notn2429;
or (n2429,s0n2429,s1n2429);
not(notn2429,n930);
and (s0n2429,notn2429,1'b0);
and (s1n2429,n930,n2364);
xor (n2430,n2431,n2361);
xor (n2431,n2275,n2359);
and (n2432,n2430,n2433);
or (n2433,n2434,n2438,n2478);
and (n2434,n2435,n2436);
wire s0n2435,s1n2435,notn2435;
or (n2435,s0n2435,s1n2435);
not(notn2435,n930);
and (s0n2435,notn2435,1'b0);
and (s1n2435,n930,n2370);
xor (n2436,n2437,n2367);
xor (n2437,n2363,n2365);
and (n2438,n2436,n2439);
or (n2439,n2440,n2444,n2477);
and (n2440,n2441,n2442);
wire s0n2441,s1n2441,notn2441;
or (n2441,s0n2441,s1n2441);
not(notn2441,n930);
and (s0n2441,notn2441,1'b0);
and (s1n2441,n930,n2377);
xor (n2442,n2443,n2374);
xor (n2443,n2369,n2372);
and (n2444,n2442,n2445);
or (n2445,n2446,n2450,n2476);
and (n2446,n2447,n2448);
wire s0n2447,s1n2447,notn2447;
or (n2447,s0n2447,s1n2447);
not(notn2447,n930);
and (s0n2447,notn2447,1'b0);
and (s1n2447,n930,n2383);
xor (n2448,n2449,n2380);
xor (n2449,n2376,n2378);
and (n2450,n2448,n2451);
or (n2451,n2452,n2456,n2475);
and (n2452,n2453,n2454);
wire s0n2453,s1n2453,notn2453;
or (n2453,s0n2453,s1n2453);
not(notn2453,n930);
and (s0n2453,notn2453,1'b0);
and (s1n2453,n930,n2389);
xor (n2454,n2455,n2386);
xor (n2455,n2382,n2384);
and (n2456,n2454,n2457);
or (n2457,n2458,n2462,n2474);
and (n2458,n2459,n2460);
wire s0n2459,s1n2459,notn2459;
or (n2459,s0n2459,s1n2459);
not(notn2459,n930);
and (s0n2459,notn2459,1'b0);
and (s1n2459,n930,n2395);
xor (n2460,n2461,n2392);
xor (n2461,n2388,n2390);
and (n2462,n2460,n2463);
or (n2463,n2464,n2468,n2473);
and (n2464,n2465,n2466);
wire s0n2465,s1n2465,notn2465;
or (n2465,s0n2465,s1n2465);
not(notn2465,n930);
and (s0n2465,notn2465,1'b0);
and (s1n2465,n930,n2401);
xor (n2466,n2467,n2398);
xor (n2467,n2394,n2396);
and (n2468,n2466,n2469);
and (n2469,n2470,n2471);
wire s0n2470,s1n2470,notn2470;
or (n2470,s0n2470,s1n2470);
not(notn2470,n930);
and (s0n2470,notn2470,1'b0);
and (s1n2470,n930,n2406);
xor (n2471,n2472,n2404);
xor (n2472,n2400,n2402);
and (n2473,n2465,n2469);
and (n2474,n2459,n2463);
and (n2475,n2453,n2457);
and (n2476,n2447,n2451);
and (n2477,n2441,n2445);
and (n2478,n2435,n2439);
and (n2479,n2429,n2433);
and (n2480,n2423,n2427);
and (n2481,n2418,n2421);
and (n2482,n2078,n2416);
or (n2483,n2484,n2489,n2577);
and (n2484,n2485,n2487);
xor (n2485,n2486,n2009);
xor (n2486,n1684,n1885);
xor (n2487,n2488,n2416);
xor (n2488,n2078,n2264);
and (n2489,n2487,n2490);
or (n2490,n2491,n2496,n2576);
and (n2491,n2492,n2494);
xor (n2492,n2493,n2014);
xor (n2493,n2011,n2012);
xor (n2494,n2495,n2421);
xor (n2495,n2418,n2419);
and (n2496,n2494,n2497);
or (n2497,n2498,n2503,n2575);
and (n2498,n2499,n2501);
xor (n2499,n2500,n2020);
xor (n2500,n2016,n2017);
xor (n2501,n2502,n2427);
xor (n2502,n2423,n2424);
and (n2503,n2501,n2504);
or (n2504,n2505,n2510,n2574);
and (n2505,n2506,n2508);
xor (n2506,n2507,n2026);
xor (n2507,n2022,n2023);
xor (n2508,n2509,n2433);
xor (n2509,n2429,n2430);
and (n2510,n2508,n2511);
or (n2511,n2512,n2517,n2573);
and (n2512,n2513,n2515);
xor (n2513,n2514,n2032);
xor (n2514,n2028,n2029);
xor (n2515,n2516,n2439);
xor (n2516,n2435,n2436);
and (n2517,n2515,n2518);
or (n2518,n2519,n2524,n2572);
and (n2519,n2520,n2522);
xor (n2520,n2521,n2038);
xor (n2521,n2034,n2035);
xor (n2522,n2523,n2445);
xor (n2523,n2441,n2442);
and (n2524,n2522,n2525);
or (n2525,n2526,n2531,n2571);
and (n2526,n2527,n2529);
xor (n2527,n2528,n2044);
xor (n2528,n2040,n2041);
xor (n2529,n2530,n2451);
xor (n2530,n2447,n2448);
and (n2531,n2529,n2532);
or (n2532,n2533,n2538,n2570);
and (n2533,n2534,n2536);
xor (n2534,n2535,n2050);
xor (n2535,n2046,n2047);
xor (n2536,n2537,n2457);
xor (n2537,n2453,n2454);
and (n2538,n2536,n2539);
or (n2539,n2540,n2545,n2569);
and (n2540,n2541,n2543);
xor (n2541,n2542,n2056);
xor (n2542,n2052,n2053);
xor (n2543,n2544,n2463);
xor (n2544,n2459,n2460);
and (n2545,n2543,n2546);
or (n2546,n2547,n2552,n2568);
and (n2547,n2548,n2550);
xor (n2548,n2549,n2062);
xor (n2549,n2058,n2059);
xor (n2550,n2551,n2469);
xor (n2551,n2465,n2466);
and (n2552,n2550,n2553);
or (n2553,n2554,n2557,n2567);
and (n2554,n2555,n2556);
xor (n2555,n2063,n2064);
xor (n2556,n2470,n2471);
and (n2557,n2556,n2558);
or (n2558,n2559,n2562,n2566);
and (n2559,n2560,n2561);
xor (n2560,n1998,n2000);
xor (n2561,n2405,n2407);
and (n2562,n2561,n2563);
and (n2563,n2564,n2565);
wire s0n2564,s1n2564,notn2564;
or (n2564,s0n2564,s1n2564);
not(notn2564,n1027);
and (s0n2564,notn2564,1'b0);
and (s1n2564,n1027,n1999);
wire s0n2565,s1n2565,notn2565;
or (n2565,s0n2565,s1n2565);
not(notn2565,n1027);
and (s0n2565,notn2565,1'b0);
and (s1n2565,n1027,n2406);
and (n2566,n2560,n2563);
and (n2567,n2555,n2558);
and (n2568,n2548,n2553);
and (n2569,n2541,n2546);
and (n2570,n2534,n2539);
and (n2571,n2527,n2532);
and (n2572,n2520,n2525);
and (n2573,n2513,n2518);
and (n2574,n2506,n2511);
and (n2575,n2499,n2504);
and (n2576,n2492,n2497);
and (n2577,n2485,n2490);
or (n2578,n2579,n2584,n2676);
and (n2579,n2580,n2582);
xor (n2580,n2581,n1592);
xor (n2581,n1587,n1589);
xor (n2582,n2583,n2490);
xor (n2583,n2485,n2487);
and (n2584,n2582,n2585);
or (n2585,n2586,n2591,n2675);
and (n2586,n2587,n2589);
xor (n2587,n2588,n1599);
xor (n2588,n1594,n1596);
xor (n2589,n2590,n2497);
xor (n2590,n2492,n2494);
and (n2591,n2589,n2592);
or (n2592,n2593,n2598,n2674);
and (n2593,n2594,n2596);
xor (n2594,n2595,n1606);
xor (n2595,n1601,n1603);
xor (n2596,n2597,n2504);
xor (n2597,n2499,n2501);
and (n2598,n2596,n2599);
or (n2599,n2600,n2605,n2673);
and (n2600,n2601,n2603);
xor (n2601,n2602,n1613);
xor (n2602,n1608,n1610);
xor (n2603,n2604,n2511);
xor (n2604,n2506,n2508);
and (n2605,n2603,n2606);
or (n2606,n2607,n2612,n2672);
and (n2607,n2608,n2610);
xor (n2608,n2609,n1620);
xor (n2609,n1615,n1617);
xor (n2610,n2611,n2518);
xor (n2611,n2513,n2515);
and (n2612,n2610,n2613);
or (n2613,n2614,n2619,n2671);
and (n2614,n2615,n2617);
xor (n2615,n2616,n1627);
xor (n2616,n1622,n1624);
xor (n2617,n2618,n2525);
xor (n2618,n2520,n2522);
and (n2619,n2617,n2620);
or (n2620,n2621,n2626,n2670);
and (n2621,n2622,n2624);
xor (n2622,n2623,n1634);
xor (n2623,n1629,n1631);
xor (n2624,n2625,n2532);
xor (n2625,n2527,n2529);
and (n2626,n2624,n2627);
or (n2627,n2628,n2633,n2669);
and (n2628,n2629,n2631);
xor (n2629,n2630,n1641);
xor (n2630,n1636,n1638);
xor (n2631,n2632,n2539);
xor (n2632,n2534,n2536);
and (n2633,n2631,n2634);
or (n2634,n2635,n2640,n2668);
and (n2635,n2636,n2638);
xor (n2636,n2637,n1648);
xor (n2637,n1643,n1645);
xor (n2638,n2639,n2546);
xor (n2639,n2541,n2543);
and (n2640,n2638,n2641);
or (n2641,n2642,n2647,n2667);
and (n2642,n2643,n2645);
xor (n2643,n2644,n1655);
xor (n2644,n1650,n1652);
xor (n2645,n2646,n2553);
xor (n2646,n2548,n2550);
and (n2647,n2645,n2648);
or (n2648,n2649,n2654,n2666);
and (n2649,n2650,n2652);
xor (n2650,n2651,n1660);
xor (n2651,n1657,n1658);
xor (n2652,n2653,n2558);
xor (n2653,n2555,n2556);
and (n2654,n2652,n2655);
or (n2655,n2656,n2661,n2665);
and (n2656,n2657,n2659);
xor (n2657,n2658,n1665);
xor (n2658,n1662,n1663);
xor (n2659,n2660,n2563);
xor (n2660,n2560,n2561);
and (n2661,n2659,n2662);
and (n2662,n2663,n2664);
xor (n2663,n1666,n1667);
xor (n2664,n2564,n2565);
and (n2665,n2657,n2662);
and (n2666,n2650,n2655);
and (n2667,n2643,n2648);
and (n2668,n2636,n2641);
and (n2669,n2629,n2634);
and (n2670,n2622,n2627);
and (n2671,n2615,n2620);
and (n2672,n2608,n2613);
and (n2673,n2601,n2606);
and (n2674,n2594,n2599);
and (n2675,n2587,n2592);
and (n2676,n2580,n2585);
and (n2677,n2678,n2680);
xor (n2678,n2679,n2585);
xor (n2679,n2580,n2582);
and (n2680,n2681,n2683);
xor (n2681,n2682,n2592);
xor (n2682,n2587,n2589);
and (n2683,n2684,n2686);
xor (n2684,n2685,n2599);
xor (n2685,n2594,n2596);
and (n2686,n2687,n2689);
xor (n2687,n2688,n2606);
xor (n2688,n2601,n2603);
and (n2689,n2690,n2692);
xor (n2690,n2691,n2613);
xor (n2691,n2608,n2610);
and (n2692,n2693,n2695);
xor (n2693,n2694,n2620);
xor (n2694,n2615,n2617);
and (n2695,n2696,n2698);
xor (n2696,n2697,n2627);
xor (n2697,n2622,n2624);
xor (n2698,n2699,n2634);
xor (n2699,n2629,n2631);
wire s0n2700,s1n2700,notn2700;
or (n2700,s0n2700,s1n2700);
not(notn2700,n2755);
and (s0n2700,notn2700,n2701);
and (s1n2700,n2755,n2707);
wire s0n2701,s1n2701,notn2701;
or (n2701,s0n2701,s1n2701);
not(notn2701,n2705);
and (s0n2701,notn2701,1'b0);
and (s1n2701,n2705,n2702);
wire s0n2702,s1n2702,notn2702;
or (n2702,s0n2702,s1n2702);
not(notn2702,n577);
and (s0n2702,notn2702,n562);
and (s1n2702,n577,n2703);
wire s0n2703,s1n2703,notn2703;
or (n2703,s0n2703,s1n2703);
not(notn2703,n2704);
and (s0n2703,notn2703,1'b0);
and (s1n2703,n2704,n21);
or (n2704,n558,n559,n560,n561);
and (n2705,n2706,n928);
and (n2706,n40,n592);
or (n2707,1'b0,n2708,n2720,n2732,n2744);
and (n2708,n2709,n2718);
or (n2709,1'b0,n2710,n2712,n2714,n2716);
and (n2710,n2711,n556);
and (n2712,n2713,n567);
and (n2714,n2715,n571);
and (n2716,n2717,n573);
and (n2718,n590,n2719);
and (n2719,n576,n27);
and (n2720,n2721,n2730);
or (n2721,1'b0,n2722,n2724,n2726,n2728);
and (n2722,n2723,n556);
and (n2724,n2725,n567);
and (n2726,n2727,n571);
and (n2728,n2729,n573);
and (n2730,n590,n2731);
and (n2731,n576,n32);
and (n2732,n2733,n2742);
or (n2733,1'b0,n2734,n2736,n2738,n2740);
and (n2734,n2735,n556);
and (n2736,n2737,n567);
and (n2738,n2739,n571);
and (n2740,n2741,n573);
and (n2742,n590,n2743);
and (n2743,n576,n36);
and (n2744,n2745,n2752);
or (n2745,1'b0,n2746,n2748,n2750,n2751);
and (n2746,n2747,n556);
and (n2748,n2749,n567);
and (n2750,n1251,n571);
and (n2751,n564,n573);
and (n2752,n590,n2753);
or (n2753,n577,n2754);
and (n2754,n576,n39);
and (n2755,n590,n2756);
nor (n2756,n2757,n2800,n2826,n2852);
wire s0n2757,s1n2757,notn2757;
or (n2757,s0n2757,s1n2757);
not(notn2757,n590);
and (s0n2757,notn2757,1'b0);
and (s1n2757,n590,n2758);
wire s0n2758,s1n2758,notn2758;
or (n2758,s0n2758,s1n2758);
not(notn2758,n590);
and (s0n2758,notn2758,n1027);
and (s1n2758,n590,n2759);
wire s0n2759,s1n2759,notn2759;
or (n2759,s0n2759,s1n2759);
not(notn2759,n648);
and (s0n2759,notn2759,n2760);
and (s1n2759,n648,n1065);
wire s0n2760,s1n2760,notn2760;
or (n2760,s0n2760,s1n2760);
not(notn2760,n577);
and (s0n2760,notn2760,n2761);
and (s1n2760,n577,n2766);
or (n2761,n2762,n2763,n2764,n2765);
and (n2762,n1032,n580);
and (n2763,n1043,n584);
and (n2764,n1054,n587);
and (n2765,n1065,n589);
or (n2766,1'b0,n2767,n2769,n2771,n2774,n2776,n2778,n2780,n2782,n2784,n2786,n2788,n2790,n2792,n2794,n2796,n2798);
and (n2767,n1035,n2768);
and (n2768,n28,n29,n581,n582,n591);
and (n2769,n1037,n2770);
and (n2770,n33,n29,n581,n582,n591);
and (n2771,n1039,n2772);
and (n2772,n28,n2773,n581,n582,n591);
not (n2773,n29);
and (n2774,n1032,n2775);
and (n2775,n33,n2773,n581,n582,n591);
and (n2776,n1046,n2777);
and (n2777,n28,n29,n585,n582,n591);
and (n2778,n1048,n2779);
and (n2779,n33,n29,n585,n582,n591);
and (n2780,n1050,n2781);
and (n2781,n28,n2773,n585,n582,n591);
and (n2782,n1043,n2783);
and (n2783,n33,n2773,n585,n582,n591);
and (n2784,n1057,n2785);
nor (n2785,n33,n2773,n585,n582,n555);
and (n2786,n1059,n2787);
nor (n2787,n28,n2773,n585,n582,n555);
and (n2788,n1061,n2789);
nor (n2789,n33,n29,n585,n582,n555);
and (n2790,n1054,n2791);
nor (n2791,n28,n29,n585,n582,n555);
and (n2792,n1068,n2793);
nor (n2793,n33,n2773,n581,n582,n555);
and (n2794,n1070,n2795);
nor (n2795,n28,n2773,n581,n582,n555);
and (n2796,n1072,n2797);
nor (n2797,n33,n29,n581,n582,n555);
and (n2798,n1065,n2799);
nor (n2799,n28,n29,n581,n582,n555);
wire s0n2800,s1n2800,notn2800;
or (n2800,s0n2800,s1n2800);
not(notn2800,n590);
and (s0n2800,notn2800,1'b0);
and (s1n2800,n590,n2801);
wire s0n2801,s1n2801,notn2801;
or (n2801,s0n2801,s1n2801);
not(notn2801,n590);
and (s0n2801,notn2801,n979);
and (s1n2801,n590,n2802);
wire s0n2802,s1n2802,notn2802;
or (n2802,s0n2802,s1n2802);
not(notn2802,n648);
and (s0n2802,notn2802,n2803);
and (s1n2802,n648,n1017);
wire s0n2803,s1n2803,notn2803;
or (n2803,s0n2803,s1n2803);
not(notn2803,n577);
and (s0n2803,notn2803,n2804);
and (s1n2803,n577,n2809);
or (n2804,n2805,n2806,n2807,n2808);
and (n2805,n984,n580);
and (n2806,n995,n584);
and (n2807,n1006,n587);
and (n2808,n1017,n589);
or (n2809,1'b0,n2810,n2811,n2812,n2813,n2814,n2815,n2816,n2817,n2818,n2819,n2820,n2821,n2822,n2823,n2824,n2825);
and (n2810,n987,n2768);
and (n2811,n989,n2770);
and (n2812,n991,n2772);
and (n2813,n984,n2775);
and (n2814,n998,n2777);
and (n2815,n1000,n2779);
and (n2816,n1002,n2781);
and (n2817,n995,n2783);
and (n2818,n1009,n2785);
and (n2819,n1011,n2787);
and (n2820,n1013,n2789);
and (n2821,n1006,n2791);
and (n2822,n1020,n2793);
and (n2823,n1022,n2795);
and (n2824,n1024,n2797);
and (n2825,n1017,n2799);
wire s0n2826,s1n2826,notn2826;
or (n2826,s0n2826,s1n2826);
not(notn2826,n590);
and (s0n2826,notn2826,1'b0);
and (s1n2826,n590,n2827);
wire s0n2827,s1n2827,notn2827;
or (n2827,s0n2827,s1n2827);
not(notn2827,n590);
and (s0n2827,notn2827,n699);
and (s1n2827,n590,n2828);
wire s0n2828,s1n2828,notn2828;
or (n2828,s0n2828,s1n2828);
not(notn2828,n648);
and (s0n2828,notn2828,n2829);
and (s1n2828,n648,n737);
wire s0n2829,s1n2829,notn2829;
or (n2829,s0n2829,s1n2829);
not(notn2829,n577);
and (s0n2829,notn2829,n2830);
and (s1n2829,n577,n2835);
or (n2830,n2831,n2832,n2833,n2834);
and (n2831,n704,n580);
and (n2832,n715,n584);
and (n2833,n726,n587);
and (n2834,n737,n589);
or (n2835,1'b0,n2836,n2837,n2838,n2839,n2840,n2841,n2842,n2843,n2844,n2845,n2846,n2847,n2848,n2849,n2850,n2851);
and (n2836,n707,n2768);
and (n2837,n709,n2770);
and (n2838,n711,n2772);
and (n2839,n704,n2775);
and (n2840,n718,n2777);
and (n2841,n720,n2779);
and (n2842,n722,n2781);
and (n2843,n715,n2783);
and (n2844,n729,n2785);
and (n2845,n731,n2787);
and (n2846,n733,n2789);
and (n2847,n726,n2791);
and (n2848,n740,n2793);
and (n2849,n742,n2795);
and (n2850,n744,n2797);
and (n2851,n737,n2799);
wire s0n2852,s1n2852,notn2852;
or (n2852,s0n2852,s1n2852);
not(notn2852,n590);
and (s0n2852,notn2852,1'b0);
and (s1n2852,n590,n2853);
wire s0n2853,s1n2853,notn2853;
or (n2853,s0n2853,s1n2853);
not(notn2853,n590);
and (s0n2853,notn2853,n651);
and (s1n2853,n590,n2854);
wire s0n2854,s1n2854,notn2854;
or (n2854,s0n2854,s1n2854);
not(notn2854,n648);
and (s0n2854,notn2854,n2855);
and (s1n2854,n648,n689);
wire s0n2855,s1n2855,notn2855;
or (n2855,s0n2855,s1n2855);
not(notn2855,n577);
and (s0n2855,notn2855,n2856);
and (s1n2855,n577,n2861);
or (n2856,n2857,n2858,n2859,n2860);
and (n2857,n656,n580);
and (n2858,n667,n584);
and (n2859,n678,n587);
and (n2860,n689,n589);
or (n2861,1'b0,n2862,n2863,n2864,n2865,n2866,n2867,n2868,n2869,n2870,n2871,n2872,n2873,n2874,n2875,n2876,n2877);
and (n2862,n659,n2768);
and (n2863,n661,n2770);
and (n2864,n663,n2772);
and (n2865,n656,n2775);
and (n2866,n670,n2777);
and (n2867,n672,n2779);
and (n2868,n674,n2781);
and (n2869,n667,n2783);
and (n2870,n681,n2785);
and (n2871,n683,n2787);
and (n2872,n685,n2789);
and (n2873,n678,n2791);
and (n2874,n692,n2793);
and (n2875,n694,n2795);
and (n2876,n696,n2797);
and (n2877,n689,n2799);
or (n2878,n2879,n2882,n2700);
and (n2879,n2880,n8688);
wire s0n2880,s1n2880,notn2880;
or (n2880,s0n2880,s1n2880);
not(notn2880,n4969);
and (s0n2880,notn2880,1'b0);
and (s1n2880,n4969,n2881);
or (n2881,1'b0,n2882,n8675,n8685,n8686,n8687);
and (n2882,n2883,n2907);
wire s0n2883,s1n2883,notn2883;
or (n2883,s0n2883,s1n2883);
not(notn2883,n2902);
and (s0n2883,notn2883,1'b0);
and (s1n2883,n2902,n2884);
xor (n2884,n2885,n8653);
or (n2885,n2886,n7879,n8652);
and (n2886,n2887,n4950);
or (n2887,1'b0,n2888,n2899,n2910,n4886);
and (n2888,n2889,n2893);
wire s0n2889,s1n2889,notn2889;
or (n2889,s0n2889,s1n2889);
not(notn2889,n2891);
and (s0n2889,notn2889,1'b0);
and (s1n2889,n2891,n2890);
and (n2891,n2892,n2704);
nand (n2892,n558,n568,n560,n574);
or (n2893,n2894,n2897);
nor (n2894,n2895,n2800,n2826,n2896);
not (n2895,n2757);
not (n2896,n2852);
and (n2897,n2757,n2800,n2898,n2852);
not (n2898,n2826);
and (n2899,n2900,n2907);
wire s0n2900,s1n2900,notn2900;
or (n2900,s0n2900,s1n2900);
not(notn2900,n2902);
and (s0n2900,notn2900,1'b0);
and (s1n2900,n2902,n2901);
or (n2902,n2903,n556);
or (n2903,n2904,n571);
or (n2904,n2905,n2906);
and (n2905,n558,n559,n560,n574);
not (n2906,n2892);
or (n2907,n2908,n2909);
and (n2908,n2895,n2800,n2826,n2896);
and (n2909,n2895,n2800,n2826,n2852);
and (n2910,n2911,n4883);
wire s0n2911,s1n2911,notn2911;
or (n2911,s0n2911,s1n2911);
not(notn2911,n4878);
and (s0n2911,notn2911,n2912);
and (s1n2911,n4878,1'b0);
wire s0n2912,s1n2912,notn2912;
or (n2912,s0n2912,s1n2912);
not(notn2912,n4873);
and (s0n2912,notn2912,n2913);
and (s1n2912,n4873,1'b1);
wire s0n2913,s1n2913,notn2913;
or (n2913,s0n2913,s1n2913);
not(notn2913,n4861);
and (s0n2913,notn2913,1'b0);
and (s1n2913,n4861,n2914);
xor (n2914,n2915,n4838);
xor (n2915,n2916,n4785);
xor (n2916,n2917,n4377);
xor (n2917,n2918,n4375);
xor (n2918,n2919,n4345);
not (n2919,n2920);
or (n2920,n2921,n3776);
or (n2921,n2922,n3049,n3775);
and (n2922,n2923,n3018);
or (n2923,1'b0,n2924,n2978,n2992,n3006);
and (n2924,n2925,n2718);
or (n2925,1'b0,n2926,n2952,n2960,n2969);
and (n2926,n2927,n2932);
wire s0n2927,s1n2927,notn2927;
or (n2927,s0n2927,s1n2927);
not(notn2927,n2929);
and (s0n2927,notn2927,n2711);
and (s1n2927,n2929,n2928);
or (n2929,n2930,n2931);
and (n2930,n2757,n2800,n2826,n2896);
and (n2931,n2757,n2800,n2826,n2852);
or (n2932,n2933,n2951);
or (n2933,n2934,n2947);
and (n2934,n2935,n556);
or (n2935,n2936,n2931);
or (n2936,n2937,n2930);
or (n2937,n2938,n2946);
or (n2938,n2939,n2945);
or (n2939,n2940,n2944);
or (n2940,n2941,n2942);
nor (n2941,n2757,n2800,n2826,n2896);
and (n2942,n2895,n2943,n2826,n2896);
not (n2943,n2800);
and (n2944,n2895,n2943,n2826,n2852);
and (n2945,n2757,n2943,n2826,n2896);
and (n2946,n2757,n2943,n2826,n2852);
and (n2947,n2948,n567);
or (n2948,n2949,n2897);
or (n2949,n2950,n2894);
nor (n2950,n2757,n2943,n2826,n2896);
and (n2951,n2907,n567);
and (n2952,n2953,n2955);
wire s0n2953,s1n2953,notn2953;
or (n2953,s0n2953,s1n2953);
not(notn2953,n2929);
and (s0n2953,notn2953,n2713);
and (s1n2953,n2929,n2954);
or (n2955,n2956,n2959);
or (n2956,n2957,n2958);
and (n2957,n2935,n567);
and (n2958,n2948,n571);
and (n2959,n2907,n573);
and (n2960,n2961,n2963);
wire s0n2961,s1n2961,notn2961;
or (n2961,s0n2961,s1n2961);
not(notn2961,n2929);
and (s0n2961,notn2961,n2715);
and (s1n2961,n2929,n2962);
or (n2963,n2964,n2967);
or (n2964,n2965,n2966);
and (n2965,n2935,n571);
and (n2966,n2948,n573);
and (n2967,n2907,n2968);
and (n2968,n557,n559,n560,n574);
and (n2969,n2970,n2972);
wire s0n2970,s1n2970,notn2970;
or (n2970,s0n2970,s1n2970);
not(notn2970,n2929);
and (s0n2970,notn2970,n2717);
and (s1n2970,n2929,n2971);
or (n2972,n2973,n2976);
or (n2973,n2974,n2975);
and (n2974,n2935,n573);
and (n2975,n2948,n2906);
and (n2976,n2907,n2977);
nor (n2977,n558,n559,n560,n574);
and (n2978,n2979,n2730);
or (n2979,1'b0,n2980,n2983,n2986,n2989);
and (n2980,n2981,n2932);
wire s0n2981,s1n2981,notn2981;
or (n2981,s0n2981,s1n2981);
not(notn2981,n2929);
and (s0n2981,notn2981,n2723);
and (s1n2981,n2929,n2982);
and (n2983,n2984,n2955);
wire s0n2984,s1n2984,notn2984;
or (n2984,s0n2984,s1n2984);
not(notn2984,n2929);
and (s0n2984,notn2984,n2725);
and (s1n2984,n2929,n2985);
and (n2986,n2987,n2963);
wire s0n2987,s1n2987,notn2987;
or (n2987,s0n2987,s1n2987);
not(notn2987,n2929);
and (s0n2987,notn2987,n2727);
and (s1n2987,n2929,n2988);
and (n2989,n2990,n2972);
wire s0n2990,s1n2990,notn2990;
or (n2990,s0n2990,s1n2990);
not(notn2990,n2929);
and (s0n2990,notn2990,n2729);
and (s1n2990,n2929,n2991);
and (n2992,n2993,n2742);
or (n2993,1'b0,n2994,n2997,n3000,n3003);
and (n2994,n2995,n2932);
wire s0n2995,s1n2995,notn2995;
or (n2995,s0n2995,s1n2995);
not(notn2995,n2929);
and (s0n2995,notn2995,n2735);
and (s1n2995,n2929,n2996);
and (n2997,n2998,n2955);
wire s0n2998,s1n2998,notn2998;
or (n2998,s0n2998,s1n2998);
not(notn2998,n2929);
and (s0n2998,notn2998,n2737);
and (s1n2998,n2929,n2999);
and (n3000,n3001,n2963);
wire s0n3001,s1n3001,notn3001;
or (n3001,s0n3001,s1n3001);
not(notn3001,n2929);
and (s0n3001,notn3001,n2739);
and (s1n3001,n2929,n3002);
and (n3003,n3004,n2972);
wire s0n3004,s1n3004,notn3004;
or (n3004,s0n3004,s1n3004);
not(notn3004,n2929);
and (s0n3004,notn3004,n2741);
and (s1n3004,n2929,n3005);
and (n3006,n3007,n2752);
or (n3007,1'b0,n3008,n3011,n3014,n3016);
and (n3008,n3009,n2932);
wire s0n3009,s1n3009,notn3009;
or (n3009,s0n3009,s1n3009);
not(notn3009,n2929);
and (s0n3009,notn3009,n2747);
and (s1n3009,n2929,n3010);
and (n3011,n3012,n2955);
wire s0n3012,s1n3012,notn3012;
or (n3012,s0n3012,s1n3012);
not(notn3012,n2929);
and (s0n3012,notn3012,n2749);
and (s1n3012,n2929,n3013);
and (n3014,n3015,n2963);
wire s0n3015,s1n3015,notn3015;
or (n3015,s0n3015,s1n3015);
not(notn3015,n2929);
and (s0n3015,notn3015,n1251);
and (s1n3015,n2929,n2087);
and (n3016,n3017,n2972);
wire s0n3017,s1n3017,notn3017;
or (n3017,s0n3017,s1n3017);
not(notn3017,n2929);
and (s0n3017,notn3017,n564);
and (s1n3017,n2929,n1692);
or (n3018,1'b0,n3019,n3028,n3034,n3043);
and (n3019,n3020,n2718);
or (n3020,1'b0,n3021,n3025,n3026,n3027);
and (n3021,n3022,n2932);
wire s0n3022,s1n3022,notn3022;
or (n3022,s0n3022,s1n3022);
not(notn3022,n2929);
and (s0n3022,notn3022,n3023);
and (s1n3022,n2929,n3024);
and (n3025,n2927,n2955);
and (n3026,n2953,n2963);
and (n3027,n2961,n2972);
and (n3028,n3029,n2730);
or (n3029,1'b0,n3030,n3031,n3032,n3033);
and (n3030,n2970,n2932);
and (n3031,n2981,n2955);
and (n3032,n2984,n2963);
and (n3033,n2987,n2972);
and (n3034,n3035,n2742);
or (n3035,1'b0,n3036,n3040,n3041,n3042);
and (n3036,n3037,n2932);
wire s0n3037,s1n3037,notn3037;
or (n3037,s0n3037,s1n3037);
not(notn3037,n2929);
and (s0n3037,notn3037,n3038);
and (s1n3037,n2929,n3039);
and (n3040,n2995,n2955);
and (n3041,n2998,n2963);
and (n3042,n3001,n2972);
and (n3043,n3044,n2752);
or (n3044,1'b0,n3045,n3046,n3047,n3048);
and (n3045,n3004,n2932);
and (n3046,n3009,n2955);
and (n3047,n3012,n2963);
and (n3048,n3015,n2972);
and (n3049,n3018,n3050);
or (n3050,n3051,n3152,n3774);
and (n3051,n3052,n3121);
or (n3052,1'b0,n3053,n3071,n3089,n3107);
and (n3053,n3054,n2718);
or (n3054,1'b0,n3055,n3059,n3063,n3067);
and (n3055,n3056,n2932);
wire s0n3056,s1n3056,notn3056;
or (n3056,s0n3056,s1n3056);
not(notn3056,n2929);
and (s0n3056,notn3056,n3057);
and (s1n3056,n2929,n3058);
and (n3059,n3060,n2955);
wire s0n3060,s1n3060,notn3060;
or (n3060,s0n3060,s1n3060);
not(notn3060,n2929);
and (s0n3060,notn3060,n3061);
and (s1n3060,n2929,n3062);
and (n3063,n3064,n2963);
wire s0n3064,s1n3064,notn3064;
or (n3064,s0n3064,s1n3064);
not(notn3064,n2929);
and (s0n3064,notn3064,n3065);
and (s1n3064,n2929,n3066);
and (n3067,n3068,n2972);
wire s0n3068,s1n3068,notn3068;
or (n3068,s0n3068,s1n3068);
not(notn3068,n2929);
and (s0n3068,notn3068,n3069);
and (s1n3068,n2929,n3070);
and (n3071,n3072,n2730);
or (n3072,1'b0,n3073,n3077,n3081,n3085);
and (n3073,n3074,n2932);
wire s0n3074,s1n3074,notn3074;
or (n3074,s0n3074,s1n3074);
not(notn3074,n2929);
and (s0n3074,notn3074,n3075);
and (s1n3074,n2929,n3076);
and (n3077,n3078,n2955);
wire s0n3078,s1n3078,notn3078;
or (n3078,s0n3078,s1n3078);
not(notn3078,n2929);
and (s0n3078,notn3078,n3079);
and (s1n3078,n2929,n3080);
and (n3081,n3082,n2963);
wire s0n3082,s1n3082,notn3082;
or (n3082,s0n3082,s1n3082);
not(notn3082,n2929);
and (s0n3082,notn3082,n3083);
and (s1n3082,n2929,n3084);
and (n3085,n3086,n2972);
wire s0n3086,s1n3086,notn3086;
or (n3086,s0n3086,s1n3086);
not(notn3086,n2929);
and (s0n3086,notn3086,n3087);
and (s1n3086,n2929,n3088);
and (n3089,n3090,n2742);
or (n3090,1'b0,n3091,n3095,n3099,n3103);
and (n3091,n3092,n2932);
wire s0n3092,s1n3092,notn3092;
or (n3092,s0n3092,s1n3092);
not(notn3092,n2929);
and (s0n3092,notn3092,n3093);
and (s1n3092,n2929,n3094);
and (n3095,n3096,n2955);
wire s0n3096,s1n3096,notn3096;
or (n3096,s0n3096,s1n3096);
not(notn3096,n2929);
and (s0n3096,notn3096,n3097);
and (s1n3096,n2929,n3098);
and (n3099,n3100,n2963);
wire s0n3100,s1n3100,notn3100;
or (n3100,s0n3100,s1n3100);
not(notn3100,n2929);
and (s0n3100,notn3100,n3101);
and (s1n3100,n2929,n3102);
and (n3103,n3104,n2972);
wire s0n3104,s1n3104,notn3104;
or (n3104,s0n3104,s1n3104);
not(notn3104,n2929);
and (s0n3104,notn3104,n3105);
and (s1n3104,n2929,n3106);
and (n3107,n3108,n2752);
or (n3108,1'b0,n3109,n3113,n3117,n3119);
and (n3109,n3110,n2932);
wire s0n3110,s1n3110,notn3110;
or (n3110,s0n3110,s1n3110);
not(notn3110,n2929);
and (s0n3110,notn3110,n3111);
and (s1n3110,n2929,n3112);
and (n3113,n3114,n2955);
wire s0n3114,s1n3114,notn3114;
or (n3114,s0n3114,s1n3114);
not(notn3114,n2929);
and (s0n3114,notn3114,n3115);
and (s1n3114,n2929,n3116);
and (n3117,n3118,n2963);
wire s0n3118,s1n3118,notn3118;
or (n3118,s0n3118,s1n3118);
not(notn3118,n2929);
and (s0n3118,notn3118,n1267);
and (s1n3118,n2929,n2103);
and (n3119,n3120,n2972);
wire s0n3120,s1n3120,notn3120;
or (n3120,s0n3120,s1n3120);
not(notn3120,n2929);
and (s0n3120,notn3120,n755);
and (s1n3120,n2929,n1708);
or (n3121,1'b0,n3122,n3131,n3137,n3146);
and (n3122,n3123,n2718);
or (n3123,1'b0,n3124,n3128,n3129,n3130);
and (n3124,n3125,n2932);
wire s0n3125,s1n3125,notn3125;
or (n3125,s0n3125,s1n3125);
not(notn3125,n2929);
and (s0n3125,notn3125,n3126);
and (s1n3125,n2929,n3127);
and (n3128,n3056,n2955);
and (n3129,n3060,n2963);
and (n3130,n3064,n2972);
and (n3131,n3132,n2730);
or (n3132,1'b0,n3133,n3134,n3135,n3136);
and (n3133,n3068,n2932);
and (n3134,n3074,n2955);
and (n3135,n3078,n2963);
and (n3136,n3082,n2972);
and (n3137,n3138,n2742);
or (n3138,1'b0,n3139,n3143,n3144,n3145);
and (n3139,n3140,n2932);
wire s0n3140,s1n3140,notn3140;
or (n3140,s0n3140,s1n3140);
not(notn3140,n2929);
and (s0n3140,notn3140,n3141);
and (s1n3140,n2929,n3142);
and (n3143,n3092,n2955);
and (n3144,n3096,n2963);
and (n3145,n3100,n2972);
and (n3146,n3147,n2752);
or (n3147,1'b0,n3148,n3149,n3150,n3151);
and (n3148,n3104,n2932);
and (n3149,n3110,n2955);
and (n3150,n3114,n2963);
and (n3151,n3118,n2972);
and (n3152,n3121,n3153);
or (n3153,n3154,n3255,n3773);
and (n3154,n3155,n3224);
or (n3155,1'b0,n3156,n3174,n3192,n3210);
and (n3156,n3157,n2718);
or (n3157,1'b0,n3158,n3162,n3166,n3170);
and (n3158,n3159,n2932);
wire s0n3159,s1n3159,notn3159;
or (n3159,s0n3159,s1n3159);
not(notn3159,n2929);
and (s0n3159,notn3159,n3160);
and (s1n3159,n2929,n3161);
and (n3162,n3163,n2955);
wire s0n3163,s1n3163,notn3163;
or (n3163,s0n3163,s1n3163);
not(notn3163,n2929);
and (s0n3163,notn3163,n3164);
and (s1n3163,n2929,n3165);
and (n3166,n3167,n2963);
wire s0n3167,s1n3167,notn3167;
or (n3167,s0n3167,s1n3167);
not(notn3167,n2929);
and (s0n3167,notn3167,n3168);
and (s1n3167,n2929,n3169);
and (n3170,n3171,n2972);
wire s0n3171,s1n3171,notn3171;
or (n3171,s0n3171,s1n3171);
not(notn3171,n2929);
and (s0n3171,notn3171,n3172);
and (s1n3171,n2929,n3173);
and (n3174,n3175,n2730);
or (n3175,1'b0,n3176,n3180,n3184,n3188);
and (n3176,n3177,n2932);
wire s0n3177,s1n3177,notn3177;
or (n3177,s0n3177,s1n3177);
not(notn3177,n2929);
and (s0n3177,notn3177,n3178);
and (s1n3177,n2929,n3179);
and (n3180,n3181,n2955);
wire s0n3181,s1n3181,notn3181;
or (n3181,s0n3181,s1n3181);
not(notn3181,n2929);
and (s0n3181,notn3181,n3182);
and (s1n3181,n2929,n3183);
and (n3184,n3185,n2963);
wire s0n3185,s1n3185,notn3185;
or (n3185,s0n3185,s1n3185);
not(notn3185,n2929);
and (s0n3185,notn3185,n3186);
and (s1n3185,n2929,n3187);
and (n3188,n3189,n2972);
wire s0n3189,s1n3189,notn3189;
or (n3189,s0n3189,s1n3189);
not(notn3189,n2929);
and (s0n3189,notn3189,n3190);
and (s1n3189,n2929,n3191);
and (n3192,n3193,n2742);
or (n3193,1'b0,n3194,n3198,n3202,n3206);
and (n3194,n3195,n2932);
wire s0n3195,s1n3195,notn3195;
or (n3195,s0n3195,s1n3195);
not(notn3195,n2929);
and (s0n3195,notn3195,n3196);
and (s1n3195,n2929,n3197);
and (n3198,n3199,n2955);
wire s0n3199,s1n3199,notn3199;
or (n3199,s0n3199,s1n3199);
not(notn3199,n2929);
and (s0n3199,notn3199,n3200);
and (s1n3199,n2929,n3201);
and (n3202,n3203,n2963);
wire s0n3203,s1n3203,notn3203;
or (n3203,s0n3203,s1n3203);
not(notn3203,n2929);
and (s0n3203,notn3203,n3204);
and (s1n3203,n2929,n3205);
and (n3206,n3207,n2972);
wire s0n3207,s1n3207,notn3207;
or (n3207,s0n3207,s1n3207);
not(notn3207,n2929);
and (s0n3207,notn3207,n3208);
and (s1n3207,n2929,n3209);
and (n3210,n3211,n2752);
or (n3211,1'b0,n3212,n3216,n3220,n3222);
and (n3212,n3213,n2932);
wire s0n3213,s1n3213,notn3213;
or (n3213,s0n3213,s1n3213);
not(notn3213,n2929);
and (s0n3213,notn3213,n3214);
and (s1n3213,n2929,n3215);
and (n3216,n3217,n2955);
wire s0n3217,s1n3217,notn3217;
or (n3217,s0n3217,s1n3217);
not(notn3217,n2929);
and (s0n3217,notn3217,n3218);
and (s1n3217,n2929,n3219);
and (n3220,n3221,n2963);
wire s0n3221,s1n3221,notn3221;
or (n3221,s0n3221,s1n3221);
not(notn3221,n2929);
and (s0n3221,notn3221,n1283);
and (s1n3221,n2929,n2119);
and (n3222,n3223,n2972);
wire s0n3223,s1n3223,notn3223;
or (n3223,s0n3223,s1n3223);
not(notn3223,n2929);
and (s0n3223,notn3223,n779);
and (s1n3223,n2929,n1727);
or (n3224,1'b0,n3225,n3234,n3240,n3249);
and (n3225,n3226,n2718);
or (n3226,1'b0,n3227,n3231,n3232,n3233);
and (n3227,n3228,n2932);
wire s0n3228,s1n3228,notn3228;
or (n3228,s0n3228,s1n3228);
not(notn3228,n2929);
and (s0n3228,notn3228,n3229);
and (s1n3228,n2929,n3230);
and (n3231,n3159,n2955);
and (n3232,n3163,n2963);
and (n3233,n3167,n2972);
and (n3234,n3235,n2730);
or (n3235,1'b0,n3236,n3237,n3238,n3239);
and (n3236,n3171,n2932);
and (n3237,n3177,n2955);
and (n3238,n3181,n2963);
and (n3239,n3185,n2972);
and (n3240,n3241,n2742);
or (n3241,1'b0,n3242,n3246,n3247,n3248);
and (n3242,n3243,n2932);
wire s0n3243,s1n3243,notn3243;
or (n3243,s0n3243,s1n3243);
not(notn3243,n2929);
and (s0n3243,notn3243,n3244);
and (s1n3243,n2929,n3245);
and (n3246,n3195,n2955);
and (n3247,n3199,n2963);
and (n3248,n3203,n2972);
and (n3249,n3250,n2752);
or (n3250,1'b0,n3251,n3252,n3253,n3254);
and (n3251,n3207,n2932);
and (n3252,n3213,n2955);
and (n3253,n3217,n2963);
and (n3254,n3221,n2972);
and (n3255,n3224,n3256);
or (n3256,n3257,n3358,n3772);
and (n3257,n3258,n3327);
or (n3258,1'b0,n3259,n3277,n3295,n3313);
and (n3259,n3260,n2718);
or (n3260,1'b0,n3261,n3265,n3269,n3273);
and (n3261,n3262,n2932);
wire s0n3262,s1n3262,notn3262;
or (n3262,s0n3262,s1n3262);
not(notn3262,n2929);
and (s0n3262,notn3262,n3263);
and (s1n3262,n2929,n3264);
and (n3265,n3266,n2955);
wire s0n3266,s1n3266,notn3266;
or (n3266,s0n3266,s1n3266);
not(notn3266,n2929);
and (s0n3266,notn3266,n3267);
and (s1n3266,n2929,n3268);
and (n3269,n3270,n2963);
wire s0n3270,s1n3270,notn3270;
or (n3270,s0n3270,s1n3270);
not(notn3270,n2929);
and (s0n3270,notn3270,n3271);
and (s1n3270,n2929,n3272);
and (n3273,n3274,n2972);
wire s0n3274,s1n3274,notn3274;
or (n3274,s0n3274,s1n3274);
not(notn3274,n2929);
and (s0n3274,notn3274,n3275);
and (s1n3274,n2929,n3276);
and (n3277,n3278,n2730);
or (n3278,1'b0,n3279,n3283,n3287,n3291);
and (n3279,n3280,n2932);
wire s0n3280,s1n3280,notn3280;
or (n3280,s0n3280,s1n3280);
not(notn3280,n2929);
and (s0n3280,notn3280,n3281);
and (s1n3280,n2929,n3282);
and (n3283,n3284,n2955);
wire s0n3284,s1n3284,notn3284;
or (n3284,s0n3284,s1n3284);
not(notn3284,n2929);
and (s0n3284,notn3284,n3285);
and (s1n3284,n2929,n3286);
and (n3287,n3288,n2963);
wire s0n3288,s1n3288,notn3288;
or (n3288,s0n3288,s1n3288);
not(notn3288,n2929);
and (s0n3288,notn3288,n3289);
and (s1n3288,n2929,n3290);
and (n3291,n3292,n2972);
wire s0n3292,s1n3292,notn3292;
or (n3292,s0n3292,s1n3292);
not(notn3292,n2929);
and (s0n3292,notn3292,n3293);
and (s1n3292,n2929,n3294);
and (n3295,n3296,n2742);
or (n3296,1'b0,n3297,n3301,n3305,n3309);
and (n3297,n3298,n2932);
wire s0n3298,s1n3298,notn3298;
or (n3298,s0n3298,s1n3298);
not(notn3298,n2929);
and (s0n3298,notn3298,n3299);
and (s1n3298,n2929,n3300);
and (n3301,n3302,n2955);
wire s0n3302,s1n3302,notn3302;
or (n3302,s0n3302,s1n3302);
not(notn3302,n2929);
and (s0n3302,notn3302,n3303);
and (s1n3302,n2929,n3304);
and (n3305,n3306,n2963);
wire s0n3306,s1n3306,notn3306;
or (n3306,s0n3306,s1n3306);
not(notn3306,n2929);
and (s0n3306,notn3306,n3307);
and (s1n3306,n2929,n3308);
and (n3309,n3310,n2972);
wire s0n3310,s1n3310,notn3310;
or (n3310,s0n3310,s1n3310);
not(notn3310,n2929);
and (s0n3310,notn3310,n3311);
and (s1n3310,n2929,n3312);
and (n3313,n3314,n2752);
or (n3314,1'b0,n3315,n3319,n3323,n3325);
and (n3315,n3316,n2932);
wire s0n3316,s1n3316,notn3316;
or (n3316,s0n3316,s1n3316);
not(notn3316,n2929);
and (s0n3316,notn3316,n3317);
and (s1n3316,n2929,n3318);
and (n3319,n3320,n2955);
wire s0n3320,s1n3320,notn3320;
or (n3320,s0n3320,s1n3320);
not(notn3320,n2929);
and (s0n3320,notn3320,n3321);
and (s1n3320,n2929,n3322);
and (n3323,n3324,n2963);
wire s0n3324,s1n3324,notn3324;
or (n3324,s0n3324,s1n3324);
not(notn3324,n2929);
and (s0n3324,notn3324,n1299);
and (s1n3324,n2929,n2135);
and (n3325,n3326,n2972);
wire s0n3326,s1n3326,notn3326;
or (n3326,s0n3326,s1n3326);
not(notn3326,n2929);
and (s0n3326,notn3326,n795);
and (s1n3326,n2929,n1753);
or (n3327,1'b0,n3328,n3337,n3343,n3352);
and (n3328,n3329,n2718);
or (n3329,1'b0,n3330,n3334,n3335,n3336);
and (n3330,n3331,n2932);
wire s0n3331,s1n3331,notn3331;
or (n3331,s0n3331,s1n3331);
not(notn3331,n2929);
and (s0n3331,notn3331,n3332);
and (s1n3331,n2929,n3333);
and (n3334,n3262,n2955);
and (n3335,n3266,n2963);
and (n3336,n3270,n2972);
and (n3337,n3338,n2730);
or (n3338,1'b0,n3339,n3340,n3341,n3342);
and (n3339,n3274,n2932);
and (n3340,n3280,n2955);
and (n3341,n3284,n2963);
and (n3342,n3288,n2972);
and (n3343,n3344,n2742);
or (n3344,1'b0,n3345,n3349,n3350,n3351);
and (n3345,n3346,n2932);
wire s0n3346,s1n3346,notn3346;
or (n3346,s0n3346,s1n3346);
not(notn3346,n2929);
and (s0n3346,notn3346,n3347);
and (s1n3346,n2929,n3348);
and (n3349,n3298,n2955);
and (n3350,n3302,n2963);
and (n3351,n3306,n2972);
and (n3352,n3353,n2752);
or (n3353,1'b0,n3354,n3355,n3356,n3357);
and (n3354,n3310,n2932);
and (n3355,n3316,n2955);
and (n3356,n3320,n2963);
and (n3357,n3324,n2972);
and (n3358,n3327,n3359);
or (n3359,n3360,n3461,n3771);
and (n3360,n3361,n3430);
or (n3361,1'b0,n3362,n3380,n3398,n3416);
and (n3362,n3363,n2718);
or (n3363,1'b0,n3364,n3368,n3372,n3376);
and (n3364,n3365,n2932);
wire s0n3365,s1n3365,notn3365;
or (n3365,s0n3365,s1n3365);
not(notn3365,n2929);
and (s0n3365,notn3365,n3366);
and (s1n3365,n2929,n3367);
and (n3368,n3369,n2955);
wire s0n3369,s1n3369,notn3369;
or (n3369,s0n3369,s1n3369);
not(notn3369,n2929);
and (s0n3369,notn3369,n3370);
and (s1n3369,n2929,n3371);
and (n3372,n3373,n2963);
wire s0n3373,s1n3373,notn3373;
or (n3373,s0n3373,s1n3373);
not(notn3373,n2929);
and (s0n3373,notn3373,n3374);
and (s1n3373,n2929,n3375);
and (n3376,n3377,n2972);
wire s0n3377,s1n3377,notn3377;
or (n3377,s0n3377,s1n3377);
not(notn3377,n2929);
and (s0n3377,notn3377,n3378);
and (s1n3377,n2929,n3379);
and (n3380,n3381,n2730);
or (n3381,1'b0,n3382,n3386,n3390,n3394);
and (n3382,n3383,n2932);
wire s0n3383,s1n3383,notn3383;
or (n3383,s0n3383,s1n3383);
not(notn3383,n2929);
and (s0n3383,notn3383,n3384);
and (s1n3383,n2929,n3385);
and (n3386,n3387,n2955);
wire s0n3387,s1n3387,notn3387;
or (n3387,s0n3387,s1n3387);
not(notn3387,n2929);
and (s0n3387,notn3387,n3388);
and (s1n3387,n2929,n3389);
and (n3390,n3391,n2963);
wire s0n3391,s1n3391,notn3391;
or (n3391,s0n3391,s1n3391);
not(notn3391,n2929);
and (s0n3391,notn3391,n3392);
and (s1n3391,n2929,n3393);
and (n3394,n3395,n2972);
wire s0n3395,s1n3395,notn3395;
or (n3395,s0n3395,s1n3395);
not(notn3395,n2929);
and (s0n3395,notn3395,n3396);
and (s1n3395,n2929,n3397);
and (n3398,n3399,n2742);
or (n3399,1'b0,n3400,n3404,n3408,n3412);
and (n3400,n3401,n2932);
wire s0n3401,s1n3401,notn3401;
or (n3401,s0n3401,s1n3401);
not(notn3401,n2929);
and (s0n3401,notn3401,n3402);
and (s1n3401,n2929,n3403);
and (n3404,n3405,n2955);
wire s0n3405,s1n3405,notn3405;
or (n3405,s0n3405,s1n3405);
not(notn3405,n2929);
and (s0n3405,notn3405,n3406);
and (s1n3405,n2929,n3407);
and (n3408,n3409,n2963);
wire s0n3409,s1n3409,notn3409;
or (n3409,s0n3409,s1n3409);
not(notn3409,n2929);
and (s0n3409,notn3409,n3410);
and (s1n3409,n2929,n3411);
and (n3412,n3413,n2972);
wire s0n3413,s1n3413,notn3413;
or (n3413,s0n3413,s1n3413);
not(notn3413,n2929);
and (s0n3413,notn3413,n3414);
and (s1n3413,n2929,n3415);
and (n3416,n3417,n2752);
or (n3417,1'b0,n3418,n3422,n3426,n3428);
and (n3418,n3419,n2932);
wire s0n3419,s1n3419,notn3419;
or (n3419,s0n3419,s1n3419);
not(notn3419,n2929);
and (s0n3419,notn3419,n3420);
and (s1n3419,n2929,n3421);
and (n3422,n3423,n2955);
wire s0n3423,s1n3423,notn3423;
or (n3423,s0n3423,s1n3423);
not(notn3423,n2929);
and (s0n3423,notn3423,n3424);
and (s1n3423,n2929,n3425);
and (n3426,n3427,n2963);
wire s0n3427,s1n3427,notn3427;
or (n3427,s0n3427,s1n3427);
not(notn3427,n2929);
and (s0n3427,notn3427,n1315);
and (s1n3427,n2929,n2151);
and (n3428,n3429,n2972);
wire s0n3429,s1n3429,notn3429;
or (n3429,s0n3429,s1n3429);
not(notn3429,n2929);
and (s0n3429,notn3429,n811);
and (s1n3429,n2929,n1769);
or (n3430,1'b0,n3431,n3440,n3446,n3455);
and (n3431,n3432,n2718);
or (n3432,1'b0,n3433,n3437,n3438,n3439);
and (n3433,n3434,n2932);
wire s0n3434,s1n3434,notn3434;
or (n3434,s0n3434,s1n3434);
not(notn3434,n2929);
and (s0n3434,notn3434,n3435);
and (s1n3434,n2929,n3436);
and (n3437,n3365,n2955);
and (n3438,n3369,n2963);
and (n3439,n3373,n2972);
and (n3440,n3441,n2730);
or (n3441,1'b0,n3442,n3443,n3444,n3445);
and (n3442,n3377,n2932);
and (n3443,n3383,n2955);
and (n3444,n3387,n2963);
and (n3445,n3391,n2972);
and (n3446,n3447,n2742);
or (n3447,1'b0,n3448,n3452,n3453,n3454);
and (n3448,n3449,n2932);
wire s0n3449,s1n3449,notn3449;
or (n3449,s0n3449,s1n3449);
not(notn3449,n2929);
and (s0n3449,notn3449,n3450);
and (s1n3449,n2929,n3451);
and (n3452,n3401,n2955);
and (n3453,n3405,n2963);
and (n3454,n3409,n2972);
and (n3455,n3456,n2752);
or (n3456,1'b0,n3457,n3458,n3459,n3460);
and (n3457,n3413,n2932);
and (n3458,n3419,n2955);
and (n3459,n3423,n2963);
and (n3460,n3427,n2972);
and (n3461,n3430,n3462);
or (n3462,n3463,n3564,n3770);
and (n3463,n3464,n3533);
or (n3464,1'b0,n3465,n3483,n3501,n3519);
and (n3465,n3466,n2718);
or (n3466,1'b0,n3467,n3471,n3475,n3479);
and (n3467,n3468,n2932);
wire s0n3468,s1n3468,notn3468;
or (n3468,s0n3468,s1n3468);
not(notn3468,n2929);
and (s0n3468,notn3468,n3469);
and (s1n3468,n2929,n3470);
and (n3471,n3472,n2955);
wire s0n3472,s1n3472,notn3472;
or (n3472,s0n3472,s1n3472);
not(notn3472,n2929);
and (s0n3472,notn3472,n3473);
and (s1n3472,n2929,n3474);
and (n3475,n3476,n2963);
wire s0n3476,s1n3476,notn3476;
or (n3476,s0n3476,s1n3476);
not(notn3476,n2929);
and (s0n3476,notn3476,n3477);
and (s1n3476,n2929,n3478);
and (n3479,n3480,n2972);
wire s0n3480,s1n3480,notn3480;
or (n3480,s0n3480,s1n3480);
not(notn3480,n2929);
and (s0n3480,notn3480,n3481);
and (s1n3480,n2929,n3482);
and (n3483,n3484,n2730);
or (n3484,1'b0,n3485,n3489,n3493,n3497);
and (n3485,n3486,n2932);
wire s0n3486,s1n3486,notn3486;
or (n3486,s0n3486,s1n3486);
not(notn3486,n2929);
and (s0n3486,notn3486,n3487);
and (s1n3486,n2929,n3488);
and (n3489,n3490,n2955);
wire s0n3490,s1n3490,notn3490;
or (n3490,s0n3490,s1n3490);
not(notn3490,n2929);
and (s0n3490,notn3490,n3491);
and (s1n3490,n2929,n3492);
and (n3493,n3494,n2963);
wire s0n3494,s1n3494,notn3494;
or (n3494,s0n3494,s1n3494);
not(notn3494,n2929);
and (s0n3494,notn3494,n3495);
and (s1n3494,n2929,n3496);
and (n3497,n3498,n2972);
wire s0n3498,s1n3498,notn3498;
or (n3498,s0n3498,s1n3498);
not(notn3498,n2929);
and (s0n3498,notn3498,n3499);
and (s1n3498,n2929,n3500);
and (n3501,n3502,n2742);
or (n3502,1'b0,n3503,n3507,n3511,n3515);
and (n3503,n3504,n2932);
wire s0n3504,s1n3504,notn3504;
or (n3504,s0n3504,s1n3504);
not(notn3504,n2929);
and (s0n3504,notn3504,n3505);
and (s1n3504,n2929,n3506);
and (n3507,n3508,n2955);
wire s0n3508,s1n3508,notn3508;
or (n3508,s0n3508,s1n3508);
not(notn3508,n2929);
and (s0n3508,notn3508,n3509);
and (s1n3508,n2929,n3510);
and (n3511,n3512,n2963);
wire s0n3512,s1n3512,notn3512;
or (n3512,s0n3512,s1n3512);
not(notn3512,n2929);
and (s0n3512,notn3512,n3513);
and (s1n3512,n2929,n3514);
and (n3515,n3516,n2972);
wire s0n3516,s1n3516,notn3516;
or (n3516,s0n3516,s1n3516);
not(notn3516,n2929);
and (s0n3516,notn3516,n3517);
and (s1n3516,n2929,n3518);
and (n3519,n3520,n2752);
or (n3520,1'b0,n3521,n3525,n3529,n3531);
and (n3521,n3522,n2932);
wire s0n3522,s1n3522,notn3522;
or (n3522,s0n3522,s1n3522);
not(notn3522,n2929);
and (s0n3522,notn3522,n3523);
and (s1n3522,n2929,n3524);
and (n3525,n3526,n2955);
wire s0n3526,s1n3526,notn3526;
or (n3526,s0n3526,s1n3526);
not(notn3526,n2929);
and (s0n3526,notn3526,n3527);
and (s1n3526,n2929,n3528);
and (n3529,n3530,n2963);
wire s0n3530,s1n3530,notn3530;
or (n3530,s0n3530,s1n3530);
not(notn3530,n2929);
and (s0n3530,notn3530,n1331);
and (s1n3530,n2929,n2167);
and (n3531,n3532,n2972);
wire s0n3532,s1n3532,notn3532;
or (n3532,s0n3532,s1n3532);
not(notn3532,n2929);
and (s0n3532,notn3532,n827);
and (s1n3532,n2929,n1790);
or (n3533,1'b0,n3534,n3543,n3549,n3558);
and (n3534,n3535,n2718);
or (n3535,1'b0,n3536,n3540,n3541,n3542);
and (n3536,n3537,n2932);
wire s0n3537,s1n3537,notn3537;
or (n3537,s0n3537,s1n3537);
not(notn3537,n2929);
and (s0n3537,notn3537,n3538);
and (s1n3537,n2929,n3539);
and (n3540,n3468,n2955);
and (n3541,n3472,n2963);
and (n3542,n3476,n2972);
and (n3543,n3544,n2730);
or (n3544,1'b0,n3545,n3546,n3547,n3548);
and (n3545,n3480,n2932);
and (n3546,n3486,n2955);
and (n3547,n3490,n2963);
and (n3548,n3494,n2972);
and (n3549,n3550,n2742);
or (n3550,1'b0,n3551,n3555,n3556,n3557);
and (n3551,n3552,n2932);
wire s0n3552,s1n3552,notn3552;
or (n3552,s0n3552,s1n3552);
not(notn3552,n2929);
and (s0n3552,notn3552,n3553);
and (s1n3552,n2929,n3554);
and (n3555,n3504,n2955);
and (n3556,n3508,n2963);
and (n3557,n3512,n2972);
and (n3558,n3559,n2752);
or (n3559,1'b0,n3560,n3561,n3562,n3563);
and (n3560,n3516,n2932);
and (n3561,n3522,n2955);
and (n3562,n3526,n2963);
and (n3563,n3530,n2972);
and (n3564,n3533,n3565);
or (n3565,n3566,n3667,n3769);
and (n3566,n3567,n3636);
or (n3567,1'b0,n3568,n3586,n3604,n3622);
and (n3568,n3569,n2718);
or (n3569,1'b0,n3570,n3574,n3578,n3582);
and (n3570,n3571,n2932);
wire s0n3571,s1n3571,notn3571;
or (n3571,s0n3571,s1n3571);
not(notn3571,n2929);
and (s0n3571,notn3571,n3572);
and (s1n3571,n2929,n3573);
and (n3574,n3575,n2955);
wire s0n3575,s1n3575,notn3575;
or (n3575,s0n3575,s1n3575);
not(notn3575,n2929);
and (s0n3575,notn3575,n3576);
and (s1n3575,n2929,n3577);
and (n3578,n3579,n2963);
wire s0n3579,s1n3579,notn3579;
or (n3579,s0n3579,s1n3579);
not(notn3579,n2929);
and (s0n3579,notn3579,n3580);
and (s1n3579,n2929,n3581);
and (n3582,n3583,n2972);
wire s0n3583,s1n3583,notn3583;
or (n3583,s0n3583,s1n3583);
not(notn3583,n2929);
and (s0n3583,notn3583,n3584);
and (s1n3583,n2929,n3585);
and (n3586,n3587,n2730);
or (n3587,1'b0,n3588,n3592,n3596,n3600);
and (n3588,n3589,n2932);
wire s0n3589,s1n3589,notn3589;
or (n3589,s0n3589,s1n3589);
not(notn3589,n2929);
and (s0n3589,notn3589,n3590);
and (s1n3589,n2929,n3591);
and (n3592,n3593,n2955);
wire s0n3593,s1n3593,notn3593;
or (n3593,s0n3593,s1n3593);
not(notn3593,n2929);
and (s0n3593,notn3593,n3594);
and (s1n3593,n2929,n3595);
and (n3596,n3597,n2963);
wire s0n3597,s1n3597,notn3597;
or (n3597,s0n3597,s1n3597);
not(notn3597,n2929);
and (s0n3597,notn3597,n3598);
and (s1n3597,n2929,n3599);
and (n3600,n3601,n2972);
wire s0n3601,s1n3601,notn3601;
or (n3601,s0n3601,s1n3601);
not(notn3601,n2929);
and (s0n3601,notn3601,n3602);
and (s1n3601,n2929,n3603);
and (n3604,n3605,n2742);
or (n3605,1'b0,n3606,n3610,n3614,n3618);
and (n3606,n3607,n2932);
wire s0n3607,s1n3607,notn3607;
or (n3607,s0n3607,s1n3607);
not(notn3607,n2929);
and (s0n3607,notn3607,n3608);
and (s1n3607,n2929,n3609);
and (n3610,n3611,n2955);
wire s0n3611,s1n3611,notn3611;
or (n3611,s0n3611,s1n3611);
not(notn3611,n2929);
and (s0n3611,notn3611,n3612);
and (s1n3611,n2929,n3613);
and (n3614,n3615,n2963);
wire s0n3615,s1n3615,notn3615;
or (n3615,s0n3615,s1n3615);
not(notn3615,n2929);
and (s0n3615,notn3615,n3616);
and (s1n3615,n2929,n3617);
and (n3618,n3619,n2972);
wire s0n3619,s1n3619,notn3619;
or (n3619,s0n3619,s1n3619);
not(notn3619,n2929);
and (s0n3619,notn3619,n3620);
and (s1n3619,n2929,n3621);
and (n3622,n3623,n2752);
or (n3623,1'b0,n3624,n3628,n3632,n3634);
and (n3624,n3625,n2932);
wire s0n3625,s1n3625,notn3625;
or (n3625,s0n3625,s1n3625);
not(notn3625,n2929);
and (s0n3625,notn3625,n3626);
and (s1n3625,n2929,n3627);
and (n3628,n3629,n2955);
wire s0n3629,s1n3629,notn3629;
or (n3629,s0n3629,s1n3629);
not(notn3629,n2929);
and (s0n3629,notn3629,n3630);
and (s1n3629,n2929,n3631);
and (n3632,n3633,n2963);
wire s0n3633,s1n3633,notn3633;
or (n3633,s0n3633,s1n3633);
not(notn3633,n2929);
and (s0n3633,notn3633,n1347);
and (s1n3633,n2929,n2184);
and (n3634,n3635,n2972);
wire s0n3635,s1n3635,notn3635;
or (n3635,s0n3635,s1n3635);
not(notn3635,n2929);
and (s0n3635,notn3635,n843);
and (s1n3635,n2929,n1820);
or (n3636,1'b0,n3637,n3646,n3652,n3661);
and (n3637,n3638,n2718);
or (n3638,1'b0,n3639,n3643,n3644,n3645);
and (n3639,n3640,n2932);
wire s0n3640,s1n3640,notn3640;
or (n3640,s0n3640,s1n3640);
not(notn3640,n2929);
and (s0n3640,notn3640,n3641);
and (s1n3640,n2929,n3642);
and (n3643,n3571,n2955);
and (n3644,n3575,n2963);
and (n3645,n3579,n2972);
and (n3646,n3647,n2730);
or (n3647,1'b0,n3648,n3649,n3650,n3651);
and (n3648,n3583,n2932);
and (n3649,n3589,n2955);
and (n3650,n3593,n2963);
and (n3651,n3597,n2972);
and (n3652,n3653,n2742);
or (n3653,1'b0,n3654,n3658,n3659,n3660);
and (n3654,n3655,n2932);
wire s0n3655,s1n3655,notn3655;
or (n3655,s0n3655,s1n3655);
not(notn3655,n2929);
and (s0n3655,notn3655,n3656);
and (s1n3655,n2929,n3657);
and (n3658,n3607,n2955);
and (n3659,n3611,n2963);
and (n3660,n3615,n2972);
and (n3661,n3662,n2752);
or (n3662,1'b0,n3663,n3664,n3665,n3666);
and (n3663,n3619,n2932);
and (n3664,n3625,n2955);
and (n3665,n3629,n2963);
and (n3666,n3633,n2972);
and (n3667,n3636,n3668);
and (n3668,n3669,n3738);
or (n3669,1'b0,n3670,n3688,n3706,n3724);
and (n3670,n3671,n2718);
or (n3671,1'b0,n3672,n3676,n3680,n3684);
and (n3672,n3673,n2932);
wire s0n3673,s1n3673,notn3673;
or (n3673,s0n3673,s1n3673);
not(notn3673,n2929);
and (s0n3673,notn3673,n3674);
and (s1n3673,n2929,n3675);
and (n3676,n3677,n2955);
wire s0n3677,s1n3677,notn3677;
or (n3677,s0n3677,s1n3677);
not(notn3677,n2929);
and (s0n3677,notn3677,n3678);
and (s1n3677,n2929,n3679);
and (n3680,n3681,n2963);
wire s0n3681,s1n3681,notn3681;
or (n3681,s0n3681,s1n3681);
not(notn3681,n2929);
and (s0n3681,notn3681,n3682);
and (s1n3681,n2929,n3683);
and (n3684,n3685,n2972);
wire s0n3685,s1n3685,notn3685;
or (n3685,s0n3685,s1n3685);
not(notn3685,n2929);
and (s0n3685,notn3685,n3686);
and (s1n3685,n2929,n3687);
and (n3688,n3689,n2730);
or (n3689,1'b0,n3690,n3694,n3698,n3702);
and (n3690,n3691,n2932);
wire s0n3691,s1n3691,notn3691;
or (n3691,s0n3691,s1n3691);
not(notn3691,n2929);
and (s0n3691,notn3691,n3692);
and (s1n3691,n2929,n3693);
and (n3694,n3695,n2955);
wire s0n3695,s1n3695,notn3695;
or (n3695,s0n3695,s1n3695);
not(notn3695,n2929);
and (s0n3695,notn3695,n3696);
and (s1n3695,n2929,n3697);
and (n3698,n3699,n2963);
wire s0n3699,s1n3699,notn3699;
or (n3699,s0n3699,s1n3699);
not(notn3699,n2929);
and (s0n3699,notn3699,n3700);
and (s1n3699,n2929,n3701);
and (n3702,n3703,n2972);
wire s0n3703,s1n3703,notn3703;
or (n3703,s0n3703,s1n3703);
not(notn3703,n2929);
and (s0n3703,notn3703,n3704);
and (s1n3703,n2929,n3705);
and (n3706,n3707,n2742);
or (n3707,1'b0,n3708,n3712,n3716,n3720);
and (n3708,n3709,n2932);
wire s0n3709,s1n3709,notn3709;
or (n3709,s0n3709,s1n3709);
not(notn3709,n2929);
and (s0n3709,notn3709,n3710);
and (s1n3709,n2929,n3711);
and (n3712,n3713,n2955);
wire s0n3713,s1n3713,notn3713;
or (n3713,s0n3713,s1n3713);
not(notn3713,n2929);
and (s0n3713,notn3713,n3714);
and (s1n3713,n2929,n3715);
and (n3716,n3717,n2963);
wire s0n3717,s1n3717,notn3717;
or (n3717,s0n3717,s1n3717);
not(notn3717,n2929);
and (s0n3717,notn3717,n3718);
and (s1n3717,n2929,n3719);
and (n3720,n3721,n2972);
wire s0n3721,s1n3721,notn3721;
or (n3721,s0n3721,s1n3721);
not(notn3721,n2929);
and (s0n3721,notn3721,n3722);
and (s1n3721,n2929,n3723);
and (n3724,n3725,n2752);
or (n3725,1'b0,n3726,n3730,n3734,n3736);
and (n3726,n3727,n2932);
wire s0n3727,s1n3727,notn3727;
or (n3727,s0n3727,s1n3727);
not(notn3727,n2929);
and (s0n3727,notn3727,n3728);
and (s1n3727,n2929,n3729);
and (n3730,n3731,n2955);
wire s0n3731,s1n3731,notn3731;
or (n3731,s0n3731,s1n3731);
not(notn3731,n2929);
and (s0n3731,notn3731,n3732);
and (s1n3731,n2929,n3733);
and (n3734,n3735,n2963);
wire s0n3735,s1n3735,notn3735;
or (n3735,s0n3735,s1n3735);
not(notn3735,n2929);
and (s0n3735,notn3735,n1362);
and (s1n3735,n2929,n2199);
and (n3736,n3737,n2972);
wire s0n3737,s1n3737,notn3737;
or (n3737,s0n3737,s1n3737);
not(notn3737,n2929);
and (s0n3737,notn3737,n858);
and (s1n3737,n2929,n1843);
or (n3738,1'b0,n3739,n3748,n3754,n3763);
and (n3739,n3740,n2718);
or (n3740,1'b0,n3741,n3745,n3746,n3747);
and (n3741,n3742,n2932);
wire s0n3742,s1n3742,notn3742;
or (n3742,s0n3742,s1n3742);
not(notn3742,n2929);
and (s0n3742,notn3742,n3743);
and (s1n3742,n2929,n3744);
and (n3745,n3673,n2955);
and (n3746,n3677,n2963);
and (n3747,n3681,n2972);
and (n3748,n3749,n2730);
or (n3749,1'b0,n3750,n3751,n3752,n3753);
and (n3750,n3685,n2932);
and (n3751,n3691,n2955);
and (n3752,n3695,n2963);
and (n3753,n3699,n2972);
and (n3754,n3755,n2742);
or (n3755,1'b0,n3756,n3760,n3761,n3762);
and (n3756,n3757,n2932);
wire s0n3757,s1n3757,notn3757;
or (n3757,s0n3757,s1n3757);
not(notn3757,n2929);
and (s0n3757,notn3757,n3758);
and (s1n3757,n2929,n3759);
and (n3760,n3709,n2955);
and (n3761,n3713,n2963);
and (n3762,n3717,n2972);
and (n3763,n3764,n2752);
or (n3764,1'b0,n3765,n3766,n3767,n3768);
and (n3765,n3721,n2932);
and (n3766,n3727,n2955);
and (n3767,n3731,n2963);
and (n3768,n3735,n2972);
and (n3769,n3567,n3668);
and (n3770,n3464,n3565);
and (n3771,n3361,n3462);
and (n3772,n3258,n3359);
and (n3773,n3155,n3256);
and (n3774,n3052,n3153);
and (n3775,n2923,n3050);
or (n3776,n3777,n3779);
xor (n3777,n3778,n3050);
xor (n3778,n2923,n3018);
or (n3779,n3780,n4293,n4344);
and (n3780,n3781,n3783);
xor (n3781,n3782,n3153);
xor (n3782,n3052,n3121);
not (n3783,n3784);
or (n3784,n3785,n3846,n4292);
and (n3785,n3786,n3815);
or (n3786,1'b0,n3787,n3793,n3802,n3808);
and (n3787,n3788,n2718);
or (n3788,1'b0,n3789,n3790,n3791,n3792);
and (n3789,n2953,n2932);
and (n3790,n2961,n2955);
and (n3791,n2970,n2963);
and (n3792,n2981,n2972);
and (n3793,n3794,n2730);
or (n3794,1'b0,n3795,n3796,n3797,n3798);
and (n3795,n2984,n2932);
and (n3796,n2987,n2955);
and (n3797,n2990,n2963);
and (n3798,n3799,n2972);
wire s0n3799,s1n3799,notn3799;
or (n3799,s0n3799,s1n3799);
not(notn3799,n2929);
and (s0n3799,notn3799,n3800);
and (s1n3799,n2929,n3801);
and (n3802,n3803,n2742);
or (n3803,1'b0,n3804,n3805,n3806,n3807);
and (n3804,n2998,n2932);
and (n3805,n3001,n2955);
and (n3806,n3004,n2963);
and (n3807,n3009,n2972);
and (n3808,n3809,n2752);
or (n3809,1'b0,n3810,n3811,n3812,n3813);
and (n3810,n3012,n2932);
and (n3811,n3015,n2955);
and (n3812,n3017,n2963);
and (n3813,n3814,n2972);
wire s0n3814,s1n3814,notn3814;
or (n3814,s0n3814,s1n3814);
not(notn3814,n2929);
and (s0n3814,notn3814,n1253);
and (s1n3814,n2929,n2089);
or (n3815,1'b0,n3816,n3825,n3831,n3840);
and (n3816,n3817,n2718);
or (n3817,1'b0,n3818,n3822,n3823,n3824);
and (n3818,n3819,n2932);
wire s0n3819,s1n3819,notn3819;
or (n3819,s0n3819,s1n3819);
not(notn3819,n2929);
and (s0n3819,notn3819,n3820);
and (s1n3819,n2929,n3821);
and (n3822,n3022,n2955);
and (n3823,n2927,n2963);
and (n3824,n2953,n2972);
and (n3825,n3826,n2730);
or (n3826,1'b0,n3827,n3828,n3829,n3830);
and (n3827,n2961,n2932);
and (n3828,n2970,n2955);
and (n3829,n2981,n2963);
and (n3830,n2984,n2972);
and (n3831,n3832,n2742);
or (n3832,1'b0,n3833,n3837,n3838,n3839);
and (n3833,n3834,n2932);
wire s0n3834,s1n3834,notn3834;
or (n3834,s0n3834,s1n3834);
not(notn3834,n2929);
and (s0n3834,notn3834,n3835);
and (s1n3834,n2929,n3836);
and (n3837,n3037,n2955);
and (n3838,n2995,n2963);
and (n3839,n2998,n2972);
and (n3840,n3841,n2752);
or (n3841,1'b0,n3842,n3843,n3844,n3845);
and (n3842,n3001,n2932);
and (n3843,n3004,n2955);
and (n3844,n3009,n2963);
and (n3845,n3012,n2972);
and (n3846,n3815,n3847);
or (n3847,n3848,n3909,n4291);
and (n3848,n3849,n3878);
or (n3849,1'b0,n3850,n3856,n3865,n3871);
and (n3850,n3851,n2718);
or (n3851,1'b0,n3852,n3853,n3854,n3855);
and (n3852,n3060,n2932);
and (n3853,n3064,n2955);
and (n3854,n3068,n2963);
and (n3855,n3074,n2972);
and (n3856,n3857,n2730);
or (n3857,1'b0,n3858,n3859,n3860,n3861);
and (n3858,n3078,n2932);
and (n3859,n3082,n2955);
and (n3860,n3086,n2963);
and (n3861,n3862,n2972);
wire s0n3862,s1n3862,notn3862;
or (n3862,s0n3862,s1n3862);
not(notn3862,n2929);
and (s0n3862,notn3862,n3863);
and (s1n3862,n2929,n3864);
and (n3865,n3866,n2742);
or (n3866,1'b0,n3867,n3868,n3869,n3870);
and (n3867,n3096,n2932);
and (n3868,n3100,n2955);
and (n3869,n3104,n2963);
and (n3870,n3110,n2972);
and (n3871,n3872,n2752);
or (n3872,1'b0,n3873,n3874,n3875,n3876);
and (n3873,n3114,n2932);
and (n3874,n3118,n2955);
and (n3875,n3120,n2963);
and (n3876,n3877,n2972);
wire s0n3877,s1n3877,notn3877;
or (n3877,s0n3877,s1n3877);
not(notn3877,n2929);
and (s0n3877,notn3877,n1269);
and (s1n3877,n2929,n2105);
or (n3878,1'b0,n3879,n3888,n3894,n3903);
and (n3879,n3880,n2718);
or (n3880,1'b0,n3881,n3885,n3886,n3887);
and (n3881,n3882,n2932);
wire s0n3882,s1n3882,notn3882;
or (n3882,s0n3882,s1n3882);
not(notn3882,n2929);
and (s0n3882,notn3882,n3883);
and (s1n3882,n2929,n3884);
and (n3885,n3125,n2955);
and (n3886,n3056,n2963);
and (n3887,n3060,n2972);
and (n3888,n3889,n2730);
or (n3889,1'b0,n3890,n3891,n3892,n3893);
and (n3890,n3064,n2932);
and (n3891,n3068,n2955);
and (n3892,n3074,n2963);
and (n3893,n3078,n2972);
and (n3894,n3895,n2742);
or (n3895,1'b0,n3896,n3900,n3901,n3902);
and (n3896,n3897,n2932);
wire s0n3897,s1n3897,notn3897;
or (n3897,s0n3897,s1n3897);
not(notn3897,n2929);
and (s0n3897,notn3897,n3898);
and (s1n3897,n2929,n3899);
and (n3900,n3140,n2955);
and (n3901,n3092,n2963);
and (n3902,n3096,n2972);
and (n3903,n3904,n2752);
or (n3904,1'b0,n3905,n3906,n3907,n3908);
and (n3905,n3100,n2932);
and (n3906,n3104,n2955);
and (n3907,n3110,n2963);
and (n3908,n3114,n2972);
and (n3909,n3878,n3910);
or (n3910,n3911,n3972,n4290);
and (n3911,n3912,n3941);
or (n3912,1'b0,n3913,n3919,n3928,n3934);
and (n3913,n3914,n2718);
or (n3914,1'b0,n3915,n3916,n3917,n3918);
and (n3915,n3163,n2932);
and (n3916,n3167,n2955);
and (n3917,n3171,n2963);
and (n3918,n3177,n2972);
and (n3919,n3920,n2730);
or (n3920,1'b0,n3921,n3922,n3923,n3924);
and (n3921,n3181,n2932);
and (n3922,n3185,n2955);
and (n3923,n3189,n2963);
and (n3924,n3925,n2972);
wire s0n3925,s1n3925,notn3925;
or (n3925,s0n3925,s1n3925);
not(notn3925,n2929);
and (s0n3925,notn3925,n3926);
and (s1n3925,n2929,n3927);
and (n3928,n3929,n2742);
or (n3929,1'b0,n3930,n3931,n3932,n3933);
and (n3930,n3199,n2932);
and (n3931,n3203,n2955);
and (n3932,n3207,n2963);
and (n3933,n3213,n2972);
and (n3934,n3935,n2752);
or (n3935,1'b0,n3936,n3937,n3938,n3939);
and (n3936,n3217,n2932);
and (n3937,n3221,n2955);
and (n3938,n3223,n2963);
and (n3939,n3940,n2972);
wire s0n3940,s1n3940,notn3940;
or (n3940,s0n3940,s1n3940);
not(notn3940,n2929);
and (s0n3940,notn3940,n1285);
and (s1n3940,n2929,n2121);
or (n3941,1'b0,n3942,n3951,n3957,n3966);
and (n3942,n3943,n2718);
or (n3943,1'b0,n3944,n3948,n3949,n3950);
and (n3944,n3945,n2932);
wire s0n3945,s1n3945,notn3945;
or (n3945,s0n3945,s1n3945);
not(notn3945,n2929);
and (s0n3945,notn3945,n3946);
and (s1n3945,n2929,n3947);
and (n3948,n3228,n2955);
and (n3949,n3159,n2963);
and (n3950,n3163,n2972);
and (n3951,n3952,n2730);
or (n3952,1'b0,n3953,n3954,n3955,n3956);
and (n3953,n3167,n2932);
and (n3954,n3171,n2955);
and (n3955,n3177,n2963);
and (n3956,n3181,n2972);
and (n3957,n3958,n2742);
or (n3958,1'b0,n3959,n3963,n3964,n3965);
and (n3959,n3960,n2932);
wire s0n3960,s1n3960,notn3960;
or (n3960,s0n3960,s1n3960);
not(notn3960,n2929);
and (s0n3960,notn3960,n3961);
and (s1n3960,n2929,n3962);
and (n3963,n3243,n2955);
and (n3964,n3195,n2963);
and (n3965,n3199,n2972);
and (n3966,n3967,n2752);
or (n3967,1'b0,n3968,n3969,n3970,n3971);
and (n3968,n3203,n2932);
and (n3969,n3207,n2955);
and (n3970,n3213,n2963);
and (n3971,n3217,n2972);
and (n3972,n3941,n3973);
or (n3973,n3974,n4035,n4289);
and (n3974,n3975,n4004);
or (n3975,1'b0,n3976,n3982,n3991,n3997);
and (n3976,n3977,n2718);
or (n3977,1'b0,n3978,n3979,n3980,n3981);
and (n3978,n3266,n2932);
and (n3979,n3270,n2955);
and (n3980,n3274,n2963);
and (n3981,n3280,n2972);
and (n3982,n3983,n2730);
or (n3983,1'b0,n3984,n3985,n3986,n3987);
and (n3984,n3284,n2932);
and (n3985,n3288,n2955);
and (n3986,n3292,n2963);
and (n3987,n3988,n2972);
wire s0n3988,s1n3988,notn3988;
or (n3988,s0n3988,s1n3988);
not(notn3988,n2929);
and (s0n3988,notn3988,n3989);
and (s1n3988,n2929,n3990);
and (n3991,n3992,n2742);
or (n3992,1'b0,n3993,n3994,n3995,n3996);
and (n3993,n3302,n2932);
and (n3994,n3306,n2955);
and (n3995,n3310,n2963);
and (n3996,n3316,n2972);
and (n3997,n3998,n2752);
or (n3998,1'b0,n3999,n4000,n4001,n4002);
and (n3999,n3320,n2932);
and (n4000,n3324,n2955);
and (n4001,n3326,n2963);
and (n4002,n4003,n2972);
wire s0n4003,s1n4003,notn4003;
or (n4003,s0n4003,s1n4003);
not(notn4003,n2929);
and (s0n4003,notn4003,n1301);
and (s1n4003,n2929,n2137);
or (n4004,1'b0,n4005,n4014,n4020,n4029);
and (n4005,n4006,n2718);
or (n4006,1'b0,n4007,n4011,n4012,n4013);
and (n4007,n4008,n2932);
wire s0n4008,s1n4008,notn4008;
or (n4008,s0n4008,s1n4008);
not(notn4008,n2929);
and (s0n4008,notn4008,n4009);
and (s1n4008,n2929,n4010);
and (n4011,n3331,n2955);
and (n4012,n3262,n2963);
and (n4013,n3266,n2972);
and (n4014,n4015,n2730);
or (n4015,1'b0,n4016,n4017,n4018,n4019);
and (n4016,n3270,n2932);
and (n4017,n3274,n2955);
and (n4018,n3280,n2963);
and (n4019,n3284,n2972);
and (n4020,n4021,n2742);
or (n4021,1'b0,n4022,n4026,n4027,n4028);
and (n4022,n4023,n2932);
wire s0n4023,s1n4023,notn4023;
or (n4023,s0n4023,s1n4023);
not(notn4023,n2929);
and (s0n4023,notn4023,n4024);
and (s1n4023,n2929,n4025);
and (n4026,n3346,n2955);
and (n4027,n3298,n2963);
and (n4028,n3302,n2972);
and (n4029,n4030,n2752);
or (n4030,1'b0,n4031,n4032,n4033,n4034);
and (n4031,n3306,n2932);
and (n4032,n3310,n2955);
and (n4033,n3316,n2963);
and (n4034,n3320,n2972);
and (n4035,n4004,n4036);
or (n4036,n4037,n4098,n4288);
and (n4037,n4038,n4067);
or (n4038,1'b0,n4039,n4045,n4054,n4060);
and (n4039,n4040,n2718);
or (n4040,1'b0,n4041,n4042,n4043,n4044);
and (n4041,n3369,n2932);
and (n4042,n3373,n2955);
and (n4043,n3377,n2963);
and (n4044,n3383,n2972);
and (n4045,n4046,n2730);
or (n4046,1'b0,n4047,n4048,n4049,n4050);
and (n4047,n3387,n2932);
and (n4048,n3391,n2955);
and (n4049,n3395,n2963);
and (n4050,n4051,n2972);
wire s0n4051,s1n4051,notn4051;
or (n4051,s0n4051,s1n4051);
not(notn4051,n2929);
and (s0n4051,notn4051,n4052);
and (s1n4051,n2929,n4053);
and (n4054,n4055,n2742);
or (n4055,1'b0,n4056,n4057,n4058,n4059);
and (n4056,n3405,n2932);
and (n4057,n3409,n2955);
and (n4058,n3413,n2963);
and (n4059,n3419,n2972);
and (n4060,n4061,n2752);
or (n4061,1'b0,n4062,n4063,n4064,n4065);
and (n4062,n3423,n2932);
and (n4063,n3427,n2955);
and (n4064,n3429,n2963);
and (n4065,n4066,n2972);
wire s0n4066,s1n4066,notn4066;
or (n4066,s0n4066,s1n4066);
not(notn4066,n2929);
and (s0n4066,notn4066,n1317);
and (s1n4066,n2929,n2153);
or (n4067,1'b0,n4068,n4077,n4083,n4092);
and (n4068,n4069,n2718);
or (n4069,1'b0,n4070,n4074,n4075,n4076);
and (n4070,n4071,n2932);
wire s0n4071,s1n4071,notn4071;
or (n4071,s0n4071,s1n4071);
not(notn4071,n2929);
and (s0n4071,notn4071,n4072);
and (s1n4071,n2929,n4073);
and (n4074,n3434,n2955);
and (n4075,n3365,n2963);
and (n4076,n3369,n2972);
and (n4077,n4078,n2730);
or (n4078,1'b0,n4079,n4080,n4081,n4082);
and (n4079,n3373,n2932);
and (n4080,n3377,n2955);
and (n4081,n3383,n2963);
and (n4082,n3387,n2972);
and (n4083,n4084,n2742);
or (n4084,1'b0,n4085,n4089,n4090,n4091);
and (n4085,n4086,n2932);
wire s0n4086,s1n4086,notn4086;
or (n4086,s0n4086,s1n4086);
not(notn4086,n2929);
and (s0n4086,notn4086,n4087);
and (s1n4086,n2929,n4088);
and (n4089,n3449,n2955);
and (n4090,n3401,n2963);
and (n4091,n3405,n2972);
and (n4092,n4093,n2752);
or (n4093,1'b0,n4094,n4095,n4096,n4097);
and (n4094,n3409,n2932);
and (n4095,n3413,n2955);
and (n4096,n3419,n2963);
and (n4097,n3423,n2972);
and (n4098,n4067,n4099);
or (n4099,n4100,n4161,n4287);
and (n4100,n4101,n4130);
or (n4101,1'b0,n4102,n4108,n4117,n4123);
and (n4102,n4103,n2718);
or (n4103,1'b0,n4104,n4105,n4106,n4107);
and (n4104,n3472,n2932);
and (n4105,n3476,n2955);
and (n4106,n3480,n2963);
and (n4107,n3486,n2972);
and (n4108,n4109,n2730);
or (n4109,1'b0,n4110,n4111,n4112,n4113);
and (n4110,n3490,n2932);
and (n4111,n3494,n2955);
and (n4112,n3498,n2963);
and (n4113,n4114,n2972);
wire s0n4114,s1n4114,notn4114;
or (n4114,s0n4114,s1n4114);
not(notn4114,n2929);
and (s0n4114,notn4114,n4115);
and (s1n4114,n2929,n4116);
and (n4117,n4118,n2742);
or (n4118,1'b0,n4119,n4120,n4121,n4122);
and (n4119,n3508,n2932);
and (n4120,n3512,n2955);
and (n4121,n3516,n2963);
and (n4122,n3522,n2972);
and (n4123,n4124,n2752);
or (n4124,1'b0,n4125,n4126,n4127,n4128);
and (n4125,n3526,n2932);
and (n4126,n3530,n2955);
and (n4127,n3532,n2963);
and (n4128,n4129,n2972);
wire s0n4129,s1n4129,notn4129;
or (n4129,s0n4129,s1n4129);
not(notn4129,n2929);
and (s0n4129,notn4129,n1333);
and (s1n4129,n2929,n2169);
or (n4130,1'b0,n4131,n4140,n4146,n4155);
and (n4131,n4132,n2718);
or (n4132,1'b0,n4133,n4137,n4138,n4139);
and (n4133,n4134,n2932);
wire s0n4134,s1n4134,notn4134;
or (n4134,s0n4134,s1n4134);
not(notn4134,n2929);
and (s0n4134,notn4134,n4135);
and (s1n4134,n2929,n4136);
and (n4137,n3537,n2955);
and (n4138,n3468,n2963);
and (n4139,n3472,n2972);
and (n4140,n4141,n2730);
or (n4141,1'b0,n4142,n4143,n4144,n4145);
and (n4142,n3476,n2932);
and (n4143,n3480,n2955);
and (n4144,n3486,n2963);
and (n4145,n3490,n2972);
and (n4146,n4147,n2742);
or (n4147,1'b0,n4148,n4152,n4153,n4154);
and (n4148,n4149,n2932);
wire s0n4149,s1n4149,notn4149;
or (n4149,s0n4149,s1n4149);
not(notn4149,n2929);
and (s0n4149,notn4149,n4150);
and (s1n4149,n2929,n4151);
and (n4152,n3552,n2955);
and (n4153,n3504,n2963);
and (n4154,n3508,n2972);
and (n4155,n4156,n2752);
or (n4156,1'b0,n4157,n4158,n4159,n4160);
and (n4157,n3512,n2932);
and (n4158,n3516,n2955);
and (n4159,n3522,n2963);
and (n4160,n3526,n2972);
and (n4161,n4130,n4162);
or (n4162,n4163,n4224,n4286);
and (n4163,n4164,n4193);
or (n4164,1'b0,n4165,n4171,n4180,n4186);
and (n4165,n4166,n2718);
or (n4166,1'b0,n4167,n4168,n4169,n4170);
and (n4167,n3575,n2932);
and (n4168,n3579,n2955);
and (n4169,n3583,n2963);
and (n4170,n3589,n2972);
and (n4171,n4172,n2730);
or (n4172,1'b0,n4173,n4174,n4175,n4176);
and (n4173,n3593,n2932);
and (n4174,n3597,n2955);
and (n4175,n3601,n2963);
and (n4176,n4177,n2972);
wire s0n4177,s1n4177,notn4177;
or (n4177,s0n4177,s1n4177);
not(notn4177,n2929);
and (s0n4177,notn4177,n4178);
and (s1n4177,n2929,n4179);
and (n4180,n4181,n2742);
or (n4181,1'b0,n4182,n4183,n4184,n4185);
and (n4182,n3611,n2932);
and (n4183,n3615,n2955);
and (n4184,n3619,n2963);
and (n4185,n3625,n2972);
and (n4186,n4187,n2752);
or (n4187,1'b0,n4188,n4189,n4190,n4191);
and (n4188,n3629,n2932);
and (n4189,n3633,n2955);
and (n4190,n3635,n2963);
and (n4191,n4192,n2972);
wire s0n4192,s1n4192,notn4192;
or (n4192,s0n4192,s1n4192);
not(notn4192,n2929);
and (s0n4192,notn4192,n1349);
and (s1n4192,n2929,n2186);
or (n4193,1'b0,n4194,n4203,n4209,n4218);
and (n4194,n4195,n2718);
or (n4195,1'b0,n4196,n4200,n4201,n4202);
and (n4196,n4197,n2932);
wire s0n4197,s1n4197,notn4197;
or (n4197,s0n4197,s1n4197);
not(notn4197,n2929);
and (s0n4197,notn4197,n4198);
and (s1n4197,n2929,n4199);
and (n4200,n3640,n2955);
and (n4201,n3571,n2963);
and (n4202,n3575,n2972);
and (n4203,n4204,n2730);
or (n4204,1'b0,n4205,n4206,n4207,n4208);
and (n4205,n3579,n2932);
and (n4206,n3583,n2955);
and (n4207,n3589,n2963);
and (n4208,n3593,n2972);
and (n4209,n4210,n2742);
or (n4210,1'b0,n4211,n4215,n4216,n4217);
and (n4211,n4212,n2932);
wire s0n4212,s1n4212,notn4212;
or (n4212,s0n4212,s1n4212);
not(notn4212,n2929);
and (s0n4212,notn4212,n4213);
and (s1n4212,n2929,n4214);
and (n4215,n3655,n2955);
and (n4216,n3607,n2963);
and (n4217,n3611,n2972);
and (n4218,n4219,n2752);
or (n4219,1'b0,n4220,n4221,n4222,n4223);
and (n4220,n3615,n2932);
and (n4221,n3619,n2955);
and (n4222,n3625,n2963);
and (n4223,n3629,n2972);
and (n4224,n4193,n4225);
and (n4225,n4226,n4255);
or (n4226,1'b0,n4227,n4233,n4242,n4248);
and (n4227,n4228,n2718);
or (n4228,1'b0,n4229,n4230,n4231,n4232);
and (n4229,n3677,n2932);
and (n4230,n3681,n2955);
and (n4231,n3685,n2963);
and (n4232,n3691,n2972);
and (n4233,n4234,n2730);
or (n4234,1'b0,n4235,n4236,n4237,n4238);
and (n4235,n3695,n2932);
and (n4236,n3699,n2955);
and (n4237,n3703,n2963);
and (n4238,n4239,n2972);
wire s0n4239,s1n4239,notn4239;
or (n4239,s0n4239,s1n4239);
not(notn4239,n2929);
and (s0n4239,notn4239,n4240);
and (s1n4239,n2929,n4241);
and (n4242,n4243,n2742);
or (n4243,1'b0,n4244,n4245,n4246,n4247);
and (n4244,n3713,n2932);
and (n4245,n3717,n2955);
and (n4246,n3721,n2963);
and (n4247,n3727,n2972);
and (n4248,n4249,n2752);
or (n4249,1'b0,n4250,n4251,n4252,n4253);
and (n4250,n3731,n2932);
and (n4251,n3735,n2955);
and (n4252,n3737,n2963);
and (n4253,n4254,n2972);
wire s0n4254,s1n4254,notn4254;
or (n4254,s0n4254,s1n4254);
not(notn4254,n2929);
and (s0n4254,notn4254,n1364);
and (s1n4254,n2929,n2201);
or (n4255,1'b0,n4256,n4265,n4271,n4280);
and (n4256,n4257,n2718);
or (n4257,1'b0,n4258,n4262,n4263,n4264);
and (n4258,n4259,n2932);
wire s0n4259,s1n4259,notn4259;
or (n4259,s0n4259,s1n4259);
not(notn4259,n2929);
and (s0n4259,notn4259,n4260);
and (s1n4259,n2929,n4261);
and (n4262,n3742,n2955);
and (n4263,n3673,n2963);
and (n4264,n3677,n2972);
and (n4265,n4266,n2730);
or (n4266,1'b0,n4267,n4268,n4269,n4270);
and (n4267,n3681,n2932);
and (n4268,n3685,n2955);
and (n4269,n3691,n2963);
and (n4270,n3695,n2972);
and (n4271,n4272,n2742);
or (n4272,1'b0,n4273,n4277,n4278,n4279);
and (n4273,n4274,n2932);
wire s0n4274,s1n4274,notn4274;
or (n4274,s0n4274,s1n4274);
not(notn4274,n2929);
and (s0n4274,notn4274,n4275);
and (s1n4274,n2929,n4276);
and (n4277,n3757,n2955);
and (n4278,n3709,n2963);
and (n4279,n3713,n2972);
and (n4280,n4281,n2752);
or (n4281,1'b0,n4282,n4283,n4284,n4285);
and (n4282,n3717,n2932);
and (n4283,n3721,n2955);
and (n4284,n3727,n2963);
and (n4285,n3731,n2972);
and (n4286,n4164,n4225);
and (n4287,n4101,n4162);
and (n4288,n4038,n4099);
and (n4289,n3975,n4036);
and (n4290,n3912,n3973);
and (n4291,n3849,n3910);
and (n4292,n3786,n3847);
and (n4293,n3783,n4294);
or (n4294,n4295,n4301,n4343);
and (n4295,n4296,n4298);
xor (n4296,n4297,n3256);
xor (n4297,n3155,n3224);
not (n4298,n4299);
xor (n4299,n4300,n3847);
xor (n4300,n3786,n3815);
and (n4301,n4298,n4302);
or (n4302,n4303,n4309,n4342);
and (n4303,n4304,n4306);
xor (n4304,n4305,n3359);
xor (n4305,n3258,n3327);
not (n4306,n4307);
xor (n4307,n4308,n3910);
xor (n4308,n3849,n3878);
and (n4309,n4306,n4310);
or (n4310,n4311,n4317,n4341);
and (n4311,n4312,n4314);
xor (n4312,n4313,n3462);
xor (n4313,n3361,n3430);
not (n4314,n4315);
xor (n4315,n4316,n3973);
xor (n4316,n3912,n3941);
and (n4317,n4314,n4318);
or (n4318,n4319,n4325,n4340);
and (n4319,n4320,n4322);
xor (n4320,n4321,n3565);
xor (n4321,n3464,n3533);
not (n4322,n4323);
xor (n4323,n4324,n4036);
xor (n4324,n3975,n4004);
and (n4325,n4322,n4326);
or (n4326,n4327,n4333,n4339);
and (n4327,n4328,n4330);
xor (n4328,n4329,n3668);
xor (n4329,n3567,n3636);
not (n4330,n4331);
xor (n4331,n4332,n4099);
xor (n4332,n4038,n4067);
and (n4333,n4330,n4334);
and (n4334,n4335,n4336);
xor (n4335,n3669,n3738);
not (n4336,n4337);
xor (n4337,n4338,n4162);
xor (n4338,n4101,n4130);
and (n4339,n4328,n4334);
and (n4340,n4320,n4326);
and (n4341,n4312,n4318);
and (n4342,n4304,n4310);
and (n4343,n4296,n4302);
and (n4344,n3781,n4294);
and (n4345,n4346,n4347);
xnor (n4346,n2921,n3776);
and (n4347,n4348,n4349);
xnor (n4348,n3777,n3779);
and (n4349,n4350,n4352);
xor (n4350,n4351,n4294);
xor (n4351,n3781,n3783);
and (n4352,n4353,n4355);
xor (n4353,n4354,n4302);
xor (n4354,n4296,n4298);
and (n4355,n4356,n4358);
xor (n4356,n4357,n4310);
xor (n4357,n4304,n4306);
and (n4358,n4359,n4361);
xor (n4359,n4360,n4318);
xor (n4360,n4312,n4314);
and (n4361,n4362,n4364);
xor (n4362,n4363,n4326);
xor (n4363,n4320,n4322);
and (n4364,n4365,n4367);
xor (n4365,n4366,n4334);
xor (n4366,n4328,n4330);
and (n4367,n4368,n4369);
xor (n4368,n4335,n4336);
and (n4369,n4370,n4373);
not (n4370,n4371);
xor (n4371,n4372,n4225);
xor (n4372,n4164,n4193);
not (n4373,n4374);
xor (n4374,n4226,n4255);
and (n4375,n2918,n4376);
and (n4376,n4377,n4378);
xor (n4377,n4346,n4347);
and (n4378,n4379,n4380);
xor (n4379,n4348,n4349);
or (n4380,n4381,n4732,n4784);
and (n4381,n4382,n4731);
or (n4382,n4383,n4424,n4730);
and (n4383,n4384,n4403);
or (n4384,1'b0,n4385,n4386,n4395,n4396);
and (n4385,n3826,n2718);
and (n4386,n4387,n2730);
or (n4387,1'b0,n4388,n4389,n4390,n4391);
and (n4388,n2987,n2932);
and (n4389,n2990,n2955);
and (n4390,n3799,n2963);
and (n4391,n4392,n2972);
wire s0n4392,s1n4392,notn4392;
or (n4392,s0n4392,s1n4392);
not(notn4392,n2929);
and (s0n4392,notn4392,n4393);
and (s1n4392,n2929,n4394);
and (n4395,n3841,n2742);
and (n4396,n4397,n2752);
or (n4397,1'b0,n4398,n4399,n4400,n4401);
and (n4398,n3015,n2932);
and (n4399,n3017,n2955);
and (n4400,n3814,n2963);
and (n4401,n4402,n2972);
wire s0n4402,s1n4402,notn4402;
or (n4402,s0n4402,s1n4402);
not(notn4402,n2929);
and (s0n4402,notn4402,n566);
and (s1n4402,n2929,n1694);
or (n4403,1'b0,n4404,n4413,n4414,n4423);
and (n4404,n4405,n2718);
or (n4405,1'b0,n4406,n4410,n4411,n4412);
and (n4406,n4407,n2932);
wire s0n4407,s1n4407,notn4407;
or (n4407,s0n4407,s1n4407);
not(notn4407,n2929);
and (s0n4407,notn4407,n4408);
and (s1n4407,n2929,n4409);
and (n4410,n3819,n2955);
and (n4411,n3022,n2963);
and (n4412,n2927,n2972);
and (n4413,n3788,n2730);
and (n4414,n4415,n2742);
or (n4415,1'b0,n4416,n4420,n4421,n4422);
and (n4416,n4417,n2932);
wire s0n4417,s1n4417,notn4417;
or (n4417,s0n4417,s1n4417);
not(notn4417,n2929);
and (s0n4417,notn4417,n4418);
and (s1n4417,n2929,n4419);
and (n4420,n3834,n2955);
and (n4421,n3037,n2963);
and (n4422,n2995,n2972);
and (n4423,n3803,n2752);
and (n4424,n4403,n4425);
or (n4425,n4426,n4467,n4729);
and (n4426,n4427,n4446);
or (n4427,1'b0,n4428,n4429,n4438,n4439);
and (n4428,n3889,n2718);
and (n4429,n4430,n2730);
or (n4430,1'b0,n4431,n4432,n4433,n4434);
and (n4431,n3082,n2932);
and (n4432,n3086,n2955);
and (n4433,n3862,n2963);
and (n4434,n4435,n2972);
wire s0n4435,s1n4435,notn4435;
or (n4435,s0n4435,s1n4435);
not(notn4435,n2929);
and (s0n4435,notn4435,n4436);
and (s1n4435,n2929,n4437);
and (n4438,n3904,n2742);
and (n4439,n4440,n2752);
or (n4440,1'b0,n4441,n4442,n4443,n4444);
and (n4441,n3118,n2932);
and (n4442,n3120,n2955);
and (n4443,n3877,n2963);
and (n4444,n4445,n2972);
wire s0n4445,s1n4445,notn4445;
or (n4445,s0n4445,s1n4445);
not(notn4445,n2929);
and (s0n4445,notn4445,n757);
and (s1n4445,n2929,n1710);
or (n4446,1'b0,n4447,n4456,n4457,n4466);
and (n4447,n4448,n2718);
or (n4448,1'b0,n4449,n4453,n4454,n4455);
and (n4449,n4450,n2932);
wire s0n4450,s1n4450,notn4450;
or (n4450,s0n4450,s1n4450);
not(notn4450,n2929);
and (s0n4450,notn4450,n4451);
and (s1n4450,n2929,n4452);
and (n4453,n3882,n2955);
and (n4454,n3125,n2963);
and (n4455,n3056,n2972);
and (n4456,n3851,n2730);
and (n4457,n4458,n2742);
or (n4458,1'b0,n4459,n4463,n4464,n4465);
and (n4459,n4460,n2932);
wire s0n4460,s1n4460,notn4460;
or (n4460,s0n4460,s1n4460);
not(notn4460,n2929);
and (s0n4460,notn4460,n4461);
and (s1n4460,n2929,n4462);
and (n4463,n3897,n2955);
and (n4464,n3140,n2963);
and (n4465,n3092,n2972);
and (n4466,n3866,n2752);
and (n4467,n4446,n4468);
or (n4468,n4469,n4510,n4728);
and (n4469,n4470,n4489);
or (n4470,1'b0,n4471,n4472,n4481,n4482);
and (n4471,n3952,n2718);
and (n4472,n4473,n2730);
or (n4473,1'b0,n4474,n4475,n4476,n4477);
and (n4474,n3185,n2932);
and (n4475,n3189,n2955);
and (n4476,n3925,n2963);
and (n4477,n4478,n2972);
wire s0n4478,s1n4478,notn4478;
or (n4478,s0n4478,s1n4478);
not(notn4478,n2929);
and (s0n4478,notn4478,n4479);
and (s1n4478,n2929,n4480);
and (n4481,n3967,n2742);
and (n4482,n4483,n2752);
or (n4483,1'b0,n4484,n4485,n4486,n4487);
and (n4484,n3221,n2932);
and (n4485,n3223,n2955);
and (n4486,n3940,n2963);
and (n4487,n4488,n2972);
wire s0n4488,s1n4488,notn4488;
or (n4488,s0n4488,s1n4488);
not(notn4488,n2929);
and (s0n4488,notn4488,n781);
and (s1n4488,n2929,n1729);
or (n4489,1'b0,n4490,n4499,n4500,n4509);
and (n4490,n4491,n2718);
or (n4491,1'b0,n4492,n4496,n4497,n4498);
and (n4492,n4493,n2932);
wire s0n4493,s1n4493,notn4493;
or (n4493,s0n4493,s1n4493);
not(notn4493,n2929);
and (s0n4493,notn4493,n4494);
and (s1n4493,n2929,n4495);
and (n4496,n3945,n2955);
and (n4497,n3228,n2963);
and (n4498,n3159,n2972);
and (n4499,n3914,n2730);
and (n4500,n4501,n2742);
or (n4501,1'b0,n4502,n4506,n4507,n4508);
and (n4502,n4503,n2932);
wire s0n4503,s1n4503,notn4503;
or (n4503,s0n4503,s1n4503);
not(notn4503,n2929);
and (s0n4503,notn4503,n4504);
and (s1n4503,n2929,n4505);
and (n4506,n3960,n2955);
and (n4507,n3243,n2963);
and (n4508,n3195,n2972);
and (n4509,n3929,n2752);
and (n4510,n4489,n4511);
or (n4511,n4512,n4553,n4727);
and (n4512,n4513,n4532);
or (n4513,1'b0,n4514,n4515,n4524,n4525);
and (n4514,n4015,n2718);
and (n4515,n4516,n2730);
or (n4516,1'b0,n4517,n4518,n4519,n4520);
and (n4517,n3288,n2932);
and (n4518,n3292,n2955);
and (n4519,n3988,n2963);
and (n4520,n4521,n2972);
wire s0n4521,s1n4521,notn4521;
or (n4521,s0n4521,s1n4521);
not(notn4521,n2929);
and (s0n4521,notn4521,n4522);
and (s1n4521,n2929,n4523);
and (n4524,n4030,n2742);
and (n4525,n4526,n2752);
or (n4526,1'b0,n4527,n4528,n4529,n4530);
and (n4527,n3324,n2932);
and (n4528,n3326,n2955);
and (n4529,n4003,n2963);
and (n4530,n4531,n2972);
wire s0n4531,s1n4531,notn4531;
or (n4531,s0n4531,s1n4531);
not(notn4531,n2929);
and (s0n4531,notn4531,n797);
and (s1n4531,n2929,n1755);
or (n4532,1'b0,n4533,n4542,n4543,n4552);
and (n4533,n4534,n2718);
or (n4534,1'b0,n4535,n4539,n4540,n4541);
and (n4535,n4536,n2932);
wire s0n4536,s1n4536,notn4536;
or (n4536,s0n4536,s1n4536);
not(notn4536,n2929);
and (s0n4536,notn4536,n4537);
and (s1n4536,n2929,n4538);
and (n4539,n4008,n2955);
and (n4540,n3331,n2963);
and (n4541,n3262,n2972);
and (n4542,n3977,n2730);
and (n4543,n4544,n2742);
or (n4544,1'b0,n4545,n4549,n4550,n4551);
and (n4545,n4546,n2932);
wire s0n4546,s1n4546,notn4546;
or (n4546,s0n4546,s1n4546);
not(notn4546,n2929);
and (s0n4546,notn4546,n4547);
and (s1n4546,n2929,n4548);
and (n4549,n4023,n2955);
and (n4550,n3346,n2963);
and (n4551,n3298,n2972);
and (n4552,n3992,n2752);
and (n4553,n4532,n4554);
or (n4554,n4555,n4596,n4726);
and (n4555,n4556,n4575);
or (n4556,1'b0,n4557,n4558,n4567,n4568);
and (n4557,n4078,n2718);
and (n4558,n4559,n2730);
or (n4559,1'b0,n4560,n4561,n4562,n4563);
and (n4560,n3391,n2932);
and (n4561,n3395,n2955);
and (n4562,n4051,n2963);
and (n4563,n4564,n2972);
wire s0n4564,s1n4564,notn4564;
or (n4564,s0n4564,s1n4564);
not(notn4564,n2929);
and (s0n4564,notn4564,n4565);
and (s1n4564,n2929,n4566);
and (n4567,n4093,n2742);
and (n4568,n4569,n2752);
or (n4569,1'b0,n4570,n4571,n4572,n4573);
and (n4570,n3427,n2932);
and (n4571,n3429,n2955);
and (n4572,n4066,n2963);
and (n4573,n4574,n2972);
wire s0n4574,s1n4574,notn4574;
or (n4574,s0n4574,s1n4574);
not(notn4574,n2929);
and (s0n4574,notn4574,n813);
and (s1n4574,n2929,n1771);
or (n4575,1'b0,n4576,n4585,n4586,n4595);
and (n4576,n4577,n2718);
or (n4577,1'b0,n4578,n4582,n4583,n4584);
and (n4578,n4579,n2932);
wire s0n4579,s1n4579,notn4579;
or (n4579,s0n4579,s1n4579);
not(notn4579,n2929);
and (s0n4579,notn4579,n4580);
and (s1n4579,n2929,n4581);
and (n4582,n4071,n2955);
and (n4583,n3434,n2963);
and (n4584,n3365,n2972);
and (n4585,n4040,n2730);
and (n4586,n4587,n2742);
or (n4587,1'b0,n4588,n4592,n4593,n4594);
and (n4588,n4589,n2932);
wire s0n4589,s1n4589,notn4589;
or (n4589,s0n4589,s1n4589);
not(notn4589,n2929);
and (s0n4589,notn4589,n4590);
and (s1n4589,n2929,n4591);
and (n4592,n4086,n2955);
and (n4593,n3449,n2963);
and (n4594,n3401,n2972);
and (n4595,n4055,n2752);
and (n4596,n4575,n4597);
or (n4597,n4598,n4639,n4725);
and (n4598,n4599,n4618);
or (n4599,1'b0,n4600,n4601,n4610,n4611);
and (n4600,n4141,n2718);
and (n4601,n4602,n2730);
or (n4602,1'b0,n4603,n4604,n4605,n4606);
and (n4603,n3494,n2932);
and (n4604,n3498,n2955);
and (n4605,n4114,n2963);
and (n4606,n4607,n2972);
wire s0n4607,s1n4607,notn4607;
or (n4607,s0n4607,s1n4607);
not(notn4607,n2929);
and (s0n4607,notn4607,n4608);
and (s1n4607,n2929,n4609);
and (n4610,n4156,n2742);
and (n4611,n4612,n2752);
or (n4612,1'b0,n4613,n4614,n4615,n4616);
and (n4613,n3530,n2932);
and (n4614,n3532,n2955);
and (n4615,n4129,n2963);
and (n4616,n4617,n2972);
wire s0n4617,s1n4617,notn4617;
or (n4617,s0n4617,s1n4617);
not(notn4617,n2929);
and (s0n4617,notn4617,n829);
and (s1n4617,n2929,n1792);
or (n4618,1'b0,n4619,n4628,n4629,n4638);
and (n4619,n4620,n2718);
or (n4620,1'b0,n4621,n4625,n4626,n4627);
and (n4621,n4622,n2932);
wire s0n4622,s1n4622,notn4622;
or (n4622,s0n4622,s1n4622);
not(notn4622,n2929);
and (s0n4622,notn4622,n4623);
and (s1n4622,n2929,n4624);
and (n4625,n4134,n2955);
and (n4626,n3537,n2963);
and (n4627,n3468,n2972);
and (n4628,n4103,n2730);
and (n4629,n4630,n2742);
or (n4630,1'b0,n4631,n4635,n4636,n4637);
and (n4631,n4632,n2932);
wire s0n4632,s1n4632,notn4632;
or (n4632,s0n4632,s1n4632);
not(notn4632,n2929);
and (s0n4632,notn4632,n4633);
and (s1n4632,n2929,n4634);
and (n4635,n4149,n2955);
and (n4636,n3552,n2963);
and (n4637,n3504,n2972);
and (n4638,n4118,n2752);
and (n4639,n4618,n4640);
or (n4640,n4641,n4682,n4724);
and (n4641,n4642,n4661);
or (n4642,1'b0,n4643,n4644,n4653,n4654);
and (n4643,n4204,n2718);
and (n4644,n4645,n2730);
or (n4645,1'b0,n4646,n4647,n4648,n4649);
and (n4646,n3597,n2932);
and (n4647,n3601,n2955);
and (n4648,n4177,n2963);
and (n4649,n4650,n2972);
wire s0n4650,s1n4650,notn4650;
or (n4650,s0n4650,s1n4650);
not(notn4650,n2929);
and (s0n4650,notn4650,n4651);
and (s1n4650,n2929,n4652);
and (n4653,n4219,n2742);
and (n4654,n4655,n2752);
or (n4655,1'b0,n4656,n4657,n4658,n4659);
and (n4656,n3633,n2932);
and (n4657,n3635,n2955);
and (n4658,n4192,n2963);
and (n4659,n4660,n2972);
wire s0n4660,s1n4660,notn4660;
or (n4660,s0n4660,s1n4660);
not(notn4660,n2929);
and (s0n4660,notn4660,n845);
and (s1n4660,n2929,n1822);
or (n4661,1'b0,n4662,n4671,n4672,n4681);
and (n4662,n4663,n2718);
or (n4663,1'b0,n4664,n4668,n4669,n4670);
and (n4664,n4665,n2932);
wire s0n4665,s1n4665,notn4665;
or (n4665,s0n4665,s1n4665);
not(notn4665,n2929);
and (s0n4665,notn4665,n4666);
and (s1n4665,n2929,n4667);
and (n4668,n4197,n2955);
and (n4669,n3640,n2963);
and (n4670,n3571,n2972);
and (n4671,n4166,n2730);
and (n4672,n4673,n2742);
or (n4673,1'b0,n4674,n4678,n4679,n4680);
and (n4674,n4675,n2932);
wire s0n4675,s1n4675,notn4675;
or (n4675,s0n4675,s1n4675);
not(notn4675,n2929);
and (s0n4675,notn4675,n4676);
and (s1n4675,n2929,n4677);
and (n4678,n4212,n2955);
and (n4679,n3655,n2963);
and (n4680,n3607,n2972);
and (n4681,n4181,n2752);
and (n4682,n4661,n4683);
and (n4683,n4684,n4703);
or (n4684,1'b0,n4685,n4686,n4695,n4696);
and (n4685,n4266,n2718);
and (n4686,n4687,n2730);
or (n4687,1'b0,n4688,n4689,n4690,n4691);
and (n4688,n3699,n2932);
and (n4689,n3703,n2955);
and (n4690,n4239,n2963);
and (n4691,n4692,n2972);
wire s0n4692,s1n4692,notn4692;
or (n4692,s0n4692,s1n4692);
not(notn4692,n2929);
and (s0n4692,notn4692,n4693);
and (s1n4692,n2929,n4694);
and (n4695,n4281,n2742);
and (n4696,n4697,n2752);
or (n4697,1'b0,n4698,n4699,n4700,n4701);
and (n4698,n3735,n2932);
and (n4699,n3737,n2955);
and (n4700,n4254,n2963);
and (n4701,n4702,n2972);
wire s0n4702,s1n4702,notn4702;
or (n4702,s0n4702,s1n4702);
not(notn4702,n2929);
and (s0n4702,notn4702,n860);
and (s1n4702,n2929,n1845);
or (n4703,1'b0,n4704,n4713,n4714,n4723);
and (n4704,n4705,n2718);
or (n4705,1'b0,n4706,n4710,n4711,n4712);
and (n4706,n4707,n2932);
wire s0n4707,s1n4707,notn4707;
or (n4707,s0n4707,s1n4707);
not(notn4707,n2929);
and (s0n4707,notn4707,n4708);
and (s1n4707,n2929,n4709);
and (n4710,n4259,n2955);
and (n4711,n3742,n2963);
and (n4712,n3673,n2972);
and (n4713,n4228,n2730);
and (n4714,n4715,n2742);
or (n4715,1'b0,n4716,n4720,n4721,n4722);
and (n4716,n4717,n2932);
wire s0n4717,s1n4717,notn4717;
or (n4717,s0n4717,s1n4717);
not(notn4717,n2929);
and (s0n4717,notn4717,n4718);
and (s1n4717,n2929,n4719);
and (n4720,n4274,n2955);
and (n4721,n3757,n2963);
and (n4722,n3709,n2972);
and (n4723,n4243,n2752);
and (n4724,n4642,n4683);
and (n4725,n4599,n4640);
and (n4726,n4556,n4597);
and (n4727,n4513,n4554);
and (n4728,n4470,n4511);
and (n4729,n4427,n4468);
and (n4730,n4384,n4425);
xor (n4731,n4350,n4352);
and (n4732,n4731,n4733);
or (n4733,n4734,n4738,n4783);
and (n4734,n4735,n4737);
xor (n4735,n4736,n4425);
xor (n4736,n4384,n4403);
xor (n4737,n4353,n4355);
and (n4738,n4737,n4739);
or (n4739,n4740,n4744,n4782);
and (n4740,n4741,n4743);
xor (n4741,n4742,n4468);
xor (n4742,n4427,n4446);
xor (n4743,n4356,n4358);
and (n4744,n4743,n4745);
or (n4745,n4746,n4750,n4781);
and (n4746,n4747,n4749);
xor (n4747,n4748,n4511);
xor (n4748,n4470,n4489);
xor (n4749,n4359,n4361);
and (n4750,n4749,n4751);
or (n4751,n4752,n4756,n4780);
and (n4752,n4753,n4755);
xor (n4753,n4754,n4554);
xor (n4754,n4513,n4532);
xor (n4755,n4362,n4364);
and (n4756,n4755,n4757);
or (n4757,n4758,n4762,n4779);
and (n4758,n4759,n4761);
xor (n4759,n4760,n4597);
xor (n4760,n4556,n4575);
xor (n4761,n4365,n4367);
and (n4762,n4761,n4763);
or (n4763,n4764,n4768,n4778);
and (n4764,n4765,n4767);
xor (n4765,n4766,n4640);
xor (n4766,n4599,n4618);
xor (n4767,n4368,n4369);
and (n4768,n4767,n4769);
or (n4769,n4770,n4774,n4777);
and (n4770,n4771,n4773);
xor (n4771,n4772,n4683);
xor (n4772,n4642,n4661);
xor (n4773,n4370,n4373);
and (n4774,n4773,n4775);
and (n4775,n4776,n4374);
xor (n4776,n4684,n4703);
and (n4777,n4771,n4775);
and (n4778,n4765,n4769);
and (n4779,n4759,n4763);
and (n4780,n4753,n4757);
and (n4781,n4747,n4751);
and (n4782,n4741,n4745);
and (n4783,n4735,n4739);
and (n4784,n4382,n4733);
or (n4785,n4786,n4787,n4837);
xor (n4786,n2918,n4376);
and (n4787,n4379,n4788);
or (n4788,n4789,n4791,n4836);
and (n4789,n4790,n4731);
xor (n4790,n4377,n4378);
and (n4791,n4731,n4792);
or (n4792,n4793,n4795,n4835);
and (n4793,n4794,n4737);
xor (n4794,n4379,n4380);
and (n4795,n4737,n4796);
or (n4796,n4797,n4800,n4834);
and (n4797,n4798,n4743);
xor (n4798,n4799,n4733);
xor (n4799,n4382,n4731);
and (n4800,n4743,n4801);
or (n4801,n4802,n4805,n4833);
and (n4802,n4803,n4749);
xor (n4803,n4804,n4739);
xor (n4804,n4735,n4737);
and (n4805,n4749,n4806);
or (n4806,n4807,n4810,n4832);
and (n4807,n4808,n4755);
xor (n4808,n4809,n4745);
xor (n4809,n4741,n4743);
and (n4810,n4755,n4811);
or (n4811,n4812,n4815,n4831);
and (n4812,n4813,n4761);
xor (n4813,n4814,n4751);
xor (n4814,n4747,n4749);
and (n4815,n4761,n4816);
or (n4816,n4817,n4820,n4830);
and (n4817,n4818,n4767);
xor (n4818,n4819,n4757);
xor (n4819,n4753,n4755);
and (n4820,n4767,n4821);
or (n4821,n4822,n4825,n4829);
and (n4822,n4823,n4773);
xor (n4823,n4824,n4763);
xor (n4824,n4759,n4761);
and (n4825,n4773,n4826);
and (n4826,n4827,n4374);
xor (n4827,n4828,n4769);
xor (n4828,n4765,n4767);
and (n4829,n4823,n4826);
and (n4830,n4818,n4821);
and (n4831,n4813,n4816);
and (n4832,n4808,n4811);
and (n4833,n4803,n4806);
and (n4834,n4798,n4801);
and (n4835,n4794,n4796);
and (n4836,n4790,n4792);
and (n4837,n4786,n4788);
and (n4838,n4839,n4841);
xor (n4839,n4840,n4788);
xor (n4840,n4786,n4379);
and (n4841,n4842,n4844);
xor (n4842,n4843,n4792);
xor (n4843,n4790,n4731);
and (n4844,n4845,n4847);
xor (n4845,n4846,n4796);
xor (n4846,n4794,n4737);
and (n4847,n4848,n4850);
xor (n4848,n4849,n4801);
xor (n4849,n4798,n4743);
and (n4850,n4851,n4853);
xor (n4851,n4852,n4806);
xor (n4852,n4803,n4749);
and (n4853,n4854,n4856);
xor (n4854,n4855,n4811);
xor (n4855,n4808,n4755);
and (n4856,n4857,n4859);
xor (n4857,n4858,n4816);
xor (n4858,n4813,n4761);
xor (n4859,n4860,n4821);
xor (n4860,n4818,n4767);
and (n4861,n4862,n4872);
and (n4862,n4863,n4871);
and (n4863,n4864,n4870);
and (n4864,n4865,n4869);
and (n4865,n4866,n4868);
and (n4866,n2704,n4867);
not (n4867,n2756);
not (n4868,n2908);
not (n4869,n2950);
not (n4870,n2909);
or (n4871,n2895,n2800,n2826,n2852);
nand (n4872,n2757,n2800,n2898,n2896);
wire s0n4873,s1n4873,notn4873;
or (n4873,s0n4873,s1n4873);
not(notn4873,n4861);
and (s0n4873,notn4873,1'b0);
and (s1n4873,n4861,n4874);
xor (n4874,n4875,n4877);
xor (n4875,n4375,n4876);
and (n4876,n4377,n4785);
and (n4877,n2915,n4838);
wire s0n4878,s1n4878,notn4878;
or (n4878,s0n4878,s1n4878);
not(notn4878,n4861);
and (s0n4878,notn4878,1'b0);
and (s1n4878,n4861,n4879);
xor (n4879,n4880,n4882);
xor (n4880,n4375,n4881);
and (n4881,n2918,n4876);
and (n4882,n4875,n4877);
or (n4883,n4884,n2931);
or (n4884,n4885,n2930);
or (n4885,n2945,n2946);
or (n4886,1'b0,n4887,n4905,n4920,n4935);
and (n4887,n4888,n2718);
or (n4888,1'b0,n4889,n4896,n4902);
and (n4889,n4890,n4895);
or (n4890,1'b0,n4891,n4892,n4893,n4894);
and (n4891,n2928,n556);
and (n4892,n2954,n567);
and (n4893,n2962,n571);
and (n4894,n2971,n573);
not (n4895,n4872);
and (n4896,n4897,n2944);
or (n4897,1'b0,n4898,n4899,n4900,n4901);
and (n4898,n3023,n556);
and (n4899,n2711,n567);
and (n4900,n2713,n571);
and (n4901,n2715,n573);
and (n4902,n2709,n4903);
or (n4903,n2942,n4904);
not (n4904,n4871);
and (n4905,n4906,n2730);
or (n4906,1'b0,n4907,n4913,n4919);
and (n4907,n4908,n4895);
or (n4908,1'b0,n4909,n4910,n4911,n4912);
and (n4909,n2982,n556);
and (n4910,n2985,n567);
and (n4911,n2988,n571);
and (n4912,n2991,n573);
and (n4913,n4914,n2944);
or (n4914,1'b0,n4915,n4916,n4917,n4918);
and (n4915,n2717,n556);
and (n4916,n2723,n567);
and (n4917,n2725,n571);
and (n4918,n2727,n573);
and (n4919,n2721,n4903);
and (n4920,n4921,n2742);
or (n4921,1'b0,n4922,n4928,n4934);
and (n4922,n4923,n4895);
or (n4923,1'b0,n4924,n4925,n4926,n4927);
and (n4924,n2996,n556);
and (n4925,n2999,n567);
and (n4926,n3002,n571);
and (n4927,n3005,n573);
and (n4928,n4929,n2944);
or (n4929,1'b0,n4930,n4931,n4932,n4933);
and (n4930,n3038,n556);
and (n4931,n2735,n567);
and (n4932,n2737,n571);
and (n4933,n2739,n573);
and (n4934,n2733,n4903);
and (n4935,n4936,n2752);
or (n4936,1'b0,n4937,n4943,n4949);
and (n4937,n4938,n4895);
or (n4938,1'b0,n4939,n4940,n4941,n4942);
and (n4939,n3010,n556);
and (n4940,n3013,n567);
and (n4941,n2087,n571);
and (n4942,n1692,n573);
and (n4943,n4944,n2944);
or (n4944,1'b0,n4945,n4946,n4947,n4948);
and (n4945,n2741,n556);
and (n4946,n2747,n567);
and (n4947,n2749,n571);
and (n4948,n1251,n573);
and (n4949,n2745,n4903);
or (n4950,1'b0,n4951,n7872,n7874,n7877);
and (n4951,n4952,n2893);
wire s0n4952,s1n4952,notn4952;
or (n4952,s0n4952,s1n4952);
not(notn4952,n2891);
and (s0n4952,notn4952,1'b0);
and (s1n4952,n2891,n4953);
wire s0n4953,s1n4953,notn4953;
or (n4953,s0n4953,s1n4953);
not(notn4953,n7861);
and (s0n4953,notn4953,n4954);
and (s1n4953,n7861,1'b0);
wire s0n4954,s1n4954,notn4954;
or (n4954,s0n4954,s1n4954);
not(notn4954,n7846);
and (s0n4954,notn4954,n4955);
and (s1n4954,n7846,1'b1);
wire s0n4955,s1n4955,notn4955;
or (n4955,s0n4955,s1n4955);
not(notn4955,n4966);
and (s0n4955,notn4955,n4956);
and (s1n4955,n4966,n7635);
wire s0n4956,s1n4956,notn4956;
or (n4956,s0n4956,s1n4956);
not(notn4956,n4966);
and (s0n4956,notn4956,n4957);
and (s1n4956,n4966,n7632);
xor (n4957,n4958,n7609);
xor (n4958,n4959,n7552);
xor (n4959,n4960,n7483);
xor (n4960,n4961,n7473);
xor (n4961,n4962,n6014);
xor (n4962,n4963,n4976);
xor (n4963,n4964,n4974);
wire s0n4964,s1n4964,notn4964;
or (n4964,s0n4964,s1n4964);
not(notn4964,n4966);
and (s0n4964,notn4964,1'b0);
and (s1n4964,n4966,n4965);
or (n4966,n4967,n4973);
or (n4967,n4968,n4972);
and (n4968,n2950,n4969);
or (n4969,n4970,n556);
or (n4970,n4971,n567);
or (n4971,n573,n571);
and (n4972,n2893,n4969);
and (n4973,n2907,n2902);
wire s0n4974,s1n4974,notn4974;
or (n4974,s0n4974,s1n4974);
not(notn4974,n4966);
and (s0n4974,notn4974,1'b0);
and (s1n4974,n4966,n4975);
or (n4976,n4977,n4982,n6013);
and (n4977,n4978,n4980);
wire s0n4978,s1n4978,notn4978;
or (n4978,s0n4978,s1n4978);
not(notn4978,n4966);
and (s0n4978,notn4978,1'b0);
and (s1n4978,n4966,n4979);
wire s0n4980,s1n4980,notn4980;
or (n4980,s0n4980,s1n4980);
not(notn4980,n4966);
and (s0n4980,notn4980,1'b0);
and (s1n4980,n4966,n4981);
and (n4982,n4980,n4983);
or (n4983,n4984,n4989,n6012);
and (n4984,n4985,n4987);
wire s0n4985,s1n4985,notn4985;
or (n4985,s0n4985,s1n4985);
not(notn4985,n4966);
and (s0n4985,notn4985,1'b0);
and (s1n4985,n4966,n4986);
wire s0n4987,s1n4987,notn4987;
or (n4987,s0n4987,s1n4987);
not(notn4987,n4966);
and (s0n4987,notn4987,1'b0);
and (s1n4987,n4966,n4988);
and (n4989,n4987,n4990);
or (n4990,n4991,n4996,n6011);
and (n4991,n4992,n4994);
wire s0n4992,s1n4992,notn4992;
or (n4992,s0n4992,s1n4992);
not(notn4992,n4966);
and (s0n4992,notn4992,1'b0);
and (s1n4992,n4966,n4993);
wire s0n4994,s1n4994,notn4994;
or (n4994,s0n4994,s1n4994);
not(notn4994,n4966);
and (s0n4994,notn4994,1'b0);
and (s1n4994,n4966,n4995);
and (n4996,n4994,n4997);
or (n4997,n4998,n5003,n6010);
and (n4998,n4999,n5001);
wire s0n4999,s1n4999,notn4999;
or (n4999,s0n4999,s1n4999);
not(notn4999,n4966);
and (s0n4999,notn4999,1'b0);
and (s1n4999,n4966,n5000);
wire s0n5001,s1n5001,notn5001;
or (n5001,s0n5001,s1n5001);
not(notn5001,n4966);
and (s0n5001,notn5001,1'b0);
and (s1n5001,n4966,n5002);
and (n5003,n5001,n5004);
or (n5004,n5005,n5143,n6009);
and (n5005,n5006,n5082);
wire s0n5006,s1n5006,notn5006;
or (n5006,s0n5006,s1n5006);
not(notn5006,n4966);
and (s0n5006,notn5006,n5007);
and (s1n5006,n4966,n5081);
or (n5007,1'b0,n5008,n5040,n5054,n5069);
and (n5008,n5009,n2718);
or (n5009,1'b0,n5010,n5025,n5030,n5035);
and (n5010,n5011,n5016);
wire s0n5011,s1n5011,notn5011;
or (n5011,s0n5011,s1n5011);
not(notn5011,n5014);
and (s0n5011,notn5011,n5012);
and (s1n5011,n5014,n5013);
or (n5014,n5015,n2909);
or (n5015,n2946,n2931);
or (n5016,n5017,n2951);
and (n5017,n5018,n556);
or (n5018,n5019,n2931);
or (n5019,n5020,n2930);
or (n5020,n5021,n2946);
or (n5021,n5022,n2945);
or (n5022,n5023,n4895);
or (n5023,n5024,n4904);
nor (n5024,n2757,n2943,n2826,n2852);
and (n5025,n5026,n5028);
wire s0n5026,s1n5026,notn5026;
or (n5026,s0n5026,s1n5026);
not(notn5026,n5014);
and (s0n5026,notn5026,n5027);
and (s1n5026,n5014,n5012);
or (n5028,n5029,n2959);
and (n5029,n5018,n567);
and (n5030,n5031,n5033);
wire s0n5031,s1n5031,notn5031;
or (n5031,s0n5031,s1n5031);
not(notn5031,n5014);
and (s0n5031,notn5031,n5032);
and (s1n5031,n5014,n5027);
or (n5033,n5034,n2967);
and (n5034,n5018,n571);
and (n5035,n5036,n5038);
wire s0n5036,s1n5036,notn5036;
or (n5036,s0n5036,s1n5036);
not(notn5036,n5014);
and (s0n5036,notn5036,n5037);
and (s1n5036,n5014,n5032);
or (n5038,n5039,n2976);
and (n5039,n5018,n573);
and (n5040,n5041,n2730);
or (n5041,1'b0,n5042,n5045,n5048,n5051);
and (n5042,n5043,n5016);
wire s0n5043,s1n5043,notn5043;
or (n5043,s0n5043,s1n5043);
not(notn5043,n5014);
and (s0n5043,notn5043,n5044);
and (s1n5043,n5014,n5037);
and (n5045,n5046,n5028);
wire s0n5046,s1n5046,notn5046;
or (n5046,s0n5046,s1n5046);
not(notn5046,n5014);
and (s0n5046,notn5046,n5047);
and (s1n5046,n5014,n5044);
and (n5048,n5049,n5033);
wire s0n5049,s1n5049,notn5049;
or (n5049,s0n5049,s1n5049);
not(notn5049,n5014);
and (s0n5049,notn5049,n5050);
and (s1n5049,n5014,n5047);
and (n5051,n5052,n5038);
wire s0n5052,s1n5052,notn5052;
or (n5052,s0n5052,s1n5052);
not(notn5052,n5014);
and (s0n5052,notn5052,n5053);
and (s1n5052,n5014,n5050);
and (n5054,n5055,n2742);
or (n5055,1'b0,n5056,n5060,n5063,n5066);
and (n5056,n5057,n5016);
wire s0n5057,s1n5057,notn5057;
or (n5057,s0n5057,s1n5057);
not(notn5057,n5014);
and (s0n5057,notn5057,n5058);
and (s1n5057,n5014,n5059);
and (n5060,n5061,n5028);
wire s0n5061,s1n5061,notn5061;
or (n5061,s0n5061,s1n5061);
not(notn5061,n5014);
and (s0n5061,notn5061,n5062);
and (s1n5061,n5014,n5058);
and (n5063,n5064,n5033);
wire s0n5064,s1n5064,notn5064;
or (n5064,s0n5064,s1n5064);
not(notn5064,n5014);
and (s0n5064,notn5064,n5065);
and (s1n5064,n5014,n5062);
and (n5066,n5067,n5038);
wire s0n5067,s1n5067,notn5067;
or (n5067,s0n5067,s1n5067);
not(notn5067,n5014);
and (s0n5067,notn5067,n5068);
and (s1n5067,n5014,n5065);
and (n5069,n5070,n2752);
or (n5070,1'b0,n5071,n5074,n5077,n5079);
and (n5071,n5072,n5016);
wire s0n5072,s1n5072,notn5072;
or (n5072,s0n5072,s1n5072);
not(notn5072,n5014);
and (s0n5072,notn5072,n5073);
and (s1n5072,n5014,n5068);
and (n5074,n5075,n5028);
wire s0n5075,s1n5075,notn5075;
or (n5075,s0n5075,s1n5075);
not(notn5075,n5014);
and (s0n5075,notn5075,n5076);
and (s1n5075,n5014,n5073);
and (n5077,n5078,n5033);
wire s0n5078,s1n5078,notn5078;
or (n5078,s0n5078,s1n5078);
not(notn5078,n5014);
and (s0n5078,notn5078,n1255);
and (s1n5078,n5014,n5076);
and (n5079,n5080,n5038);
wire s0n5080,s1n5080,notn5080;
or (n5080,s0n5080,s1n5080);
not(notn5080,n5014);
and (s0n5080,notn5080,n570);
and (s1n5080,n5014,n1255);
wire s0n5082,s1n5082,notn5082;
or (n5082,s0n5082,s1n5082);
not(notn5082,n4966);
and (s0n5082,notn5082,n5083);
and (s1n5082,n4966,n5142);
or (n5083,1'b0,n5084,n5099,n5113,n5128);
and (n5084,n5085,n2718);
or (n5085,1'b0,n5086,n5090,n5093,n5096);
and (n5086,n5087,n5016);
wire s0n5087,s1n5087,notn5087;
or (n5087,s0n5087,s1n5087);
not(notn5087,n5014);
and (s0n5087,notn5087,n5088);
and (s1n5087,n5014,n5089);
and (n5090,n5091,n5028);
wire s0n5091,s1n5091,notn5091;
or (n5091,s0n5091,s1n5091);
not(notn5091,n5014);
and (s0n5091,notn5091,n5092);
and (s1n5091,n5014,n5088);
and (n5093,n5094,n5033);
wire s0n5094,s1n5094,notn5094;
or (n5094,s0n5094,s1n5094);
not(notn5094,n5014);
and (s0n5094,notn5094,n5095);
and (s1n5094,n5014,n5092);
and (n5096,n5097,n5038);
wire s0n5097,s1n5097,notn5097;
or (n5097,s0n5097,s1n5097);
not(notn5097,n5014);
and (s0n5097,notn5097,n5098);
and (s1n5097,n5014,n5095);
and (n5099,n5100,n2730);
or (n5100,1'b0,n5101,n5104,n5107,n5110);
and (n5101,n5102,n5016);
wire s0n5102,s1n5102,notn5102;
or (n5102,s0n5102,s1n5102);
not(notn5102,n5014);
and (s0n5102,notn5102,n5103);
and (s1n5102,n5014,n5098);
and (n5104,n5105,n5028);
wire s0n5105,s1n5105,notn5105;
or (n5105,s0n5105,s1n5105);
not(notn5105,n5014);
and (s0n5105,notn5105,n5106);
and (s1n5105,n5014,n5103);
and (n5107,n5108,n5033);
wire s0n5108,s1n5108,notn5108;
or (n5108,s0n5108,s1n5108);
not(notn5108,n5014);
and (s0n5108,notn5108,n5109);
and (s1n5108,n5014,n5106);
and (n5110,n5111,n5038);
wire s0n5111,s1n5111,notn5111;
or (n5111,s0n5111,s1n5111);
not(notn5111,n5014);
and (s0n5111,notn5111,n5112);
and (s1n5111,n5014,n5109);
and (n5113,n5114,n2742);
or (n5114,1'b0,n5115,n5119,n5122,n5125);
and (n5115,n5116,n5016);
wire s0n5116,s1n5116,notn5116;
or (n5116,s0n5116,s1n5116);
not(notn5116,n5014);
and (s0n5116,notn5116,n5117);
and (s1n5116,n5014,n5118);
and (n5119,n5120,n5028);
wire s0n5120,s1n5120,notn5120;
or (n5120,s0n5120,s1n5120);
not(notn5120,n5014);
and (s0n5120,notn5120,n5121);
and (s1n5120,n5014,n5117);
and (n5122,n5123,n5033);
wire s0n5123,s1n5123,notn5123;
or (n5123,s0n5123,s1n5123);
not(notn5123,n5014);
and (s0n5123,notn5123,n5124);
and (s1n5123,n5014,n5121);
and (n5125,n5126,n5038);
wire s0n5126,s1n5126,notn5126;
or (n5126,s0n5126,s1n5126);
not(notn5126,n5014);
and (s0n5126,notn5126,n5127);
and (s1n5126,n5014,n5124);
and (n5128,n5129,n2752);
or (n5129,1'b0,n5130,n5133,n5136,n5139);
and (n5130,n5131,n5016);
wire s0n5131,s1n5131,notn5131;
or (n5131,s0n5131,s1n5131);
not(notn5131,n5014);
and (s0n5131,notn5131,n5132);
and (s1n5131,n5014,n5127);
and (n5133,n5134,n5028);
wire s0n5134,s1n5134,notn5134;
or (n5134,s0n5134,s1n5134);
not(notn5134,n5014);
and (s0n5134,notn5134,n5135);
and (s1n5134,n5014,n5132);
and (n5136,n5137,n5033);
wire s0n5137,s1n5137,notn5137;
or (n5137,s0n5137,s1n5137);
not(notn5137,n5014);
and (s0n5137,notn5137,n5138);
and (s1n5137,n5014,n5135);
and (n5139,n5140,n5038);
wire s0n5140,s1n5140,notn5140;
or (n5140,s0n5140,s1n5140);
not(notn5140,n5014);
and (s0n5140,notn5140,n5141);
and (s1n5140,n5014,n5138);
and (n5143,n5082,n5144);
or (n5144,n5145,n5266,n6008);
and (n5145,n5146,n5205);
wire s0n5146,s1n5146,notn5146;
or (n5146,s0n5146,s1n5146);
not(notn5146,n4966);
and (s0n5146,notn5146,n5147);
and (s1n5146,n4966,n5204);
or (n5147,1'b0,n5148,n5163,n5177,n5192);
and (n5148,n5149,n2718);
or (n5149,1'b0,n5150,n5154,n5157,n5160);
and (n5150,n5151,n5016);
wire s0n5151,s1n5151,notn5151;
or (n5151,s0n5151,s1n5151);
not(notn5151,n5014);
and (s0n5151,notn5151,n5152);
and (s1n5151,n5014,n5153);
and (n5154,n5155,n5028);
wire s0n5155,s1n5155,notn5155;
or (n5155,s0n5155,s1n5155);
not(notn5155,n5014);
and (s0n5155,notn5155,n5156);
and (s1n5155,n5014,n5152);
and (n5157,n5158,n5033);
wire s0n5158,s1n5158,notn5158;
or (n5158,s0n5158,s1n5158);
not(notn5158,n5014);
and (s0n5158,notn5158,n5159);
and (s1n5158,n5014,n5156);
and (n5160,n5161,n5038);
wire s0n5161,s1n5161,notn5161;
or (n5161,s0n5161,s1n5161);
not(notn5161,n5014);
and (s0n5161,notn5161,n5162);
and (s1n5161,n5014,n5159);
and (n5163,n5164,n2730);
or (n5164,1'b0,n5165,n5168,n5171,n5174);
and (n5165,n5166,n5016);
wire s0n5166,s1n5166,notn5166;
or (n5166,s0n5166,s1n5166);
not(notn5166,n5014);
and (s0n5166,notn5166,n5167);
and (s1n5166,n5014,n5162);
and (n5168,n5169,n5028);
wire s0n5169,s1n5169,notn5169;
or (n5169,s0n5169,s1n5169);
not(notn5169,n5014);
and (s0n5169,notn5169,n5170);
and (s1n5169,n5014,n5167);
and (n5171,n5172,n5033);
wire s0n5172,s1n5172,notn5172;
or (n5172,s0n5172,s1n5172);
not(notn5172,n5014);
and (s0n5172,notn5172,n5173);
and (s1n5172,n5014,n5170);
and (n5174,n5175,n5038);
wire s0n5175,s1n5175,notn5175;
or (n5175,s0n5175,s1n5175);
not(notn5175,n5014);
and (s0n5175,notn5175,n5176);
and (s1n5175,n5014,n5173);
and (n5177,n5178,n2742);
or (n5178,1'b0,n5179,n5183,n5186,n5189);
and (n5179,n5180,n5016);
wire s0n5180,s1n5180,notn5180;
or (n5180,s0n5180,s1n5180);
not(notn5180,n5014);
and (s0n5180,notn5180,n5181);
and (s1n5180,n5014,n5182);
and (n5183,n5184,n5028);
wire s0n5184,s1n5184,notn5184;
or (n5184,s0n5184,s1n5184);
not(notn5184,n5014);
and (s0n5184,notn5184,n5185);
and (s1n5184,n5014,n5181);
and (n5186,n5187,n5033);
wire s0n5187,s1n5187,notn5187;
or (n5187,s0n5187,s1n5187);
not(notn5187,n5014);
and (s0n5187,notn5187,n5188);
and (s1n5187,n5014,n5185);
and (n5189,n5190,n5038);
wire s0n5190,s1n5190,notn5190;
or (n5190,s0n5190,s1n5190);
not(notn5190,n5014);
and (s0n5190,notn5190,n5191);
and (s1n5190,n5014,n5188);
and (n5192,n5193,n2752);
or (n5193,1'b0,n5194,n5197,n5200,n5202);
and (n5194,n5195,n5016);
wire s0n5195,s1n5195,notn5195;
or (n5195,s0n5195,s1n5195);
not(notn5195,n5014);
and (s0n5195,notn5195,n5196);
and (s1n5195,n5014,n5191);
and (n5197,n5198,n5028);
wire s0n5198,s1n5198,notn5198;
or (n5198,s0n5198,s1n5198);
not(notn5198,n5014);
and (s0n5198,notn5198,n5199);
and (s1n5198,n5014,n5196);
and (n5200,n5201,n5033);
wire s0n5201,s1n5201,notn5201;
or (n5201,s0n5201,s1n5201);
not(notn5201,n5014);
and (s0n5201,notn5201,n1271);
and (s1n5201,n5014,n5199);
and (n5202,n5203,n5038);
wire s0n5203,s1n5203,notn5203;
or (n5203,s0n5203,s1n5203);
not(notn5203,n5014);
and (s0n5203,notn5203,n759);
and (s1n5203,n5014,n1271);
wire s0n5205,s1n5205,notn5205;
or (n5205,s0n5205,s1n5205);
not(notn5205,n4966);
and (s0n5205,notn5205,n5206);
and (s1n5205,n4966,n5265);
or (n5206,1'b0,n5207,n5222,n5236,n5251);
and (n5207,n5208,n2718);
or (n5208,1'b0,n5209,n5213,n5216,n5219);
and (n5209,n5210,n5016);
wire s0n5210,s1n5210,notn5210;
or (n5210,s0n5210,s1n5210);
not(notn5210,n5014);
and (s0n5210,notn5210,n5211);
and (s1n5210,n5014,n5212);
and (n5213,n5214,n5028);
wire s0n5214,s1n5214,notn5214;
or (n5214,s0n5214,s1n5214);
not(notn5214,n5014);
and (s0n5214,notn5214,n5215);
and (s1n5214,n5014,n5211);
and (n5216,n5217,n5033);
wire s0n5217,s1n5217,notn5217;
or (n5217,s0n5217,s1n5217);
not(notn5217,n5014);
and (s0n5217,notn5217,n5218);
and (s1n5217,n5014,n5215);
and (n5219,n5220,n5038);
wire s0n5220,s1n5220,notn5220;
or (n5220,s0n5220,s1n5220);
not(notn5220,n5014);
and (s0n5220,notn5220,n5221);
and (s1n5220,n5014,n5218);
and (n5222,n5223,n2730);
or (n5223,1'b0,n5224,n5227,n5230,n5233);
and (n5224,n5225,n5016);
wire s0n5225,s1n5225,notn5225;
or (n5225,s0n5225,s1n5225);
not(notn5225,n5014);
and (s0n5225,notn5225,n5226);
and (s1n5225,n5014,n5221);
and (n5227,n5228,n5028);
wire s0n5228,s1n5228,notn5228;
or (n5228,s0n5228,s1n5228);
not(notn5228,n5014);
and (s0n5228,notn5228,n5229);
and (s1n5228,n5014,n5226);
and (n5230,n5231,n5033);
wire s0n5231,s1n5231,notn5231;
or (n5231,s0n5231,s1n5231);
not(notn5231,n5014);
and (s0n5231,notn5231,n5232);
and (s1n5231,n5014,n5229);
and (n5233,n5234,n5038);
wire s0n5234,s1n5234,notn5234;
or (n5234,s0n5234,s1n5234);
not(notn5234,n5014);
and (s0n5234,notn5234,n5235);
and (s1n5234,n5014,n5232);
and (n5236,n5237,n2742);
or (n5237,1'b0,n5238,n5242,n5245,n5248);
and (n5238,n5239,n5016);
wire s0n5239,s1n5239,notn5239;
or (n5239,s0n5239,s1n5239);
not(notn5239,n5014);
and (s0n5239,notn5239,n5240);
and (s1n5239,n5014,n5241);
and (n5242,n5243,n5028);
wire s0n5243,s1n5243,notn5243;
or (n5243,s0n5243,s1n5243);
not(notn5243,n5014);
and (s0n5243,notn5243,n5244);
and (s1n5243,n5014,n5240);
and (n5245,n5246,n5033);
wire s0n5246,s1n5246,notn5246;
or (n5246,s0n5246,s1n5246);
not(notn5246,n5014);
and (s0n5246,notn5246,n5247);
and (s1n5246,n5014,n5244);
and (n5248,n5249,n5038);
wire s0n5249,s1n5249,notn5249;
or (n5249,s0n5249,s1n5249);
not(notn5249,n5014);
and (s0n5249,notn5249,n5250);
and (s1n5249,n5014,n5247);
and (n5251,n5252,n2752);
or (n5252,1'b0,n5253,n5256,n5259,n5262);
and (n5253,n5254,n5016);
wire s0n5254,s1n5254,notn5254;
or (n5254,s0n5254,s1n5254);
not(notn5254,n5014);
and (s0n5254,notn5254,n5255);
and (s1n5254,n5014,n5250);
and (n5256,n5257,n5028);
wire s0n5257,s1n5257,notn5257;
or (n5257,s0n5257,s1n5257);
not(notn5257,n5014);
and (s0n5257,notn5257,n5258);
and (s1n5257,n5014,n5255);
and (n5259,n5260,n5033);
wire s0n5260,s1n5260,notn5260;
or (n5260,s0n5260,s1n5260);
not(notn5260,n5014);
and (s0n5260,notn5260,n5261);
and (s1n5260,n5014,n5258);
and (n5262,n5263,n5038);
wire s0n5263,s1n5263,notn5263;
or (n5263,s0n5263,s1n5263);
not(notn5263,n5014);
and (s0n5263,notn5263,n5264);
and (s1n5263,n5014,n5261);
and (n5266,n5205,n5267);
or (n5267,n5268,n5389,n6007);
and (n5268,n5269,n5328);
wire s0n5269,s1n5269,notn5269;
or (n5269,s0n5269,s1n5269);
not(notn5269,n4966);
and (s0n5269,notn5269,n5270);
and (s1n5269,n4966,n5327);
or (n5270,1'b0,n5271,n5286,n5300,n5315);
and (n5271,n5272,n2718);
or (n5272,1'b0,n5273,n5277,n5280,n5283);
and (n5273,n5274,n5016);
wire s0n5274,s1n5274,notn5274;
or (n5274,s0n5274,s1n5274);
not(notn5274,n5014);
and (s0n5274,notn5274,n5275);
and (s1n5274,n5014,n5276);
and (n5277,n5278,n5028);
wire s0n5278,s1n5278,notn5278;
or (n5278,s0n5278,s1n5278);
not(notn5278,n5014);
and (s0n5278,notn5278,n5279);
and (s1n5278,n5014,n5275);
and (n5280,n5281,n5033);
wire s0n5281,s1n5281,notn5281;
or (n5281,s0n5281,s1n5281);
not(notn5281,n5014);
and (s0n5281,notn5281,n5282);
and (s1n5281,n5014,n5279);
and (n5283,n5284,n5038);
wire s0n5284,s1n5284,notn5284;
or (n5284,s0n5284,s1n5284);
not(notn5284,n5014);
and (s0n5284,notn5284,n5285);
and (s1n5284,n5014,n5282);
and (n5286,n5287,n2730);
or (n5287,1'b0,n5288,n5291,n5294,n5297);
and (n5288,n5289,n5016);
wire s0n5289,s1n5289,notn5289;
or (n5289,s0n5289,s1n5289);
not(notn5289,n5014);
and (s0n5289,notn5289,n5290);
and (s1n5289,n5014,n5285);
and (n5291,n5292,n5028);
wire s0n5292,s1n5292,notn5292;
or (n5292,s0n5292,s1n5292);
not(notn5292,n5014);
and (s0n5292,notn5292,n5293);
and (s1n5292,n5014,n5290);
and (n5294,n5295,n5033);
wire s0n5295,s1n5295,notn5295;
or (n5295,s0n5295,s1n5295);
not(notn5295,n5014);
and (s0n5295,notn5295,n5296);
and (s1n5295,n5014,n5293);
and (n5297,n5298,n5038);
wire s0n5298,s1n5298,notn5298;
or (n5298,s0n5298,s1n5298);
not(notn5298,n5014);
and (s0n5298,notn5298,n5299);
and (s1n5298,n5014,n5296);
and (n5300,n5301,n2742);
or (n5301,1'b0,n5302,n5306,n5309,n5312);
and (n5302,n5303,n5016);
wire s0n5303,s1n5303,notn5303;
or (n5303,s0n5303,s1n5303);
not(notn5303,n5014);
and (s0n5303,notn5303,n5304);
and (s1n5303,n5014,n5305);
and (n5306,n5307,n5028);
wire s0n5307,s1n5307,notn5307;
or (n5307,s0n5307,s1n5307);
not(notn5307,n5014);
and (s0n5307,notn5307,n5308);
and (s1n5307,n5014,n5304);
and (n5309,n5310,n5033);
wire s0n5310,s1n5310,notn5310;
or (n5310,s0n5310,s1n5310);
not(notn5310,n5014);
and (s0n5310,notn5310,n5311);
and (s1n5310,n5014,n5308);
and (n5312,n5313,n5038);
wire s0n5313,s1n5313,notn5313;
or (n5313,s0n5313,s1n5313);
not(notn5313,n5014);
and (s0n5313,notn5313,n5314);
and (s1n5313,n5014,n5311);
and (n5315,n5316,n2752);
or (n5316,1'b0,n5317,n5320,n5323,n5325);
and (n5317,n5318,n5016);
wire s0n5318,s1n5318,notn5318;
or (n5318,s0n5318,s1n5318);
not(notn5318,n5014);
and (s0n5318,notn5318,n5319);
and (s1n5318,n5014,n5314);
and (n5320,n5321,n5028);
wire s0n5321,s1n5321,notn5321;
or (n5321,s0n5321,s1n5321);
not(notn5321,n5014);
and (s0n5321,notn5321,n5322);
and (s1n5321,n5014,n5319);
and (n5323,n5324,n5033);
wire s0n5324,s1n5324,notn5324;
or (n5324,s0n5324,s1n5324);
not(notn5324,n5014);
and (s0n5324,notn5324,n1287);
and (s1n5324,n5014,n5322);
and (n5325,n5326,n5038);
wire s0n5326,s1n5326,notn5326;
or (n5326,s0n5326,s1n5326);
not(notn5326,n5014);
and (s0n5326,notn5326,n783);
and (s1n5326,n5014,n1287);
wire s0n5328,s1n5328,notn5328;
or (n5328,s0n5328,s1n5328);
not(notn5328,n4966);
and (s0n5328,notn5328,n5329);
and (s1n5328,n4966,n5388);
or (n5329,1'b0,n5330,n5345,n5359,n5374);
and (n5330,n5331,n2718);
or (n5331,1'b0,n5332,n5336,n5339,n5342);
and (n5332,n5333,n5016);
wire s0n5333,s1n5333,notn5333;
or (n5333,s0n5333,s1n5333);
not(notn5333,n5014);
and (s0n5333,notn5333,n5334);
and (s1n5333,n5014,n5335);
and (n5336,n5337,n5028);
wire s0n5337,s1n5337,notn5337;
or (n5337,s0n5337,s1n5337);
not(notn5337,n5014);
and (s0n5337,notn5337,n5338);
and (s1n5337,n5014,n5334);
and (n5339,n5340,n5033);
wire s0n5340,s1n5340,notn5340;
or (n5340,s0n5340,s1n5340);
not(notn5340,n5014);
and (s0n5340,notn5340,n5341);
and (s1n5340,n5014,n5338);
and (n5342,n5343,n5038);
wire s0n5343,s1n5343,notn5343;
or (n5343,s0n5343,s1n5343);
not(notn5343,n5014);
and (s0n5343,notn5343,n5344);
and (s1n5343,n5014,n5341);
and (n5345,n5346,n2730);
or (n5346,1'b0,n5347,n5350,n5353,n5356);
and (n5347,n5348,n5016);
wire s0n5348,s1n5348,notn5348;
or (n5348,s0n5348,s1n5348);
not(notn5348,n5014);
and (s0n5348,notn5348,n5349);
and (s1n5348,n5014,n5344);
and (n5350,n5351,n5028);
wire s0n5351,s1n5351,notn5351;
or (n5351,s0n5351,s1n5351);
not(notn5351,n5014);
and (s0n5351,notn5351,n5352);
and (s1n5351,n5014,n5349);
and (n5353,n5354,n5033);
wire s0n5354,s1n5354,notn5354;
or (n5354,s0n5354,s1n5354);
not(notn5354,n5014);
and (s0n5354,notn5354,n5355);
and (s1n5354,n5014,n5352);
and (n5356,n5357,n5038);
wire s0n5357,s1n5357,notn5357;
or (n5357,s0n5357,s1n5357);
not(notn5357,n5014);
and (s0n5357,notn5357,n5358);
and (s1n5357,n5014,n5355);
and (n5359,n5360,n2742);
or (n5360,1'b0,n5361,n5365,n5368,n5371);
and (n5361,n5362,n5016);
wire s0n5362,s1n5362,notn5362;
or (n5362,s0n5362,s1n5362);
not(notn5362,n5014);
and (s0n5362,notn5362,n5363);
and (s1n5362,n5014,n5364);
and (n5365,n5366,n5028);
wire s0n5366,s1n5366,notn5366;
or (n5366,s0n5366,s1n5366);
not(notn5366,n5014);
and (s0n5366,notn5366,n5367);
and (s1n5366,n5014,n5363);
and (n5368,n5369,n5033);
wire s0n5369,s1n5369,notn5369;
or (n5369,s0n5369,s1n5369);
not(notn5369,n5014);
and (s0n5369,notn5369,n5370);
and (s1n5369,n5014,n5367);
and (n5371,n5372,n5038);
wire s0n5372,s1n5372,notn5372;
or (n5372,s0n5372,s1n5372);
not(notn5372,n5014);
and (s0n5372,notn5372,n5373);
and (s1n5372,n5014,n5370);
and (n5374,n5375,n2752);
or (n5375,1'b0,n5376,n5379,n5382,n5385);
and (n5376,n5377,n5016);
wire s0n5377,s1n5377,notn5377;
or (n5377,s0n5377,s1n5377);
not(notn5377,n5014);
and (s0n5377,notn5377,n5378);
and (s1n5377,n5014,n5373);
and (n5379,n5380,n5028);
wire s0n5380,s1n5380,notn5380;
or (n5380,s0n5380,s1n5380);
not(notn5380,n5014);
and (s0n5380,notn5380,n5381);
and (s1n5380,n5014,n5378);
and (n5382,n5383,n5033);
wire s0n5383,s1n5383,notn5383;
or (n5383,s0n5383,s1n5383);
not(notn5383,n5014);
and (s0n5383,notn5383,n5384);
and (s1n5383,n5014,n5381);
and (n5385,n5386,n5038);
wire s0n5386,s1n5386,notn5386;
or (n5386,s0n5386,s1n5386);
not(notn5386,n5014);
and (s0n5386,notn5386,n5387);
and (s1n5386,n5014,n5384);
and (n5389,n5328,n5390);
or (n5390,n5391,n5512,n6006);
and (n5391,n5392,n5451);
wire s0n5392,s1n5392,notn5392;
or (n5392,s0n5392,s1n5392);
not(notn5392,n4966);
and (s0n5392,notn5392,n5393);
and (s1n5392,n4966,n5450);
or (n5393,1'b0,n5394,n5409,n5423,n5438);
and (n5394,n5395,n2718);
or (n5395,1'b0,n5396,n5400,n5403,n5406);
and (n5396,n5397,n5016);
wire s0n5397,s1n5397,notn5397;
or (n5397,s0n5397,s1n5397);
not(notn5397,n5014);
and (s0n5397,notn5397,n5398);
and (s1n5397,n5014,n5399);
and (n5400,n5401,n5028);
wire s0n5401,s1n5401,notn5401;
or (n5401,s0n5401,s1n5401);
not(notn5401,n5014);
and (s0n5401,notn5401,n5402);
and (s1n5401,n5014,n5398);
and (n5403,n5404,n5033);
wire s0n5404,s1n5404,notn5404;
or (n5404,s0n5404,s1n5404);
not(notn5404,n5014);
and (s0n5404,notn5404,n5405);
and (s1n5404,n5014,n5402);
and (n5406,n5407,n5038);
wire s0n5407,s1n5407,notn5407;
or (n5407,s0n5407,s1n5407);
not(notn5407,n5014);
and (s0n5407,notn5407,n5408);
and (s1n5407,n5014,n5405);
and (n5409,n5410,n2730);
or (n5410,1'b0,n5411,n5414,n5417,n5420);
and (n5411,n5412,n5016);
wire s0n5412,s1n5412,notn5412;
or (n5412,s0n5412,s1n5412);
not(notn5412,n5014);
and (s0n5412,notn5412,n5413);
and (s1n5412,n5014,n5408);
and (n5414,n5415,n5028);
wire s0n5415,s1n5415,notn5415;
or (n5415,s0n5415,s1n5415);
not(notn5415,n5014);
and (s0n5415,notn5415,n5416);
and (s1n5415,n5014,n5413);
and (n5417,n5418,n5033);
wire s0n5418,s1n5418,notn5418;
or (n5418,s0n5418,s1n5418);
not(notn5418,n5014);
and (s0n5418,notn5418,n5419);
and (s1n5418,n5014,n5416);
and (n5420,n5421,n5038);
wire s0n5421,s1n5421,notn5421;
or (n5421,s0n5421,s1n5421);
not(notn5421,n5014);
and (s0n5421,notn5421,n5422);
and (s1n5421,n5014,n5419);
and (n5423,n5424,n2742);
or (n5424,1'b0,n5425,n5429,n5432,n5435);
and (n5425,n5426,n5016);
wire s0n5426,s1n5426,notn5426;
or (n5426,s0n5426,s1n5426);
not(notn5426,n5014);
and (s0n5426,notn5426,n5427);
and (s1n5426,n5014,n5428);
and (n5429,n5430,n5028);
wire s0n5430,s1n5430,notn5430;
or (n5430,s0n5430,s1n5430);
not(notn5430,n5014);
and (s0n5430,notn5430,n5431);
and (s1n5430,n5014,n5427);
and (n5432,n5433,n5033);
wire s0n5433,s1n5433,notn5433;
or (n5433,s0n5433,s1n5433);
not(notn5433,n5014);
and (s0n5433,notn5433,n5434);
and (s1n5433,n5014,n5431);
and (n5435,n5436,n5038);
wire s0n5436,s1n5436,notn5436;
or (n5436,s0n5436,s1n5436);
not(notn5436,n5014);
and (s0n5436,notn5436,n5437);
and (s1n5436,n5014,n5434);
and (n5438,n5439,n2752);
or (n5439,1'b0,n5440,n5443,n5446,n5448);
and (n5440,n5441,n5016);
wire s0n5441,s1n5441,notn5441;
or (n5441,s0n5441,s1n5441);
not(notn5441,n5014);
and (s0n5441,notn5441,n5442);
and (s1n5441,n5014,n5437);
and (n5443,n5444,n5028);
wire s0n5444,s1n5444,notn5444;
or (n5444,s0n5444,s1n5444);
not(notn5444,n5014);
and (s0n5444,notn5444,n5445);
and (s1n5444,n5014,n5442);
and (n5446,n5447,n5033);
wire s0n5447,s1n5447,notn5447;
or (n5447,s0n5447,s1n5447);
not(notn5447,n5014);
and (s0n5447,notn5447,n1303);
and (s1n5447,n5014,n5445);
and (n5448,n5449,n5038);
wire s0n5449,s1n5449,notn5449;
or (n5449,s0n5449,s1n5449);
not(notn5449,n5014);
and (s0n5449,notn5449,n799);
and (s1n5449,n5014,n1303);
wire s0n5451,s1n5451,notn5451;
or (n5451,s0n5451,s1n5451);
not(notn5451,n4966);
and (s0n5451,notn5451,n5452);
and (s1n5451,n4966,n5511);
or (n5452,1'b0,n5453,n5468,n5482,n5497);
and (n5453,n5454,n2718);
or (n5454,1'b0,n5455,n5459,n5462,n5465);
and (n5455,n5456,n5016);
wire s0n5456,s1n5456,notn5456;
or (n5456,s0n5456,s1n5456);
not(notn5456,n5014);
and (s0n5456,notn5456,n5457);
and (s1n5456,n5014,n5458);
and (n5459,n5460,n5028);
wire s0n5460,s1n5460,notn5460;
or (n5460,s0n5460,s1n5460);
not(notn5460,n5014);
and (s0n5460,notn5460,n5461);
and (s1n5460,n5014,n5457);
and (n5462,n5463,n5033);
wire s0n5463,s1n5463,notn5463;
or (n5463,s0n5463,s1n5463);
not(notn5463,n5014);
and (s0n5463,notn5463,n5464);
and (s1n5463,n5014,n5461);
and (n5465,n5466,n5038);
wire s0n5466,s1n5466,notn5466;
or (n5466,s0n5466,s1n5466);
not(notn5466,n5014);
and (s0n5466,notn5466,n5467);
and (s1n5466,n5014,n5464);
and (n5468,n5469,n2730);
or (n5469,1'b0,n5470,n5473,n5476,n5479);
and (n5470,n5471,n5016);
wire s0n5471,s1n5471,notn5471;
or (n5471,s0n5471,s1n5471);
not(notn5471,n5014);
and (s0n5471,notn5471,n5472);
and (s1n5471,n5014,n5467);
and (n5473,n5474,n5028);
wire s0n5474,s1n5474,notn5474;
or (n5474,s0n5474,s1n5474);
not(notn5474,n5014);
and (s0n5474,notn5474,n5475);
and (s1n5474,n5014,n5472);
and (n5476,n5477,n5033);
wire s0n5477,s1n5477,notn5477;
or (n5477,s0n5477,s1n5477);
not(notn5477,n5014);
and (s0n5477,notn5477,n5478);
and (s1n5477,n5014,n5475);
and (n5479,n5480,n5038);
wire s0n5480,s1n5480,notn5480;
or (n5480,s0n5480,s1n5480);
not(notn5480,n5014);
and (s0n5480,notn5480,n5481);
and (s1n5480,n5014,n5478);
and (n5482,n5483,n2742);
or (n5483,1'b0,n5484,n5488,n5491,n5494);
and (n5484,n5485,n5016);
wire s0n5485,s1n5485,notn5485;
or (n5485,s0n5485,s1n5485);
not(notn5485,n5014);
and (s0n5485,notn5485,n5486);
and (s1n5485,n5014,n5487);
and (n5488,n5489,n5028);
wire s0n5489,s1n5489,notn5489;
or (n5489,s0n5489,s1n5489);
not(notn5489,n5014);
and (s0n5489,notn5489,n5490);
and (s1n5489,n5014,n5486);
and (n5491,n5492,n5033);
wire s0n5492,s1n5492,notn5492;
or (n5492,s0n5492,s1n5492);
not(notn5492,n5014);
and (s0n5492,notn5492,n5493);
and (s1n5492,n5014,n5490);
and (n5494,n5495,n5038);
wire s0n5495,s1n5495,notn5495;
or (n5495,s0n5495,s1n5495);
not(notn5495,n5014);
and (s0n5495,notn5495,n5496);
and (s1n5495,n5014,n5493);
and (n5497,n5498,n2752);
or (n5498,1'b0,n5499,n5502,n5505,n5508);
and (n5499,n5500,n5016);
wire s0n5500,s1n5500,notn5500;
or (n5500,s0n5500,s1n5500);
not(notn5500,n5014);
and (s0n5500,notn5500,n5501);
and (s1n5500,n5014,n5496);
and (n5502,n5503,n5028);
wire s0n5503,s1n5503,notn5503;
or (n5503,s0n5503,s1n5503);
not(notn5503,n5014);
and (s0n5503,notn5503,n5504);
and (s1n5503,n5014,n5501);
and (n5505,n5506,n5033);
wire s0n5506,s1n5506,notn5506;
or (n5506,s0n5506,s1n5506);
not(notn5506,n5014);
and (s0n5506,notn5506,n5507);
and (s1n5506,n5014,n5504);
and (n5508,n5509,n5038);
wire s0n5509,s1n5509,notn5509;
or (n5509,s0n5509,s1n5509);
not(notn5509,n5014);
and (s0n5509,notn5509,n5510);
and (s1n5509,n5014,n5507);
and (n5512,n5451,n5513);
or (n5513,n5514,n5635,n6005);
and (n5514,n5515,n5574);
wire s0n5515,s1n5515,notn5515;
or (n5515,s0n5515,s1n5515);
not(notn5515,n4966);
and (s0n5515,notn5515,n5516);
and (s1n5515,n4966,n5573);
or (n5516,1'b0,n5517,n5532,n5546,n5561);
and (n5517,n5518,n2718);
or (n5518,1'b0,n5519,n5523,n5526,n5529);
and (n5519,n5520,n5016);
wire s0n5520,s1n5520,notn5520;
or (n5520,s0n5520,s1n5520);
not(notn5520,n5014);
and (s0n5520,notn5520,n5521);
and (s1n5520,n5014,n5522);
and (n5523,n5524,n5028);
wire s0n5524,s1n5524,notn5524;
or (n5524,s0n5524,s1n5524);
not(notn5524,n5014);
and (s0n5524,notn5524,n5525);
and (s1n5524,n5014,n5521);
and (n5526,n5527,n5033);
wire s0n5527,s1n5527,notn5527;
or (n5527,s0n5527,s1n5527);
not(notn5527,n5014);
and (s0n5527,notn5527,n5528);
and (s1n5527,n5014,n5525);
and (n5529,n5530,n5038);
wire s0n5530,s1n5530,notn5530;
or (n5530,s0n5530,s1n5530);
not(notn5530,n5014);
and (s0n5530,notn5530,n5531);
and (s1n5530,n5014,n5528);
and (n5532,n5533,n2730);
or (n5533,1'b0,n5534,n5537,n5540,n5543);
and (n5534,n5535,n5016);
wire s0n5535,s1n5535,notn5535;
or (n5535,s0n5535,s1n5535);
not(notn5535,n5014);
and (s0n5535,notn5535,n5536);
and (s1n5535,n5014,n5531);
and (n5537,n5538,n5028);
wire s0n5538,s1n5538,notn5538;
or (n5538,s0n5538,s1n5538);
not(notn5538,n5014);
and (s0n5538,notn5538,n5539);
and (s1n5538,n5014,n5536);
and (n5540,n5541,n5033);
wire s0n5541,s1n5541,notn5541;
or (n5541,s0n5541,s1n5541);
not(notn5541,n5014);
and (s0n5541,notn5541,n5542);
and (s1n5541,n5014,n5539);
and (n5543,n5544,n5038);
wire s0n5544,s1n5544,notn5544;
or (n5544,s0n5544,s1n5544);
not(notn5544,n5014);
and (s0n5544,notn5544,n5545);
and (s1n5544,n5014,n5542);
and (n5546,n5547,n2742);
or (n5547,1'b0,n5548,n5552,n5555,n5558);
and (n5548,n5549,n5016);
wire s0n5549,s1n5549,notn5549;
or (n5549,s0n5549,s1n5549);
not(notn5549,n5014);
and (s0n5549,notn5549,n5550);
and (s1n5549,n5014,n5551);
and (n5552,n5553,n5028);
wire s0n5553,s1n5553,notn5553;
or (n5553,s0n5553,s1n5553);
not(notn5553,n5014);
and (s0n5553,notn5553,n5554);
and (s1n5553,n5014,n5550);
and (n5555,n5556,n5033);
wire s0n5556,s1n5556,notn5556;
or (n5556,s0n5556,s1n5556);
not(notn5556,n5014);
and (s0n5556,notn5556,n5557);
and (s1n5556,n5014,n5554);
and (n5558,n5559,n5038);
wire s0n5559,s1n5559,notn5559;
or (n5559,s0n5559,s1n5559);
not(notn5559,n5014);
and (s0n5559,notn5559,n5560);
and (s1n5559,n5014,n5557);
and (n5561,n5562,n2752);
or (n5562,1'b0,n5563,n5566,n5569,n5571);
and (n5563,n5564,n5016);
wire s0n5564,s1n5564,notn5564;
or (n5564,s0n5564,s1n5564);
not(notn5564,n5014);
and (s0n5564,notn5564,n5565);
and (s1n5564,n5014,n5560);
and (n5566,n5567,n5028);
wire s0n5567,s1n5567,notn5567;
or (n5567,s0n5567,s1n5567);
not(notn5567,n5014);
and (s0n5567,notn5567,n5568);
and (s1n5567,n5014,n5565);
and (n5569,n5570,n5033);
wire s0n5570,s1n5570,notn5570;
or (n5570,s0n5570,s1n5570);
not(notn5570,n5014);
and (s0n5570,notn5570,n1319);
and (s1n5570,n5014,n5568);
and (n5571,n5572,n5038);
wire s0n5572,s1n5572,notn5572;
or (n5572,s0n5572,s1n5572);
not(notn5572,n5014);
and (s0n5572,notn5572,n815);
and (s1n5572,n5014,n1319);
wire s0n5574,s1n5574,notn5574;
or (n5574,s0n5574,s1n5574);
not(notn5574,n4966);
and (s0n5574,notn5574,n5575);
and (s1n5574,n4966,n5634);
or (n5575,1'b0,n5576,n5591,n5605,n5620);
and (n5576,n5577,n2718);
or (n5577,1'b0,n5578,n5582,n5585,n5588);
and (n5578,n5579,n5016);
wire s0n5579,s1n5579,notn5579;
or (n5579,s0n5579,s1n5579);
not(notn5579,n5014);
and (s0n5579,notn5579,n5580);
and (s1n5579,n5014,n5581);
and (n5582,n5583,n5028);
wire s0n5583,s1n5583,notn5583;
or (n5583,s0n5583,s1n5583);
not(notn5583,n5014);
and (s0n5583,notn5583,n5584);
and (s1n5583,n5014,n5580);
and (n5585,n5586,n5033);
wire s0n5586,s1n5586,notn5586;
or (n5586,s0n5586,s1n5586);
not(notn5586,n5014);
and (s0n5586,notn5586,n5587);
and (s1n5586,n5014,n5584);
and (n5588,n5589,n5038);
wire s0n5589,s1n5589,notn5589;
or (n5589,s0n5589,s1n5589);
not(notn5589,n5014);
and (s0n5589,notn5589,n5590);
and (s1n5589,n5014,n5587);
and (n5591,n5592,n2730);
or (n5592,1'b0,n5593,n5596,n5599,n5602);
and (n5593,n5594,n5016);
wire s0n5594,s1n5594,notn5594;
or (n5594,s0n5594,s1n5594);
not(notn5594,n5014);
and (s0n5594,notn5594,n5595);
and (s1n5594,n5014,n5590);
and (n5596,n5597,n5028);
wire s0n5597,s1n5597,notn5597;
or (n5597,s0n5597,s1n5597);
not(notn5597,n5014);
and (s0n5597,notn5597,n5598);
and (s1n5597,n5014,n5595);
and (n5599,n5600,n5033);
wire s0n5600,s1n5600,notn5600;
or (n5600,s0n5600,s1n5600);
not(notn5600,n5014);
and (s0n5600,notn5600,n5601);
and (s1n5600,n5014,n5598);
and (n5602,n5603,n5038);
wire s0n5603,s1n5603,notn5603;
or (n5603,s0n5603,s1n5603);
not(notn5603,n5014);
and (s0n5603,notn5603,n5604);
and (s1n5603,n5014,n5601);
and (n5605,n5606,n2742);
or (n5606,1'b0,n5607,n5611,n5614,n5617);
and (n5607,n5608,n5016);
wire s0n5608,s1n5608,notn5608;
or (n5608,s0n5608,s1n5608);
not(notn5608,n5014);
and (s0n5608,notn5608,n5609);
and (s1n5608,n5014,n5610);
and (n5611,n5612,n5028);
wire s0n5612,s1n5612,notn5612;
or (n5612,s0n5612,s1n5612);
not(notn5612,n5014);
and (s0n5612,notn5612,n5613);
and (s1n5612,n5014,n5609);
and (n5614,n5615,n5033);
wire s0n5615,s1n5615,notn5615;
or (n5615,s0n5615,s1n5615);
not(notn5615,n5014);
and (s0n5615,notn5615,n5616);
and (s1n5615,n5014,n5613);
and (n5617,n5618,n5038);
wire s0n5618,s1n5618,notn5618;
or (n5618,s0n5618,s1n5618);
not(notn5618,n5014);
and (s0n5618,notn5618,n5619);
and (s1n5618,n5014,n5616);
and (n5620,n5621,n2752);
or (n5621,1'b0,n5622,n5625,n5628,n5631);
and (n5622,n5623,n5016);
wire s0n5623,s1n5623,notn5623;
or (n5623,s0n5623,s1n5623);
not(notn5623,n5014);
and (s0n5623,notn5623,n5624);
and (s1n5623,n5014,n5619);
and (n5625,n5626,n5028);
wire s0n5626,s1n5626,notn5626;
or (n5626,s0n5626,s1n5626);
not(notn5626,n5014);
and (s0n5626,notn5626,n5627);
and (s1n5626,n5014,n5624);
and (n5628,n5629,n5033);
wire s0n5629,s1n5629,notn5629;
or (n5629,s0n5629,s1n5629);
not(notn5629,n5014);
and (s0n5629,notn5629,n5630);
and (s1n5629,n5014,n5627);
and (n5631,n5632,n5038);
wire s0n5632,s1n5632,notn5632;
or (n5632,s0n5632,s1n5632);
not(notn5632,n5014);
and (s0n5632,notn5632,n5633);
and (s1n5632,n5014,n5630);
and (n5635,n5574,n5636);
or (n5636,n5637,n5758,n6004);
and (n5637,n5638,n5697);
wire s0n5638,s1n5638,notn5638;
or (n5638,s0n5638,s1n5638);
not(notn5638,n4966);
and (s0n5638,notn5638,n5639);
and (s1n5638,n4966,n5696);
or (n5639,1'b0,n5640,n5655,n5669,n5684);
and (n5640,n5641,n2718);
or (n5641,1'b0,n5642,n5646,n5649,n5652);
and (n5642,n5643,n5016);
wire s0n5643,s1n5643,notn5643;
or (n5643,s0n5643,s1n5643);
not(notn5643,n5014);
and (s0n5643,notn5643,n5644);
and (s1n5643,n5014,n5645);
and (n5646,n5647,n5028);
wire s0n5647,s1n5647,notn5647;
or (n5647,s0n5647,s1n5647);
not(notn5647,n5014);
and (s0n5647,notn5647,n5648);
and (s1n5647,n5014,n5644);
and (n5649,n5650,n5033);
wire s0n5650,s1n5650,notn5650;
or (n5650,s0n5650,s1n5650);
not(notn5650,n5014);
and (s0n5650,notn5650,n5651);
and (s1n5650,n5014,n5648);
and (n5652,n5653,n5038);
wire s0n5653,s1n5653,notn5653;
or (n5653,s0n5653,s1n5653);
not(notn5653,n5014);
and (s0n5653,notn5653,n5654);
and (s1n5653,n5014,n5651);
and (n5655,n5656,n2730);
or (n5656,1'b0,n5657,n5660,n5663,n5666);
and (n5657,n5658,n5016);
wire s0n5658,s1n5658,notn5658;
or (n5658,s0n5658,s1n5658);
not(notn5658,n5014);
and (s0n5658,notn5658,n5659);
and (s1n5658,n5014,n5654);
and (n5660,n5661,n5028);
wire s0n5661,s1n5661,notn5661;
or (n5661,s0n5661,s1n5661);
not(notn5661,n5014);
and (s0n5661,notn5661,n5662);
and (s1n5661,n5014,n5659);
and (n5663,n5664,n5033);
wire s0n5664,s1n5664,notn5664;
or (n5664,s0n5664,s1n5664);
not(notn5664,n5014);
and (s0n5664,notn5664,n5665);
and (s1n5664,n5014,n5662);
and (n5666,n5667,n5038);
wire s0n5667,s1n5667,notn5667;
or (n5667,s0n5667,s1n5667);
not(notn5667,n5014);
and (s0n5667,notn5667,n5668);
and (s1n5667,n5014,n5665);
and (n5669,n5670,n2742);
or (n5670,1'b0,n5671,n5675,n5678,n5681);
and (n5671,n5672,n5016);
wire s0n5672,s1n5672,notn5672;
or (n5672,s0n5672,s1n5672);
not(notn5672,n5014);
and (s0n5672,notn5672,n5673);
and (s1n5672,n5014,n5674);
and (n5675,n5676,n5028);
wire s0n5676,s1n5676,notn5676;
or (n5676,s0n5676,s1n5676);
not(notn5676,n5014);
and (s0n5676,notn5676,n5677);
and (s1n5676,n5014,n5673);
and (n5678,n5679,n5033);
wire s0n5679,s1n5679,notn5679;
or (n5679,s0n5679,s1n5679);
not(notn5679,n5014);
and (s0n5679,notn5679,n5680);
and (s1n5679,n5014,n5677);
and (n5681,n5682,n5038);
wire s0n5682,s1n5682,notn5682;
or (n5682,s0n5682,s1n5682);
not(notn5682,n5014);
and (s0n5682,notn5682,n5683);
and (s1n5682,n5014,n5680);
and (n5684,n5685,n2752);
or (n5685,1'b0,n5686,n5689,n5692,n5694);
and (n5686,n5687,n5016);
wire s0n5687,s1n5687,notn5687;
or (n5687,s0n5687,s1n5687);
not(notn5687,n5014);
and (s0n5687,notn5687,n5688);
and (s1n5687,n5014,n5683);
and (n5689,n5690,n5028);
wire s0n5690,s1n5690,notn5690;
or (n5690,s0n5690,s1n5690);
not(notn5690,n5014);
and (s0n5690,notn5690,n5691);
and (s1n5690,n5014,n5688);
and (n5692,n5693,n5033);
wire s0n5693,s1n5693,notn5693;
or (n5693,s0n5693,s1n5693);
not(notn5693,n5014);
and (s0n5693,notn5693,n1335);
and (s1n5693,n5014,n5691);
and (n5694,n5695,n5038);
wire s0n5695,s1n5695,notn5695;
or (n5695,s0n5695,s1n5695);
not(notn5695,n5014);
and (s0n5695,notn5695,n831);
and (s1n5695,n5014,n1335);
wire s0n5697,s1n5697,notn5697;
or (n5697,s0n5697,s1n5697);
not(notn5697,n4966);
and (s0n5697,notn5697,n5698);
and (s1n5697,n4966,n5757);
or (n5698,1'b0,n5699,n5714,n5728,n5743);
and (n5699,n5700,n2718);
or (n5700,1'b0,n5701,n5705,n5708,n5711);
and (n5701,n5702,n5016);
wire s0n5702,s1n5702,notn5702;
or (n5702,s0n5702,s1n5702);
not(notn5702,n5014);
and (s0n5702,notn5702,n5703);
and (s1n5702,n5014,n5704);
and (n5705,n5706,n5028);
wire s0n5706,s1n5706,notn5706;
or (n5706,s0n5706,s1n5706);
not(notn5706,n5014);
and (s0n5706,notn5706,n5707);
and (s1n5706,n5014,n5703);
and (n5708,n5709,n5033);
wire s0n5709,s1n5709,notn5709;
or (n5709,s0n5709,s1n5709);
not(notn5709,n5014);
and (s0n5709,notn5709,n5710);
and (s1n5709,n5014,n5707);
and (n5711,n5712,n5038);
wire s0n5712,s1n5712,notn5712;
or (n5712,s0n5712,s1n5712);
not(notn5712,n5014);
and (s0n5712,notn5712,n5713);
and (s1n5712,n5014,n5710);
and (n5714,n5715,n2730);
or (n5715,1'b0,n5716,n5719,n5722,n5725);
and (n5716,n5717,n5016);
wire s0n5717,s1n5717,notn5717;
or (n5717,s0n5717,s1n5717);
not(notn5717,n5014);
and (s0n5717,notn5717,n5718);
and (s1n5717,n5014,n5713);
and (n5719,n5720,n5028);
wire s0n5720,s1n5720,notn5720;
or (n5720,s0n5720,s1n5720);
not(notn5720,n5014);
and (s0n5720,notn5720,n5721);
and (s1n5720,n5014,n5718);
and (n5722,n5723,n5033);
wire s0n5723,s1n5723,notn5723;
or (n5723,s0n5723,s1n5723);
not(notn5723,n5014);
and (s0n5723,notn5723,n5724);
and (s1n5723,n5014,n5721);
and (n5725,n5726,n5038);
wire s0n5726,s1n5726,notn5726;
or (n5726,s0n5726,s1n5726);
not(notn5726,n5014);
and (s0n5726,notn5726,n5727);
and (s1n5726,n5014,n5724);
and (n5728,n5729,n2742);
or (n5729,1'b0,n5730,n5734,n5737,n5740);
and (n5730,n5731,n5016);
wire s0n5731,s1n5731,notn5731;
or (n5731,s0n5731,s1n5731);
not(notn5731,n5014);
and (s0n5731,notn5731,n5732);
and (s1n5731,n5014,n5733);
and (n5734,n5735,n5028);
wire s0n5735,s1n5735,notn5735;
or (n5735,s0n5735,s1n5735);
not(notn5735,n5014);
and (s0n5735,notn5735,n5736);
and (s1n5735,n5014,n5732);
and (n5737,n5738,n5033);
wire s0n5738,s1n5738,notn5738;
or (n5738,s0n5738,s1n5738);
not(notn5738,n5014);
and (s0n5738,notn5738,n5739);
and (s1n5738,n5014,n5736);
and (n5740,n5741,n5038);
wire s0n5741,s1n5741,notn5741;
or (n5741,s0n5741,s1n5741);
not(notn5741,n5014);
and (s0n5741,notn5741,n5742);
and (s1n5741,n5014,n5739);
and (n5743,n5744,n2752);
or (n5744,1'b0,n5745,n5748,n5751,n5754);
and (n5745,n5746,n5016);
wire s0n5746,s1n5746,notn5746;
or (n5746,s0n5746,s1n5746);
not(notn5746,n5014);
and (s0n5746,notn5746,n5747);
and (s1n5746,n5014,n5742);
and (n5748,n5749,n5028);
wire s0n5749,s1n5749,notn5749;
or (n5749,s0n5749,s1n5749);
not(notn5749,n5014);
and (s0n5749,notn5749,n5750);
and (s1n5749,n5014,n5747);
and (n5751,n5752,n5033);
wire s0n5752,s1n5752,notn5752;
or (n5752,s0n5752,s1n5752);
not(notn5752,n5014);
and (s0n5752,notn5752,n5753);
and (s1n5752,n5014,n5750);
and (n5754,n5755,n5038);
wire s0n5755,s1n5755,notn5755;
or (n5755,s0n5755,s1n5755);
not(notn5755,n5014);
and (s0n5755,notn5755,n5756);
and (s1n5755,n5014,n5753);
and (n5758,n5697,n5759);
or (n5759,n5760,n5881,n6003);
and (n5760,n5761,n5820);
wire s0n5761,s1n5761,notn5761;
or (n5761,s0n5761,s1n5761);
not(notn5761,n4966);
and (s0n5761,notn5761,n5762);
and (s1n5761,n4966,n5819);
or (n5762,1'b0,n5763,n5778,n5792,n5807);
and (n5763,n5764,n2718);
or (n5764,1'b0,n5765,n5769,n5772,n5775);
and (n5765,n5766,n5016);
wire s0n5766,s1n5766,notn5766;
or (n5766,s0n5766,s1n5766);
not(notn5766,n5014);
and (s0n5766,notn5766,n5767);
and (s1n5766,n5014,n5768);
and (n5769,n5770,n5028);
wire s0n5770,s1n5770,notn5770;
or (n5770,s0n5770,s1n5770);
not(notn5770,n5014);
and (s0n5770,notn5770,n5771);
and (s1n5770,n5014,n5767);
and (n5772,n5773,n5033);
wire s0n5773,s1n5773,notn5773;
or (n5773,s0n5773,s1n5773);
not(notn5773,n5014);
and (s0n5773,notn5773,n5774);
and (s1n5773,n5014,n5771);
and (n5775,n5776,n5038);
wire s0n5776,s1n5776,notn5776;
or (n5776,s0n5776,s1n5776);
not(notn5776,n5014);
and (s0n5776,notn5776,n5777);
and (s1n5776,n5014,n5774);
and (n5778,n5779,n2730);
or (n5779,1'b0,n5780,n5783,n5786,n5789);
and (n5780,n5781,n5016);
wire s0n5781,s1n5781,notn5781;
or (n5781,s0n5781,s1n5781);
not(notn5781,n5014);
and (s0n5781,notn5781,n5782);
and (s1n5781,n5014,n5777);
and (n5783,n5784,n5028);
wire s0n5784,s1n5784,notn5784;
or (n5784,s0n5784,s1n5784);
not(notn5784,n5014);
and (s0n5784,notn5784,n5785);
and (s1n5784,n5014,n5782);
and (n5786,n5787,n5033);
wire s0n5787,s1n5787,notn5787;
or (n5787,s0n5787,s1n5787);
not(notn5787,n5014);
and (s0n5787,notn5787,n5788);
and (s1n5787,n5014,n5785);
and (n5789,n5790,n5038);
wire s0n5790,s1n5790,notn5790;
or (n5790,s0n5790,s1n5790);
not(notn5790,n5014);
and (s0n5790,notn5790,n5791);
and (s1n5790,n5014,n5788);
and (n5792,n5793,n2742);
or (n5793,1'b0,n5794,n5798,n5801,n5804);
and (n5794,n5795,n5016);
wire s0n5795,s1n5795,notn5795;
or (n5795,s0n5795,s1n5795);
not(notn5795,n5014);
and (s0n5795,notn5795,n5796);
and (s1n5795,n5014,n5797);
and (n5798,n5799,n5028);
wire s0n5799,s1n5799,notn5799;
or (n5799,s0n5799,s1n5799);
not(notn5799,n5014);
and (s0n5799,notn5799,n5800);
and (s1n5799,n5014,n5796);
and (n5801,n5802,n5033);
wire s0n5802,s1n5802,notn5802;
or (n5802,s0n5802,s1n5802);
not(notn5802,n5014);
and (s0n5802,notn5802,n5803);
and (s1n5802,n5014,n5800);
and (n5804,n5805,n5038);
wire s0n5805,s1n5805,notn5805;
or (n5805,s0n5805,s1n5805);
not(notn5805,n5014);
and (s0n5805,notn5805,n5806);
and (s1n5805,n5014,n5803);
and (n5807,n5808,n2752);
or (n5808,1'b0,n5809,n5812,n5815,n5817);
and (n5809,n5810,n5016);
wire s0n5810,s1n5810,notn5810;
or (n5810,s0n5810,s1n5810);
not(notn5810,n5014);
and (s0n5810,notn5810,n5811);
and (s1n5810,n5014,n5806);
and (n5812,n5813,n5028);
wire s0n5813,s1n5813,notn5813;
or (n5813,s0n5813,s1n5813);
not(notn5813,n5014);
and (s0n5813,notn5813,n5814);
and (s1n5813,n5014,n5811);
and (n5815,n5816,n5033);
wire s0n5816,s1n5816,notn5816;
or (n5816,s0n5816,s1n5816);
not(notn5816,n5014);
and (s0n5816,notn5816,n1351);
and (s1n5816,n5014,n5814);
and (n5817,n5818,n5038);
wire s0n5818,s1n5818,notn5818;
or (n5818,s0n5818,s1n5818);
not(notn5818,n5014);
and (s0n5818,notn5818,n847);
and (s1n5818,n5014,n1351);
wire s0n5820,s1n5820,notn5820;
or (n5820,s0n5820,s1n5820);
not(notn5820,n4966);
and (s0n5820,notn5820,n5821);
and (s1n5820,n4966,n5880);
or (n5821,1'b0,n5822,n5837,n5851,n5866);
and (n5822,n5823,n2718);
or (n5823,1'b0,n5824,n5828,n5831,n5834);
and (n5824,n5825,n5016);
wire s0n5825,s1n5825,notn5825;
or (n5825,s0n5825,s1n5825);
not(notn5825,n5014);
and (s0n5825,notn5825,n5826);
and (s1n5825,n5014,n5827);
and (n5828,n5829,n5028);
wire s0n5829,s1n5829,notn5829;
or (n5829,s0n5829,s1n5829);
not(notn5829,n5014);
and (s0n5829,notn5829,n5830);
and (s1n5829,n5014,n5826);
and (n5831,n5832,n5033);
wire s0n5832,s1n5832,notn5832;
or (n5832,s0n5832,s1n5832);
not(notn5832,n5014);
and (s0n5832,notn5832,n5833);
and (s1n5832,n5014,n5830);
and (n5834,n5835,n5038);
wire s0n5835,s1n5835,notn5835;
or (n5835,s0n5835,s1n5835);
not(notn5835,n5014);
and (s0n5835,notn5835,n5836);
and (s1n5835,n5014,n5833);
and (n5837,n5838,n2730);
or (n5838,1'b0,n5839,n5842,n5845,n5848);
and (n5839,n5840,n5016);
wire s0n5840,s1n5840,notn5840;
or (n5840,s0n5840,s1n5840);
not(notn5840,n5014);
and (s0n5840,notn5840,n5841);
and (s1n5840,n5014,n5836);
and (n5842,n5843,n5028);
wire s0n5843,s1n5843,notn5843;
or (n5843,s0n5843,s1n5843);
not(notn5843,n5014);
and (s0n5843,notn5843,n5844);
and (s1n5843,n5014,n5841);
and (n5845,n5846,n5033);
wire s0n5846,s1n5846,notn5846;
or (n5846,s0n5846,s1n5846);
not(notn5846,n5014);
and (s0n5846,notn5846,n5847);
and (s1n5846,n5014,n5844);
and (n5848,n5849,n5038);
wire s0n5849,s1n5849,notn5849;
or (n5849,s0n5849,s1n5849);
not(notn5849,n5014);
and (s0n5849,notn5849,n5850);
and (s1n5849,n5014,n5847);
and (n5851,n5852,n2742);
or (n5852,1'b0,n5853,n5857,n5860,n5863);
and (n5853,n5854,n5016);
wire s0n5854,s1n5854,notn5854;
or (n5854,s0n5854,s1n5854);
not(notn5854,n5014);
and (s0n5854,notn5854,n5855);
and (s1n5854,n5014,n5856);
and (n5857,n5858,n5028);
wire s0n5858,s1n5858,notn5858;
or (n5858,s0n5858,s1n5858);
not(notn5858,n5014);
and (s0n5858,notn5858,n5859);
and (s1n5858,n5014,n5855);
and (n5860,n5861,n5033);
wire s0n5861,s1n5861,notn5861;
or (n5861,s0n5861,s1n5861);
not(notn5861,n5014);
and (s0n5861,notn5861,n5862);
and (s1n5861,n5014,n5859);
and (n5863,n5864,n5038);
wire s0n5864,s1n5864,notn5864;
or (n5864,s0n5864,s1n5864);
not(notn5864,n5014);
and (s0n5864,notn5864,n5865);
and (s1n5864,n5014,n5862);
and (n5866,n5867,n2752);
or (n5867,1'b0,n5868,n5871,n5874,n5877);
and (n5868,n5869,n5016);
wire s0n5869,s1n5869,notn5869;
or (n5869,s0n5869,s1n5869);
not(notn5869,n5014);
and (s0n5869,notn5869,n5870);
and (s1n5869,n5014,n5865);
and (n5871,n5872,n5028);
wire s0n5872,s1n5872,notn5872;
or (n5872,s0n5872,s1n5872);
not(notn5872,n5014);
and (s0n5872,notn5872,n5873);
and (s1n5872,n5014,n5870);
and (n5874,n5875,n5033);
wire s0n5875,s1n5875,notn5875;
or (n5875,s0n5875,s1n5875);
not(notn5875,n5014);
and (s0n5875,notn5875,n5876);
and (s1n5875,n5014,n5873);
and (n5877,n5878,n5038);
wire s0n5878,s1n5878,notn5878;
or (n5878,s0n5878,s1n5878);
not(notn5878,n5014);
and (s0n5878,notn5878,n5879);
and (s1n5878,n5014,n5876);
and (n5881,n5820,n5882);
and (n5882,n5883,n5942);
wire s0n5883,s1n5883,notn5883;
or (n5883,s0n5883,s1n5883);
not(notn5883,n4966);
and (s0n5883,notn5883,n5884);
and (s1n5883,n4966,n5941);
or (n5884,1'b0,n5885,n5900,n5914,n5929);
and (n5885,n5886,n2718);
or (n5886,1'b0,n5887,n5891,n5894,n5897);
and (n5887,n5888,n5016);
wire s0n5888,s1n5888,notn5888;
or (n5888,s0n5888,s1n5888);
not(notn5888,n5014);
and (s0n5888,notn5888,n5889);
and (s1n5888,n5014,n5890);
and (n5891,n5892,n5028);
wire s0n5892,s1n5892,notn5892;
or (n5892,s0n5892,s1n5892);
not(notn5892,n5014);
and (s0n5892,notn5892,n5893);
and (s1n5892,n5014,n5889);
and (n5894,n5895,n5033);
wire s0n5895,s1n5895,notn5895;
or (n5895,s0n5895,s1n5895);
not(notn5895,n5014);
and (s0n5895,notn5895,n5896);
and (s1n5895,n5014,n5893);
and (n5897,n5898,n5038);
wire s0n5898,s1n5898,notn5898;
or (n5898,s0n5898,s1n5898);
not(notn5898,n5014);
and (s0n5898,notn5898,n5899);
and (s1n5898,n5014,n5896);
and (n5900,n5901,n2730);
or (n5901,1'b0,n5902,n5905,n5908,n5911);
and (n5902,n5903,n5016);
wire s0n5903,s1n5903,notn5903;
or (n5903,s0n5903,s1n5903);
not(notn5903,n5014);
and (s0n5903,notn5903,n5904);
and (s1n5903,n5014,n5899);
and (n5905,n5906,n5028);
wire s0n5906,s1n5906,notn5906;
or (n5906,s0n5906,s1n5906);
not(notn5906,n5014);
and (s0n5906,notn5906,n5907);
and (s1n5906,n5014,n5904);
and (n5908,n5909,n5033);
wire s0n5909,s1n5909,notn5909;
or (n5909,s0n5909,s1n5909);
not(notn5909,n5014);
and (s0n5909,notn5909,n5910);
and (s1n5909,n5014,n5907);
and (n5911,n5912,n5038);
wire s0n5912,s1n5912,notn5912;
or (n5912,s0n5912,s1n5912);
not(notn5912,n5014);
and (s0n5912,notn5912,n5913);
and (s1n5912,n5014,n5910);
and (n5914,n5915,n2742);
or (n5915,1'b0,n5916,n5920,n5923,n5926);
and (n5916,n5917,n5016);
wire s0n5917,s1n5917,notn5917;
or (n5917,s0n5917,s1n5917);
not(notn5917,n5014);
and (s0n5917,notn5917,n5918);
and (s1n5917,n5014,n5919);
and (n5920,n5921,n5028);
wire s0n5921,s1n5921,notn5921;
or (n5921,s0n5921,s1n5921);
not(notn5921,n5014);
and (s0n5921,notn5921,n5922);
and (s1n5921,n5014,n5918);
and (n5923,n5924,n5033);
wire s0n5924,s1n5924,notn5924;
or (n5924,s0n5924,s1n5924);
not(notn5924,n5014);
and (s0n5924,notn5924,n5925);
and (s1n5924,n5014,n5922);
and (n5926,n5927,n5038);
wire s0n5927,s1n5927,notn5927;
or (n5927,s0n5927,s1n5927);
not(notn5927,n5014);
and (s0n5927,notn5927,n5928);
and (s1n5927,n5014,n5925);
and (n5929,n5930,n2752);
or (n5930,1'b0,n5931,n5934,n5937,n5939);
and (n5931,n5932,n5016);
wire s0n5932,s1n5932,notn5932;
or (n5932,s0n5932,s1n5932);
not(notn5932,n5014);
and (s0n5932,notn5932,n5933);
and (s1n5932,n5014,n5928);
and (n5934,n5935,n5028);
wire s0n5935,s1n5935,notn5935;
or (n5935,s0n5935,s1n5935);
not(notn5935,n5014);
and (s0n5935,notn5935,n5936);
and (s1n5935,n5014,n5933);
and (n5937,n5938,n5033);
wire s0n5938,s1n5938,notn5938;
or (n5938,s0n5938,s1n5938);
not(notn5938,n5014);
and (s0n5938,notn5938,n1366);
and (s1n5938,n5014,n5936);
and (n5939,n5940,n5038);
wire s0n5940,s1n5940,notn5940;
or (n5940,s0n5940,s1n5940);
not(notn5940,n5014);
and (s0n5940,notn5940,n862);
and (s1n5940,n5014,n1366);
wire s0n5942,s1n5942,notn5942;
or (n5942,s0n5942,s1n5942);
not(notn5942,n4966);
and (s0n5942,notn5942,n5943);
and (s1n5942,n4966,n6002);
or (n5943,1'b0,n5944,n5959,n5973,n5988);
and (n5944,n5945,n2718);
or (n5945,1'b0,n5946,n5950,n5953,n5956);
and (n5946,n5947,n5016);
wire s0n5947,s1n5947,notn5947;
or (n5947,s0n5947,s1n5947);
not(notn5947,n5014);
and (s0n5947,notn5947,n5948);
and (s1n5947,n5014,n5949);
and (n5950,n5951,n5028);
wire s0n5951,s1n5951,notn5951;
or (n5951,s0n5951,s1n5951);
not(notn5951,n5014);
and (s0n5951,notn5951,n5952);
and (s1n5951,n5014,n5948);
and (n5953,n5954,n5033);
wire s0n5954,s1n5954,notn5954;
or (n5954,s0n5954,s1n5954);
not(notn5954,n5014);
and (s0n5954,notn5954,n5955);
and (s1n5954,n5014,n5952);
and (n5956,n5957,n5038);
wire s0n5957,s1n5957,notn5957;
or (n5957,s0n5957,s1n5957);
not(notn5957,n5014);
and (s0n5957,notn5957,n5958);
and (s1n5957,n5014,n5955);
and (n5959,n5960,n2730);
or (n5960,1'b0,n5961,n5964,n5967,n5970);
and (n5961,n5962,n5016);
wire s0n5962,s1n5962,notn5962;
or (n5962,s0n5962,s1n5962);
not(notn5962,n5014);
and (s0n5962,notn5962,n5963);
and (s1n5962,n5014,n5958);
and (n5964,n5965,n5028);
wire s0n5965,s1n5965,notn5965;
or (n5965,s0n5965,s1n5965);
not(notn5965,n5014);
and (s0n5965,notn5965,n5966);
and (s1n5965,n5014,n5963);
and (n5967,n5968,n5033);
wire s0n5968,s1n5968,notn5968;
or (n5968,s0n5968,s1n5968);
not(notn5968,n5014);
and (s0n5968,notn5968,n5969);
and (s1n5968,n5014,n5966);
and (n5970,n5971,n5038);
wire s0n5971,s1n5971,notn5971;
or (n5971,s0n5971,s1n5971);
not(notn5971,n5014);
and (s0n5971,notn5971,n5972);
and (s1n5971,n5014,n5969);
and (n5973,n5974,n2742);
or (n5974,1'b0,n5975,n5979,n5982,n5985);
and (n5975,n5976,n5016);
wire s0n5976,s1n5976,notn5976;
or (n5976,s0n5976,s1n5976);
not(notn5976,n5014);
and (s0n5976,notn5976,n5977);
and (s1n5976,n5014,n5978);
and (n5979,n5980,n5028);
wire s0n5980,s1n5980,notn5980;
or (n5980,s0n5980,s1n5980);
not(notn5980,n5014);
and (s0n5980,notn5980,n5981);
and (s1n5980,n5014,n5977);
and (n5982,n5983,n5033);
wire s0n5983,s1n5983,notn5983;
or (n5983,s0n5983,s1n5983);
not(notn5983,n5014);
and (s0n5983,notn5983,n5984);
and (s1n5983,n5014,n5981);
and (n5985,n5986,n5038);
wire s0n5986,s1n5986,notn5986;
or (n5986,s0n5986,s1n5986);
not(notn5986,n5014);
and (s0n5986,notn5986,n5987);
and (s1n5986,n5014,n5984);
and (n5988,n5989,n2752);
or (n5989,1'b0,n5990,n5993,n5996,n5999);
and (n5990,n5991,n5016);
wire s0n5991,s1n5991,notn5991;
or (n5991,s0n5991,s1n5991);
not(notn5991,n5014);
and (s0n5991,notn5991,n5992);
and (s1n5991,n5014,n5987);
and (n5993,n5994,n5028);
wire s0n5994,s1n5994,notn5994;
or (n5994,s0n5994,s1n5994);
not(notn5994,n5014);
and (s0n5994,notn5994,n5995);
and (s1n5994,n5014,n5992);
and (n5996,n5997,n5033);
wire s0n5997,s1n5997,notn5997;
or (n5997,s0n5997,s1n5997);
not(notn5997,n5014);
and (s0n5997,notn5997,n5998);
and (s1n5997,n5014,n5995);
and (n5999,n6000,n5038);
wire s0n6000,s1n6000,notn6000;
or (n6000,s0n6000,s1n6000);
not(notn6000,n5014);
and (s0n6000,notn6000,n6001);
and (s1n6000,n5014,n5998);
and (n6003,n5761,n5882);
and (n6004,n5638,n5759);
and (n6005,n5515,n5636);
and (n6006,n5392,n5513);
and (n6007,n5269,n5390);
and (n6008,n5146,n5267);
and (n6009,n5006,n5144);
and (n6010,n4999,n5004);
and (n6011,n4992,n4997);
and (n6012,n4985,n4990);
and (n6013,n4978,n4983);
xor (n6014,n6015,n7438);
xor (n6015,n6016,n7352);
xor (n6016,n6017,n6756);
xor (n6017,n6018,n6023);
xor (n6018,n6019,n6021);
wire s0n6019,s1n6019,notn6019;
or (n6019,s0n6019,s1n6019);
not(notn6019,n4966);
and (s0n6019,notn6019,1'b0);
and (s1n6019,n4966,n6020);
wire s0n6021,s1n6021,notn6021;
or (n6021,s0n6021,s1n6021);
not(notn6021,n4966);
and (s0n6021,notn6021,1'b0);
and (s1n6021,n4966,n6022);
or (n6023,n6024,n6029,n6755);
and (n6024,n6025,n6027);
wire s0n6025,s1n6025,notn6025;
or (n6025,s0n6025,s1n6025);
not(notn6025,n4966);
and (s0n6025,notn6025,1'b0);
and (s1n6025,n4966,n6026);
wire s0n6027,s1n6027,notn6027;
or (n6027,s0n6027,s1n6027);
not(notn6027,n4966);
and (s0n6027,notn6027,1'b0);
and (s1n6027,n4966,n6028);
and (n6029,n6027,n6030);
or (n6030,n6031,n6036,n6754);
and (n6031,n6032,n6034);
wire s0n6032,s1n6032,notn6032;
or (n6032,s0n6032,s1n6032);
not(notn6032,n4966);
and (s0n6032,notn6032,1'b0);
and (s1n6032,n4966,n6033);
wire s0n6034,s1n6034,notn6034;
or (n6034,s0n6034,s1n6034);
not(notn6034,n4966);
and (s0n6034,notn6034,1'b0);
and (s1n6034,n4966,n6035);
and (n6036,n6034,n6037);
or (n6037,n6038,n6125,n6753);
and (n6038,n6039,n6082);
wire s0n6039,s1n6039,notn6039;
or (n6039,s0n6039,s1n6039);
not(notn6039,n4966);
and (s0n6039,notn6039,n6040);
and (s1n6039,n4966,n6081);
or (n6040,1'b0,n6041,n6051,n6061,n6071);
and (n6041,n6042,n2718);
or (n6042,1'b0,n6043,n6045,n6047,n6049);
and (n6043,n6044,n5016);
wire s0n6044,s1n6044,notn6044;
or (n6044,s0n6044,s1n6044);
not(notn6044,n5014);
and (s0n6044,notn6044,n2711);
and (s1n6044,n5014,n3023);
and (n6045,n6046,n5028);
wire s0n6046,s1n6046,notn6046;
or (n6046,s0n6046,s1n6046);
not(notn6046,n5014);
and (s0n6046,notn6046,n2713);
and (s1n6046,n5014,n2711);
and (n6047,n6048,n5033);
wire s0n6048,s1n6048,notn6048;
or (n6048,s0n6048,s1n6048);
not(notn6048,n5014);
and (s0n6048,notn6048,n2715);
and (s1n6048,n5014,n2713);
and (n6049,n6050,n5038);
wire s0n6050,s1n6050,notn6050;
or (n6050,s0n6050,s1n6050);
not(notn6050,n5014);
and (s0n6050,notn6050,n2717);
and (s1n6050,n5014,n2715);
and (n6051,n6052,n2730);
or (n6052,1'b0,n6053,n6055,n6057,n6059);
and (n6053,n6054,n5016);
wire s0n6054,s1n6054,notn6054;
or (n6054,s0n6054,s1n6054);
not(notn6054,n5014);
and (s0n6054,notn6054,n2723);
and (s1n6054,n5014,n2717);
and (n6055,n6056,n5028);
wire s0n6056,s1n6056,notn6056;
or (n6056,s0n6056,s1n6056);
not(notn6056,n5014);
and (s0n6056,notn6056,n2725);
and (s1n6056,n5014,n2723);
and (n6057,n6058,n5033);
wire s0n6058,s1n6058,notn6058;
or (n6058,s0n6058,s1n6058);
not(notn6058,n5014);
and (s0n6058,notn6058,n2727);
and (s1n6058,n5014,n2725);
and (n6059,n6060,n5038);
wire s0n6060,s1n6060,notn6060;
or (n6060,s0n6060,s1n6060);
not(notn6060,n5014);
and (s0n6060,notn6060,n2729);
and (s1n6060,n5014,n2727);
and (n6061,n6062,n2742);
or (n6062,1'b0,n6063,n6065,n6067,n6069);
and (n6063,n6064,n5016);
wire s0n6064,s1n6064,notn6064;
or (n6064,s0n6064,s1n6064);
not(notn6064,n5014);
and (s0n6064,notn6064,n2735);
and (s1n6064,n5014,n3038);
and (n6065,n6066,n5028);
wire s0n6066,s1n6066,notn6066;
or (n6066,s0n6066,s1n6066);
not(notn6066,n5014);
and (s0n6066,notn6066,n2737);
and (s1n6066,n5014,n2735);
and (n6067,n6068,n5033);
wire s0n6068,s1n6068,notn6068;
or (n6068,s0n6068,s1n6068);
not(notn6068,n5014);
and (s0n6068,notn6068,n2739);
and (s1n6068,n5014,n2737);
and (n6069,n6070,n5038);
wire s0n6070,s1n6070,notn6070;
or (n6070,s0n6070,s1n6070);
not(notn6070,n5014);
and (s0n6070,notn6070,n2741);
and (s1n6070,n5014,n2739);
and (n6071,n6072,n2752);
or (n6072,1'b0,n6073,n6075,n6077,n6079);
and (n6073,n6074,n5016);
wire s0n6074,s1n6074,notn6074;
or (n6074,s0n6074,s1n6074);
not(notn6074,n5014);
and (s0n6074,notn6074,n2747);
and (s1n6074,n5014,n2741);
and (n6075,n6076,n5028);
wire s0n6076,s1n6076,notn6076;
or (n6076,s0n6076,s1n6076);
not(notn6076,n5014);
and (s0n6076,notn6076,n2749);
and (s1n6076,n5014,n2747);
and (n6077,n6078,n5033);
wire s0n6078,s1n6078,notn6078;
or (n6078,s0n6078,s1n6078);
not(notn6078,n5014);
and (s0n6078,notn6078,n1251);
and (s1n6078,n5014,n2749);
and (n6079,n6080,n5038);
wire s0n6080,s1n6080,notn6080;
or (n6080,s0n6080,s1n6080);
not(notn6080,n5014);
and (s0n6080,notn6080,n564);
and (s1n6080,n5014,n1251);
wire s0n6082,s1n6082,notn6082;
or (n6082,s0n6082,s1n6082);
not(notn6082,n4966);
and (s0n6082,notn6082,n6083);
and (s1n6082,n4966,n6124);
or (n6083,1'b0,n6084,n6094,n6104,n6114);
and (n6084,n6085,n2718);
or (n6085,1'b0,n6086,n6088,n6090,n6092);
and (n6086,n6087,n5016);
wire s0n6087,s1n6087,notn6087;
or (n6087,s0n6087,s1n6087);
not(notn6087,n5014);
and (s0n6087,notn6087,n2928);
and (s1n6087,n5014,n3024);
and (n6088,n6089,n5028);
wire s0n6089,s1n6089,notn6089;
or (n6089,s0n6089,s1n6089);
not(notn6089,n5014);
and (s0n6089,notn6089,n2954);
and (s1n6089,n5014,n2928);
and (n6090,n6091,n5033);
wire s0n6091,s1n6091,notn6091;
or (n6091,s0n6091,s1n6091);
not(notn6091,n5014);
and (s0n6091,notn6091,n2962);
and (s1n6091,n5014,n2954);
and (n6092,n6093,n5038);
wire s0n6093,s1n6093,notn6093;
or (n6093,s0n6093,s1n6093);
not(notn6093,n5014);
and (s0n6093,notn6093,n2971);
and (s1n6093,n5014,n2962);
and (n6094,n6095,n2730);
or (n6095,1'b0,n6096,n6098,n6100,n6102);
and (n6096,n6097,n5016);
wire s0n6097,s1n6097,notn6097;
or (n6097,s0n6097,s1n6097);
not(notn6097,n5014);
and (s0n6097,notn6097,n2982);
and (s1n6097,n5014,n2971);
and (n6098,n6099,n5028);
wire s0n6099,s1n6099,notn6099;
or (n6099,s0n6099,s1n6099);
not(notn6099,n5014);
and (s0n6099,notn6099,n2985);
and (s1n6099,n5014,n2982);
and (n6100,n6101,n5033);
wire s0n6101,s1n6101,notn6101;
or (n6101,s0n6101,s1n6101);
not(notn6101,n5014);
and (s0n6101,notn6101,n2988);
and (s1n6101,n5014,n2985);
and (n6102,n6103,n5038);
wire s0n6103,s1n6103,notn6103;
or (n6103,s0n6103,s1n6103);
not(notn6103,n5014);
and (s0n6103,notn6103,n2991);
and (s1n6103,n5014,n2988);
and (n6104,n6105,n2742);
or (n6105,1'b0,n6106,n6108,n6110,n6112);
and (n6106,n6107,n5016);
wire s0n6107,s1n6107,notn6107;
or (n6107,s0n6107,s1n6107);
not(notn6107,n5014);
and (s0n6107,notn6107,n2996);
and (s1n6107,n5014,n3039);
and (n6108,n6109,n5028);
wire s0n6109,s1n6109,notn6109;
or (n6109,s0n6109,s1n6109);
not(notn6109,n5014);
and (s0n6109,notn6109,n2999);
and (s1n6109,n5014,n2996);
and (n6110,n6111,n5033);
wire s0n6111,s1n6111,notn6111;
or (n6111,s0n6111,s1n6111);
not(notn6111,n5014);
and (s0n6111,notn6111,n3002);
and (s1n6111,n5014,n2999);
and (n6112,n6113,n5038);
wire s0n6113,s1n6113,notn6113;
or (n6113,s0n6113,s1n6113);
not(notn6113,n5014);
and (s0n6113,notn6113,n3005);
and (s1n6113,n5014,n3002);
and (n6114,n6115,n2752);
or (n6115,1'b0,n6116,n6118,n6120,n6122);
and (n6116,n6117,n5016);
wire s0n6117,s1n6117,notn6117;
or (n6117,s0n6117,s1n6117);
not(notn6117,n5014);
and (s0n6117,notn6117,n3010);
and (s1n6117,n5014,n3005);
and (n6118,n6119,n5028);
wire s0n6119,s1n6119,notn6119;
or (n6119,s0n6119,s1n6119);
not(notn6119,n5014);
and (s0n6119,notn6119,n3013);
and (s1n6119,n5014,n3010);
and (n6120,n6121,n5033);
wire s0n6121,s1n6121,notn6121;
or (n6121,s0n6121,s1n6121);
not(notn6121,n5014);
and (s0n6121,notn6121,n2087);
and (s1n6121,n5014,n3013);
and (n6122,n6123,n5038);
wire s0n6123,s1n6123,notn6123;
or (n6123,s0n6123,s1n6123);
not(notn6123,n5014);
and (s0n6123,notn6123,n1692);
and (s1n6123,n5014,n2087);
and (n6125,n6082,n6126);
or (n6126,n6127,n6214,n6752);
and (n6127,n6128,n6171);
wire s0n6128,s1n6128,notn6128;
or (n6128,s0n6128,s1n6128);
not(notn6128,n4966);
and (s0n6128,notn6128,n6129);
and (s1n6128,n4966,n6170);
or (n6129,1'b0,n6130,n6140,n6150,n6160);
and (n6130,n6131,n2718);
or (n6131,1'b0,n6132,n6134,n6136,n6138);
and (n6132,n6133,n5016);
wire s0n6133,s1n6133,notn6133;
or (n6133,s0n6133,s1n6133);
not(notn6133,n5014);
and (s0n6133,notn6133,n3057);
and (s1n6133,n5014,n3126);
and (n6134,n6135,n5028);
wire s0n6135,s1n6135,notn6135;
or (n6135,s0n6135,s1n6135);
not(notn6135,n5014);
and (s0n6135,notn6135,n3061);
and (s1n6135,n5014,n3057);
and (n6136,n6137,n5033);
wire s0n6137,s1n6137,notn6137;
or (n6137,s0n6137,s1n6137);
not(notn6137,n5014);
and (s0n6137,notn6137,n3065);
and (s1n6137,n5014,n3061);
and (n6138,n6139,n5038);
wire s0n6139,s1n6139,notn6139;
or (n6139,s0n6139,s1n6139);
not(notn6139,n5014);
and (s0n6139,notn6139,n3069);
and (s1n6139,n5014,n3065);
and (n6140,n6141,n2730);
or (n6141,1'b0,n6142,n6144,n6146,n6148);
and (n6142,n6143,n5016);
wire s0n6143,s1n6143,notn6143;
or (n6143,s0n6143,s1n6143);
not(notn6143,n5014);
and (s0n6143,notn6143,n3075);
and (s1n6143,n5014,n3069);
and (n6144,n6145,n5028);
wire s0n6145,s1n6145,notn6145;
or (n6145,s0n6145,s1n6145);
not(notn6145,n5014);
and (s0n6145,notn6145,n3079);
and (s1n6145,n5014,n3075);
and (n6146,n6147,n5033);
wire s0n6147,s1n6147,notn6147;
or (n6147,s0n6147,s1n6147);
not(notn6147,n5014);
and (s0n6147,notn6147,n3083);
and (s1n6147,n5014,n3079);
and (n6148,n6149,n5038);
wire s0n6149,s1n6149,notn6149;
or (n6149,s0n6149,s1n6149);
not(notn6149,n5014);
and (s0n6149,notn6149,n3087);
and (s1n6149,n5014,n3083);
and (n6150,n6151,n2742);
or (n6151,1'b0,n6152,n6154,n6156,n6158);
and (n6152,n6153,n5016);
wire s0n6153,s1n6153,notn6153;
or (n6153,s0n6153,s1n6153);
not(notn6153,n5014);
and (s0n6153,notn6153,n3093);
and (s1n6153,n5014,n3141);
and (n6154,n6155,n5028);
wire s0n6155,s1n6155,notn6155;
or (n6155,s0n6155,s1n6155);
not(notn6155,n5014);
and (s0n6155,notn6155,n3097);
and (s1n6155,n5014,n3093);
and (n6156,n6157,n5033);
wire s0n6157,s1n6157,notn6157;
or (n6157,s0n6157,s1n6157);
not(notn6157,n5014);
and (s0n6157,notn6157,n3101);
and (s1n6157,n5014,n3097);
and (n6158,n6159,n5038);
wire s0n6159,s1n6159,notn6159;
or (n6159,s0n6159,s1n6159);
not(notn6159,n5014);
and (s0n6159,notn6159,n3105);
and (s1n6159,n5014,n3101);
and (n6160,n6161,n2752);
or (n6161,1'b0,n6162,n6164,n6166,n6168);
and (n6162,n6163,n5016);
wire s0n6163,s1n6163,notn6163;
or (n6163,s0n6163,s1n6163);
not(notn6163,n5014);
and (s0n6163,notn6163,n3111);
and (s1n6163,n5014,n3105);
and (n6164,n6165,n5028);
wire s0n6165,s1n6165,notn6165;
or (n6165,s0n6165,s1n6165);
not(notn6165,n5014);
and (s0n6165,notn6165,n3115);
and (s1n6165,n5014,n3111);
and (n6166,n6167,n5033);
wire s0n6167,s1n6167,notn6167;
or (n6167,s0n6167,s1n6167);
not(notn6167,n5014);
and (s0n6167,notn6167,n1267);
and (s1n6167,n5014,n3115);
and (n6168,n6169,n5038);
wire s0n6169,s1n6169,notn6169;
or (n6169,s0n6169,s1n6169);
not(notn6169,n5014);
and (s0n6169,notn6169,n755);
and (s1n6169,n5014,n1267);
wire s0n6171,s1n6171,notn6171;
or (n6171,s0n6171,s1n6171);
not(notn6171,n4966);
and (s0n6171,notn6171,n6172);
and (s1n6171,n4966,n6213);
or (n6172,1'b0,n6173,n6183,n6193,n6203);
and (n6173,n6174,n2718);
or (n6174,1'b0,n6175,n6177,n6179,n6181);
and (n6175,n6176,n5016);
wire s0n6176,s1n6176,notn6176;
or (n6176,s0n6176,s1n6176);
not(notn6176,n5014);
and (s0n6176,notn6176,n3058);
and (s1n6176,n5014,n3127);
and (n6177,n6178,n5028);
wire s0n6178,s1n6178,notn6178;
or (n6178,s0n6178,s1n6178);
not(notn6178,n5014);
and (s0n6178,notn6178,n3062);
and (s1n6178,n5014,n3058);
and (n6179,n6180,n5033);
wire s0n6180,s1n6180,notn6180;
or (n6180,s0n6180,s1n6180);
not(notn6180,n5014);
and (s0n6180,notn6180,n3066);
and (s1n6180,n5014,n3062);
and (n6181,n6182,n5038);
wire s0n6182,s1n6182,notn6182;
or (n6182,s0n6182,s1n6182);
not(notn6182,n5014);
and (s0n6182,notn6182,n3070);
and (s1n6182,n5014,n3066);
and (n6183,n6184,n2730);
or (n6184,1'b0,n6185,n6187,n6189,n6191);
and (n6185,n6186,n5016);
wire s0n6186,s1n6186,notn6186;
or (n6186,s0n6186,s1n6186);
not(notn6186,n5014);
and (s0n6186,notn6186,n3076);
and (s1n6186,n5014,n3070);
and (n6187,n6188,n5028);
wire s0n6188,s1n6188,notn6188;
or (n6188,s0n6188,s1n6188);
not(notn6188,n5014);
and (s0n6188,notn6188,n3080);
and (s1n6188,n5014,n3076);
and (n6189,n6190,n5033);
wire s0n6190,s1n6190,notn6190;
or (n6190,s0n6190,s1n6190);
not(notn6190,n5014);
and (s0n6190,notn6190,n3084);
and (s1n6190,n5014,n3080);
and (n6191,n6192,n5038);
wire s0n6192,s1n6192,notn6192;
or (n6192,s0n6192,s1n6192);
not(notn6192,n5014);
and (s0n6192,notn6192,n3088);
and (s1n6192,n5014,n3084);
and (n6193,n6194,n2742);
or (n6194,1'b0,n6195,n6197,n6199,n6201);
and (n6195,n6196,n5016);
wire s0n6196,s1n6196,notn6196;
or (n6196,s0n6196,s1n6196);
not(notn6196,n5014);
and (s0n6196,notn6196,n3094);
and (s1n6196,n5014,n3142);
and (n6197,n6198,n5028);
wire s0n6198,s1n6198,notn6198;
or (n6198,s0n6198,s1n6198);
not(notn6198,n5014);
and (s0n6198,notn6198,n3098);
and (s1n6198,n5014,n3094);
and (n6199,n6200,n5033);
wire s0n6200,s1n6200,notn6200;
or (n6200,s0n6200,s1n6200);
not(notn6200,n5014);
and (s0n6200,notn6200,n3102);
and (s1n6200,n5014,n3098);
and (n6201,n6202,n5038);
wire s0n6202,s1n6202,notn6202;
or (n6202,s0n6202,s1n6202);
not(notn6202,n5014);
and (s0n6202,notn6202,n3106);
and (s1n6202,n5014,n3102);
and (n6203,n6204,n2752);
or (n6204,1'b0,n6205,n6207,n6209,n6211);
and (n6205,n6206,n5016);
wire s0n6206,s1n6206,notn6206;
or (n6206,s0n6206,s1n6206);
not(notn6206,n5014);
and (s0n6206,notn6206,n3112);
and (s1n6206,n5014,n3106);
and (n6207,n6208,n5028);
wire s0n6208,s1n6208,notn6208;
or (n6208,s0n6208,s1n6208);
not(notn6208,n5014);
and (s0n6208,notn6208,n3116);
and (s1n6208,n5014,n3112);
and (n6209,n6210,n5033);
wire s0n6210,s1n6210,notn6210;
or (n6210,s0n6210,s1n6210);
not(notn6210,n5014);
and (s0n6210,notn6210,n2103);
and (s1n6210,n5014,n3116);
and (n6211,n6212,n5038);
wire s0n6212,s1n6212,notn6212;
or (n6212,s0n6212,s1n6212);
not(notn6212,n5014);
and (s0n6212,notn6212,n1708);
and (s1n6212,n5014,n2103);
and (n6214,n6171,n6215);
or (n6215,n6216,n6303,n6751);
and (n6216,n6217,n6260);
wire s0n6217,s1n6217,notn6217;
or (n6217,s0n6217,s1n6217);
not(notn6217,n4966);
and (s0n6217,notn6217,n6218);
and (s1n6217,n4966,n6259);
or (n6218,1'b0,n6219,n6229,n6239,n6249);
and (n6219,n6220,n2718);
or (n6220,1'b0,n6221,n6223,n6225,n6227);
and (n6221,n6222,n5016);
wire s0n6222,s1n6222,notn6222;
or (n6222,s0n6222,s1n6222);
not(notn6222,n5014);
and (s0n6222,notn6222,n3160);
and (s1n6222,n5014,n3229);
and (n6223,n6224,n5028);
wire s0n6224,s1n6224,notn6224;
or (n6224,s0n6224,s1n6224);
not(notn6224,n5014);
and (s0n6224,notn6224,n3164);
and (s1n6224,n5014,n3160);
and (n6225,n6226,n5033);
wire s0n6226,s1n6226,notn6226;
or (n6226,s0n6226,s1n6226);
not(notn6226,n5014);
and (s0n6226,notn6226,n3168);
and (s1n6226,n5014,n3164);
and (n6227,n6228,n5038);
wire s0n6228,s1n6228,notn6228;
or (n6228,s0n6228,s1n6228);
not(notn6228,n5014);
and (s0n6228,notn6228,n3172);
and (s1n6228,n5014,n3168);
and (n6229,n6230,n2730);
or (n6230,1'b0,n6231,n6233,n6235,n6237);
and (n6231,n6232,n5016);
wire s0n6232,s1n6232,notn6232;
or (n6232,s0n6232,s1n6232);
not(notn6232,n5014);
and (s0n6232,notn6232,n3178);
and (s1n6232,n5014,n3172);
and (n6233,n6234,n5028);
wire s0n6234,s1n6234,notn6234;
or (n6234,s0n6234,s1n6234);
not(notn6234,n5014);
and (s0n6234,notn6234,n3182);
and (s1n6234,n5014,n3178);
and (n6235,n6236,n5033);
wire s0n6236,s1n6236,notn6236;
or (n6236,s0n6236,s1n6236);
not(notn6236,n5014);
and (s0n6236,notn6236,n3186);
and (s1n6236,n5014,n3182);
and (n6237,n6238,n5038);
wire s0n6238,s1n6238,notn6238;
or (n6238,s0n6238,s1n6238);
not(notn6238,n5014);
and (s0n6238,notn6238,n3190);
and (s1n6238,n5014,n3186);
and (n6239,n6240,n2742);
or (n6240,1'b0,n6241,n6243,n6245,n6247);
and (n6241,n6242,n5016);
wire s0n6242,s1n6242,notn6242;
or (n6242,s0n6242,s1n6242);
not(notn6242,n5014);
and (s0n6242,notn6242,n3196);
and (s1n6242,n5014,n3244);
and (n6243,n6244,n5028);
wire s0n6244,s1n6244,notn6244;
or (n6244,s0n6244,s1n6244);
not(notn6244,n5014);
and (s0n6244,notn6244,n3200);
and (s1n6244,n5014,n3196);
and (n6245,n6246,n5033);
wire s0n6246,s1n6246,notn6246;
or (n6246,s0n6246,s1n6246);
not(notn6246,n5014);
and (s0n6246,notn6246,n3204);
and (s1n6246,n5014,n3200);
and (n6247,n6248,n5038);
wire s0n6248,s1n6248,notn6248;
or (n6248,s0n6248,s1n6248);
not(notn6248,n5014);
and (s0n6248,notn6248,n3208);
and (s1n6248,n5014,n3204);
and (n6249,n6250,n2752);
or (n6250,1'b0,n6251,n6253,n6255,n6257);
and (n6251,n6252,n5016);
wire s0n6252,s1n6252,notn6252;
or (n6252,s0n6252,s1n6252);
not(notn6252,n5014);
and (s0n6252,notn6252,n3214);
and (s1n6252,n5014,n3208);
and (n6253,n6254,n5028);
wire s0n6254,s1n6254,notn6254;
or (n6254,s0n6254,s1n6254);
not(notn6254,n5014);
and (s0n6254,notn6254,n3218);
and (s1n6254,n5014,n3214);
and (n6255,n6256,n5033);
wire s0n6256,s1n6256,notn6256;
or (n6256,s0n6256,s1n6256);
not(notn6256,n5014);
and (s0n6256,notn6256,n1283);
and (s1n6256,n5014,n3218);
and (n6257,n6258,n5038);
wire s0n6258,s1n6258,notn6258;
or (n6258,s0n6258,s1n6258);
not(notn6258,n5014);
and (s0n6258,notn6258,n779);
and (s1n6258,n5014,n1283);
wire s0n6260,s1n6260,notn6260;
or (n6260,s0n6260,s1n6260);
not(notn6260,n4966);
and (s0n6260,notn6260,n6261);
and (s1n6260,n4966,n6302);
or (n6261,1'b0,n6262,n6272,n6282,n6292);
and (n6262,n6263,n2718);
or (n6263,1'b0,n6264,n6266,n6268,n6270);
and (n6264,n6265,n5016);
wire s0n6265,s1n6265,notn6265;
or (n6265,s0n6265,s1n6265);
not(notn6265,n5014);
and (s0n6265,notn6265,n3161);
and (s1n6265,n5014,n3230);
and (n6266,n6267,n5028);
wire s0n6267,s1n6267,notn6267;
or (n6267,s0n6267,s1n6267);
not(notn6267,n5014);
and (s0n6267,notn6267,n3165);
and (s1n6267,n5014,n3161);
and (n6268,n6269,n5033);
wire s0n6269,s1n6269,notn6269;
or (n6269,s0n6269,s1n6269);
not(notn6269,n5014);
and (s0n6269,notn6269,n3169);
and (s1n6269,n5014,n3165);
and (n6270,n6271,n5038);
wire s0n6271,s1n6271,notn6271;
or (n6271,s0n6271,s1n6271);
not(notn6271,n5014);
and (s0n6271,notn6271,n3173);
and (s1n6271,n5014,n3169);
and (n6272,n6273,n2730);
or (n6273,1'b0,n6274,n6276,n6278,n6280);
and (n6274,n6275,n5016);
wire s0n6275,s1n6275,notn6275;
or (n6275,s0n6275,s1n6275);
not(notn6275,n5014);
and (s0n6275,notn6275,n3179);
and (s1n6275,n5014,n3173);
and (n6276,n6277,n5028);
wire s0n6277,s1n6277,notn6277;
or (n6277,s0n6277,s1n6277);
not(notn6277,n5014);
and (s0n6277,notn6277,n3183);
and (s1n6277,n5014,n3179);
and (n6278,n6279,n5033);
wire s0n6279,s1n6279,notn6279;
or (n6279,s0n6279,s1n6279);
not(notn6279,n5014);
and (s0n6279,notn6279,n3187);
and (s1n6279,n5014,n3183);
and (n6280,n6281,n5038);
wire s0n6281,s1n6281,notn6281;
or (n6281,s0n6281,s1n6281);
not(notn6281,n5014);
and (s0n6281,notn6281,n3191);
and (s1n6281,n5014,n3187);
and (n6282,n6283,n2742);
or (n6283,1'b0,n6284,n6286,n6288,n6290);
and (n6284,n6285,n5016);
wire s0n6285,s1n6285,notn6285;
or (n6285,s0n6285,s1n6285);
not(notn6285,n5014);
and (s0n6285,notn6285,n3197);
and (s1n6285,n5014,n3245);
and (n6286,n6287,n5028);
wire s0n6287,s1n6287,notn6287;
or (n6287,s0n6287,s1n6287);
not(notn6287,n5014);
and (s0n6287,notn6287,n3201);
and (s1n6287,n5014,n3197);
and (n6288,n6289,n5033);
wire s0n6289,s1n6289,notn6289;
or (n6289,s0n6289,s1n6289);
not(notn6289,n5014);
and (s0n6289,notn6289,n3205);
and (s1n6289,n5014,n3201);
and (n6290,n6291,n5038);
wire s0n6291,s1n6291,notn6291;
or (n6291,s0n6291,s1n6291);
not(notn6291,n5014);
and (s0n6291,notn6291,n3209);
and (s1n6291,n5014,n3205);
and (n6292,n6293,n2752);
or (n6293,1'b0,n6294,n6296,n6298,n6300);
and (n6294,n6295,n5016);
wire s0n6295,s1n6295,notn6295;
or (n6295,s0n6295,s1n6295);
not(notn6295,n5014);
and (s0n6295,notn6295,n3215);
and (s1n6295,n5014,n3209);
and (n6296,n6297,n5028);
wire s0n6297,s1n6297,notn6297;
or (n6297,s0n6297,s1n6297);
not(notn6297,n5014);
and (s0n6297,notn6297,n3219);
and (s1n6297,n5014,n3215);
and (n6298,n6299,n5033);
wire s0n6299,s1n6299,notn6299;
or (n6299,s0n6299,s1n6299);
not(notn6299,n5014);
and (s0n6299,notn6299,n2119);
and (s1n6299,n5014,n3219);
and (n6300,n6301,n5038);
wire s0n6301,s1n6301,notn6301;
or (n6301,s0n6301,s1n6301);
not(notn6301,n5014);
and (s0n6301,notn6301,n1727);
and (s1n6301,n5014,n2119);
and (n6303,n6260,n6304);
or (n6304,n6305,n6392,n6750);
and (n6305,n6306,n6349);
wire s0n6306,s1n6306,notn6306;
or (n6306,s0n6306,s1n6306);
not(notn6306,n4966);
and (s0n6306,notn6306,n6307);
and (s1n6306,n4966,n6348);
or (n6307,1'b0,n6308,n6318,n6328,n6338);
and (n6308,n6309,n2718);
or (n6309,1'b0,n6310,n6312,n6314,n6316);
and (n6310,n6311,n5016);
wire s0n6311,s1n6311,notn6311;
or (n6311,s0n6311,s1n6311);
not(notn6311,n5014);
and (s0n6311,notn6311,n3263);
and (s1n6311,n5014,n3332);
and (n6312,n6313,n5028);
wire s0n6313,s1n6313,notn6313;
or (n6313,s0n6313,s1n6313);
not(notn6313,n5014);
and (s0n6313,notn6313,n3267);
and (s1n6313,n5014,n3263);
and (n6314,n6315,n5033);
wire s0n6315,s1n6315,notn6315;
or (n6315,s0n6315,s1n6315);
not(notn6315,n5014);
and (s0n6315,notn6315,n3271);
and (s1n6315,n5014,n3267);
and (n6316,n6317,n5038);
wire s0n6317,s1n6317,notn6317;
or (n6317,s0n6317,s1n6317);
not(notn6317,n5014);
and (s0n6317,notn6317,n3275);
and (s1n6317,n5014,n3271);
and (n6318,n6319,n2730);
or (n6319,1'b0,n6320,n6322,n6324,n6326);
and (n6320,n6321,n5016);
wire s0n6321,s1n6321,notn6321;
or (n6321,s0n6321,s1n6321);
not(notn6321,n5014);
and (s0n6321,notn6321,n3281);
and (s1n6321,n5014,n3275);
and (n6322,n6323,n5028);
wire s0n6323,s1n6323,notn6323;
or (n6323,s0n6323,s1n6323);
not(notn6323,n5014);
and (s0n6323,notn6323,n3285);
and (s1n6323,n5014,n3281);
and (n6324,n6325,n5033);
wire s0n6325,s1n6325,notn6325;
or (n6325,s0n6325,s1n6325);
not(notn6325,n5014);
and (s0n6325,notn6325,n3289);
and (s1n6325,n5014,n3285);
and (n6326,n6327,n5038);
wire s0n6327,s1n6327,notn6327;
or (n6327,s0n6327,s1n6327);
not(notn6327,n5014);
and (s0n6327,notn6327,n3293);
and (s1n6327,n5014,n3289);
and (n6328,n6329,n2742);
or (n6329,1'b0,n6330,n6332,n6334,n6336);
and (n6330,n6331,n5016);
wire s0n6331,s1n6331,notn6331;
or (n6331,s0n6331,s1n6331);
not(notn6331,n5014);
and (s0n6331,notn6331,n3299);
and (s1n6331,n5014,n3347);
and (n6332,n6333,n5028);
wire s0n6333,s1n6333,notn6333;
or (n6333,s0n6333,s1n6333);
not(notn6333,n5014);
and (s0n6333,notn6333,n3303);
and (s1n6333,n5014,n3299);
and (n6334,n6335,n5033);
wire s0n6335,s1n6335,notn6335;
or (n6335,s0n6335,s1n6335);
not(notn6335,n5014);
and (s0n6335,notn6335,n3307);
and (s1n6335,n5014,n3303);
and (n6336,n6337,n5038);
wire s0n6337,s1n6337,notn6337;
or (n6337,s0n6337,s1n6337);
not(notn6337,n5014);
and (s0n6337,notn6337,n3311);
and (s1n6337,n5014,n3307);
and (n6338,n6339,n2752);
or (n6339,1'b0,n6340,n6342,n6344,n6346);
and (n6340,n6341,n5016);
wire s0n6341,s1n6341,notn6341;
or (n6341,s0n6341,s1n6341);
not(notn6341,n5014);
and (s0n6341,notn6341,n3317);
and (s1n6341,n5014,n3311);
and (n6342,n6343,n5028);
wire s0n6343,s1n6343,notn6343;
or (n6343,s0n6343,s1n6343);
not(notn6343,n5014);
and (s0n6343,notn6343,n3321);
and (s1n6343,n5014,n3317);
and (n6344,n6345,n5033);
wire s0n6345,s1n6345,notn6345;
or (n6345,s0n6345,s1n6345);
not(notn6345,n5014);
and (s0n6345,notn6345,n1299);
and (s1n6345,n5014,n3321);
and (n6346,n6347,n5038);
wire s0n6347,s1n6347,notn6347;
or (n6347,s0n6347,s1n6347);
not(notn6347,n5014);
and (s0n6347,notn6347,n795);
and (s1n6347,n5014,n1299);
wire s0n6349,s1n6349,notn6349;
or (n6349,s0n6349,s1n6349);
not(notn6349,n4966);
and (s0n6349,notn6349,n6350);
and (s1n6349,n4966,n6391);
or (n6350,1'b0,n6351,n6361,n6371,n6381);
and (n6351,n6352,n2718);
or (n6352,1'b0,n6353,n6355,n6357,n6359);
and (n6353,n6354,n5016);
wire s0n6354,s1n6354,notn6354;
or (n6354,s0n6354,s1n6354);
not(notn6354,n5014);
and (s0n6354,notn6354,n3264);
and (s1n6354,n5014,n3333);
and (n6355,n6356,n5028);
wire s0n6356,s1n6356,notn6356;
or (n6356,s0n6356,s1n6356);
not(notn6356,n5014);
and (s0n6356,notn6356,n3268);
and (s1n6356,n5014,n3264);
and (n6357,n6358,n5033);
wire s0n6358,s1n6358,notn6358;
or (n6358,s0n6358,s1n6358);
not(notn6358,n5014);
and (s0n6358,notn6358,n3272);
and (s1n6358,n5014,n3268);
and (n6359,n6360,n5038);
wire s0n6360,s1n6360,notn6360;
or (n6360,s0n6360,s1n6360);
not(notn6360,n5014);
and (s0n6360,notn6360,n3276);
and (s1n6360,n5014,n3272);
and (n6361,n6362,n2730);
or (n6362,1'b0,n6363,n6365,n6367,n6369);
and (n6363,n6364,n5016);
wire s0n6364,s1n6364,notn6364;
or (n6364,s0n6364,s1n6364);
not(notn6364,n5014);
and (s0n6364,notn6364,n3282);
and (s1n6364,n5014,n3276);
and (n6365,n6366,n5028);
wire s0n6366,s1n6366,notn6366;
or (n6366,s0n6366,s1n6366);
not(notn6366,n5014);
and (s0n6366,notn6366,n3286);
and (s1n6366,n5014,n3282);
and (n6367,n6368,n5033);
wire s0n6368,s1n6368,notn6368;
or (n6368,s0n6368,s1n6368);
not(notn6368,n5014);
and (s0n6368,notn6368,n3290);
and (s1n6368,n5014,n3286);
and (n6369,n6370,n5038);
wire s0n6370,s1n6370,notn6370;
or (n6370,s0n6370,s1n6370);
not(notn6370,n5014);
and (s0n6370,notn6370,n3294);
and (s1n6370,n5014,n3290);
and (n6371,n6372,n2742);
or (n6372,1'b0,n6373,n6375,n6377,n6379);
and (n6373,n6374,n5016);
wire s0n6374,s1n6374,notn6374;
or (n6374,s0n6374,s1n6374);
not(notn6374,n5014);
and (s0n6374,notn6374,n3300);
and (s1n6374,n5014,n3348);
and (n6375,n6376,n5028);
wire s0n6376,s1n6376,notn6376;
or (n6376,s0n6376,s1n6376);
not(notn6376,n5014);
and (s0n6376,notn6376,n3304);
and (s1n6376,n5014,n3300);
and (n6377,n6378,n5033);
wire s0n6378,s1n6378,notn6378;
or (n6378,s0n6378,s1n6378);
not(notn6378,n5014);
and (s0n6378,notn6378,n3308);
and (s1n6378,n5014,n3304);
and (n6379,n6380,n5038);
wire s0n6380,s1n6380,notn6380;
or (n6380,s0n6380,s1n6380);
not(notn6380,n5014);
and (s0n6380,notn6380,n3312);
and (s1n6380,n5014,n3308);
and (n6381,n6382,n2752);
or (n6382,1'b0,n6383,n6385,n6387,n6389);
and (n6383,n6384,n5016);
wire s0n6384,s1n6384,notn6384;
or (n6384,s0n6384,s1n6384);
not(notn6384,n5014);
and (s0n6384,notn6384,n3318);
and (s1n6384,n5014,n3312);
and (n6385,n6386,n5028);
wire s0n6386,s1n6386,notn6386;
or (n6386,s0n6386,s1n6386);
not(notn6386,n5014);
and (s0n6386,notn6386,n3322);
and (s1n6386,n5014,n3318);
and (n6387,n6388,n5033);
wire s0n6388,s1n6388,notn6388;
or (n6388,s0n6388,s1n6388);
not(notn6388,n5014);
and (s0n6388,notn6388,n2135);
and (s1n6388,n5014,n3322);
and (n6389,n6390,n5038);
wire s0n6390,s1n6390,notn6390;
or (n6390,s0n6390,s1n6390);
not(notn6390,n5014);
and (s0n6390,notn6390,n1753);
and (s1n6390,n5014,n2135);
and (n6392,n6349,n6393);
or (n6393,n6394,n6481,n6749);
and (n6394,n6395,n6438);
wire s0n6395,s1n6395,notn6395;
or (n6395,s0n6395,s1n6395);
not(notn6395,n4966);
and (s0n6395,notn6395,n6396);
and (s1n6395,n4966,n6437);
or (n6396,1'b0,n6397,n6407,n6417,n6427);
and (n6397,n6398,n2718);
or (n6398,1'b0,n6399,n6401,n6403,n6405);
and (n6399,n6400,n5016);
wire s0n6400,s1n6400,notn6400;
or (n6400,s0n6400,s1n6400);
not(notn6400,n5014);
and (s0n6400,notn6400,n3366);
and (s1n6400,n5014,n3435);
and (n6401,n6402,n5028);
wire s0n6402,s1n6402,notn6402;
or (n6402,s0n6402,s1n6402);
not(notn6402,n5014);
and (s0n6402,notn6402,n3370);
and (s1n6402,n5014,n3366);
and (n6403,n6404,n5033);
wire s0n6404,s1n6404,notn6404;
or (n6404,s0n6404,s1n6404);
not(notn6404,n5014);
and (s0n6404,notn6404,n3374);
and (s1n6404,n5014,n3370);
and (n6405,n6406,n5038);
wire s0n6406,s1n6406,notn6406;
or (n6406,s0n6406,s1n6406);
not(notn6406,n5014);
and (s0n6406,notn6406,n3378);
and (s1n6406,n5014,n3374);
and (n6407,n6408,n2730);
or (n6408,1'b0,n6409,n6411,n6413,n6415);
and (n6409,n6410,n5016);
wire s0n6410,s1n6410,notn6410;
or (n6410,s0n6410,s1n6410);
not(notn6410,n5014);
and (s0n6410,notn6410,n3384);
and (s1n6410,n5014,n3378);
and (n6411,n6412,n5028);
wire s0n6412,s1n6412,notn6412;
or (n6412,s0n6412,s1n6412);
not(notn6412,n5014);
and (s0n6412,notn6412,n3388);
and (s1n6412,n5014,n3384);
and (n6413,n6414,n5033);
wire s0n6414,s1n6414,notn6414;
or (n6414,s0n6414,s1n6414);
not(notn6414,n5014);
and (s0n6414,notn6414,n3392);
and (s1n6414,n5014,n3388);
and (n6415,n6416,n5038);
wire s0n6416,s1n6416,notn6416;
or (n6416,s0n6416,s1n6416);
not(notn6416,n5014);
and (s0n6416,notn6416,n3396);
and (s1n6416,n5014,n3392);
and (n6417,n6418,n2742);
or (n6418,1'b0,n6419,n6421,n6423,n6425);
and (n6419,n6420,n5016);
wire s0n6420,s1n6420,notn6420;
or (n6420,s0n6420,s1n6420);
not(notn6420,n5014);
and (s0n6420,notn6420,n3402);
and (s1n6420,n5014,n3450);
and (n6421,n6422,n5028);
wire s0n6422,s1n6422,notn6422;
or (n6422,s0n6422,s1n6422);
not(notn6422,n5014);
and (s0n6422,notn6422,n3406);
and (s1n6422,n5014,n3402);
and (n6423,n6424,n5033);
wire s0n6424,s1n6424,notn6424;
or (n6424,s0n6424,s1n6424);
not(notn6424,n5014);
and (s0n6424,notn6424,n3410);
and (s1n6424,n5014,n3406);
and (n6425,n6426,n5038);
wire s0n6426,s1n6426,notn6426;
or (n6426,s0n6426,s1n6426);
not(notn6426,n5014);
and (s0n6426,notn6426,n3414);
and (s1n6426,n5014,n3410);
and (n6427,n6428,n2752);
or (n6428,1'b0,n6429,n6431,n6433,n6435);
and (n6429,n6430,n5016);
wire s0n6430,s1n6430,notn6430;
or (n6430,s0n6430,s1n6430);
not(notn6430,n5014);
and (s0n6430,notn6430,n3420);
and (s1n6430,n5014,n3414);
and (n6431,n6432,n5028);
wire s0n6432,s1n6432,notn6432;
or (n6432,s0n6432,s1n6432);
not(notn6432,n5014);
and (s0n6432,notn6432,n3424);
and (s1n6432,n5014,n3420);
and (n6433,n6434,n5033);
wire s0n6434,s1n6434,notn6434;
or (n6434,s0n6434,s1n6434);
not(notn6434,n5014);
and (s0n6434,notn6434,n1315);
and (s1n6434,n5014,n3424);
and (n6435,n6436,n5038);
wire s0n6436,s1n6436,notn6436;
or (n6436,s0n6436,s1n6436);
not(notn6436,n5014);
and (s0n6436,notn6436,n811);
and (s1n6436,n5014,n1315);
wire s0n6438,s1n6438,notn6438;
or (n6438,s0n6438,s1n6438);
not(notn6438,n4966);
and (s0n6438,notn6438,n6439);
and (s1n6438,n4966,n6480);
or (n6439,1'b0,n6440,n6450,n6460,n6470);
and (n6440,n6441,n2718);
or (n6441,1'b0,n6442,n6444,n6446,n6448);
and (n6442,n6443,n5016);
wire s0n6443,s1n6443,notn6443;
or (n6443,s0n6443,s1n6443);
not(notn6443,n5014);
and (s0n6443,notn6443,n3367);
and (s1n6443,n5014,n3436);
and (n6444,n6445,n5028);
wire s0n6445,s1n6445,notn6445;
or (n6445,s0n6445,s1n6445);
not(notn6445,n5014);
and (s0n6445,notn6445,n3371);
and (s1n6445,n5014,n3367);
and (n6446,n6447,n5033);
wire s0n6447,s1n6447,notn6447;
or (n6447,s0n6447,s1n6447);
not(notn6447,n5014);
and (s0n6447,notn6447,n3375);
and (s1n6447,n5014,n3371);
and (n6448,n6449,n5038);
wire s0n6449,s1n6449,notn6449;
or (n6449,s0n6449,s1n6449);
not(notn6449,n5014);
and (s0n6449,notn6449,n3379);
and (s1n6449,n5014,n3375);
and (n6450,n6451,n2730);
or (n6451,1'b0,n6452,n6454,n6456,n6458);
and (n6452,n6453,n5016);
wire s0n6453,s1n6453,notn6453;
or (n6453,s0n6453,s1n6453);
not(notn6453,n5014);
and (s0n6453,notn6453,n3385);
and (s1n6453,n5014,n3379);
and (n6454,n6455,n5028);
wire s0n6455,s1n6455,notn6455;
or (n6455,s0n6455,s1n6455);
not(notn6455,n5014);
and (s0n6455,notn6455,n3389);
and (s1n6455,n5014,n3385);
and (n6456,n6457,n5033);
wire s0n6457,s1n6457,notn6457;
or (n6457,s0n6457,s1n6457);
not(notn6457,n5014);
and (s0n6457,notn6457,n3393);
and (s1n6457,n5014,n3389);
and (n6458,n6459,n5038);
wire s0n6459,s1n6459,notn6459;
or (n6459,s0n6459,s1n6459);
not(notn6459,n5014);
and (s0n6459,notn6459,n3397);
and (s1n6459,n5014,n3393);
and (n6460,n6461,n2742);
or (n6461,1'b0,n6462,n6464,n6466,n6468);
and (n6462,n6463,n5016);
wire s0n6463,s1n6463,notn6463;
or (n6463,s0n6463,s1n6463);
not(notn6463,n5014);
and (s0n6463,notn6463,n3403);
and (s1n6463,n5014,n3451);
and (n6464,n6465,n5028);
wire s0n6465,s1n6465,notn6465;
or (n6465,s0n6465,s1n6465);
not(notn6465,n5014);
and (s0n6465,notn6465,n3407);
and (s1n6465,n5014,n3403);
and (n6466,n6467,n5033);
wire s0n6467,s1n6467,notn6467;
or (n6467,s0n6467,s1n6467);
not(notn6467,n5014);
and (s0n6467,notn6467,n3411);
and (s1n6467,n5014,n3407);
and (n6468,n6469,n5038);
wire s0n6469,s1n6469,notn6469;
or (n6469,s0n6469,s1n6469);
not(notn6469,n5014);
and (s0n6469,notn6469,n3415);
and (s1n6469,n5014,n3411);
and (n6470,n6471,n2752);
or (n6471,1'b0,n6472,n6474,n6476,n6478);
and (n6472,n6473,n5016);
wire s0n6473,s1n6473,notn6473;
or (n6473,s0n6473,s1n6473);
not(notn6473,n5014);
and (s0n6473,notn6473,n3421);
and (s1n6473,n5014,n3415);
and (n6474,n6475,n5028);
wire s0n6475,s1n6475,notn6475;
or (n6475,s0n6475,s1n6475);
not(notn6475,n5014);
and (s0n6475,notn6475,n3425);
and (s1n6475,n5014,n3421);
and (n6476,n6477,n5033);
wire s0n6477,s1n6477,notn6477;
or (n6477,s0n6477,s1n6477);
not(notn6477,n5014);
and (s0n6477,notn6477,n2151);
and (s1n6477,n5014,n3425);
and (n6478,n6479,n5038);
wire s0n6479,s1n6479,notn6479;
or (n6479,s0n6479,s1n6479);
not(notn6479,n5014);
and (s0n6479,notn6479,n1769);
and (s1n6479,n5014,n2151);
and (n6481,n6438,n6482);
or (n6482,n6483,n6570,n6748);
and (n6483,n6484,n6527);
wire s0n6484,s1n6484,notn6484;
or (n6484,s0n6484,s1n6484);
not(notn6484,n4966);
and (s0n6484,notn6484,n6485);
and (s1n6484,n4966,n6526);
or (n6485,1'b0,n6486,n6496,n6506,n6516);
and (n6486,n6487,n2718);
or (n6487,1'b0,n6488,n6490,n6492,n6494);
and (n6488,n6489,n5016);
wire s0n6489,s1n6489,notn6489;
or (n6489,s0n6489,s1n6489);
not(notn6489,n5014);
and (s0n6489,notn6489,n3469);
and (s1n6489,n5014,n3538);
and (n6490,n6491,n5028);
wire s0n6491,s1n6491,notn6491;
or (n6491,s0n6491,s1n6491);
not(notn6491,n5014);
and (s0n6491,notn6491,n3473);
and (s1n6491,n5014,n3469);
and (n6492,n6493,n5033);
wire s0n6493,s1n6493,notn6493;
or (n6493,s0n6493,s1n6493);
not(notn6493,n5014);
and (s0n6493,notn6493,n3477);
and (s1n6493,n5014,n3473);
and (n6494,n6495,n5038);
wire s0n6495,s1n6495,notn6495;
or (n6495,s0n6495,s1n6495);
not(notn6495,n5014);
and (s0n6495,notn6495,n3481);
and (s1n6495,n5014,n3477);
and (n6496,n6497,n2730);
or (n6497,1'b0,n6498,n6500,n6502,n6504);
and (n6498,n6499,n5016);
wire s0n6499,s1n6499,notn6499;
or (n6499,s0n6499,s1n6499);
not(notn6499,n5014);
and (s0n6499,notn6499,n3487);
and (s1n6499,n5014,n3481);
and (n6500,n6501,n5028);
wire s0n6501,s1n6501,notn6501;
or (n6501,s0n6501,s1n6501);
not(notn6501,n5014);
and (s0n6501,notn6501,n3491);
and (s1n6501,n5014,n3487);
and (n6502,n6503,n5033);
wire s0n6503,s1n6503,notn6503;
or (n6503,s0n6503,s1n6503);
not(notn6503,n5014);
and (s0n6503,notn6503,n3495);
and (s1n6503,n5014,n3491);
and (n6504,n6505,n5038);
wire s0n6505,s1n6505,notn6505;
or (n6505,s0n6505,s1n6505);
not(notn6505,n5014);
and (s0n6505,notn6505,n3499);
and (s1n6505,n5014,n3495);
and (n6506,n6507,n2742);
or (n6507,1'b0,n6508,n6510,n6512,n6514);
and (n6508,n6509,n5016);
wire s0n6509,s1n6509,notn6509;
or (n6509,s0n6509,s1n6509);
not(notn6509,n5014);
and (s0n6509,notn6509,n3505);
and (s1n6509,n5014,n3553);
and (n6510,n6511,n5028);
wire s0n6511,s1n6511,notn6511;
or (n6511,s0n6511,s1n6511);
not(notn6511,n5014);
and (s0n6511,notn6511,n3509);
and (s1n6511,n5014,n3505);
and (n6512,n6513,n5033);
wire s0n6513,s1n6513,notn6513;
or (n6513,s0n6513,s1n6513);
not(notn6513,n5014);
and (s0n6513,notn6513,n3513);
and (s1n6513,n5014,n3509);
and (n6514,n6515,n5038);
wire s0n6515,s1n6515,notn6515;
or (n6515,s0n6515,s1n6515);
not(notn6515,n5014);
and (s0n6515,notn6515,n3517);
and (s1n6515,n5014,n3513);
and (n6516,n6517,n2752);
or (n6517,1'b0,n6518,n6520,n6522,n6524);
and (n6518,n6519,n5016);
wire s0n6519,s1n6519,notn6519;
or (n6519,s0n6519,s1n6519);
not(notn6519,n5014);
and (s0n6519,notn6519,n3523);
and (s1n6519,n5014,n3517);
and (n6520,n6521,n5028);
wire s0n6521,s1n6521,notn6521;
or (n6521,s0n6521,s1n6521);
not(notn6521,n5014);
and (s0n6521,notn6521,n3527);
and (s1n6521,n5014,n3523);
and (n6522,n6523,n5033);
wire s0n6523,s1n6523,notn6523;
or (n6523,s0n6523,s1n6523);
not(notn6523,n5014);
and (s0n6523,notn6523,n1331);
and (s1n6523,n5014,n3527);
and (n6524,n6525,n5038);
wire s0n6525,s1n6525,notn6525;
or (n6525,s0n6525,s1n6525);
not(notn6525,n5014);
and (s0n6525,notn6525,n827);
and (s1n6525,n5014,n1331);
wire s0n6527,s1n6527,notn6527;
or (n6527,s0n6527,s1n6527);
not(notn6527,n4966);
and (s0n6527,notn6527,n6528);
and (s1n6527,n4966,n6569);
or (n6528,1'b0,n6529,n6539,n6549,n6559);
and (n6529,n6530,n2718);
or (n6530,1'b0,n6531,n6533,n6535,n6537);
and (n6531,n6532,n5016);
wire s0n6532,s1n6532,notn6532;
or (n6532,s0n6532,s1n6532);
not(notn6532,n5014);
and (s0n6532,notn6532,n3470);
and (s1n6532,n5014,n3539);
and (n6533,n6534,n5028);
wire s0n6534,s1n6534,notn6534;
or (n6534,s0n6534,s1n6534);
not(notn6534,n5014);
and (s0n6534,notn6534,n3474);
and (s1n6534,n5014,n3470);
and (n6535,n6536,n5033);
wire s0n6536,s1n6536,notn6536;
or (n6536,s0n6536,s1n6536);
not(notn6536,n5014);
and (s0n6536,notn6536,n3478);
and (s1n6536,n5014,n3474);
and (n6537,n6538,n5038);
wire s0n6538,s1n6538,notn6538;
or (n6538,s0n6538,s1n6538);
not(notn6538,n5014);
and (s0n6538,notn6538,n3482);
and (s1n6538,n5014,n3478);
and (n6539,n6540,n2730);
or (n6540,1'b0,n6541,n6543,n6545,n6547);
and (n6541,n6542,n5016);
wire s0n6542,s1n6542,notn6542;
or (n6542,s0n6542,s1n6542);
not(notn6542,n5014);
and (s0n6542,notn6542,n3488);
and (s1n6542,n5014,n3482);
and (n6543,n6544,n5028);
wire s0n6544,s1n6544,notn6544;
or (n6544,s0n6544,s1n6544);
not(notn6544,n5014);
and (s0n6544,notn6544,n3492);
and (s1n6544,n5014,n3488);
and (n6545,n6546,n5033);
wire s0n6546,s1n6546,notn6546;
or (n6546,s0n6546,s1n6546);
not(notn6546,n5014);
and (s0n6546,notn6546,n3496);
and (s1n6546,n5014,n3492);
and (n6547,n6548,n5038);
wire s0n6548,s1n6548,notn6548;
or (n6548,s0n6548,s1n6548);
not(notn6548,n5014);
and (s0n6548,notn6548,n3500);
and (s1n6548,n5014,n3496);
and (n6549,n6550,n2742);
or (n6550,1'b0,n6551,n6553,n6555,n6557);
and (n6551,n6552,n5016);
wire s0n6552,s1n6552,notn6552;
or (n6552,s0n6552,s1n6552);
not(notn6552,n5014);
and (s0n6552,notn6552,n3506);
and (s1n6552,n5014,n3554);
and (n6553,n6554,n5028);
wire s0n6554,s1n6554,notn6554;
or (n6554,s0n6554,s1n6554);
not(notn6554,n5014);
and (s0n6554,notn6554,n3510);
and (s1n6554,n5014,n3506);
and (n6555,n6556,n5033);
wire s0n6556,s1n6556,notn6556;
or (n6556,s0n6556,s1n6556);
not(notn6556,n5014);
and (s0n6556,notn6556,n3514);
and (s1n6556,n5014,n3510);
and (n6557,n6558,n5038);
wire s0n6558,s1n6558,notn6558;
or (n6558,s0n6558,s1n6558);
not(notn6558,n5014);
and (s0n6558,notn6558,n3518);
and (s1n6558,n5014,n3514);
and (n6559,n6560,n2752);
or (n6560,1'b0,n6561,n6563,n6565,n6567);
and (n6561,n6562,n5016);
wire s0n6562,s1n6562,notn6562;
or (n6562,s0n6562,s1n6562);
not(notn6562,n5014);
and (s0n6562,notn6562,n3524);
and (s1n6562,n5014,n3518);
and (n6563,n6564,n5028);
wire s0n6564,s1n6564,notn6564;
or (n6564,s0n6564,s1n6564);
not(notn6564,n5014);
and (s0n6564,notn6564,n3528);
and (s1n6564,n5014,n3524);
and (n6565,n6566,n5033);
wire s0n6566,s1n6566,notn6566;
or (n6566,s0n6566,s1n6566);
not(notn6566,n5014);
and (s0n6566,notn6566,n2167);
and (s1n6566,n5014,n3528);
and (n6567,n6568,n5038);
wire s0n6568,s1n6568,notn6568;
or (n6568,s0n6568,s1n6568);
not(notn6568,n5014);
and (s0n6568,notn6568,n1790);
and (s1n6568,n5014,n2167);
and (n6570,n6527,n6571);
or (n6571,n6572,n6659,n6747);
and (n6572,n6573,n6616);
wire s0n6573,s1n6573,notn6573;
or (n6573,s0n6573,s1n6573);
not(notn6573,n4966);
and (s0n6573,notn6573,n6574);
and (s1n6573,n4966,n6615);
or (n6574,1'b0,n6575,n6585,n6595,n6605);
and (n6575,n6576,n2718);
or (n6576,1'b0,n6577,n6579,n6581,n6583);
and (n6577,n6578,n5016);
wire s0n6578,s1n6578,notn6578;
or (n6578,s0n6578,s1n6578);
not(notn6578,n5014);
and (s0n6578,notn6578,n3572);
and (s1n6578,n5014,n3641);
and (n6579,n6580,n5028);
wire s0n6580,s1n6580,notn6580;
or (n6580,s0n6580,s1n6580);
not(notn6580,n5014);
and (s0n6580,notn6580,n3576);
and (s1n6580,n5014,n3572);
and (n6581,n6582,n5033);
wire s0n6582,s1n6582,notn6582;
or (n6582,s0n6582,s1n6582);
not(notn6582,n5014);
and (s0n6582,notn6582,n3580);
and (s1n6582,n5014,n3576);
and (n6583,n6584,n5038);
wire s0n6584,s1n6584,notn6584;
or (n6584,s0n6584,s1n6584);
not(notn6584,n5014);
and (s0n6584,notn6584,n3584);
and (s1n6584,n5014,n3580);
and (n6585,n6586,n2730);
or (n6586,1'b0,n6587,n6589,n6591,n6593);
and (n6587,n6588,n5016);
wire s0n6588,s1n6588,notn6588;
or (n6588,s0n6588,s1n6588);
not(notn6588,n5014);
and (s0n6588,notn6588,n3590);
and (s1n6588,n5014,n3584);
and (n6589,n6590,n5028);
wire s0n6590,s1n6590,notn6590;
or (n6590,s0n6590,s1n6590);
not(notn6590,n5014);
and (s0n6590,notn6590,n3594);
and (s1n6590,n5014,n3590);
and (n6591,n6592,n5033);
wire s0n6592,s1n6592,notn6592;
or (n6592,s0n6592,s1n6592);
not(notn6592,n5014);
and (s0n6592,notn6592,n3598);
and (s1n6592,n5014,n3594);
and (n6593,n6594,n5038);
wire s0n6594,s1n6594,notn6594;
or (n6594,s0n6594,s1n6594);
not(notn6594,n5014);
and (s0n6594,notn6594,n3602);
and (s1n6594,n5014,n3598);
and (n6595,n6596,n2742);
or (n6596,1'b0,n6597,n6599,n6601,n6603);
and (n6597,n6598,n5016);
wire s0n6598,s1n6598,notn6598;
or (n6598,s0n6598,s1n6598);
not(notn6598,n5014);
and (s0n6598,notn6598,n3608);
and (s1n6598,n5014,n3656);
and (n6599,n6600,n5028);
wire s0n6600,s1n6600,notn6600;
or (n6600,s0n6600,s1n6600);
not(notn6600,n5014);
and (s0n6600,notn6600,n3612);
and (s1n6600,n5014,n3608);
and (n6601,n6602,n5033);
wire s0n6602,s1n6602,notn6602;
or (n6602,s0n6602,s1n6602);
not(notn6602,n5014);
and (s0n6602,notn6602,n3616);
and (s1n6602,n5014,n3612);
and (n6603,n6604,n5038);
wire s0n6604,s1n6604,notn6604;
or (n6604,s0n6604,s1n6604);
not(notn6604,n5014);
and (s0n6604,notn6604,n3620);
and (s1n6604,n5014,n3616);
and (n6605,n6606,n2752);
or (n6606,1'b0,n6607,n6609,n6611,n6613);
and (n6607,n6608,n5016);
wire s0n6608,s1n6608,notn6608;
or (n6608,s0n6608,s1n6608);
not(notn6608,n5014);
and (s0n6608,notn6608,n3626);
and (s1n6608,n5014,n3620);
and (n6609,n6610,n5028);
wire s0n6610,s1n6610,notn6610;
or (n6610,s0n6610,s1n6610);
not(notn6610,n5014);
and (s0n6610,notn6610,n3630);
and (s1n6610,n5014,n3626);
and (n6611,n6612,n5033);
wire s0n6612,s1n6612,notn6612;
or (n6612,s0n6612,s1n6612);
not(notn6612,n5014);
and (s0n6612,notn6612,n1347);
and (s1n6612,n5014,n3630);
and (n6613,n6614,n5038);
wire s0n6614,s1n6614,notn6614;
or (n6614,s0n6614,s1n6614);
not(notn6614,n5014);
and (s0n6614,notn6614,n843);
and (s1n6614,n5014,n1347);
wire s0n6616,s1n6616,notn6616;
or (n6616,s0n6616,s1n6616);
not(notn6616,n4966);
and (s0n6616,notn6616,n6617);
and (s1n6616,n4966,n6658);
or (n6617,1'b0,n6618,n6628,n6638,n6648);
and (n6618,n6619,n2718);
or (n6619,1'b0,n6620,n6622,n6624,n6626);
and (n6620,n6621,n5016);
wire s0n6621,s1n6621,notn6621;
or (n6621,s0n6621,s1n6621);
not(notn6621,n5014);
and (s0n6621,notn6621,n3573);
and (s1n6621,n5014,n3642);
and (n6622,n6623,n5028);
wire s0n6623,s1n6623,notn6623;
or (n6623,s0n6623,s1n6623);
not(notn6623,n5014);
and (s0n6623,notn6623,n3577);
and (s1n6623,n5014,n3573);
and (n6624,n6625,n5033);
wire s0n6625,s1n6625,notn6625;
or (n6625,s0n6625,s1n6625);
not(notn6625,n5014);
and (s0n6625,notn6625,n3581);
and (s1n6625,n5014,n3577);
and (n6626,n6627,n5038);
wire s0n6627,s1n6627,notn6627;
or (n6627,s0n6627,s1n6627);
not(notn6627,n5014);
and (s0n6627,notn6627,n3585);
and (s1n6627,n5014,n3581);
and (n6628,n6629,n2730);
or (n6629,1'b0,n6630,n6632,n6634,n6636);
and (n6630,n6631,n5016);
wire s0n6631,s1n6631,notn6631;
or (n6631,s0n6631,s1n6631);
not(notn6631,n5014);
and (s0n6631,notn6631,n3591);
and (s1n6631,n5014,n3585);
and (n6632,n6633,n5028);
wire s0n6633,s1n6633,notn6633;
or (n6633,s0n6633,s1n6633);
not(notn6633,n5014);
and (s0n6633,notn6633,n3595);
and (s1n6633,n5014,n3591);
and (n6634,n6635,n5033);
wire s0n6635,s1n6635,notn6635;
or (n6635,s0n6635,s1n6635);
not(notn6635,n5014);
and (s0n6635,notn6635,n3599);
and (s1n6635,n5014,n3595);
and (n6636,n6637,n5038);
wire s0n6637,s1n6637,notn6637;
or (n6637,s0n6637,s1n6637);
not(notn6637,n5014);
and (s0n6637,notn6637,n3603);
and (s1n6637,n5014,n3599);
and (n6638,n6639,n2742);
or (n6639,1'b0,n6640,n6642,n6644,n6646);
and (n6640,n6641,n5016);
wire s0n6641,s1n6641,notn6641;
or (n6641,s0n6641,s1n6641);
not(notn6641,n5014);
and (s0n6641,notn6641,n3609);
and (s1n6641,n5014,n3657);
and (n6642,n6643,n5028);
wire s0n6643,s1n6643,notn6643;
or (n6643,s0n6643,s1n6643);
not(notn6643,n5014);
and (s0n6643,notn6643,n3613);
and (s1n6643,n5014,n3609);
and (n6644,n6645,n5033);
wire s0n6645,s1n6645,notn6645;
or (n6645,s0n6645,s1n6645);
not(notn6645,n5014);
and (s0n6645,notn6645,n3617);
and (s1n6645,n5014,n3613);
and (n6646,n6647,n5038);
wire s0n6647,s1n6647,notn6647;
or (n6647,s0n6647,s1n6647);
not(notn6647,n5014);
and (s0n6647,notn6647,n3621);
and (s1n6647,n5014,n3617);
and (n6648,n6649,n2752);
or (n6649,1'b0,n6650,n6652,n6654,n6656);
and (n6650,n6651,n5016);
wire s0n6651,s1n6651,notn6651;
or (n6651,s0n6651,s1n6651);
not(notn6651,n5014);
and (s0n6651,notn6651,n3627);
and (s1n6651,n5014,n3621);
and (n6652,n6653,n5028);
wire s0n6653,s1n6653,notn6653;
or (n6653,s0n6653,s1n6653);
not(notn6653,n5014);
and (s0n6653,notn6653,n3631);
and (s1n6653,n5014,n3627);
and (n6654,n6655,n5033);
wire s0n6655,s1n6655,notn6655;
or (n6655,s0n6655,s1n6655);
not(notn6655,n5014);
and (s0n6655,notn6655,n2184);
and (s1n6655,n5014,n3631);
and (n6656,n6657,n5038);
wire s0n6657,s1n6657,notn6657;
or (n6657,s0n6657,s1n6657);
not(notn6657,n5014);
and (s0n6657,notn6657,n1820);
and (s1n6657,n5014,n2184);
and (n6659,n6616,n6660);
and (n6660,n6661,n6704);
wire s0n6661,s1n6661,notn6661;
or (n6661,s0n6661,s1n6661);
not(notn6661,n4966);
and (s0n6661,notn6661,n6662);
and (s1n6661,n4966,n6703);
or (n6662,1'b0,n6663,n6673,n6683,n6693);
and (n6663,n6664,n2718);
or (n6664,1'b0,n6665,n6667,n6669,n6671);
and (n6665,n6666,n5016);
wire s0n6666,s1n6666,notn6666;
or (n6666,s0n6666,s1n6666);
not(notn6666,n5014);
and (s0n6666,notn6666,n3674);
and (s1n6666,n5014,n3743);
and (n6667,n6668,n5028);
wire s0n6668,s1n6668,notn6668;
or (n6668,s0n6668,s1n6668);
not(notn6668,n5014);
and (s0n6668,notn6668,n3678);
and (s1n6668,n5014,n3674);
and (n6669,n6670,n5033);
wire s0n6670,s1n6670,notn6670;
or (n6670,s0n6670,s1n6670);
not(notn6670,n5014);
and (s0n6670,notn6670,n3682);
and (s1n6670,n5014,n3678);
and (n6671,n6672,n5038);
wire s0n6672,s1n6672,notn6672;
or (n6672,s0n6672,s1n6672);
not(notn6672,n5014);
and (s0n6672,notn6672,n3686);
and (s1n6672,n5014,n3682);
and (n6673,n6674,n2730);
or (n6674,1'b0,n6675,n6677,n6679,n6681);
and (n6675,n6676,n5016);
wire s0n6676,s1n6676,notn6676;
or (n6676,s0n6676,s1n6676);
not(notn6676,n5014);
and (s0n6676,notn6676,n3692);
and (s1n6676,n5014,n3686);
and (n6677,n6678,n5028);
wire s0n6678,s1n6678,notn6678;
or (n6678,s0n6678,s1n6678);
not(notn6678,n5014);
and (s0n6678,notn6678,n3696);
and (s1n6678,n5014,n3692);
and (n6679,n6680,n5033);
wire s0n6680,s1n6680,notn6680;
or (n6680,s0n6680,s1n6680);
not(notn6680,n5014);
and (s0n6680,notn6680,n3700);
and (s1n6680,n5014,n3696);
and (n6681,n6682,n5038);
wire s0n6682,s1n6682,notn6682;
or (n6682,s0n6682,s1n6682);
not(notn6682,n5014);
and (s0n6682,notn6682,n3704);
and (s1n6682,n5014,n3700);
and (n6683,n6684,n2742);
or (n6684,1'b0,n6685,n6687,n6689,n6691);
and (n6685,n6686,n5016);
wire s0n6686,s1n6686,notn6686;
or (n6686,s0n6686,s1n6686);
not(notn6686,n5014);
and (s0n6686,notn6686,n3710);
and (s1n6686,n5014,n3758);
and (n6687,n6688,n5028);
wire s0n6688,s1n6688,notn6688;
or (n6688,s0n6688,s1n6688);
not(notn6688,n5014);
and (s0n6688,notn6688,n3714);
and (s1n6688,n5014,n3710);
and (n6689,n6690,n5033);
wire s0n6690,s1n6690,notn6690;
or (n6690,s0n6690,s1n6690);
not(notn6690,n5014);
and (s0n6690,notn6690,n3718);
and (s1n6690,n5014,n3714);
and (n6691,n6692,n5038);
wire s0n6692,s1n6692,notn6692;
or (n6692,s0n6692,s1n6692);
not(notn6692,n5014);
and (s0n6692,notn6692,n3722);
and (s1n6692,n5014,n3718);
and (n6693,n6694,n2752);
or (n6694,1'b0,n6695,n6697,n6699,n6701);
and (n6695,n6696,n5016);
wire s0n6696,s1n6696,notn6696;
or (n6696,s0n6696,s1n6696);
not(notn6696,n5014);
and (s0n6696,notn6696,n3728);
and (s1n6696,n5014,n3722);
and (n6697,n6698,n5028);
wire s0n6698,s1n6698,notn6698;
or (n6698,s0n6698,s1n6698);
not(notn6698,n5014);
and (s0n6698,notn6698,n3732);
and (s1n6698,n5014,n3728);
and (n6699,n6700,n5033);
wire s0n6700,s1n6700,notn6700;
or (n6700,s0n6700,s1n6700);
not(notn6700,n5014);
and (s0n6700,notn6700,n1362);
and (s1n6700,n5014,n3732);
and (n6701,n6702,n5038);
wire s0n6702,s1n6702,notn6702;
or (n6702,s0n6702,s1n6702);
not(notn6702,n5014);
and (s0n6702,notn6702,n858);
and (s1n6702,n5014,n1362);
wire s0n6704,s1n6704,notn6704;
or (n6704,s0n6704,s1n6704);
not(notn6704,n4966);
and (s0n6704,notn6704,n6705);
and (s1n6704,n4966,n6746);
or (n6705,1'b0,n6706,n6716,n6726,n6736);
and (n6706,n6707,n2718);
or (n6707,1'b0,n6708,n6710,n6712,n6714);
and (n6708,n6709,n5016);
wire s0n6709,s1n6709,notn6709;
or (n6709,s0n6709,s1n6709);
not(notn6709,n5014);
and (s0n6709,notn6709,n3675);
and (s1n6709,n5014,n3744);
and (n6710,n6711,n5028);
wire s0n6711,s1n6711,notn6711;
or (n6711,s0n6711,s1n6711);
not(notn6711,n5014);
and (s0n6711,notn6711,n3679);
and (s1n6711,n5014,n3675);
and (n6712,n6713,n5033);
wire s0n6713,s1n6713,notn6713;
or (n6713,s0n6713,s1n6713);
not(notn6713,n5014);
and (s0n6713,notn6713,n3683);
and (s1n6713,n5014,n3679);
and (n6714,n6715,n5038);
wire s0n6715,s1n6715,notn6715;
or (n6715,s0n6715,s1n6715);
not(notn6715,n5014);
and (s0n6715,notn6715,n3687);
and (s1n6715,n5014,n3683);
and (n6716,n6717,n2730);
or (n6717,1'b0,n6718,n6720,n6722,n6724);
and (n6718,n6719,n5016);
wire s0n6719,s1n6719,notn6719;
or (n6719,s0n6719,s1n6719);
not(notn6719,n5014);
and (s0n6719,notn6719,n3693);
and (s1n6719,n5014,n3687);
and (n6720,n6721,n5028);
wire s0n6721,s1n6721,notn6721;
or (n6721,s0n6721,s1n6721);
not(notn6721,n5014);
and (s0n6721,notn6721,n3697);
and (s1n6721,n5014,n3693);
and (n6722,n6723,n5033);
wire s0n6723,s1n6723,notn6723;
or (n6723,s0n6723,s1n6723);
not(notn6723,n5014);
and (s0n6723,notn6723,n3701);
and (s1n6723,n5014,n3697);
and (n6724,n6725,n5038);
wire s0n6725,s1n6725,notn6725;
or (n6725,s0n6725,s1n6725);
not(notn6725,n5014);
and (s0n6725,notn6725,n3705);
and (s1n6725,n5014,n3701);
and (n6726,n6727,n2742);
or (n6727,1'b0,n6728,n6730,n6732,n6734);
and (n6728,n6729,n5016);
wire s0n6729,s1n6729,notn6729;
or (n6729,s0n6729,s1n6729);
not(notn6729,n5014);
and (s0n6729,notn6729,n3711);
and (s1n6729,n5014,n3759);
and (n6730,n6731,n5028);
wire s0n6731,s1n6731,notn6731;
or (n6731,s0n6731,s1n6731);
not(notn6731,n5014);
and (s0n6731,notn6731,n3715);
and (s1n6731,n5014,n3711);
and (n6732,n6733,n5033);
wire s0n6733,s1n6733,notn6733;
or (n6733,s0n6733,s1n6733);
not(notn6733,n5014);
and (s0n6733,notn6733,n3719);
and (s1n6733,n5014,n3715);
and (n6734,n6735,n5038);
wire s0n6735,s1n6735,notn6735;
or (n6735,s0n6735,s1n6735);
not(notn6735,n5014);
and (s0n6735,notn6735,n3723);
and (s1n6735,n5014,n3719);
and (n6736,n6737,n2752);
or (n6737,1'b0,n6738,n6740,n6742,n6744);
and (n6738,n6739,n5016);
wire s0n6739,s1n6739,notn6739;
or (n6739,s0n6739,s1n6739);
not(notn6739,n5014);
and (s0n6739,notn6739,n3729);
and (s1n6739,n5014,n3723);
and (n6740,n6741,n5028);
wire s0n6741,s1n6741,notn6741;
or (n6741,s0n6741,s1n6741);
not(notn6741,n5014);
and (s0n6741,notn6741,n3733);
and (s1n6741,n5014,n3729);
and (n6742,n6743,n5033);
wire s0n6743,s1n6743,notn6743;
or (n6743,s0n6743,s1n6743);
not(notn6743,n5014);
and (s0n6743,notn6743,n2199);
and (s1n6743,n5014,n3733);
and (n6744,n6745,n5038);
wire s0n6745,s1n6745,notn6745;
or (n6745,s0n6745,s1n6745);
not(notn6745,n5014);
and (s0n6745,notn6745,n1843);
and (s1n6745,n5014,n2199);
and (n6747,n6573,n6660);
and (n6748,n6484,n6571);
and (n6749,n6395,n6482);
and (n6750,n6306,n6393);
and (n6751,n6217,n6304);
and (n6752,n6128,n6215);
and (n6753,n6039,n6126);
and (n6754,n6032,n6037);
and (n6755,n6025,n6030);
not (n6756,n6757);
xor (n6757,n6758,n6763);
xor (n6758,n6759,n6761);
wire s0n6759,s1n6759,notn6759;
or (n6759,s0n6759,s1n6759);
not(notn6759,n4966);
and (s0n6759,notn6759,1'b0);
and (s1n6759,n4966,n6760);
wire s0n6761,s1n6761,notn6761;
or (n6761,s0n6761,s1n6761);
not(notn6761,n4966);
and (s0n6761,notn6761,1'b0);
and (s1n6761,n4966,n6762);
or (n6763,n6764,n6769,n7351);
and (n6764,n6765,n6767);
wire s0n6765,s1n6765,notn6765;
or (n6765,s0n6765,s1n6765);
not(notn6765,n4966);
and (s0n6765,notn6765,1'b0);
and (s1n6765,n4966,n6766);
wire s0n6767,s1n6767,notn6767;
or (n6767,s0n6767,s1n6767);
not(notn6767,n4966);
and (s0n6767,notn6767,1'b0);
and (s1n6767,n4966,n6768);
and (n6769,n6767,n6770);
or (n6770,n6771,n6776,n7350);
and (n6771,n6772,n6774);
wire s0n6772,s1n6772,notn6772;
or (n6772,s0n6772,s1n6772);
not(notn6772,n4966);
and (s0n6772,notn6772,1'b0);
and (s1n6772,n4966,n6773);
wire s0n6774,s1n6774,notn6774;
or (n6774,s0n6774,s1n6774);
not(notn6774,n4966);
and (s0n6774,notn6774,1'b0);
and (s1n6774,n4966,n6775);
and (n6776,n6774,n6777);
or (n6777,n6778,n6783,n7349);
and (n6778,n6779,n6781);
wire s0n6779,s1n6779,notn6779;
or (n6779,s0n6779,s1n6779);
not(notn6779,n4966);
and (s0n6779,notn6779,1'b0);
and (s1n6779,n4966,n6780);
wire s0n6781,s1n6781,notn6781;
or (n6781,s0n6781,s1n6781);
not(notn6781,n4966);
and (s0n6781,notn6781,1'b0);
and (s1n6781,n4966,n6782);
and (n6783,n6781,n6784);
or (n6784,n6785,n6790,n7348);
and (n6785,n6786,n6788);
wire s0n6786,s1n6786,notn6786;
or (n6786,s0n6786,s1n6786);
not(notn6786,n4966);
and (s0n6786,notn6786,1'b0);
and (s1n6786,n4966,n6787);
wire s0n6788,s1n6788,notn6788;
or (n6788,s0n6788,s1n6788);
not(notn6788,n4966);
and (s0n6788,notn6788,1'b0);
and (s1n6788,n4966,n6789);
and (n6790,n6788,n6791);
or (n6791,n6792,n6859,n7347);
and (n6792,n6793,n6825);
wire s0n6793,s1n6793,notn6793;
or (n6793,s0n6793,s1n6793);
not(notn6793,n4966);
and (s0n6793,notn6793,n6794);
and (s1n6793,n4966,n6824);
or (n6794,1'b0,n6795,n6796,n6797,n6812);
and (n6795,n5114,n2718);
and (n6796,n5129,n2730);
and (n6797,n6798,n2742);
or (n6798,1'b0,n6799,n6803,n6806,n6809);
and (n6799,n6800,n5016);
wire s0n6800,s1n6800,notn6800;
or (n6800,s0n6800,s1n6800);
not(notn6800,n5014);
and (s0n6800,notn6800,n6801);
and (s1n6800,n5014,n6802);
and (n6803,n6804,n5028);
wire s0n6804,s1n6804,notn6804;
or (n6804,s0n6804,s1n6804);
not(notn6804,n5014);
and (s0n6804,notn6804,n6805);
and (s1n6804,n5014,n6801);
and (n6806,n6807,n5033);
wire s0n6807,s1n6807,notn6807;
or (n6807,s0n6807,s1n6807);
not(notn6807,n5014);
and (s0n6807,notn6807,n6808);
and (s1n6807,n5014,n6805);
and (n6809,n6810,n5038);
wire s0n6810,s1n6810,notn6810;
or (n6810,s0n6810,s1n6810);
not(notn6810,n5014);
and (s0n6810,notn6810,n6811);
and (s1n6810,n5014,n6808);
and (n6812,n6813,n2752);
or (n6813,1'b0,n6814,n6817,n6820,n6822);
and (n6814,n6815,n5016);
wire s0n6815,s1n6815,notn6815;
or (n6815,s0n6815,s1n6815);
not(notn6815,n5014);
and (s0n6815,notn6815,n6816);
and (s1n6815,n5014,n6811);
and (n6817,n6818,n5028);
wire s0n6818,s1n6818,notn6818;
or (n6818,s0n6818,s1n6818);
not(notn6818,n5014);
and (s0n6818,notn6818,n6819);
and (s1n6818,n5014,n6816);
and (n6820,n6821,n5033);
wire s0n6821,s1n6821,notn6821;
or (n6821,s0n6821,s1n6821);
not(notn6821,n5014);
and (s0n6821,notn6821,n2091);
and (s1n6821,n5014,n6819);
and (n6822,n6823,n5038);
wire s0n6823,s1n6823,notn6823;
or (n6823,s0n6823,s1n6823);
not(notn6823,n5014);
and (s0n6823,notn6823,n1696);
and (s1n6823,n5014,n2091);
wire s0n6825,s1n6825,notn6825;
or (n6825,s0n6825,s1n6825);
not(notn6825,n4966);
and (s0n6825,notn6825,n6826);
and (s1n6825,n4966,n6858);
or (n6826,1'b0,n6827,n6842,n6856,n6857);
and (n6827,n6828,n2718);
or (n6828,1'b0,n6829,n6833,n6836,n6839);
and (n6829,n6830,n5016);
wire s0n6830,s1n6830,notn6830;
or (n6830,s0n6830,s1n6830);
not(notn6830,n5014);
and (s0n6830,notn6830,n6831);
and (s1n6830,n5014,n6832);
and (n6833,n6834,n5028);
wire s0n6834,s1n6834,notn6834;
or (n6834,s0n6834,s1n6834);
not(notn6834,n5014);
and (s0n6834,notn6834,n6835);
and (s1n6834,n5014,n6831);
and (n6836,n6837,n5033);
wire s0n6837,s1n6837,notn6837;
or (n6837,s0n6837,s1n6837);
not(notn6837,n5014);
and (s0n6837,notn6837,n6838);
and (s1n6837,n5014,n6835);
and (n6839,n6840,n5038);
wire s0n6840,s1n6840,notn6840;
or (n6840,s0n6840,s1n6840);
not(notn6840,n5014);
and (s0n6840,notn6840,n6841);
and (s1n6840,n5014,n6838);
and (n6842,n6843,n2730);
or (n6843,1'b0,n6844,n6847,n6850,n6853);
and (n6844,n6845,n5016);
wire s0n6845,s1n6845,notn6845;
or (n6845,s0n6845,s1n6845);
not(notn6845,n5014);
and (s0n6845,notn6845,n6846);
and (s1n6845,n5014,n6841);
and (n6847,n6848,n5028);
wire s0n6848,s1n6848,notn6848;
or (n6848,s0n6848,s1n6848);
not(notn6848,n5014);
and (s0n6848,notn6848,n6849);
and (s1n6848,n5014,n6846);
and (n6850,n6851,n5033);
wire s0n6851,s1n6851,notn6851;
or (n6851,s0n6851,s1n6851);
not(notn6851,n5014);
and (s0n6851,notn6851,n6852);
and (s1n6851,n5014,n6849);
and (n6853,n6854,n5038);
wire s0n6854,s1n6854,notn6854;
or (n6854,s0n6854,s1n6854);
not(notn6854,n5014);
and (s0n6854,notn6854,n6855);
and (s1n6854,n5014,n6852);
and (n6856,n5009,n2742);
and (n6857,n5041,n2752);
and (n6859,n6825,n6860);
or (n6860,n6861,n6928,n7346);
and (n6861,n6862,n6894);
wire s0n6862,s1n6862,notn6862;
or (n6862,s0n6862,s1n6862);
not(notn6862,n4966);
and (s0n6862,notn6862,n6863);
and (s1n6862,n4966,n6893);
or (n6863,1'b0,n6864,n6865,n6866,n6881);
and (n6864,n5237,n2718);
and (n6865,n5252,n2730);
and (n6866,n6867,n2742);
or (n6867,1'b0,n6868,n6872,n6875,n6878);
and (n6868,n6869,n5016);
wire s0n6869,s1n6869,notn6869;
or (n6869,s0n6869,s1n6869);
not(notn6869,n5014);
and (s0n6869,notn6869,n6870);
and (s1n6869,n5014,n6871);
and (n6872,n6873,n5028);
wire s0n6873,s1n6873,notn6873;
or (n6873,s0n6873,s1n6873);
not(notn6873,n5014);
and (s0n6873,notn6873,n6874);
and (s1n6873,n5014,n6870);
and (n6875,n6876,n5033);
wire s0n6876,s1n6876,notn6876;
or (n6876,s0n6876,s1n6876);
not(notn6876,n5014);
and (s0n6876,notn6876,n6877);
and (s1n6876,n5014,n6874);
and (n6878,n6879,n5038);
wire s0n6879,s1n6879,notn6879;
or (n6879,s0n6879,s1n6879);
not(notn6879,n5014);
and (s0n6879,notn6879,n6880);
and (s1n6879,n5014,n6877);
and (n6881,n6882,n2752);
or (n6882,1'b0,n6883,n6886,n6889,n6891);
and (n6883,n6884,n5016);
wire s0n6884,s1n6884,notn6884;
or (n6884,s0n6884,s1n6884);
not(notn6884,n5014);
and (s0n6884,notn6884,n6885);
and (s1n6884,n5014,n6880);
and (n6886,n6887,n5028);
wire s0n6887,s1n6887,notn6887;
or (n6887,s0n6887,s1n6887);
not(notn6887,n5014);
and (s0n6887,notn6887,n6888);
and (s1n6887,n5014,n6885);
and (n6889,n6890,n5033);
wire s0n6890,s1n6890,notn6890;
or (n6890,s0n6890,s1n6890);
not(notn6890,n5014);
and (s0n6890,notn6890,n2107);
and (s1n6890,n5014,n6888);
and (n6891,n6892,n5038);
wire s0n6892,s1n6892,notn6892;
or (n6892,s0n6892,s1n6892);
not(notn6892,n5014);
and (s0n6892,notn6892,n1712);
and (s1n6892,n5014,n2107);
wire s0n6894,s1n6894,notn6894;
or (n6894,s0n6894,s1n6894);
not(notn6894,n4966);
and (s0n6894,notn6894,n6895);
and (s1n6894,n4966,n6927);
or (n6895,1'b0,n6896,n6911,n6925,n6926);
and (n6896,n6897,n2718);
or (n6897,1'b0,n6898,n6902,n6905,n6908);
and (n6898,n6899,n5016);
wire s0n6899,s1n6899,notn6899;
or (n6899,s0n6899,s1n6899);
not(notn6899,n5014);
and (s0n6899,notn6899,n6900);
and (s1n6899,n5014,n6901);
and (n6902,n6903,n5028);
wire s0n6903,s1n6903,notn6903;
or (n6903,s0n6903,s1n6903);
not(notn6903,n5014);
and (s0n6903,notn6903,n6904);
and (s1n6903,n5014,n6900);
and (n6905,n6906,n5033);
wire s0n6906,s1n6906,notn6906;
or (n6906,s0n6906,s1n6906);
not(notn6906,n5014);
and (s0n6906,notn6906,n6907);
and (s1n6906,n5014,n6904);
and (n6908,n6909,n5038);
wire s0n6909,s1n6909,notn6909;
or (n6909,s0n6909,s1n6909);
not(notn6909,n5014);
and (s0n6909,notn6909,n6910);
and (s1n6909,n5014,n6907);
and (n6911,n6912,n2730);
or (n6912,1'b0,n6913,n6916,n6919,n6922);
and (n6913,n6914,n5016);
wire s0n6914,s1n6914,notn6914;
or (n6914,s0n6914,s1n6914);
not(notn6914,n5014);
and (s0n6914,notn6914,n6915);
and (s1n6914,n5014,n6910);
and (n6916,n6917,n5028);
wire s0n6917,s1n6917,notn6917;
or (n6917,s0n6917,s1n6917);
not(notn6917,n5014);
and (s0n6917,notn6917,n6918);
and (s1n6917,n5014,n6915);
and (n6919,n6920,n5033);
wire s0n6920,s1n6920,notn6920;
or (n6920,s0n6920,s1n6920);
not(notn6920,n5014);
and (s0n6920,notn6920,n6921);
and (s1n6920,n5014,n6918);
and (n6922,n6923,n5038);
wire s0n6923,s1n6923,notn6923;
or (n6923,s0n6923,s1n6923);
not(notn6923,n5014);
and (s0n6923,notn6923,n6924);
and (s1n6923,n5014,n6921);
and (n6925,n5149,n2742);
and (n6926,n5164,n2752);
and (n6928,n6894,n6929);
or (n6929,n6930,n6997,n7345);
and (n6930,n6931,n6963);
wire s0n6931,s1n6931,notn6931;
or (n6931,s0n6931,s1n6931);
not(notn6931,n4966);
and (s0n6931,notn6931,n6932);
and (s1n6931,n4966,n6962);
or (n6932,1'b0,n6933,n6934,n6935,n6950);
and (n6933,n5360,n2718);
and (n6934,n5375,n2730);
and (n6935,n6936,n2742);
or (n6936,1'b0,n6937,n6941,n6944,n6947);
and (n6937,n6938,n5016);
wire s0n6938,s1n6938,notn6938;
or (n6938,s0n6938,s1n6938);
not(notn6938,n5014);
and (s0n6938,notn6938,n6939);
and (s1n6938,n5014,n6940);
and (n6941,n6942,n5028);
wire s0n6942,s1n6942,notn6942;
or (n6942,s0n6942,s1n6942);
not(notn6942,n5014);
and (s0n6942,notn6942,n6943);
and (s1n6942,n5014,n6939);
and (n6944,n6945,n5033);
wire s0n6945,s1n6945,notn6945;
or (n6945,s0n6945,s1n6945);
not(notn6945,n5014);
and (s0n6945,notn6945,n6946);
and (s1n6945,n5014,n6943);
and (n6947,n6948,n5038);
wire s0n6948,s1n6948,notn6948;
or (n6948,s0n6948,s1n6948);
not(notn6948,n5014);
and (s0n6948,notn6948,n6949);
and (s1n6948,n5014,n6946);
and (n6950,n6951,n2752);
or (n6951,1'b0,n6952,n6955,n6958,n6960);
and (n6952,n6953,n5016);
wire s0n6953,s1n6953,notn6953;
or (n6953,s0n6953,s1n6953);
not(notn6953,n5014);
and (s0n6953,notn6953,n6954);
and (s1n6953,n5014,n6949);
and (n6955,n6956,n5028);
wire s0n6956,s1n6956,notn6956;
or (n6956,s0n6956,s1n6956);
not(notn6956,n5014);
and (s0n6956,notn6956,n6957);
and (s1n6956,n5014,n6954);
and (n6958,n6959,n5033);
wire s0n6959,s1n6959,notn6959;
or (n6959,s0n6959,s1n6959);
not(notn6959,n5014);
and (s0n6959,notn6959,n2123);
and (s1n6959,n5014,n6957);
and (n6960,n6961,n5038);
wire s0n6961,s1n6961,notn6961;
or (n6961,s0n6961,s1n6961);
not(notn6961,n5014);
and (s0n6961,notn6961,n1731);
and (s1n6961,n5014,n2123);
wire s0n6963,s1n6963,notn6963;
or (n6963,s0n6963,s1n6963);
not(notn6963,n4966);
and (s0n6963,notn6963,n6964);
and (s1n6963,n4966,n6996);
or (n6964,1'b0,n6965,n6980,n6994,n6995);
and (n6965,n6966,n2718);
or (n6966,1'b0,n6967,n6971,n6974,n6977);
and (n6967,n6968,n5016);
wire s0n6968,s1n6968,notn6968;
or (n6968,s0n6968,s1n6968);
not(notn6968,n5014);
and (s0n6968,notn6968,n6969);
and (s1n6968,n5014,n6970);
and (n6971,n6972,n5028);
wire s0n6972,s1n6972,notn6972;
or (n6972,s0n6972,s1n6972);
not(notn6972,n5014);
and (s0n6972,notn6972,n6973);
and (s1n6972,n5014,n6969);
and (n6974,n6975,n5033);
wire s0n6975,s1n6975,notn6975;
or (n6975,s0n6975,s1n6975);
not(notn6975,n5014);
and (s0n6975,notn6975,n6976);
and (s1n6975,n5014,n6973);
and (n6977,n6978,n5038);
wire s0n6978,s1n6978,notn6978;
or (n6978,s0n6978,s1n6978);
not(notn6978,n5014);
and (s0n6978,notn6978,n6979);
and (s1n6978,n5014,n6976);
and (n6980,n6981,n2730);
or (n6981,1'b0,n6982,n6985,n6988,n6991);
and (n6982,n6983,n5016);
wire s0n6983,s1n6983,notn6983;
or (n6983,s0n6983,s1n6983);
not(notn6983,n5014);
and (s0n6983,notn6983,n6984);
and (s1n6983,n5014,n6979);
and (n6985,n6986,n5028);
wire s0n6986,s1n6986,notn6986;
or (n6986,s0n6986,s1n6986);
not(notn6986,n5014);
and (s0n6986,notn6986,n6987);
and (s1n6986,n5014,n6984);
and (n6988,n6989,n5033);
wire s0n6989,s1n6989,notn6989;
or (n6989,s0n6989,s1n6989);
not(notn6989,n5014);
and (s0n6989,notn6989,n6990);
and (s1n6989,n5014,n6987);
and (n6991,n6992,n5038);
wire s0n6992,s1n6992,notn6992;
or (n6992,s0n6992,s1n6992);
not(notn6992,n5014);
and (s0n6992,notn6992,n6993);
and (s1n6992,n5014,n6990);
and (n6994,n5272,n2742);
and (n6995,n5287,n2752);
and (n6997,n6963,n6998);
or (n6998,n6999,n7066,n7344);
and (n6999,n7000,n7032);
wire s0n7000,s1n7000,notn7000;
or (n7000,s0n7000,s1n7000);
not(notn7000,n4966);
and (s0n7000,notn7000,n7001);
and (s1n7000,n4966,n7031);
or (n7001,1'b0,n7002,n7003,n7004,n7019);
and (n7002,n5483,n2718);
and (n7003,n5498,n2730);
and (n7004,n7005,n2742);
or (n7005,1'b0,n7006,n7010,n7013,n7016);
and (n7006,n7007,n5016);
wire s0n7007,s1n7007,notn7007;
or (n7007,s0n7007,s1n7007);
not(notn7007,n5014);
and (s0n7007,notn7007,n7008);
and (s1n7007,n5014,n7009);
and (n7010,n7011,n5028);
wire s0n7011,s1n7011,notn7011;
or (n7011,s0n7011,s1n7011);
not(notn7011,n5014);
and (s0n7011,notn7011,n7012);
and (s1n7011,n5014,n7008);
and (n7013,n7014,n5033);
wire s0n7014,s1n7014,notn7014;
or (n7014,s0n7014,s1n7014);
not(notn7014,n5014);
and (s0n7014,notn7014,n7015);
and (s1n7014,n5014,n7012);
and (n7016,n7017,n5038);
wire s0n7017,s1n7017,notn7017;
or (n7017,s0n7017,s1n7017);
not(notn7017,n5014);
and (s0n7017,notn7017,n7018);
and (s1n7017,n5014,n7015);
and (n7019,n7020,n2752);
or (n7020,1'b0,n7021,n7024,n7027,n7029);
and (n7021,n7022,n5016);
wire s0n7022,s1n7022,notn7022;
or (n7022,s0n7022,s1n7022);
not(notn7022,n5014);
and (s0n7022,notn7022,n7023);
and (s1n7022,n5014,n7018);
and (n7024,n7025,n5028);
wire s0n7025,s1n7025,notn7025;
or (n7025,s0n7025,s1n7025);
not(notn7025,n5014);
and (s0n7025,notn7025,n7026);
and (s1n7025,n5014,n7023);
and (n7027,n7028,n5033);
wire s0n7028,s1n7028,notn7028;
or (n7028,s0n7028,s1n7028);
not(notn7028,n5014);
and (s0n7028,notn7028,n2139);
and (s1n7028,n5014,n7026);
and (n7029,n7030,n5038);
wire s0n7030,s1n7030,notn7030;
or (n7030,s0n7030,s1n7030);
not(notn7030,n5014);
and (s0n7030,notn7030,n1757);
and (s1n7030,n5014,n2139);
wire s0n7032,s1n7032,notn7032;
or (n7032,s0n7032,s1n7032);
not(notn7032,n4966);
and (s0n7032,notn7032,n7033);
and (s1n7032,n4966,n7065);
or (n7033,1'b0,n7034,n7049,n7063,n7064);
and (n7034,n7035,n2718);
or (n7035,1'b0,n7036,n7040,n7043,n7046);
and (n7036,n7037,n5016);
wire s0n7037,s1n7037,notn7037;
or (n7037,s0n7037,s1n7037);
not(notn7037,n5014);
and (s0n7037,notn7037,n7038);
and (s1n7037,n5014,n7039);
and (n7040,n7041,n5028);
wire s0n7041,s1n7041,notn7041;
or (n7041,s0n7041,s1n7041);
not(notn7041,n5014);
and (s0n7041,notn7041,n7042);
and (s1n7041,n5014,n7038);
and (n7043,n7044,n5033);
wire s0n7044,s1n7044,notn7044;
or (n7044,s0n7044,s1n7044);
not(notn7044,n5014);
and (s0n7044,notn7044,n7045);
and (s1n7044,n5014,n7042);
and (n7046,n7047,n5038);
wire s0n7047,s1n7047,notn7047;
or (n7047,s0n7047,s1n7047);
not(notn7047,n5014);
and (s0n7047,notn7047,n7048);
and (s1n7047,n5014,n7045);
and (n7049,n7050,n2730);
or (n7050,1'b0,n7051,n7054,n7057,n7060);
and (n7051,n7052,n5016);
wire s0n7052,s1n7052,notn7052;
or (n7052,s0n7052,s1n7052);
not(notn7052,n5014);
and (s0n7052,notn7052,n7053);
and (s1n7052,n5014,n7048);
and (n7054,n7055,n5028);
wire s0n7055,s1n7055,notn7055;
or (n7055,s0n7055,s1n7055);
not(notn7055,n5014);
and (s0n7055,notn7055,n7056);
and (s1n7055,n5014,n7053);
and (n7057,n7058,n5033);
wire s0n7058,s1n7058,notn7058;
or (n7058,s0n7058,s1n7058);
not(notn7058,n5014);
and (s0n7058,notn7058,n7059);
and (s1n7058,n5014,n7056);
and (n7060,n7061,n5038);
wire s0n7061,s1n7061,notn7061;
or (n7061,s0n7061,s1n7061);
not(notn7061,n5014);
and (s0n7061,notn7061,n7062);
and (s1n7061,n5014,n7059);
and (n7063,n5395,n2742);
and (n7064,n5410,n2752);
and (n7066,n7032,n7067);
or (n7067,n7068,n7135,n7343);
and (n7068,n7069,n7101);
wire s0n7069,s1n7069,notn7069;
or (n7069,s0n7069,s1n7069);
not(notn7069,n4966);
and (s0n7069,notn7069,n7070);
and (s1n7069,n4966,n7100);
or (n7070,1'b0,n7071,n7072,n7073,n7088);
and (n7071,n5606,n2718);
and (n7072,n5621,n2730);
and (n7073,n7074,n2742);
or (n7074,1'b0,n7075,n7079,n7082,n7085);
and (n7075,n7076,n5016);
wire s0n7076,s1n7076,notn7076;
or (n7076,s0n7076,s1n7076);
not(notn7076,n5014);
and (s0n7076,notn7076,n7077);
and (s1n7076,n5014,n7078);
and (n7079,n7080,n5028);
wire s0n7080,s1n7080,notn7080;
or (n7080,s0n7080,s1n7080);
not(notn7080,n5014);
and (s0n7080,notn7080,n7081);
and (s1n7080,n5014,n7077);
and (n7082,n7083,n5033);
wire s0n7083,s1n7083,notn7083;
or (n7083,s0n7083,s1n7083);
not(notn7083,n5014);
and (s0n7083,notn7083,n7084);
and (s1n7083,n5014,n7081);
and (n7085,n7086,n5038);
wire s0n7086,s1n7086,notn7086;
or (n7086,s0n7086,s1n7086);
not(notn7086,n5014);
and (s0n7086,notn7086,n7087);
and (s1n7086,n5014,n7084);
and (n7088,n7089,n2752);
or (n7089,1'b0,n7090,n7093,n7096,n7098);
and (n7090,n7091,n5016);
wire s0n7091,s1n7091,notn7091;
or (n7091,s0n7091,s1n7091);
not(notn7091,n5014);
and (s0n7091,notn7091,n7092);
and (s1n7091,n5014,n7087);
and (n7093,n7094,n5028);
wire s0n7094,s1n7094,notn7094;
or (n7094,s0n7094,s1n7094);
not(notn7094,n5014);
and (s0n7094,notn7094,n7095);
and (s1n7094,n5014,n7092);
and (n7096,n7097,n5033);
wire s0n7097,s1n7097,notn7097;
or (n7097,s0n7097,s1n7097);
not(notn7097,n5014);
and (s0n7097,notn7097,n2155);
and (s1n7097,n5014,n7095);
and (n7098,n7099,n5038);
wire s0n7099,s1n7099,notn7099;
or (n7099,s0n7099,s1n7099);
not(notn7099,n5014);
and (s0n7099,notn7099,n1773);
and (s1n7099,n5014,n2155);
wire s0n7101,s1n7101,notn7101;
or (n7101,s0n7101,s1n7101);
not(notn7101,n4966);
and (s0n7101,notn7101,n7102);
and (s1n7101,n4966,n7134);
or (n7102,1'b0,n7103,n7118,n7132,n7133);
and (n7103,n7104,n2718);
or (n7104,1'b0,n7105,n7109,n7112,n7115);
and (n7105,n7106,n5016);
wire s0n7106,s1n7106,notn7106;
or (n7106,s0n7106,s1n7106);
not(notn7106,n5014);
and (s0n7106,notn7106,n7107);
and (s1n7106,n5014,n7108);
and (n7109,n7110,n5028);
wire s0n7110,s1n7110,notn7110;
or (n7110,s0n7110,s1n7110);
not(notn7110,n5014);
and (s0n7110,notn7110,n7111);
and (s1n7110,n5014,n7107);
and (n7112,n7113,n5033);
wire s0n7113,s1n7113,notn7113;
or (n7113,s0n7113,s1n7113);
not(notn7113,n5014);
and (s0n7113,notn7113,n7114);
and (s1n7113,n5014,n7111);
and (n7115,n7116,n5038);
wire s0n7116,s1n7116,notn7116;
or (n7116,s0n7116,s1n7116);
not(notn7116,n5014);
and (s0n7116,notn7116,n7117);
and (s1n7116,n5014,n7114);
and (n7118,n7119,n2730);
or (n7119,1'b0,n7120,n7123,n7126,n7129);
and (n7120,n7121,n5016);
wire s0n7121,s1n7121,notn7121;
or (n7121,s0n7121,s1n7121);
not(notn7121,n5014);
and (s0n7121,notn7121,n7122);
and (s1n7121,n5014,n7117);
and (n7123,n7124,n5028);
wire s0n7124,s1n7124,notn7124;
or (n7124,s0n7124,s1n7124);
not(notn7124,n5014);
and (s0n7124,notn7124,n7125);
and (s1n7124,n5014,n7122);
and (n7126,n7127,n5033);
wire s0n7127,s1n7127,notn7127;
or (n7127,s0n7127,s1n7127);
not(notn7127,n5014);
and (s0n7127,notn7127,n7128);
and (s1n7127,n5014,n7125);
and (n7129,n7130,n5038);
wire s0n7130,s1n7130,notn7130;
or (n7130,s0n7130,s1n7130);
not(notn7130,n5014);
and (s0n7130,notn7130,n7131);
and (s1n7130,n5014,n7128);
and (n7132,n5518,n2742);
and (n7133,n5533,n2752);
and (n7135,n7101,n7136);
or (n7136,n7137,n7204,n7342);
and (n7137,n7138,n7170);
wire s0n7138,s1n7138,notn7138;
or (n7138,s0n7138,s1n7138);
not(notn7138,n4966);
and (s0n7138,notn7138,n7139);
and (s1n7138,n4966,n7169);
or (n7139,1'b0,n7140,n7141,n7142,n7157);
and (n7140,n5729,n2718);
and (n7141,n5744,n2730);
and (n7142,n7143,n2742);
or (n7143,1'b0,n7144,n7148,n7151,n7154);
and (n7144,n7145,n5016);
wire s0n7145,s1n7145,notn7145;
or (n7145,s0n7145,s1n7145);
not(notn7145,n5014);
and (s0n7145,notn7145,n7146);
and (s1n7145,n5014,n7147);
and (n7148,n7149,n5028);
wire s0n7149,s1n7149,notn7149;
or (n7149,s0n7149,s1n7149);
not(notn7149,n5014);
and (s0n7149,notn7149,n7150);
and (s1n7149,n5014,n7146);
and (n7151,n7152,n5033);
wire s0n7152,s1n7152,notn7152;
or (n7152,s0n7152,s1n7152);
not(notn7152,n5014);
and (s0n7152,notn7152,n7153);
and (s1n7152,n5014,n7150);
and (n7154,n7155,n5038);
wire s0n7155,s1n7155,notn7155;
or (n7155,s0n7155,s1n7155);
not(notn7155,n5014);
and (s0n7155,notn7155,n7156);
and (s1n7155,n5014,n7153);
and (n7157,n7158,n2752);
or (n7158,1'b0,n7159,n7162,n7165,n7167);
and (n7159,n7160,n5016);
wire s0n7160,s1n7160,notn7160;
or (n7160,s0n7160,s1n7160);
not(notn7160,n5014);
and (s0n7160,notn7160,n7161);
and (s1n7160,n5014,n7156);
and (n7162,n7163,n5028);
wire s0n7163,s1n7163,notn7163;
or (n7163,s0n7163,s1n7163);
not(notn7163,n5014);
and (s0n7163,notn7163,n7164);
and (s1n7163,n5014,n7161);
and (n7165,n7166,n5033);
wire s0n7166,s1n7166,notn7166;
or (n7166,s0n7166,s1n7166);
not(notn7166,n5014);
and (s0n7166,notn7166,n2171);
and (s1n7166,n5014,n7164);
and (n7167,n7168,n5038);
wire s0n7168,s1n7168,notn7168;
or (n7168,s0n7168,s1n7168);
not(notn7168,n5014);
and (s0n7168,notn7168,n1794);
and (s1n7168,n5014,n2171);
wire s0n7170,s1n7170,notn7170;
or (n7170,s0n7170,s1n7170);
not(notn7170,n4966);
and (s0n7170,notn7170,n7171);
and (s1n7170,n4966,n7203);
or (n7171,1'b0,n7172,n7187,n7201,n7202);
and (n7172,n7173,n2718);
or (n7173,1'b0,n7174,n7178,n7181,n7184);
and (n7174,n7175,n5016);
wire s0n7175,s1n7175,notn7175;
or (n7175,s0n7175,s1n7175);
not(notn7175,n5014);
and (s0n7175,notn7175,n7176);
and (s1n7175,n5014,n7177);
and (n7178,n7179,n5028);
wire s0n7179,s1n7179,notn7179;
or (n7179,s0n7179,s1n7179);
not(notn7179,n5014);
and (s0n7179,notn7179,n7180);
and (s1n7179,n5014,n7176);
and (n7181,n7182,n5033);
wire s0n7182,s1n7182,notn7182;
or (n7182,s0n7182,s1n7182);
not(notn7182,n5014);
and (s0n7182,notn7182,n7183);
and (s1n7182,n5014,n7180);
and (n7184,n7185,n5038);
wire s0n7185,s1n7185,notn7185;
or (n7185,s0n7185,s1n7185);
not(notn7185,n5014);
and (s0n7185,notn7185,n7186);
and (s1n7185,n5014,n7183);
and (n7187,n7188,n2730);
or (n7188,1'b0,n7189,n7192,n7195,n7198);
and (n7189,n7190,n5016);
wire s0n7190,s1n7190,notn7190;
or (n7190,s0n7190,s1n7190);
not(notn7190,n5014);
and (s0n7190,notn7190,n7191);
and (s1n7190,n5014,n7186);
and (n7192,n7193,n5028);
wire s0n7193,s1n7193,notn7193;
or (n7193,s0n7193,s1n7193);
not(notn7193,n5014);
and (s0n7193,notn7193,n7194);
and (s1n7193,n5014,n7191);
and (n7195,n7196,n5033);
wire s0n7196,s1n7196,notn7196;
or (n7196,s0n7196,s1n7196);
not(notn7196,n5014);
and (s0n7196,notn7196,n7197);
and (s1n7196,n5014,n7194);
and (n7198,n7199,n5038);
wire s0n7199,s1n7199,notn7199;
or (n7199,s0n7199,s1n7199);
not(notn7199,n5014);
and (s0n7199,notn7199,n7200);
and (s1n7199,n5014,n7197);
and (n7201,n5641,n2742);
and (n7202,n5656,n2752);
and (n7204,n7170,n7205);
or (n7205,n7206,n7273,n7341);
and (n7206,n7207,n7239);
wire s0n7207,s1n7207,notn7207;
or (n7207,s0n7207,s1n7207);
not(notn7207,n4966);
and (s0n7207,notn7207,n7208);
and (s1n7207,n4966,n7238);
or (n7208,1'b0,n7209,n7210,n7211,n7226);
and (n7209,n5852,n2718);
and (n7210,n5867,n2730);
and (n7211,n7212,n2742);
or (n7212,1'b0,n7213,n7217,n7220,n7223);
and (n7213,n7214,n5016);
wire s0n7214,s1n7214,notn7214;
or (n7214,s0n7214,s1n7214);
not(notn7214,n5014);
and (s0n7214,notn7214,n7215);
and (s1n7214,n5014,n7216);
and (n7217,n7218,n5028);
wire s0n7218,s1n7218,notn7218;
or (n7218,s0n7218,s1n7218);
not(notn7218,n5014);
and (s0n7218,notn7218,n7219);
and (s1n7218,n5014,n7215);
and (n7220,n7221,n5033);
wire s0n7221,s1n7221,notn7221;
or (n7221,s0n7221,s1n7221);
not(notn7221,n5014);
and (s0n7221,notn7221,n7222);
and (s1n7221,n5014,n7219);
and (n7223,n7224,n5038);
wire s0n7224,s1n7224,notn7224;
or (n7224,s0n7224,s1n7224);
not(notn7224,n5014);
and (s0n7224,notn7224,n7225);
and (s1n7224,n5014,n7222);
and (n7226,n7227,n2752);
or (n7227,1'b0,n7228,n7231,n7234,n7236);
and (n7228,n7229,n5016);
wire s0n7229,s1n7229,notn7229;
or (n7229,s0n7229,s1n7229);
not(notn7229,n5014);
and (s0n7229,notn7229,n7230);
and (s1n7229,n5014,n7225);
and (n7231,n7232,n5028);
wire s0n7232,s1n7232,notn7232;
or (n7232,s0n7232,s1n7232);
not(notn7232,n5014);
and (s0n7232,notn7232,n7233);
and (s1n7232,n5014,n7230);
and (n7234,n7235,n5033);
wire s0n7235,s1n7235,notn7235;
or (n7235,s0n7235,s1n7235);
not(notn7235,n5014);
and (s0n7235,notn7235,n2188);
and (s1n7235,n5014,n7233);
and (n7236,n7237,n5038);
wire s0n7237,s1n7237,notn7237;
or (n7237,s0n7237,s1n7237);
not(notn7237,n5014);
and (s0n7237,notn7237,n1824);
and (s1n7237,n5014,n2188);
wire s0n7239,s1n7239,notn7239;
or (n7239,s0n7239,s1n7239);
not(notn7239,n4966);
and (s0n7239,notn7239,n7240);
and (s1n7239,n4966,n7272);
or (n7240,1'b0,n7241,n7256,n7270,n7271);
and (n7241,n7242,n2718);
or (n7242,1'b0,n7243,n7247,n7250,n7253);
and (n7243,n7244,n5016);
wire s0n7244,s1n7244,notn7244;
or (n7244,s0n7244,s1n7244);
not(notn7244,n5014);
and (s0n7244,notn7244,n7245);
and (s1n7244,n5014,n7246);
and (n7247,n7248,n5028);
wire s0n7248,s1n7248,notn7248;
or (n7248,s0n7248,s1n7248);
not(notn7248,n5014);
and (s0n7248,notn7248,n7249);
and (s1n7248,n5014,n7245);
and (n7250,n7251,n5033);
wire s0n7251,s1n7251,notn7251;
or (n7251,s0n7251,s1n7251);
not(notn7251,n5014);
and (s0n7251,notn7251,n7252);
and (s1n7251,n5014,n7249);
and (n7253,n7254,n5038);
wire s0n7254,s1n7254,notn7254;
or (n7254,s0n7254,s1n7254);
not(notn7254,n5014);
and (s0n7254,notn7254,n7255);
and (s1n7254,n5014,n7252);
and (n7256,n7257,n2730);
or (n7257,1'b0,n7258,n7261,n7264,n7267);
and (n7258,n7259,n5016);
wire s0n7259,s1n7259,notn7259;
or (n7259,s0n7259,s1n7259);
not(notn7259,n5014);
and (s0n7259,notn7259,n7260);
and (s1n7259,n5014,n7255);
and (n7261,n7262,n5028);
wire s0n7262,s1n7262,notn7262;
or (n7262,s0n7262,s1n7262);
not(notn7262,n5014);
and (s0n7262,notn7262,n7263);
and (s1n7262,n5014,n7260);
and (n7264,n7265,n5033);
wire s0n7265,s1n7265,notn7265;
or (n7265,s0n7265,s1n7265);
not(notn7265,n5014);
and (s0n7265,notn7265,n7266);
and (s1n7265,n5014,n7263);
and (n7267,n7268,n5038);
wire s0n7268,s1n7268,notn7268;
or (n7268,s0n7268,s1n7268);
not(notn7268,n5014);
and (s0n7268,notn7268,n7269);
and (s1n7268,n5014,n7266);
and (n7270,n5764,n2742);
and (n7271,n5779,n2752);
and (n7273,n7239,n7274);
and (n7274,n7275,n7307);
wire s0n7275,s1n7275,notn7275;
or (n7275,s0n7275,s1n7275);
not(notn7275,n4966);
and (s0n7275,notn7275,n7276);
and (s1n7275,n4966,n7306);
or (n7276,1'b0,n7277,n7278,n7279,n7294);
and (n7277,n5974,n2718);
and (n7278,n5989,n2730);
and (n7279,n7280,n2742);
or (n7280,1'b0,n7281,n7285,n7288,n7291);
and (n7281,n7282,n5016);
wire s0n7282,s1n7282,notn7282;
or (n7282,s0n7282,s1n7282);
not(notn7282,n5014);
and (s0n7282,notn7282,n7283);
and (s1n7282,n5014,n7284);
and (n7285,n7286,n5028);
wire s0n7286,s1n7286,notn7286;
or (n7286,s0n7286,s1n7286);
not(notn7286,n5014);
and (s0n7286,notn7286,n7287);
and (s1n7286,n5014,n7283);
and (n7288,n7289,n5033);
wire s0n7289,s1n7289,notn7289;
or (n7289,s0n7289,s1n7289);
not(notn7289,n5014);
and (s0n7289,notn7289,n7290);
and (s1n7289,n5014,n7287);
and (n7291,n7292,n5038);
wire s0n7292,s1n7292,notn7292;
or (n7292,s0n7292,s1n7292);
not(notn7292,n5014);
and (s0n7292,notn7292,n7293);
and (s1n7292,n5014,n7290);
and (n7294,n7295,n2752);
or (n7295,1'b0,n7296,n7299,n7302,n7304);
and (n7296,n7297,n5016);
wire s0n7297,s1n7297,notn7297;
or (n7297,s0n7297,s1n7297);
not(notn7297,n5014);
and (s0n7297,notn7297,n7298);
and (s1n7297,n5014,n7293);
and (n7299,n7300,n5028);
wire s0n7300,s1n7300,notn7300;
or (n7300,s0n7300,s1n7300);
not(notn7300,n5014);
and (s0n7300,notn7300,n7301);
and (s1n7300,n5014,n7298);
and (n7302,n7303,n5033);
wire s0n7303,s1n7303,notn7303;
or (n7303,s0n7303,s1n7303);
not(notn7303,n5014);
and (s0n7303,notn7303,n2203);
and (s1n7303,n5014,n7301);
and (n7304,n7305,n5038);
wire s0n7305,s1n7305,notn7305;
or (n7305,s0n7305,s1n7305);
not(notn7305,n5014);
and (s0n7305,notn7305,n1847);
and (s1n7305,n5014,n2203);
wire s0n7307,s1n7307,notn7307;
or (n7307,s0n7307,s1n7307);
not(notn7307,n4966);
and (s0n7307,notn7307,n7308);
and (s1n7307,n4966,n7340);
or (n7308,1'b0,n7309,n7324,n7338,n7339);
and (n7309,n7310,n2718);
or (n7310,1'b0,n7311,n7315,n7318,n7321);
and (n7311,n7312,n5016);
wire s0n7312,s1n7312,notn7312;
or (n7312,s0n7312,s1n7312);
not(notn7312,n5014);
and (s0n7312,notn7312,n7313);
and (s1n7312,n5014,n7314);
and (n7315,n7316,n5028);
wire s0n7316,s1n7316,notn7316;
or (n7316,s0n7316,s1n7316);
not(notn7316,n5014);
and (s0n7316,notn7316,n7317);
and (s1n7316,n5014,n7313);
and (n7318,n7319,n5033);
wire s0n7319,s1n7319,notn7319;
or (n7319,s0n7319,s1n7319);
not(notn7319,n5014);
and (s0n7319,notn7319,n7320);
and (s1n7319,n5014,n7317);
and (n7321,n7322,n5038);
wire s0n7322,s1n7322,notn7322;
or (n7322,s0n7322,s1n7322);
not(notn7322,n5014);
and (s0n7322,notn7322,n7323);
and (s1n7322,n5014,n7320);
and (n7324,n7325,n2730);
or (n7325,1'b0,n7326,n7329,n7332,n7335);
and (n7326,n7327,n5016);
wire s0n7327,s1n7327,notn7327;
or (n7327,s0n7327,s1n7327);
not(notn7327,n5014);
and (s0n7327,notn7327,n7328);
and (s1n7327,n5014,n7323);
and (n7329,n7330,n5028);
wire s0n7330,s1n7330,notn7330;
or (n7330,s0n7330,s1n7330);
not(notn7330,n5014);
and (s0n7330,notn7330,n7331);
and (s1n7330,n5014,n7328);
and (n7332,n7333,n5033);
wire s0n7333,s1n7333,notn7333;
or (n7333,s0n7333,s1n7333);
not(notn7333,n5014);
and (s0n7333,notn7333,n7334);
and (s1n7333,n5014,n7331);
and (n7335,n7336,n5038);
wire s0n7336,s1n7336,notn7336;
or (n7336,s0n7336,s1n7336);
not(notn7336,n5014);
and (s0n7336,notn7336,n7337);
and (s1n7336,n5014,n7334);
and (n7338,n5886,n2742);
and (n7339,n5901,n2752);
and (n7341,n7207,n7274);
and (n7342,n7138,n7205);
and (n7343,n7069,n7136);
and (n7344,n7000,n7067);
and (n7345,n6931,n6998);
and (n7346,n6862,n6929);
and (n7347,n6793,n6860);
and (n7348,n6786,n6791);
and (n7349,n6779,n6784);
and (n7350,n6772,n6777);
and (n7351,n6765,n6770);
or (n7352,n7353,n7359,n7437);
and (n7353,n7354,n7356);
xor (n7354,n7355,n6030);
xor (n7355,n6025,n6027);
not (n7356,n7357);
xor (n7357,n7358,n6770);
xor (n7358,n6765,n6767);
and (n7359,n7356,n7360);
or (n7360,n7361,n7367,n7436);
and (n7361,n7362,n7364);
xor (n7362,n7363,n6037);
xor (n7363,n6032,n6034);
not (n7364,n7365);
xor (n7365,n7366,n6777);
xor (n7366,n6772,n6774);
and (n7367,n7364,n7368);
or (n7368,n7369,n7375,n7435);
and (n7369,n7370,n7372);
xor (n7370,n7371,n6126);
xor (n7371,n6039,n6082);
not (n7372,n7373);
xor (n7373,n7374,n6784);
xor (n7374,n6779,n6781);
and (n7375,n7372,n7376);
or (n7376,n7377,n7383,n7434);
and (n7377,n7378,n7380);
xor (n7378,n7379,n6215);
xor (n7379,n6128,n6171);
not (n7380,n7381);
xor (n7381,n7382,n6791);
xor (n7382,n6786,n6788);
and (n7383,n7380,n7384);
or (n7384,n7385,n7391,n7433);
and (n7385,n7386,n7388);
xor (n7386,n7387,n6304);
xor (n7387,n6217,n6260);
not (n7388,n7389);
xor (n7389,n7390,n6860);
xor (n7390,n6793,n6825);
and (n7391,n7388,n7392);
or (n7392,n7393,n7399,n7432);
and (n7393,n7394,n7396);
xor (n7394,n7395,n6393);
xor (n7395,n6306,n6349);
not (n7396,n7397);
xor (n7397,n7398,n6929);
xor (n7398,n6862,n6894);
and (n7399,n7396,n7400);
or (n7400,n7401,n7407,n7431);
and (n7401,n7402,n7404);
xor (n7402,n7403,n6482);
xor (n7403,n6395,n6438);
not (n7404,n7405);
xor (n7405,n7406,n6998);
xor (n7406,n6931,n6963);
and (n7407,n7404,n7408);
or (n7408,n7409,n7415,n7430);
and (n7409,n7410,n7412);
xor (n7410,n7411,n6571);
xor (n7411,n6484,n6527);
not (n7412,n7413);
xor (n7413,n7414,n7067);
xor (n7414,n7000,n7032);
and (n7415,n7412,n7416);
or (n7416,n7417,n7423,n7429);
and (n7417,n7418,n7420);
xor (n7418,n7419,n6660);
xor (n7419,n6573,n6616);
not (n7420,n7421);
xor (n7421,n7422,n7136);
xor (n7422,n7069,n7101);
and (n7423,n7420,n7424);
and (n7424,n7425,n7426);
xor (n7425,n6661,n6704);
not (n7426,n7427);
xor (n7427,n7428,n7205);
xor (n7428,n7138,n7170);
and (n7429,n7418,n7424);
and (n7430,n7410,n7416);
and (n7431,n7402,n7408);
and (n7432,n7394,n7400);
and (n7433,n7386,n7392);
and (n7434,n7378,n7384);
and (n7435,n7370,n7376);
and (n7436,n7362,n7368);
and (n7437,n7354,n7360);
and (n7438,n7439,n7441);
xor (n7439,n7440,n7360);
xor (n7440,n7354,n7356);
and (n7441,n7442,n7444);
xor (n7442,n7443,n7368);
xor (n7443,n7362,n7364);
and (n7444,n7445,n7447);
xor (n7445,n7446,n7376);
xor (n7446,n7370,n7372);
and (n7447,n7448,n7450);
xor (n7448,n7449,n7384);
xor (n7449,n7378,n7380);
and (n7450,n7451,n7453);
xor (n7451,n7452,n7392);
xor (n7452,n7386,n7388);
and (n7453,n7454,n7456);
xor (n7454,n7455,n7400);
xor (n7455,n7394,n7396);
and (n7456,n7457,n7459);
xor (n7457,n7458,n7408);
xor (n7458,n7402,n7404);
and (n7459,n7460,n7462);
xor (n7460,n7461,n7416);
xor (n7461,n7410,n7412);
and (n7462,n7463,n7465);
xor (n7463,n7464,n7424);
xor (n7464,n7418,n7420);
and (n7465,n7466,n7467);
xor (n7466,n7425,n7426);
and (n7467,n7468,n7471);
not (n7468,n7469);
xor (n7469,n7470,n7274);
xor (n7470,n7207,n7239);
not (n7471,n7472);
xor (n7472,n7275,n7307);
or (n7473,n7474,n7478,n7551);
and (n7474,n7475,n7477);
xor (n7475,n7476,n4983);
xor (n7476,n4978,n4980);
xor (n7477,n7439,n7441);
and (n7478,n7477,n7479);
or (n7479,n7480,n7484,n7550);
and (n7480,n7481,n7483);
xor (n7481,n7482,n4990);
xor (n7482,n4985,n4987);
xor (n7483,n7442,n7444);
and (n7484,n7483,n7485);
or (n7485,n7486,n7490,n7549);
and (n7486,n7487,n7489);
xor (n7487,n7488,n4997);
xor (n7488,n4992,n4994);
xor (n7489,n7445,n7447);
and (n7490,n7489,n7491);
or (n7491,n7492,n7496,n7548);
and (n7492,n7493,n7495);
xor (n7493,n7494,n5004);
xor (n7494,n4999,n5001);
xor (n7495,n7448,n7450);
and (n7496,n7495,n7497);
or (n7497,n7498,n7502,n7547);
and (n7498,n7499,n7501);
xor (n7499,n7500,n5144);
xor (n7500,n5006,n5082);
xor (n7501,n7451,n7453);
and (n7502,n7501,n7503);
or (n7503,n7504,n7508,n7546);
and (n7504,n7505,n7507);
xor (n7505,n7506,n5267);
xor (n7506,n5146,n5205);
xor (n7507,n7454,n7456);
and (n7508,n7507,n7509);
or (n7509,n7510,n7514,n7545);
and (n7510,n7511,n7513);
xor (n7511,n7512,n5390);
xor (n7512,n5269,n5328);
xor (n7513,n7457,n7459);
and (n7514,n7513,n7515);
or (n7515,n7516,n7520,n7544);
and (n7516,n7517,n7519);
xor (n7517,n7518,n5513);
xor (n7518,n5392,n5451);
xor (n7519,n7460,n7462);
and (n7520,n7519,n7521);
or (n7521,n7522,n7526,n7543);
and (n7522,n7523,n7525);
xor (n7523,n7524,n5636);
xor (n7524,n5515,n5574);
xor (n7525,n7463,n7465);
and (n7526,n7525,n7527);
or (n7527,n7528,n7532,n7542);
and (n7528,n7529,n7531);
xor (n7529,n7530,n5759);
xor (n7530,n5638,n5697);
xor (n7531,n7466,n7467);
and (n7532,n7531,n7533);
or (n7533,n7534,n7538,n7541);
and (n7534,n7535,n7537);
xor (n7535,n7536,n5882);
xor (n7536,n5761,n5820);
xor (n7537,n7468,n7471);
and (n7538,n7537,n7539);
and (n7539,n7540,n7472);
xor (n7540,n5883,n5942);
and (n7541,n7535,n7539);
and (n7542,n7529,n7533);
and (n7543,n7523,n7527);
and (n7544,n7517,n7521);
and (n7545,n7511,n7515);
and (n7546,n7505,n7509);
and (n7547,n7499,n7503);
and (n7548,n7493,n7497);
and (n7549,n7487,n7491);
and (n7550,n7481,n7485);
and (n7551,n7475,n7479);
or (n7552,n7553,n7556,n7608);
and (n7553,n7554,n7489);
xor (n7554,n7555,n7479);
xor (n7555,n7475,n7477);
and (n7556,n7489,n7557);
or (n7557,n7558,n7561,n7607);
and (n7558,n7559,n7495);
xor (n7559,n7560,n7485);
xor (n7560,n7481,n7483);
and (n7561,n7495,n7562);
or (n7562,n7563,n7566,n7606);
and (n7563,n7564,n7501);
xor (n7564,n7565,n7491);
xor (n7565,n7487,n7489);
and (n7566,n7501,n7567);
or (n7567,n7568,n7571,n7605);
and (n7568,n7569,n7507);
xor (n7569,n7570,n7497);
xor (n7570,n7493,n7495);
and (n7571,n7507,n7572);
or (n7572,n7573,n7576,n7604);
and (n7573,n7574,n7513);
xor (n7574,n7575,n7503);
xor (n7575,n7499,n7501);
and (n7576,n7513,n7577);
or (n7577,n7578,n7581,n7603);
and (n7578,n7579,n7519);
xor (n7579,n7580,n7509);
xor (n7580,n7505,n7507);
and (n7581,n7519,n7582);
or (n7582,n7583,n7586,n7602);
and (n7583,n7584,n7525);
xor (n7584,n7585,n7515);
xor (n7585,n7511,n7513);
and (n7586,n7525,n7587);
or (n7587,n7588,n7591,n7601);
and (n7588,n7589,n7531);
xor (n7589,n7590,n7521);
xor (n7590,n7517,n7519);
and (n7591,n7531,n7592);
or (n7592,n7593,n7596,n7600);
and (n7593,n7594,n7537);
xor (n7594,n7595,n7527);
xor (n7595,n7523,n7525);
and (n7596,n7537,n7597);
and (n7597,n7598,n7472);
xor (n7598,n7599,n7533);
xor (n7599,n7529,n7531);
and (n7600,n7594,n7597);
and (n7601,n7589,n7592);
and (n7602,n7584,n7587);
and (n7603,n7579,n7582);
and (n7604,n7574,n7577);
and (n7605,n7569,n7572);
and (n7606,n7564,n7567);
and (n7607,n7559,n7562);
and (n7608,n7554,n7557);
and (n7609,n7610,n7612);
xor (n7610,n7611,n7557);
xor (n7611,n7554,n7489);
and (n7612,n7613,n7615);
xor (n7613,n7614,n7562);
xor (n7614,n7559,n7495);
and (n7615,n7616,n7618);
xor (n7616,n7617,n7567);
xor (n7617,n7564,n7501);
and (n7618,n7619,n7621);
xor (n7619,n7620,n7572);
xor (n7620,n7569,n7507);
and (n7621,n7622,n7624);
xor (n7622,n7623,n7577);
xor (n7623,n7574,n7513);
and (n7624,n7625,n7627);
xor (n7625,n7626,n7582);
xor (n7626,n7579,n7519);
and (n7627,n7628,n7630);
xor (n7628,n7629,n7587);
xor (n7629,n7584,n7525);
xor (n7630,n7631,n7592);
xor (n7631,n7589,n7531);
xor (n7632,n4958,n7633);
and (n7633,n7610,n7634);
and (n7634,n7613,n7616);
wire s0n7635,s1n7635,notn7635;
or (n7635,s0n7635,s1n7635);
not(notn7635,n4966);
and (s0n7635,notn7635,n7636);
and (s1n7635,n4966,n7840);
xor (n7636,n7637,n7827);
xor (n7637,n7638,n7799);
xor (n7638,n7639,n7778);
xor (n7639,n7640,n7772);
xor (n7640,n7641,n7663);
xor (n7641,n7642,n7647);
xor (n7642,n7643,n7645);
wire s0n7643,s1n7643,notn7643;
or (n7643,s0n7643,s1n7643);
not(notn7643,n4966);
and (s0n7643,notn7643,1'b0);
and (s1n7643,n4966,n7644);
wire s0n7645,s1n7645,notn7645;
or (n7645,s0n7645,s1n7645);
not(notn7645,n4966);
and (s0n7645,notn7645,1'b0);
and (s1n7645,n4966,n7646);
or (n7647,n7648,n7649,n7662);
and (n7648,n7643,n7645);
and (n7649,n7645,n7650);
or (n7650,n7651,n7656,n7661);
and (n7651,n7652,n7654);
wire s0n7652,s1n7652,notn7652;
or (n7652,s0n7652,s1n7652);
not(notn7652,n4966);
and (s0n7652,notn7652,1'b0);
and (s1n7652,n4966,n7653);
wire s0n7654,s1n7654,notn7654;
or (n7654,s0n7654,s1n7654);
not(notn7654,n4966);
and (s0n7654,notn7654,1'b0);
and (s1n7654,n4966,n7655);
and (n7656,n7654,n7657);
or (n7657,n7658,n7659,n7660);
and (n7658,n4964,n4974);
and (n7659,n4974,n4976);
and (n7660,n4964,n4976);
and (n7661,n7652,n7657);
and (n7662,n7643,n7650);
xor (n7663,n7664,n7759);
xor (n7664,n7665,n7727);
xor (n7665,n7666,n7704);
xor (n7666,n7667,n7672);
xor (n7667,n7668,n7670);
wire s0n7668,s1n7668,notn7668;
or (n7668,s0n7668,s1n7668);
not(notn7668,n4966);
and (s0n7668,notn7668,1'b0);
and (s1n7668,n4966,n7669);
wire s0n7670,s1n7670,notn7670;
or (n7670,s0n7670,s1n7670);
not(notn7670,n4966);
and (s0n7670,notn7670,1'b0);
and (s1n7670,n4966,n7671);
or (n7672,n7673,n7674,n7703);
and (n7673,n7668,n7670);
and (n7674,n7670,n7675);
or (n7675,n7676,n7681,n7702);
and (n7676,n7677,n7679);
wire s0n7677,s1n7677,notn7677;
or (n7677,s0n7677,s1n7677);
not(notn7677,n4966);
and (s0n7677,notn7677,1'b0);
and (s1n7677,n4966,n7678);
wire s0n7679,s1n7679,notn7679;
or (n7679,s0n7679,s1n7679);
not(notn7679,n4966);
and (s0n7679,notn7679,1'b0);
and (s1n7679,n4966,n7680);
and (n7681,n7679,n7682);
or (n7682,n7683,n7688,n7701);
and (n7683,n7684,n7686);
wire s0n7684,s1n7684,notn7684;
or (n7684,s0n7684,s1n7684);
not(notn7684,n4966);
and (s0n7684,notn7684,1'b0);
and (s1n7684,n4966,n7685);
wire s0n7686,s1n7686,notn7686;
or (n7686,s0n7686,s1n7686);
not(notn7686,n4966);
and (s0n7686,notn7686,1'b0);
and (s1n7686,n4966,n7687);
and (n7688,n7686,n7689);
or (n7689,n7690,n7695,n7700);
and (n7690,n7691,n7693);
wire s0n7691,s1n7691,notn7691;
or (n7691,s0n7691,s1n7691);
not(notn7691,n4966);
and (s0n7691,notn7691,1'b0);
and (s1n7691,n4966,n7692);
wire s0n7693,s1n7693,notn7693;
or (n7693,s0n7693,s1n7693);
not(notn7693,n4966);
and (s0n7693,notn7693,1'b0);
and (s1n7693,n4966,n7694);
and (n7695,n7693,n7696);
or (n7696,n7697,n7698,n7699);
and (n7697,n6019,n6021);
and (n7698,n6021,n6023);
and (n7699,n6019,n6023);
and (n7700,n7691,n7696);
and (n7701,n7684,n7689);
and (n7702,n7677,n7682);
and (n7703,n7668,n7675);
not (n7704,n7705);
xor (n7705,n7706,n7711);
xor (n7706,n7707,n7709);
wire s0n7707,s1n7707,notn7707;
or (n7707,s0n7707,s1n7707);
not(notn7707,n4966);
and (s0n7707,notn7707,1'b0);
and (s1n7707,n4966,n7708);
wire s0n7709,s1n7709,notn7709;
or (n7709,s0n7709,s1n7709);
not(notn7709,n4966);
and (s0n7709,notn7709,1'b0);
and (s1n7709,n4966,n7710);
or (n7711,n7712,n7713,n7726);
and (n7712,n7707,n7709);
and (n7713,n7709,n7714);
or (n7714,n7715,n7720,n7725);
and (n7715,n7716,n7718);
wire s0n7716,s1n7716,notn7716;
or (n7716,s0n7716,s1n7716);
not(notn7716,n4966);
and (s0n7716,notn7716,1'b0);
and (s1n7716,n4966,n7717);
wire s0n7718,s1n7718,notn7718;
or (n7718,s0n7718,s1n7718);
not(notn7718,n4966);
and (s0n7718,notn7718,1'b0);
and (s1n7718,n4966,n7719);
and (n7720,n7718,n7721);
or (n7721,n7722,n7723,n7724);
and (n7722,n6759,n6761);
and (n7723,n6761,n6763);
and (n7724,n6759,n6763);
and (n7725,n7716,n7721);
and (n7726,n7707,n7714);
or (n7727,n7728,n7730,n7758);
and (n7728,n7729,n7704);
xor (n7729,n7667,n7675);
and (n7730,n7704,n7731);
or (n7731,n7732,n7735,n7757);
and (n7732,n7733,n7704);
xor (n7733,n7734,n7682);
xor (n7734,n7677,n7679);
and (n7735,n7704,n7736);
or (n7736,n7737,n7742,n7756);
and (n7737,n7738,n7740);
xor (n7738,n7739,n7689);
xor (n7739,n7684,n7686);
not (n7740,n7741);
xor (n7741,n7706,n7714);
and (n7742,n7740,n7743);
or (n7743,n7744,n7750,n7755);
and (n7744,n7745,n7747);
xor (n7745,n7746,n7696);
xor (n7746,n7691,n7693);
not (n7747,n7748);
xor (n7748,n7749,n7721);
xor (n7749,n7716,n7718);
and (n7750,n7747,n7751);
or (n7751,n7752,n7753,n7754);
and (n7752,n6017,n6756);
and (n7753,n6756,n7352);
and (n7754,n6017,n7352);
and (n7755,n7745,n7751);
and (n7756,n7738,n7743);
and (n7757,n7733,n7736);
and (n7758,n7729,n7731);
and (n7759,n7760,n7762);
xor (n7760,n7761,n7731);
xor (n7761,n7729,n7704);
and (n7762,n7763,n7765);
xor (n7763,n7764,n7736);
xor (n7764,n7733,n7704);
and (n7765,n7766,n7768);
xor (n7766,n7767,n7743);
xor (n7767,n7738,n7740);
and (n7768,n7769,n7771);
xor (n7769,n7770,n7751);
xor (n7770,n7745,n7747);
and (n7771,n6015,n7438);
or (n7772,n7773,n7775,n7798);
and (n7773,n7641,n7774);
xor (n7774,n7760,n7762);
and (n7775,n7774,n7776);
or (n7776,n7777,n7779,n7797);
and (n7777,n7641,n7778);
xor (n7778,n7763,n7765);
and (n7779,n7778,n7780);
or (n7780,n7781,n7784,n7796);
and (n7781,n7782,n7783);
xor (n7782,n7642,n7650);
xor (n7783,n7766,n7768);
and (n7784,n7783,n7785);
or (n7785,n7786,n7790,n7795);
and (n7786,n7787,n7789);
xor (n7787,n7788,n7657);
xor (n7788,n7652,n7654);
xor (n7789,n7769,n7771);
and (n7790,n7789,n7791);
or (n7791,n7792,n7793,n7794);
and (n7792,n4962,n6014);
and (n7793,n6014,n7473);
and (n7794,n4962,n7473);
and (n7795,n7787,n7791);
and (n7796,n7782,n7785);
and (n7797,n7641,n7780);
and (n7798,n7641,n7776);
or (n7799,n7800,n7803,n7826);
and (n7800,n7801,n7783);
xor (n7801,n7802,n7776);
xor (n7802,n7641,n7774);
and (n7803,n7783,n7804);
or (n7804,n7805,n7808,n7825);
and (n7805,n7806,n7789);
xor (n7806,n7807,n7780);
xor (n7807,n7641,n7778);
and (n7808,n7789,n7809);
or (n7809,n7810,n7813,n7824);
and (n7810,n7811,n6014);
xor (n7811,n7812,n7785);
xor (n7812,n7782,n7783);
and (n7813,n6014,n7814);
or (n7814,n7815,n7818,n7823);
and (n7815,n7816,n7477);
xor (n7816,n7817,n7791);
xor (n7817,n7787,n7789);
and (n7818,n7477,n7819);
or (n7819,n7820,n7821,n7822);
and (n7820,n4960,n7483);
and (n7821,n7483,n7552);
and (n7822,n4960,n7552);
and (n7823,n7816,n7819);
and (n7824,n7811,n7814);
and (n7825,n7806,n7809);
and (n7826,n7801,n7804);
and (n7827,n7828,n7830);
xor (n7828,n7829,n7804);
xor (n7829,n7801,n7783);
and (n7830,n7831,n7833);
xor (n7831,n7832,n7809);
xor (n7832,n7806,n7789);
and (n7833,n7834,n7836);
xor (n7834,n7835,n7814);
xor (n7835,n7811,n6014);
and (n7836,n7837,n7839);
xor (n7837,n7838,n7819);
xor (n7838,n7816,n7477);
and (n7839,n4958,n7609);
xor (n7840,n7637,n7841);
and (n7841,n7828,n7842);
and (n7842,n7831,n7843);
and (n7843,n7834,n7844);
and (n7844,n7837,n7845);
and (n7845,n4958,n7633);
wire s0n7846,s1n7846,notn7846;
or (n7846,s0n7846,s1n7846);
not(notn7846,n4966);
and (s0n7846,notn7846,n7847);
and (s1n7846,n4966,n7850);
wire s0n7847,s1n7847,notn7847;
or (n7847,s0n7847,s1n7847);
not(notn7847,n4966);
and (s0n7847,notn7847,n7848);
and (s1n7847,n4966,n7849);
xor (n7848,n7837,n7839);
xor (n7849,n7837,n7845);
wire s0n7850,s1n7850,notn7850;
or (n7850,s0n7850,s1n7850);
not(notn7850,n4966);
and (s0n7850,notn7850,n7851);
and (s1n7850,n4966,n7859);
xor (n7851,n7852,n7858);
xor (n7852,n7853,n7854);
xor (n7853,n7639,n7774);
or (n7854,n7855,n7856,n7857);
and (n7855,n7639,n7778);
and (n7856,n7778,n7799);
and (n7857,n7639,n7799);
and (n7858,n7637,n7827);
xor (n7859,n7852,n7860);
and (n7860,n7637,n7841);
wire s0n7861,s1n7861,notn7861;
or (n7861,s0n7861,s1n7861);
not(notn7861,n4966);
and (s0n7861,notn7861,n7862);
and (s1n7861,n4966,n7870);
xor (n7862,n7863,n7869);
xor (n7863,n7864,n7865);
xor (n7864,n7639,n7663);
or (n7865,n7866,n7867,n7868);
and (n7866,n7639,n7774);
and (n7867,n7774,n7854);
and (n7868,n7639,n7854);
and (n7869,n7852,n7858);
xor (n7870,n7863,n7871);
and (n7871,n7852,n7860);
and (n7872,n7873,n2907);
wire s0n7873,s1n7873,notn7873;
or (n7873,s0n7873,s1n7873);
not(notn7873,n2902);
and (s0n7873,notn7873,1'b0);
and (s1n7873,n2902,n4953);
and (n7874,n4953,n7875);
or (n7875,n7876,n4883);
or (n7876,n4904,n4895);
and (n7877,n2911,n7878);
or (n7878,n2942,n2944);
and (n7879,n4950,n7880);
or (n7880,n7881,n7991,n8651);
and (n7881,n7882,n7975);
or (n7882,1'b0,n7883,n7886,n7889,n7894);
and (n7883,n7884,n2893);
wire s0n7884,s1n7884,notn7884;
or (n7884,s0n7884,s1n7884);
not(notn7884,n2891);
and (s0n7884,notn7884,1'b0);
and (s1n7884,n2891,n7885);
and (n7886,n7887,n2907);
wire s0n7887,s1n7887,notn7887;
or (n7887,s0n7887,s1n7887);
not(notn7887,n2902);
and (s0n7887,notn7887,1'b0);
and (s1n7887,n2902,n7888);
and (n7889,n7890,n4883);
wire s0n7890,s1n7890,notn7890;
or (n7890,s0n7890,s1n7890);
not(notn7890,n4878);
and (s0n7890,notn7890,n7891);
and (s1n7890,n4878,1'b0);
wire s0n7891,s1n7891,notn7891;
or (n7891,s0n7891,s1n7891);
not(notn7891,n4873);
and (s0n7891,notn7891,n7892);
and (s1n7891,n4873,1'b1);
wire s0n7892,s1n7892,notn7892;
or (n7892,s0n7892,s1n7892);
not(notn7892,n4861);
and (s0n7892,notn7892,1'b0);
and (s1n7892,n4861,n7893);
xor (n7893,n4839,n4841);
or (n7894,1'b0,n7895,n7915,n7935,n7955);
and (n7895,n7896,n2718);
or (n7896,1'b0,n7897,n7903,n7909);
and (n7897,n7898,n4895);
or (n7898,1'b0,n7899,n7900,n7901,n7902);
and (n7899,n3058,n556);
and (n7900,n3062,n567);
and (n7901,n3066,n571);
and (n7902,n3070,n573);
and (n7903,n7904,n2944);
or (n7904,1'b0,n7905,n7906,n7907,n7908);
and (n7905,n3126,n556);
and (n7906,n3057,n567);
and (n7907,n3061,n571);
and (n7908,n3065,n573);
and (n7909,n7910,n4903);
or (n7910,1'b0,n7911,n7912,n7913,n7914);
and (n7911,n3057,n556);
and (n7912,n3061,n567);
and (n7913,n3065,n571);
and (n7914,n3069,n573);
and (n7915,n7916,n2730);
or (n7916,1'b0,n7917,n7923,n7929);
and (n7917,n7918,n4895);
or (n7918,1'b0,n7919,n7920,n7921,n7922);
and (n7919,n3076,n556);
and (n7920,n3080,n567);
and (n7921,n3084,n571);
and (n7922,n3088,n573);
and (n7923,n7924,n2944);
or (n7924,1'b0,n7925,n7926,n7927,n7928);
and (n7925,n3069,n556);
and (n7926,n3075,n567);
and (n7927,n3079,n571);
and (n7928,n3083,n573);
and (n7929,n7930,n4903);
or (n7930,1'b0,n7931,n7932,n7933,n7934);
and (n7931,n3075,n556);
and (n7932,n3079,n567);
and (n7933,n3083,n571);
and (n7934,n3087,n573);
and (n7935,n7936,n2742);
or (n7936,1'b0,n7937,n7943,n7949);
and (n7937,n7938,n4895);
or (n7938,1'b0,n7939,n7940,n7941,n7942);
and (n7939,n3094,n556);
and (n7940,n3098,n567);
and (n7941,n3102,n571);
and (n7942,n3106,n573);
and (n7943,n7944,n2944);
or (n7944,1'b0,n7945,n7946,n7947,n7948);
and (n7945,n3141,n556);
and (n7946,n3093,n567);
and (n7947,n3097,n571);
and (n7948,n3101,n573);
and (n7949,n7950,n4903);
or (n7950,1'b0,n7951,n7952,n7953,n7954);
and (n7951,n3093,n556);
and (n7952,n3097,n567);
and (n7953,n3101,n571);
and (n7954,n3105,n573);
and (n7955,n7956,n2752);
or (n7956,1'b0,n7957,n7963,n7969);
and (n7957,n7958,n4895);
or (n7958,1'b0,n7959,n7960,n7961,n7962);
and (n7959,n3112,n556);
and (n7960,n3116,n567);
and (n7961,n2103,n571);
and (n7962,n1708,n573);
and (n7963,n7964,n2944);
or (n7964,1'b0,n7965,n7966,n7967,n7968);
and (n7965,n3105,n556);
and (n7966,n3111,n567);
and (n7967,n3115,n571);
and (n7968,n1267,n573);
and (n7969,n7970,n4903);
or (n7970,1'b0,n7971,n7972,n7973,n7974);
and (n7971,n3111,n556);
and (n7972,n3115,n567);
and (n7973,n1267,n571);
and (n7974,n755,n573);
or (n7975,1'b0,n7976,n7987,n7989,n7990);
and (n7976,n7977,n2893);
wire s0n7977,s1n7977,notn7977;
or (n7977,s0n7977,s1n7977);
not(notn7977,n2891);
and (s0n7977,notn7977,1'b0);
and (s1n7977,n2891,n7978);
wire s0n7978,s1n7978,notn7978;
or (n7978,s0n7978,s1n7978);
not(notn7978,n7861);
and (s0n7978,notn7978,n7979);
and (s1n7978,n7861,1'b0);
wire s0n7979,s1n7979,notn7979;
or (n7979,s0n7979,s1n7979);
not(notn7979,n7846);
and (s0n7979,notn7979,n7980);
and (s1n7979,n7846,1'b1);
wire s0n7980,s1n7980,notn7980;
or (n7980,s0n7980,s1n7980);
not(notn7980,n4966);
and (s0n7980,notn7980,n7981);
and (s1n7980,n4966,n7984);
wire s0n7981,s1n7981,notn7981;
or (n7981,s0n7981,s1n7981);
not(notn7981,n4966);
and (s0n7981,notn7981,n7982);
and (s1n7981,n4966,n7983);
xor (n7982,n7610,n7612);
xor (n7983,n7610,n7634);
wire s0n7984,s1n7984,notn7984;
or (n7984,s0n7984,s1n7984);
not(notn7984,n4966);
and (s0n7984,notn7984,n7985);
and (s1n7984,n4966,n7986);
xor (n7985,n7828,n7830);
xor (n7986,n7828,n7842);
and (n7987,n7988,n2907);
wire s0n7988,s1n7988,notn7988;
or (n7988,s0n7988,s1n7988);
not(notn7988,n2902);
and (s0n7988,notn7988,1'b0);
and (s1n7988,n2902,n7978);
and (n7989,n7978,n7875);
and (n7990,n7890,n7878);
and (n7991,n7975,n7992);
or (n7992,n7993,n8103,n8650);
and (n7993,n7994,n8087);
or (n7994,1'b0,n7995,n7998,n8001,n8006);
and (n7995,n7996,n2893);
wire s0n7996,s1n7996,notn7996;
or (n7996,s0n7996,s1n7996);
not(notn7996,n2891);
and (s0n7996,notn7996,1'b0);
and (s1n7996,n2891,n7997);
and (n7998,n7999,n2907);
wire s0n7999,s1n7999,notn7999;
or (n7999,s0n7999,s1n7999);
not(notn7999,n2902);
and (s0n7999,notn7999,1'b0);
and (s1n7999,n2902,n8000);
and (n8001,n8002,n4883);
wire s0n8002,s1n8002,notn8002;
or (n8002,s0n8002,s1n8002);
not(notn8002,n4878);
and (s0n8002,notn8002,n8003);
and (s1n8002,n4878,1'b0);
wire s0n8003,s1n8003,notn8003;
or (n8003,s0n8003,s1n8003);
not(notn8003,n4873);
and (s0n8003,notn8003,n8004);
and (s1n8003,n4873,1'b1);
wire s0n8004,s1n8004,notn8004;
or (n8004,s0n8004,s1n8004);
not(notn8004,n4861);
and (s0n8004,notn8004,1'b0);
and (s1n8004,n4861,n8005);
xor (n8005,n4842,n4844);
or (n8006,1'b0,n8007,n8027,n8047,n8067);
and (n8007,n8008,n2718);
or (n8008,1'b0,n8009,n8015,n8021);
and (n8009,n8010,n4895);
or (n8010,1'b0,n8011,n8012,n8013,n8014);
and (n8011,n3161,n556);
and (n8012,n3165,n567);
and (n8013,n3169,n571);
and (n8014,n3173,n573);
and (n8015,n8016,n2944);
or (n8016,1'b0,n8017,n8018,n8019,n8020);
and (n8017,n3229,n556);
and (n8018,n3160,n567);
and (n8019,n3164,n571);
and (n8020,n3168,n573);
and (n8021,n8022,n4903);
or (n8022,1'b0,n8023,n8024,n8025,n8026);
and (n8023,n3160,n556);
and (n8024,n3164,n567);
and (n8025,n3168,n571);
and (n8026,n3172,n573);
and (n8027,n8028,n2730);
or (n8028,1'b0,n8029,n8035,n8041);
and (n8029,n8030,n4895);
or (n8030,1'b0,n8031,n8032,n8033,n8034);
and (n8031,n3179,n556);
and (n8032,n3183,n567);
and (n8033,n3187,n571);
and (n8034,n3191,n573);
and (n8035,n8036,n2944);
or (n8036,1'b0,n8037,n8038,n8039,n8040);
and (n8037,n3172,n556);
and (n8038,n3178,n567);
and (n8039,n3182,n571);
and (n8040,n3186,n573);
and (n8041,n8042,n4903);
or (n8042,1'b0,n8043,n8044,n8045,n8046);
and (n8043,n3178,n556);
and (n8044,n3182,n567);
and (n8045,n3186,n571);
and (n8046,n3190,n573);
and (n8047,n8048,n2742);
or (n8048,1'b0,n8049,n8055,n8061);
and (n8049,n8050,n4895);
or (n8050,1'b0,n8051,n8052,n8053,n8054);
and (n8051,n3197,n556);
and (n8052,n3201,n567);
and (n8053,n3205,n571);
and (n8054,n3209,n573);
and (n8055,n8056,n2944);
or (n8056,1'b0,n8057,n8058,n8059,n8060);
and (n8057,n3244,n556);
and (n8058,n3196,n567);
and (n8059,n3200,n571);
and (n8060,n3204,n573);
and (n8061,n8062,n4903);
or (n8062,1'b0,n8063,n8064,n8065,n8066);
and (n8063,n3196,n556);
and (n8064,n3200,n567);
and (n8065,n3204,n571);
and (n8066,n3208,n573);
and (n8067,n8068,n2752);
or (n8068,1'b0,n8069,n8075,n8081);
and (n8069,n8070,n4895);
or (n8070,1'b0,n8071,n8072,n8073,n8074);
and (n8071,n3215,n556);
and (n8072,n3219,n567);
and (n8073,n2119,n571);
and (n8074,n1727,n573);
and (n8075,n8076,n2944);
or (n8076,1'b0,n8077,n8078,n8079,n8080);
and (n8077,n3208,n556);
and (n8078,n3214,n567);
and (n8079,n3218,n571);
and (n8080,n1283,n573);
and (n8081,n8082,n4903);
or (n8082,1'b0,n8083,n8084,n8085,n8086);
and (n8083,n3214,n556);
and (n8084,n3218,n567);
and (n8085,n1283,n571);
and (n8086,n779,n573);
or (n8087,1'b0,n8088,n8099,n8101,n8102);
and (n8088,n8089,n2893);
wire s0n8089,s1n8089,notn8089;
or (n8089,s0n8089,s1n8089);
not(notn8089,n2891);
and (s0n8089,notn8089,1'b0);
and (s1n8089,n2891,n8090);
wire s0n8090,s1n8090,notn8090;
or (n8090,s0n8090,s1n8090);
not(notn8090,n7861);
and (s0n8090,notn8090,n8091);
and (s1n8090,n7861,1'b0);
wire s0n8091,s1n8091,notn8091;
or (n8091,s0n8091,s1n8091);
not(notn8091,n7846);
and (s0n8091,notn8091,n8092);
and (s1n8091,n7846,1'b1);
wire s0n8092,s1n8092,notn8092;
or (n8092,s0n8092,s1n8092);
not(notn8092,n4966);
and (s0n8092,notn8092,n8093);
and (s1n8092,n4966,n8096);
wire s0n8093,s1n8093,notn8093;
or (n8093,s0n8093,s1n8093);
not(notn8093,n4966);
and (s0n8093,notn8093,n8094);
and (s1n8093,n4966,n8095);
xor (n8094,n7613,n7615);
xor (n8095,n7613,n7616);
wire s0n8096,s1n8096,notn8096;
or (n8096,s0n8096,s1n8096);
not(notn8096,n4966);
and (s0n8096,notn8096,n8097);
and (s1n8096,n4966,n8098);
xor (n8097,n7831,n7833);
xor (n8098,n7831,n7843);
and (n8099,n8100,n2907);
wire s0n8100,s1n8100,notn8100;
or (n8100,s0n8100,s1n8100);
not(notn8100,n2902);
and (s0n8100,notn8100,1'b0);
and (s1n8100,n2902,n8090);
and (n8101,n8090,n7875);
and (n8102,n8002,n7878);
and (n8103,n8087,n8104);
or (n8104,n8105,n8215,n8649);
and (n8105,n8106,n8199);
or (n8106,1'b0,n8107,n8110,n8113,n8118);
and (n8107,n8108,n2893);
wire s0n8108,s1n8108,notn8108;
or (n8108,s0n8108,s1n8108);
not(notn8108,n2891);
and (s0n8108,notn8108,1'b0);
and (s1n8108,n2891,n8109);
and (n8110,n8111,n2907);
wire s0n8111,s1n8111,notn8111;
or (n8111,s0n8111,s1n8111);
not(notn8111,n2902);
and (s0n8111,notn8111,1'b0);
and (s1n8111,n2902,n8112);
and (n8113,n8114,n4883);
wire s0n8114,s1n8114,notn8114;
or (n8114,s0n8114,s1n8114);
not(notn8114,n4878);
and (s0n8114,notn8114,n8115);
and (s1n8114,n4878,1'b0);
wire s0n8115,s1n8115,notn8115;
or (n8115,s0n8115,s1n8115);
not(notn8115,n4873);
and (s0n8115,notn8115,n8116);
and (s1n8115,n4873,1'b1);
wire s0n8116,s1n8116,notn8116;
or (n8116,s0n8116,s1n8116);
not(notn8116,n4861);
and (s0n8116,notn8116,1'b0);
and (s1n8116,n4861,n8117);
xor (n8117,n4845,n4847);
or (n8118,1'b0,n8119,n8139,n8159,n8179);
and (n8119,n8120,n2718);
or (n8120,1'b0,n8121,n8127,n8133);
and (n8121,n8122,n4895);
or (n8122,1'b0,n8123,n8124,n8125,n8126);
and (n8123,n3264,n556);
and (n8124,n3268,n567);
and (n8125,n3272,n571);
and (n8126,n3276,n573);
and (n8127,n8128,n2944);
or (n8128,1'b0,n8129,n8130,n8131,n8132);
and (n8129,n3332,n556);
and (n8130,n3263,n567);
and (n8131,n3267,n571);
and (n8132,n3271,n573);
and (n8133,n8134,n4903);
or (n8134,1'b0,n8135,n8136,n8137,n8138);
and (n8135,n3263,n556);
and (n8136,n3267,n567);
and (n8137,n3271,n571);
and (n8138,n3275,n573);
and (n8139,n8140,n2730);
or (n8140,1'b0,n8141,n8147,n8153);
and (n8141,n8142,n4895);
or (n8142,1'b0,n8143,n8144,n8145,n8146);
and (n8143,n3282,n556);
and (n8144,n3286,n567);
and (n8145,n3290,n571);
and (n8146,n3294,n573);
and (n8147,n8148,n2944);
or (n8148,1'b0,n8149,n8150,n8151,n8152);
and (n8149,n3275,n556);
and (n8150,n3281,n567);
and (n8151,n3285,n571);
and (n8152,n3289,n573);
and (n8153,n8154,n4903);
or (n8154,1'b0,n8155,n8156,n8157,n8158);
and (n8155,n3281,n556);
and (n8156,n3285,n567);
and (n8157,n3289,n571);
and (n8158,n3293,n573);
and (n8159,n8160,n2742);
or (n8160,1'b0,n8161,n8167,n8173);
and (n8161,n8162,n4895);
or (n8162,1'b0,n8163,n8164,n8165,n8166);
and (n8163,n3300,n556);
and (n8164,n3304,n567);
and (n8165,n3308,n571);
and (n8166,n3312,n573);
and (n8167,n8168,n2944);
or (n8168,1'b0,n8169,n8170,n8171,n8172);
and (n8169,n3347,n556);
and (n8170,n3299,n567);
and (n8171,n3303,n571);
and (n8172,n3307,n573);
and (n8173,n8174,n4903);
or (n8174,1'b0,n8175,n8176,n8177,n8178);
and (n8175,n3299,n556);
and (n8176,n3303,n567);
and (n8177,n3307,n571);
and (n8178,n3311,n573);
and (n8179,n8180,n2752);
or (n8180,1'b0,n8181,n8187,n8193);
and (n8181,n8182,n4895);
or (n8182,1'b0,n8183,n8184,n8185,n8186);
and (n8183,n3318,n556);
and (n8184,n3322,n567);
and (n8185,n2135,n571);
and (n8186,n1753,n573);
and (n8187,n8188,n2944);
or (n8188,1'b0,n8189,n8190,n8191,n8192);
and (n8189,n3311,n556);
and (n8190,n3317,n567);
and (n8191,n3321,n571);
and (n8192,n1299,n573);
and (n8193,n8194,n4903);
or (n8194,1'b0,n8195,n8196,n8197,n8198);
and (n8195,n3317,n556);
and (n8196,n3321,n567);
and (n8197,n1299,n571);
and (n8198,n795,n573);
or (n8199,1'b0,n8200,n8211,n8213,n8214);
and (n8200,n8201,n2893);
wire s0n8201,s1n8201,notn8201;
or (n8201,s0n8201,s1n8201);
not(notn8201,n2891);
and (s0n8201,notn8201,1'b0);
and (s1n8201,n2891,n8202);
wire s0n8202,s1n8202,notn8202;
or (n8202,s0n8202,s1n8202);
not(notn8202,n7861);
and (s0n8202,notn8202,n8203);
and (s1n8202,n7861,1'b0);
wire s0n8203,s1n8203,notn8203;
or (n8203,s0n8203,s1n8203);
not(notn8203,n7846);
and (s0n8203,notn8203,n8204);
and (s1n8203,n7846,1'b1);
wire s0n8204,s1n8204,notn8204;
or (n8204,s0n8204,s1n8204);
not(notn8204,n4966);
and (s0n8204,notn8204,n8205);
and (s1n8204,n4966,n8208);
wire s0n8205,s1n8205,notn8205;
or (n8205,s0n8205,s1n8205);
not(notn8205,n4966);
and (s0n8205,notn8205,n8206);
and (s1n8205,n4966,n8207);
xor (n8206,n7616,n7618);
not (n8207,n7616);
wire s0n8208,s1n8208,notn8208;
or (n8208,s0n8208,s1n8208);
not(notn8208,n4966);
and (s0n8208,notn8208,n8209);
and (s1n8208,n4966,n8210);
xor (n8209,n7834,n7836);
xor (n8210,n7834,n7844);
and (n8211,n8212,n2907);
wire s0n8212,s1n8212,notn8212;
or (n8212,s0n8212,s1n8212);
not(notn8212,n2902);
and (s0n8212,notn8212,1'b0);
and (s1n8212,n2902,n8202);
and (n8213,n8202,n7875);
and (n8214,n8114,n7878);
and (n8215,n8199,n8216);
or (n8216,n8217,n8323,n8648);
and (n8217,n8218,n8311);
or (n8218,1'b0,n8219,n8222,n8225,n8230);
and (n8219,n8220,n2893);
wire s0n8220,s1n8220,notn8220;
or (n8220,s0n8220,s1n8220);
not(notn8220,n2891);
and (s0n8220,notn8220,1'b0);
and (s1n8220,n2891,n8221);
and (n8222,n8223,n2907);
wire s0n8223,s1n8223,notn8223;
or (n8223,s0n8223,s1n8223);
not(notn8223,n2902);
and (s0n8223,notn8223,1'b0);
and (s1n8223,n2902,n8224);
and (n8225,n8226,n4883);
wire s0n8226,s1n8226,notn8226;
or (n8226,s0n8226,s1n8226);
not(notn8226,n4878);
and (s0n8226,notn8226,n8227);
and (s1n8226,n4878,1'b0);
wire s0n8227,s1n8227,notn8227;
or (n8227,s0n8227,s1n8227);
not(notn8227,n4873);
and (s0n8227,notn8227,n8228);
and (s1n8227,n4873,1'b1);
wire s0n8228,s1n8228,notn8228;
or (n8228,s0n8228,s1n8228);
not(notn8228,n4861);
and (s0n8228,notn8228,1'b0);
and (s1n8228,n4861,n8229);
xor (n8229,n4848,n4850);
or (n8230,1'b0,n8231,n8251,n8271,n8291);
and (n8231,n8232,n2718);
or (n8232,1'b0,n8233,n8239,n8245);
and (n8233,n8234,n4895);
or (n8234,1'b0,n8235,n8236,n8237,n8238);
and (n8235,n3367,n556);
and (n8236,n3371,n567);
and (n8237,n3375,n571);
and (n8238,n3379,n573);
and (n8239,n8240,n2944);
or (n8240,1'b0,n8241,n8242,n8243,n8244);
and (n8241,n3435,n556);
and (n8242,n3366,n567);
and (n8243,n3370,n571);
and (n8244,n3374,n573);
and (n8245,n8246,n4903);
or (n8246,1'b0,n8247,n8248,n8249,n8250);
and (n8247,n3366,n556);
and (n8248,n3370,n567);
and (n8249,n3374,n571);
and (n8250,n3378,n573);
and (n8251,n8252,n2730);
or (n8252,1'b0,n8253,n8259,n8265);
and (n8253,n8254,n4895);
or (n8254,1'b0,n8255,n8256,n8257,n8258);
and (n8255,n3385,n556);
and (n8256,n3389,n567);
and (n8257,n3393,n571);
and (n8258,n3397,n573);
and (n8259,n8260,n2944);
or (n8260,1'b0,n8261,n8262,n8263,n8264);
and (n8261,n3378,n556);
and (n8262,n3384,n567);
and (n8263,n3388,n571);
and (n8264,n3392,n573);
and (n8265,n8266,n4903);
or (n8266,1'b0,n8267,n8268,n8269,n8270);
and (n8267,n3384,n556);
and (n8268,n3388,n567);
and (n8269,n3392,n571);
and (n8270,n3396,n573);
and (n8271,n8272,n2742);
or (n8272,1'b0,n8273,n8279,n8285);
and (n8273,n8274,n4895);
or (n8274,1'b0,n8275,n8276,n8277,n8278);
and (n8275,n3403,n556);
and (n8276,n3407,n567);
and (n8277,n3411,n571);
and (n8278,n3415,n573);
and (n8279,n8280,n2944);
or (n8280,1'b0,n8281,n8282,n8283,n8284);
and (n8281,n3450,n556);
and (n8282,n3402,n567);
and (n8283,n3406,n571);
and (n8284,n3410,n573);
and (n8285,n8286,n4903);
or (n8286,1'b0,n8287,n8288,n8289,n8290);
and (n8287,n3402,n556);
and (n8288,n3406,n567);
and (n8289,n3410,n571);
and (n8290,n3414,n573);
and (n8291,n8292,n2752);
or (n8292,1'b0,n8293,n8299,n8305);
and (n8293,n8294,n4895);
or (n8294,1'b0,n8295,n8296,n8297,n8298);
and (n8295,n3421,n556);
and (n8296,n3425,n567);
and (n8297,n2151,n571);
and (n8298,n1769,n573);
and (n8299,n8300,n2944);
or (n8300,1'b0,n8301,n8302,n8303,n8304);
and (n8301,n3414,n556);
and (n8302,n3420,n567);
and (n8303,n3424,n571);
and (n8304,n1315,n573);
and (n8305,n8306,n4903);
or (n8306,1'b0,n8307,n8308,n8309,n8310);
and (n8307,n3420,n556);
and (n8308,n3424,n567);
and (n8309,n1315,n571);
and (n8310,n811,n573);
or (n8311,1'b0,n8312,n8319,n8321,n8322);
and (n8312,n8313,n2893);
wire s0n8313,s1n8313,notn8313;
or (n8313,s0n8313,s1n8313);
not(notn8313,n2891);
and (s0n8313,notn8313,1'b0);
and (s1n8313,n2891,n8314);
wire s0n8314,s1n8314,notn8314;
or (n8314,s0n8314,s1n8314);
not(notn8314,n7861);
and (s0n8314,notn8314,n8315);
and (s1n8314,n7861,1'b0);
wire s0n8315,s1n8315,notn8315;
or (n8315,s0n8315,s1n8315);
not(notn8315,n7846);
and (s0n8315,notn8315,n8316);
and (s1n8315,n7846,1'b1);
wire s0n8316,s1n8316,notn8316;
or (n8316,s0n8316,s1n8316);
not(notn8316,n4966);
and (s0n8316,notn8316,n8317);
and (s1n8316,n4966,n7847);
wire s0n8317,s1n8317,notn8317;
or (n8317,s0n8317,s1n8317);
not(notn8317,n4966);
and (s0n8317,notn8317,n8318);
and (s1n8317,n4966,n7619);
xor (n8318,n7619,n7621);
and (n8319,n8320,n2907);
wire s0n8320,s1n8320,notn8320;
or (n8320,s0n8320,s1n8320);
not(notn8320,n2902);
and (s0n8320,notn8320,1'b0);
and (s1n8320,n2902,n8314);
and (n8321,n8314,n7875);
and (n8322,n8226,n7878);
and (n8323,n8311,n8324);
or (n8324,n8325,n8431,n8647);
and (n8325,n8326,n8419);
or (n8326,1'b0,n8327,n8330,n8333,n8338);
and (n8327,n8328,n2893);
wire s0n8328,s1n8328,notn8328;
or (n8328,s0n8328,s1n8328);
not(notn8328,n2891);
and (s0n8328,notn8328,1'b0);
and (s1n8328,n2891,n8329);
and (n8330,n8331,n2907);
wire s0n8331,s1n8331,notn8331;
or (n8331,s0n8331,s1n8331);
not(notn8331,n2902);
and (s0n8331,notn8331,1'b0);
and (s1n8331,n2902,n8332);
and (n8333,n8334,n4883);
wire s0n8334,s1n8334,notn8334;
or (n8334,s0n8334,s1n8334);
not(notn8334,n4878);
and (s0n8334,notn8334,n8335);
and (s1n8334,n4878,1'b0);
wire s0n8335,s1n8335,notn8335;
or (n8335,s0n8335,s1n8335);
not(notn8335,n4873);
and (s0n8335,notn8335,n8336);
and (s1n8335,n4873,1'b1);
wire s0n8336,s1n8336,notn8336;
or (n8336,s0n8336,s1n8336);
not(notn8336,n4861);
and (s0n8336,notn8336,1'b0);
and (s1n8336,n4861,n8337);
xor (n8337,n4851,n4853);
or (n8338,1'b0,n8339,n8359,n8379,n8399);
and (n8339,n8340,n2718);
or (n8340,1'b0,n8341,n8347,n8353);
and (n8341,n8342,n4895);
or (n8342,1'b0,n8343,n8344,n8345,n8346);
and (n8343,n3470,n556);
and (n8344,n3474,n567);
and (n8345,n3478,n571);
and (n8346,n3482,n573);
and (n8347,n8348,n2944);
or (n8348,1'b0,n8349,n8350,n8351,n8352);
and (n8349,n3538,n556);
and (n8350,n3469,n567);
and (n8351,n3473,n571);
and (n8352,n3477,n573);
and (n8353,n8354,n4903);
or (n8354,1'b0,n8355,n8356,n8357,n8358);
and (n8355,n3469,n556);
and (n8356,n3473,n567);
and (n8357,n3477,n571);
and (n8358,n3481,n573);
and (n8359,n8360,n2730);
or (n8360,1'b0,n8361,n8367,n8373);
and (n8361,n8362,n4895);
or (n8362,1'b0,n8363,n8364,n8365,n8366);
and (n8363,n3488,n556);
and (n8364,n3492,n567);
and (n8365,n3496,n571);
and (n8366,n3500,n573);
and (n8367,n8368,n2944);
or (n8368,1'b0,n8369,n8370,n8371,n8372);
and (n8369,n3481,n556);
and (n8370,n3487,n567);
and (n8371,n3491,n571);
and (n8372,n3495,n573);
and (n8373,n8374,n4903);
or (n8374,1'b0,n8375,n8376,n8377,n8378);
and (n8375,n3487,n556);
and (n8376,n3491,n567);
and (n8377,n3495,n571);
and (n8378,n3499,n573);
and (n8379,n8380,n2742);
or (n8380,1'b0,n8381,n8387,n8393);
and (n8381,n8382,n4895);
or (n8382,1'b0,n8383,n8384,n8385,n8386);
and (n8383,n3506,n556);
and (n8384,n3510,n567);
and (n8385,n3514,n571);
and (n8386,n3518,n573);
and (n8387,n8388,n2944);
or (n8388,1'b0,n8389,n8390,n8391,n8392);
and (n8389,n3553,n556);
and (n8390,n3505,n567);
and (n8391,n3509,n571);
and (n8392,n3513,n573);
and (n8393,n8394,n4903);
or (n8394,1'b0,n8395,n8396,n8397,n8398);
and (n8395,n3505,n556);
and (n8396,n3509,n567);
and (n8397,n3513,n571);
and (n8398,n3517,n573);
and (n8399,n8400,n2752);
or (n8400,1'b0,n8401,n8407,n8413);
and (n8401,n8402,n4895);
or (n8402,1'b0,n8403,n8404,n8405,n8406);
and (n8403,n3524,n556);
and (n8404,n3528,n567);
and (n8405,n2167,n571);
and (n8406,n1790,n573);
and (n8407,n8408,n2944);
or (n8408,1'b0,n8409,n8410,n8411,n8412);
and (n8409,n3517,n556);
and (n8410,n3523,n567);
and (n8411,n3527,n571);
and (n8412,n1331,n573);
and (n8413,n8414,n4903);
or (n8414,1'b0,n8415,n8416,n8417,n8418);
and (n8415,n3523,n556);
and (n8416,n3527,n567);
and (n8417,n1331,n571);
and (n8418,n827,n573);
or (n8419,1'b0,n8420,n8427,n8429,n8430);
and (n8420,n8421,n2893);
wire s0n8421,s1n8421,notn8421;
or (n8421,s0n8421,s1n8421);
not(notn8421,n2891);
and (s0n8421,notn8421,1'b0);
and (s1n8421,n2891,n8422);
wire s0n8422,s1n8422,notn8422;
or (n8422,s0n8422,s1n8422);
not(notn8422,n7861);
and (s0n8422,notn8422,n8423);
and (s1n8422,n7861,1'b0);
wire s0n8423,s1n8423,notn8423;
or (n8423,s0n8423,s1n8423);
not(notn8423,n7846);
and (s0n8423,notn8423,n8424);
and (s1n8423,n7846,1'b1);
wire s0n8424,s1n8424,notn8424;
or (n8424,s0n8424,s1n8424);
not(notn8424,n4966);
and (s0n8424,notn8424,n8425);
and (s1n8424,n4966,n4956);
wire s0n8425,s1n8425,notn8425;
or (n8425,s0n8425,s1n8425);
not(notn8425,n4966);
and (s0n8425,notn8425,n8426);
and (s1n8425,n4966,n7622);
xor (n8426,n7622,n7624);
and (n8427,n8428,n2907);
wire s0n8428,s1n8428,notn8428;
or (n8428,s0n8428,s1n8428);
not(notn8428,n2902);
and (s0n8428,notn8428,1'b0);
and (s1n8428,n2902,n8422);
and (n8429,n8422,n7875);
and (n8430,n8334,n7878);
and (n8431,n8419,n8432);
or (n8432,n8433,n8539,n8646);
and (n8433,n8434,n8527);
or (n8434,1'b0,n8435,n8438,n8441,n8446);
and (n8435,n8436,n2893);
wire s0n8436,s1n8436,notn8436;
or (n8436,s0n8436,s1n8436);
not(notn8436,n2891);
and (s0n8436,notn8436,1'b0);
and (s1n8436,n2891,n8437);
and (n8438,n8439,n2907);
wire s0n8439,s1n8439,notn8439;
or (n8439,s0n8439,s1n8439);
not(notn8439,n2902);
and (s0n8439,notn8439,1'b0);
and (s1n8439,n2902,n8440);
and (n8441,n8442,n4883);
wire s0n8442,s1n8442,notn8442;
or (n8442,s0n8442,s1n8442);
not(notn8442,n4878);
and (s0n8442,notn8442,n8443);
and (s1n8442,n4878,1'b0);
wire s0n8443,s1n8443,notn8443;
or (n8443,s0n8443,s1n8443);
not(notn8443,n4873);
and (s0n8443,notn8443,n8444);
and (s1n8443,n4873,1'b1);
wire s0n8444,s1n8444,notn8444;
or (n8444,s0n8444,s1n8444);
not(notn8444,n4861);
and (s0n8444,notn8444,1'b0);
and (s1n8444,n4861,n8445);
xor (n8445,n4854,n4856);
or (n8446,1'b0,n8447,n8467,n8487,n8507);
and (n8447,n8448,n2718);
or (n8448,1'b0,n8449,n8455,n8461);
and (n8449,n8450,n4895);
or (n8450,1'b0,n8451,n8452,n8453,n8454);
and (n8451,n3573,n556);
and (n8452,n3577,n567);
and (n8453,n3581,n571);
and (n8454,n3585,n573);
and (n8455,n8456,n2944);
or (n8456,1'b0,n8457,n8458,n8459,n8460);
and (n8457,n3641,n556);
and (n8458,n3572,n567);
and (n8459,n3576,n571);
and (n8460,n3580,n573);
and (n8461,n8462,n4903);
or (n8462,1'b0,n8463,n8464,n8465,n8466);
and (n8463,n3572,n556);
and (n8464,n3576,n567);
and (n8465,n3580,n571);
and (n8466,n3584,n573);
and (n8467,n8468,n2730);
or (n8468,1'b0,n8469,n8475,n8481);
and (n8469,n8470,n4895);
or (n8470,1'b0,n8471,n8472,n8473,n8474);
and (n8471,n3591,n556);
and (n8472,n3595,n567);
and (n8473,n3599,n571);
and (n8474,n3603,n573);
and (n8475,n8476,n2944);
or (n8476,1'b0,n8477,n8478,n8479,n8480);
and (n8477,n3584,n556);
and (n8478,n3590,n567);
and (n8479,n3594,n571);
and (n8480,n3598,n573);
and (n8481,n8482,n4903);
or (n8482,1'b0,n8483,n8484,n8485,n8486);
and (n8483,n3590,n556);
and (n8484,n3594,n567);
and (n8485,n3598,n571);
and (n8486,n3602,n573);
and (n8487,n8488,n2742);
or (n8488,1'b0,n8489,n8495,n8501);
and (n8489,n8490,n4895);
or (n8490,1'b0,n8491,n8492,n8493,n8494);
and (n8491,n3609,n556);
and (n8492,n3613,n567);
and (n8493,n3617,n571);
and (n8494,n3621,n573);
and (n8495,n8496,n2944);
or (n8496,1'b0,n8497,n8498,n8499,n8500);
and (n8497,n3656,n556);
and (n8498,n3608,n567);
and (n8499,n3612,n571);
and (n8500,n3616,n573);
and (n8501,n8502,n4903);
or (n8502,1'b0,n8503,n8504,n8505,n8506);
and (n8503,n3608,n556);
and (n8504,n3612,n567);
and (n8505,n3616,n571);
and (n8506,n3620,n573);
and (n8507,n8508,n2752);
or (n8508,1'b0,n8509,n8515,n8521);
and (n8509,n8510,n4895);
or (n8510,1'b0,n8511,n8512,n8513,n8514);
and (n8511,n3627,n556);
and (n8512,n3631,n567);
and (n8513,n2184,n571);
and (n8514,n1820,n573);
and (n8515,n8516,n2944);
or (n8516,1'b0,n8517,n8518,n8519,n8520);
and (n8517,n3620,n556);
and (n8518,n3626,n567);
and (n8519,n3630,n571);
and (n8520,n1347,n573);
and (n8521,n8522,n4903);
or (n8522,1'b0,n8523,n8524,n8525,n8526);
and (n8523,n3626,n556);
and (n8524,n3630,n567);
and (n8525,n1347,n571);
and (n8526,n843,n573);
or (n8527,1'b0,n8528,n8535,n8537,n8538);
and (n8528,n8529,n2893);
wire s0n8529,s1n8529,notn8529;
or (n8529,s0n8529,s1n8529);
not(notn8529,n2891);
and (s0n8529,notn8529,1'b0);
and (s1n8529,n2891,n8530);
wire s0n8530,s1n8530,notn8530;
or (n8530,s0n8530,s1n8530);
not(notn8530,n7861);
and (s0n8530,notn8530,n8531);
and (s1n8530,n7861,1'b0);
wire s0n8531,s1n8531,notn8531;
or (n8531,s0n8531,s1n8531);
not(notn8531,n7846);
and (s0n8531,notn8531,n8532);
and (s1n8531,n7846,1'b1);
wire s0n8532,s1n8532,notn8532;
or (n8532,s0n8532,s1n8532);
not(notn8532,n4966);
and (s0n8532,notn8532,n8533);
and (s1n8532,n4966,n7981);
wire s0n8533,s1n8533,notn8533;
or (n8533,s0n8533,s1n8533);
not(notn8533,n4966);
and (s0n8533,notn8533,n8534);
and (s1n8533,n4966,n7625);
xor (n8534,n7625,n7627);
and (n8535,n8536,n2907);
wire s0n8536,s1n8536,notn8536;
or (n8536,s0n8536,s1n8536);
not(notn8536,n2902);
and (s0n8536,notn8536,1'b0);
and (s1n8536,n2902,n8530);
and (n8537,n8530,n7875);
and (n8538,n8442,n7878);
and (n8539,n8527,n8540);
and (n8540,n8541,n8634);
or (n8541,1'b0,n8542,n8545,n8548,n8553);
and (n8542,n8543,n2893);
wire s0n8543,s1n8543,notn8543;
or (n8543,s0n8543,s1n8543);
not(notn8543,n2891);
and (s0n8543,notn8543,1'b0);
and (s1n8543,n2891,n8544);
and (n8545,n8546,n2907);
wire s0n8546,s1n8546,notn8546;
or (n8546,s0n8546,s1n8546);
not(notn8546,n2902);
and (s0n8546,notn8546,1'b0);
and (s1n8546,n2902,n8547);
and (n8548,n8549,n4883);
wire s0n8549,s1n8549,notn8549;
or (n8549,s0n8549,s1n8549);
not(notn8549,n4878);
and (s0n8549,notn8549,n8550);
and (s1n8549,n4878,1'b0);
wire s0n8550,s1n8550,notn8550;
or (n8550,s0n8550,s1n8550);
not(notn8550,n4873);
and (s0n8550,notn8550,n8551);
and (s1n8550,n4873,1'b1);
wire s0n8551,s1n8551,notn8551;
or (n8551,s0n8551,s1n8551);
not(notn8551,n4861);
and (s0n8551,notn8551,1'b0);
and (s1n8551,n4861,n8552);
xor (n8552,n4857,n4859);
or (n8553,1'b0,n8554,n8574,n8594,n8614);
and (n8554,n8555,n2718);
or (n8555,1'b0,n8556,n8562,n8568);
and (n8556,n8557,n4895);
or (n8557,1'b0,n8558,n8559,n8560,n8561);
and (n8558,n3675,n556);
and (n8559,n3679,n567);
and (n8560,n3683,n571);
and (n8561,n3687,n573);
and (n8562,n8563,n2944);
or (n8563,1'b0,n8564,n8565,n8566,n8567);
and (n8564,n3743,n556);
and (n8565,n3674,n567);
and (n8566,n3678,n571);
and (n8567,n3682,n573);
and (n8568,n8569,n4903);
or (n8569,1'b0,n8570,n8571,n8572,n8573);
and (n8570,n3674,n556);
and (n8571,n3678,n567);
and (n8572,n3682,n571);
and (n8573,n3686,n573);
and (n8574,n8575,n2730);
or (n8575,1'b0,n8576,n8582,n8588);
and (n8576,n8577,n4895);
or (n8577,1'b0,n8578,n8579,n8580,n8581);
and (n8578,n3693,n556);
and (n8579,n3697,n567);
and (n8580,n3701,n571);
and (n8581,n3705,n573);
and (n8582,n8583,n2944);
or (n8583,1'b0,n8584,n8585,n8586,n8587);
and (n8584,n3686,n556);
and (n8585,n3692,n567);
and (n8586,n3696,n571);
and (n8587,n3700,n573);
and (n8588,n8589,n4903);
or (n8589,1'b0,n8590,n8591,n8592,n8593);
and (n8590,n3692,n556);
and (n8591,n3696,n567);
and (n8592,n3700,n571);
and (n8593,n3704,n573);
and (n8594,n8595,n2742);
or (n8595,1'b0,n8596,n8602,n8608);
and (n8596,n8597,n4895);
or (n8597,1'b0,n8598,n8599,n8600,n8601);
and (n8598,n3711,n556);
and (n8599,n3715,n567);
and (n8600,n3719,n571);
and (n8601,n3723,n573);
and (n8602,n8603,n2944);
or (n8603,1'b0,n8604,n8605,n8606,n8607);
and (n8604,n3758,n556);
and (n8605,n3710,n567);
and (n8606,n3714,n571);
and (n8607,n3718,n573);
and (n8608,n8609,n4903);
or (n8609,1'b0,n8610,n8611,n8612,n8613);
and (n8610,n3710,n556);
and (n8611,n3714,n567);
and (n8612,n3718,n571);
and (n8613,n3722,n573);
and (n8614,n8615,n2752);
or (n8615,1'b0,n8616,n8622,n8628);
and (n8616,n8617,n4895);
or (n8617,1'b0,n8618,n8619,n8620,n8621);
and (n8618,n3729,n556);
and (n8619,n3733,n567);
and (n8620,n2199,n571);
and (n8621,n1843,n573);
and (n8622,n8623,n2944);
or (n8623,1'b0,n8624,n8625,n8626,n8627);
and (n8624,n3722,n556);
and (n8625,n3728,n567);
and (n8626,n3732,n571);
and (n8627,n1362,n573);
and (n8628,n8629,n4903);
or (n8629,1'b0,n8630,n8631,n8632,n8633);
and (n8630,n3728,n556);
and (n8631,n3732,n567);
and (n8632,n1362,n571);
and (n8633,n858,n573);
or (n8634,1'b0,n8635,n8642,n8644,n8645);
and (n8635,n8636,n2893);
wire s0n8636,s1n8636,notn8636;
or (n8636,s0n8636,s1n8636);
not(notn8636,n2891);
and (s0n8636,notn8636,1'b0);
and (s1n8636,n2891,n8637);
wire s0n8637,s1n8637,notn8637;
or (n8637,s0n8637,s1n8637);
not(notn8637,n7861);
and (s0n8637,notn8637,n8638);
and (s1n8637,n7861,1'b0);
wire s0n8638,s1n8638,notn8638;
or (n8638,s0n8638,s1n8638);
not(notn8638,n7846);
and (s0n8638,notn8638,n8639);
and (s1n8638,n7846,1'b1);
wire s0n8639,s1n8639,notn8639;
or (n8639,s0n8639,s1n8639);
not(notn8639,n4966);
and (s0n8639,notn8639,n8640);
and (s1n8639,n4966,n8093);
wire s0n8640,s1n8640,notn8640;
or (n8640,s0n8640,s1n8640);
not(notn8640,n4966);
and (s0n8640,notn8640,n8641);
and (s1n8640,n4966,n7628);
xor (n8641,n7628,n7630);
and (n8642,n8643,n2907);
wire s0n8643,s1n8643,notn8643;
or (n8643,s0n8643,s1n8643);
not(notn8643,n2902);
and (s0n8643,notn8643,1'b0);
and (s1n8643,n2902,n8637);
and (n8644,n8637,n7875);
and (n8645,n8549,n7878);
and (n8646,n8434,n8540);
and (n8647,n8326,n8432);
and (n8648,n8218,n8324);
and (n8649,n8106,n8216);
and (n8650,n7994,n8104);
and (n8651,n7882,n7992);
and (n8652,n2887,n7880);
and (n8653,n8654,n8656);
xor (n8654,n8655,n7880);
xor (n8655,n2887,n4950);
and (n8656,n8657,n8659);
xor (n8657,n8658,n7992);
xor (n8658,n7882,n7975);
and (n8659,n8660,n8662);
xor (n8660,n8661,n8104);
xor (n8661,n7994,n8087);
and (n8662,n8663,n8665);
xor (n8663,n8664,n8216);
xor (n8664,n8106,n8199);
and (n8665,n8666,n8668);
xor (n8666,n8667,n8324);
xor (n8667,n8218,n8311);
and (n8668,n8669,n8671);
xor (n8669,n8670,n8432);
xor (n8670,n8326,n8419);
and (n8671,n8672,n8674);
xor (n8672,n8673,n8540);
xor (n8673,n8434,n8527);
xor (n8674,n8541,n8634);
and (n8675,n8676,n8677);
wire s0n8676,s1n8676,notn8676;
or (n8676,s0n8676,s1n8676);
not(notn8676,n4969);
and (s0n8676,notn8676,1'b0);
and (s1n8676,n4969,n2884);
or (n8677,n8678,n2897);
or (n8678,n8679,n2894);
or (n8679,n8680,n2931);
or (n8680,n8681,n2930);
or (n8681,n8682,n4895);
or (n8682,n8683,n2946);
or (n8683,n8684,n2945);
or (n8684,n7878,n4904);
and (n8685,n4952,n2950);
and (n8686,n4953,n5024);
and (n8687,n2911,n2941);
nor (n8688,n2756,n2908,n2909);
and (n8689,n590,n2704);
and (n8690,n3,n8691);
not (n8691,n567);
or (n8692,n8693,n8694);
and (n8693,n7,n608);
and (n8694,n3,n8695);
not (n8695,n608);
and (n8696,n40,n2704);
wire s0n8697,s1n8697,notn8697;
or (n8697,s0n8697,s1n8697);
not(notn8697,n2907);
and (s0n8697,notn8697,n8698);
and (s1n8697,n2907,n13864);
or (n8698,n8699,n13862);
and (n8699,n8700,n573);
wire s0n8700,s1n8700,notn8700;
or (n8700,s0n8700,s1n8700);
not(notn8700,n8689);
and (s0n8700,notn8700,n8701);
and (s1n8700,n8689,n9929);
wire s0n8701,s1n8701,notn8701;
or (n8701,s0n8701,s1n8701);
not(notn8701,n2705);
and (s0n8701,notn8701,n8702);
and (s1n8701,n2705,n9900);
xor (n8702,n8703,n9877);
xor (n8703,n8704,n9779);
xor (n8704,n8705,n9079);
xor (n8705,n8706,n8987);
xor (n8706,n8707,n8847);
xor (n8707,n8708,n8709);
wire s0n8708,s1n8708,notn8708;
or (n8708,s0n8708,s1n8708);
not(notn8708,n928);
and (s0n8708,notn8708,1'b0);
and (s1n8708,n928,n1685);
or (n8709,n8710,n8761,n8846);
and (n8710,n8711,n8714);
xor (n8711,n8712,n8713);
and (n8712,n1890,n928);
wire s0n8713,s1n8713,notn8713;
or (n8713,s0n8713,s1n8713);
not(notn8713,n1081);
and (s0n8713,notn8713,1'b0);
and (s1n8713,n1081,n1685);
and (n8714,n8715,n8716);
wire s0n8715,s1n8715,notn8715;
or (n8715,s0n8715,s1n8715);
not(notn8715,n1084);
and (s0n8715,notn8715,1'b0);
and (s1n8715,n1084,n1685);
or (n8716,n8717,n8719,n8760);
and (n8717,n8718,n1891);
and (n8718,n1890,n1084);
and (n8719,n1891,n8720);
or (n8720,n8721,n8723,n8759);
and (n8721,n8722,n1948);
wire s0n8722,s1n8722,notn8722;
or (n8722,s0n8722,s1n8722);
not(notn8722,n1084);
and (s0n8722,notn8722,1'b0);
and (s1n8722,n1084,n1896);
and (n8723,n1948,n8724);
or (n8724,n8725,n8727,n8758);
and (n8725,n8726,n1956);
and (n8726,n1953,n1084);
and (n8727,n1956,n8728);
or (n8728,n8729,n8731,n8757);
and (n8729,n8730,n1963);
and (n8730,n1961,n1084);
and (n8731,n1963,n8732);
or (n8732,n8733,n8735,n8756);
and (n8733,n8734,n1970);
wire s0n8734,s1n8734,notn8734;
or (n8734,s0n8734,s1n8734);
not(notn8734,n1084);
and (s0n8734,notn8734,1'b0);
and (s1n8734,n1084,n1968);
and (n8735,n1970,n8736);
or (n8736,n8737,n8739,n8755);
and (n8737,n8738,n1977);
wire s0n8738,s1n8738,notn8738;
or (n8738,s0n8738,s1n8738);
not(notn8738,n1084);
and (s0n8738,notn8738,1'b0);
and (s1n8738,n1084,n1975);
and (n8739,n1977,n8740);
or (n8740,n8741,n8743,n8754);
and (n8741,n8742,n1983);
and (n8742,n1982,n1084);
and (n8743,n1983,n8744);
or (n8744,n8745,n8747,n8749);
and (n8745,n8746,n1989);
and (n8746,n1988,n1084);
and (n8747,n1989,n8748);
or (n8748,n8749,n8751,n8752);
and (n8749,n8750,n1995);
wire s0n8750,s1n8750,notn8750;
or (n8750,s0n8750,s1n8750);
not(notn8750,n1084);
and (s0n8750,notn8750,1'b0);
and (s1n8750,n1084,n1994);
and (n8751,n1995,n8752);
and (n8752,n8753,n2000);
wire s0n8753,s1n8753,notn8753;
or (n8753,s0n8753,s1n8753);
not(notn8753,n1084);
and (s0n8753,notn8753,1'b0);
and (s1n8753,n1084,n1999);
and (n8754,n8742,n8744);
and (n8755,n8738,n8740);
and (n8756,n8734,n8736);
and (n8757,n8730,n8732);
and (n8758,n8726,n8728);
and (n8759,n8722,n8724);
and (n8760,n8718,n8720);
and (n8761,n8714,n8762);
or (n8762,n8763,n8768,n8845);
and (n8763,n8764,n8767);
xor (n8764,n8765,n8766);
wire s0n8765,s1n8765,notn8765;
or (n8765,s0n8765,s1n8765);
not(notn8765,n928);
and (s0n8765,notn8765,1'b0);
and (s1n8765,n928,n1896);
and (n8766,n1890,n1081);
xor (n8767,n8715,n8716);
and (n8768,n8767,n8769);
or (n8769,n8770,n8776,n8844);
and (n8770,n8771,n8774);
xor (n8771,n8772,n8773);
and (n8772,n1953,n928);
wire s0n8773,s1n8773,notn8773;
or (n8773,s0n8773,s1n8773);
not(notn8773,n1081);
and (s0n8773,notn8773,1'b0);
and (s1n8773,n1081,n1896);
xor (n8774,n8775,n8720);
xor (n8775,n8718,n1891);
and (n8776,n8774,n8777);
or (n8777,n8778,n8784,n8843);
and (n8778,n8779,n8782);
xor (n8779,n8780,n8781);
and (n8780,n1961,n928);
and (n8781,n1953,n1081);
xor (n8782,n8783,n8724);
xor (n8783,n8722,n1948);
and (n8784,n8782,n8785);
or (n8785,n8786,n8792,n8842);
and (n8786,n8787,n8790);
xor (n8787,n8788,n8789);
wire s0n8788,s1n8788,notn8788;
or (n8788,s0n8788,s1n8788);
not(notn8788,n928);
and (s0n8788,notn8788,1'b0);
and (s1n8788,n928,n1968);
and (n8789,n1961,n1081);
xor (n8790,n8791,n8728);
xor (n8791,n8726,n1956);
and (n8792,n8790,n8793);
or (n8793,n8794,n8800,n8841);
and (n8794,n8795,n8798);
xor (n8795,n8796,n8797);
wire s0n8796,s1n8796,notn8796;
or (n8796,s0n8796,s1n8796);
not(notn8796,n928);
and (s0n8796,notn8796,1'b0);
and (s1n8796,n928,n1975);
wire s0n8797,s1n8797,notn8797;
or (n8797,s0n8797,s1n8797);
not(notn8797,n1081);
and (s0n8797,notn8797,1'b0);
and (s1n8797,n1081,n1968);
xor (n8798,n8799,n8732);
xor (n8799,n8730,n1963);
and (n8800,n8798,n8801);
or (n8801,n8802,n8808,n8840);
and (n8802,n8803,n8806);
xor (n8803,n8804,n8805);
and (n8804,n1982,n928);
wire s0n8805,s1n8805,notn8805;
or (n8805,s0n8805,s1n8805);
not(notn8805,n1081);
and (s0n8805,notn8805,1'b0);
and (s1n8805,n1081,n1975);
xor (n8806,n8807,n8736);
xor (n8807,n8734,n1970);
and (n8808,n8806,n8809);
or (n8809,n8810,n8816,n8839);
and (n8810,n8811,n8814);
xor (n8811,n8812,n8813);
and (n8812,n1988,n928);
and (n8813,n1982,n1081);
xor (n8814,n8815,n8740);
xor (n8815,n8738,n1977);
and (n8816,n8814,n8817);
or (n8817,n8818,n8824,n8838);
and (n8818,n8819,n8822);
xor (n8819,n8820,n8821);
wire s0n8820,s1n8820,notn8820;
or (n8820,s0n8820,s1n8820);
not(notn8820,n928);
and (s0n8820,notn8820,1'b0);
and (s1n8820,n928,n1994);
and (n8821,n1988,n1081);
xor (n8822,n8823,n8744);
xor (n8823,n8742,n1983);
and (n8824,n8822,n8825);
or (n8825,n8826,n8832,n8837);
and (n8826,n8827,n8830);
xor (n8827,n8828,n8829);
wire s0n8828,s1n8828,notn8828;
or (n8828,s0n8828,s1n8828);
not(notn8828,n928);
and (s0n8828,notn8828,1'b0);
and (s1n8828,n928,n1999);
wire s0n8829,s1n8829,notn8829;
or (n8829,s0n8829,s1n8829);
not(notn8829,n1081);
and (s0n8829,notn8829,1'b0);
and (s1n8829,n1081,n1994);
xor (n8830,n8831,n8748);
xor (n8831,n8746,n1989);
and (n8832,n8830,n8833);
and (n8833,n8834,n8835);
wire s0n8834,s1n8834,notn8834;
or (n8834,s0n8834,s1n8834);
not(notn8834,n1081);
and (s0n8834,notn8834,1'b0);
and (s1n8834,n1081,n1999);
xor (n8835,n8836,n8752);
xor (n8836,n8750,n1995);
and (n8837,n8827,n8833);
and (n8838,n8819,n8825);
and (n8839,n8811,n8817);
and (n8840,n8803,n8809);
and (n8841,n8795,n8801);
and (n8842,n8787,n8793);
and (n8843,n8779,n8785);
and (n8844,n8771,n8777);
and (n8845,n8764,n8769);
and (n8846,n8711,n8762);
xor (n8847,n8848,n8849);
wire s0n8848,s1n8848,notn8848;
or (n8848,s0n8848,s1n8848);
not(notn8848,n928);
and (s0n8848,notn8848,1'b0);
and (s1n8848,n928,n2079);
or (n8849,n8850,n8901,n8986);
and (n8850,n8851,n8854);
xor (n8851,n8852,n8853);
wire s0n8852,s1n8852,notn8852;
or (n8852,s0n8852,s1n8852);
not(notn8852,n928);
and (s0n8852,notn8852,1'b0);
and (s1n8852,n928,n2269);
wire s0n8853,s1n8853,notn8853;
or (n8853,s0n8853,s1n8853);
not(notn8853,n1081);
and (s0n8853,notn8853,1'b0);
and (s1n8853,n1081,n2079);
and (n8854,n8855,n8856);
wire s0n8855,s1n8855,notn8855;
or (n8855,s0n8855,s1n8855);
not(notn8855,n1084);
and (s0n8855,notn8855,1'b0);
and (s1n8855,n1084,n2079);
or (n8856,n8857,n8859,n8900);
and (n8857,n8858,n2271);
wire s0n8858,s1n8858,notn8858;
or (n8858,s0n8858,s1n8858);
not(notn8858,n1084);
and (s0n8858,notn8858,1'b0);
and (s1n8858,n1084,n2269);
and (n8859,n2271,n8860);
or (n8860,n8861,n8863,n8899);
and (n8861,n8862,n2359);
and (n8862,n2276,n1084);
and (n8863,n2359,n8864);
or (n8864,n8865,n8867,n8898);
and (n8865,n8866,n2365);
and (n8866,n2364,n1084);
and (n8867,n2365,n8868);
or (n8868,n8869,n8871,n8897);
and (n8869,n8870,n2372);
wire s0n8870,s1n8870,notn8870;
or (n8870,s0n8870,s1n8870);
not(notn8870,n1084);
and (s0n8870,notn8870,1'b0);
and (s1n8870,n1084,n2370);
and (n8871,n2372,n8872);
or (n8872,n8873,n8875,n8896);
and (n8873,n8874,n2378);
and (n8874,n2377,n1084);
and (n8875,n2378,n8876);
or (n8876,n8877,n8879,n8895);
and (n8877,n8878,n2384);
and (n8878,n2383,n1084);
and (n8879,n2384,n8880);
or (n8880,n8881,n8883,n8894);
and (n8881,n8882,n2390);
and (n8882,n2389,n1084);
and (n8883,n2390,n8884);
or (n8884,n8885,n8887,n8889);
and (n8885,n8886,n2396);
wire s0n8886,s1n8886,notn8886;
or (n8886,s0n8886,s1n8886);
not(notn8886,n1084);
and (s0n8886,notn8886,1'b0);
and (s1n8886,n1084,n2395);
and (n8887,n2396,n8888);
or (n8888,n8889,n8891,n8892);
and (n8889,n8890,n2402);
wire s0n8890,s1n8890,notn8890;
or (n8890,s0n8890,s1n8890);
not(notn8890,n1084);
and (s0n8890,notn8890,1'b0);
and (s1n8890,n1084,n2401);
and (n8891,n2402,n8892);
and (n8892,n8893,n2407);
wire s0n8893,s1n8893,notn8893;
or (n8893,s0n8893,s1n8893);
not(notn8893,n1084);
and (s0n8893,notn8893,1'b0);
and (s1n8893,n1084,n2406);
and (n8894,n8882,n8884);
and (n8895,n8878,n8880);
and (n8896,n8874,n8876);
and (n8897,n8870,n8872);
and (n8898,n8866,n8868);
and (n8899,n8862,n8864);
and (n8900,n8858,n8860);
and (n8901,n8854,n8902);
or (n8902,n8903,n8908,n8985);
and (n8903,n8904,n8907);
xor (n8904,n8905,n8906);
and (n8905,n2276,n928);
wire s0n8906,s1n8906,notn8906;
or (n8906,s0n8906,s1n8906);
not(notn8906,n1081);
and (s0n8906,notn8906,1'b0);
and (s1n8906,n1081,n2269);
xor (n8907,n8855,n8856);
and (n8908,n8907,n8909);
or (n8909,n8910,n8916,n8984);
and (n8910,n8911,n8914);
xor (n8911,n8912,n8913);
and (n8912,n2364,n928);
and (n8913,n2276,n1081);
xor (n8914,n8915,n8860);
xor (n8915,n8858,n2271);
and (n8916,n8914,n8917);
or (n8917,n8918,n8924,n8983);
and (n8918,n8919,n8922);
xor (n8919,n8920,n8921);
wire s0n8920,s1n8920,notn8920;
or (n8920,s0n8920,s1n8920);
not(notn8920,n928);
and (s0n8920,notn8920,1'b0);
and (s1n8920,n928,n2370);
and (n8921,n2364,n1081);
xor (n8922,n8923,n8864);
xor (n8923,n8862,n2359);
and (n8924,n8922,n8925);
or (n8925,n8926,n8932,n8982);
and (n8926,n8927,n8930);
xor (n8927,n8928,n8929);
and (n8928,n2377,n928);
wire s0n8929,s1n8929,notn8929;
or (n8929,s0n8929,s1n8929);
not(notn8929,n1081);
and (s0n8929,notn8929,1'b0);
and (s1n8929,n1081,n2370);
xor (n8930,n8931,n8868);
xor (n8931,n8866,n2365);
and (n8932,n8930,n8933);
or (n8933,n8934,n8940,n8981);
and (n8934,n8935,n8938);
xor (n8935,n8936,n8937);
and (n8936,n2383,n928);
and (n8937,n2377,n1081);
xor (n8938,n8939,n8872);
xor (n8939,n8870,n2372);
and (n8940,n8938,n8941);
or (n8941,n8942,n8948,n8980);
and (n8942,n8943,n8946);
xor (n8943,n8944,n8945);
and (n8944,n2389,n928);
and (n8945,n2383,n1081);
xor (n8946,n8947,n8876);
xor (n8947,n8874,n2378);
and (n8948,n8946,n8949);
or (n8949,n8950,n8956,n8979);
and (n8950,n8951,n8954);
xor (n8951,n8952,n8953);
wire s0n8952,s1n8952,notn8952;
or (n8952,s0n8952,s1n8952);
not(notn8952,n928);
and (s0n8952,notn8952,1'b0);
and (s1n8952,n928,n2395);
and (n8953,n2389,n1081);
xor (n8954,n8955,n8880);
xor (n8955,n8878,n2384);
and (n8956,n8954,n8957);
or (n8957,n8958,n8964,n8978);
and (n8958,n8959,n8962);
xor (n8959,n8960,n8961);
and (n8960,n928,n2401);
wire s0n8961,s1n8961,notn8961;
or (n8961,s0n8961,s1n8961);
not(notn8961,n1081);
and (s0n8961,notn8961,1'b0);
and (s1n8961,n1081,n2395);
xor (n8962,n8963,n8884);
xor (n8963,n8882,n2390);
and (n8964,n8962,n8965);
or (n8965,n8966,n8972,n8977);
and (n8966,n8967,n8970);
xor (n8967,n8968,n8969);
wire s0n8968,s1n8968,notn8968;
or (n8968,s0n8968,s1n8968);
not(notn8968,n928);
and (s0n8968,notn8968,1'b0);
and (s1n8968,n928,n2406);
and (n8969,n1081,n2401);
xor (n8970,n8971,n8888);
xor (n8971,n8886,n2396);
and (n8972,n8970,n8973);
and (n8973,n8974,n8975);
wire s0n8974,s1n8974,notn8974;
or (n8974,s0n8974,s1n8974);
not(notn8974,n1081);
and (s0n8974,notn8974,1'b0);
and (s1n8974,n1081,n2406);
xor (n8975,n8976,n8892);
xor (n8976,n8890,n2402);
and (n8977,n8967,n8973);
and (n8978,n8959,n8965);
and (n8979,n8951,n8957);
and (n8980,n8943,n8949);
and (n8981,n8935,n8941);
and (n8982,n8927,n8933);
and (n8983,n8919,n8925);
and (n8984,n8911,n8917);
and (n8985,n8904,n8909);
and (n8986,n8851,n8902);
or (n8987,n8988,n8993,n9078);
and (n8988,n8989,n8991);
xor (n8989,n8990,n8762);
xor (n8990,n8711,n8714);
xor (n8991,n8992,n8902);
xor (n8992,n8851,n8854);
and (n8993,n8991,n8994);
or (n8994,n8995,n9000,n9077);
and (n8995,n8996,n8998);
xor (n8996,n8997,n8769);
xor (n8997,n8764,n8767);
xor (n8998,n8999,n8909);
xor (n8999,n8904,n8907);
and (n9000,n8998,n9001);
or (n9001,n9002,n9007,n9076);
and (n9002,n9003,n9005);
xor (n9003,n9004,n8777);
xor (n9004,n8771,n8774);
xor (n9005,n9006,n8917);
xor (n9006,n8911,n8914);
and (n9007,n9005,n9008);
or (n9008,n9009,n9014,n9075);
and (n9009,n9010,n9012);
xor (n9010,n9011,n8785);
xor (n9011,n8779,n8782);
xor (n9012,n9013,n8925);
xor (n9013,n8919,n8922);
and (n9014,n9012,n9015);
or (n9015,n9016,n9021,n9074);
and (n9016,n9017,n9019);
xor (n9017,n9018,n8793);
xor (n9018,n8787,n8790);
xor (n9019,n9020,n8933);
xor (n9020,n8927,n8930);
and (n9021,n9019,n9022);
or (n9022,n9023,n9028,n9073);
and (n9023,n9024,n9026);
xor (n9024,n9025,n8801);
xor (n9025,n8795,n8798);
xor (n9026,n9027,n8941);
xor (n9027,n8935,n8938);
and (n9028,n9026,n9029);
or (n9029,n9030,n9035,n9072);
and (n9030,n9031,n9033);
xor (n9031,n9032,n8809);
xor (n9032,n8803,n8806);
xor (n9033,n9034,n8949);
xor (n9034,n8943,n8946);
and (n9035,n9033,n9036);
or (n9036,n9037,n9042,n9071);
and (n9037,n9038,n9040);
xor (n9038,n9039,n8817);
xor (n9039,n8811,n8814);
xor (n9040,n9041,n8957);
xor (n9041,n8951,n8954);
and (n9042,n9040,n9043);
or (n9043,n9044,n9049,n9070);
and (n9044,n9045,n9047);
xor (n9045,n9046,n8825);
xor (n9046,n8819,n8822);
xor (n9047,n9048,n8965);
xor (n9048,n8959,n8962);
and (n9049,n9047,n9050);
or (n9050,n9051,n9056,n9069);
and (n9051,n9052,n9054);
xor (n9052,n9053,n8833);
xor (n9053,n8827,n8830);
xor (n9054,n9055,n8973);
xor (n9055,n8967,n8970);
and (n9056,n9054,n9057);
or (n9057,n9058,n9061,n9068);
and (n9058,n9059,n9060);
xor (n9059,n8834,n8835);
xor (n9060,n8974,n8975);
and (n9061,n9060,n9062);
or (n9062,n9063,n9066,n9067);
and (n9063,n9064,n9065);
xor (n9064,n8753,n2000);
xor (n9065,n8893,n2407);
and (n9066,n9065,n2563);
and (n9067,n9064,n2563);
and (n9068,n9059,n9062);
and (n9069,n9052,n9057);
and (n9070,n9045,n9050);
and (n9071,n9038,n9043);
and (n9072,n9031,n9036);
and (n9073,n9024,n9029);
and (n9074,n9017,n9022);
and (n9075,n9010,n9015);
and (n9076,n9003,n9008);
and (n9077,n8996,n9001);
and (n9078,n8989,n8994);
xor (n9079,n9080,n9684);
xor (n9080,n9081,n9394);
or (n9081,n9082,n9326,n9393);
and (n9082,n9083,n9259);
and (n9083,n9084,n930);
xnor (n9084,n9085,n9095);
not (n9085,n9086);
and (n9086,n592,n9087);
wire s0n9087,s1n9087,notn9087;
or (n9087,s0n9087,s1n9087);
not(notn9087,n575);
and (s0n9087,notn9087,n9088);
and (s1n9087,n575,n9089);
wire s0n9088,s1n9088,notn9088;
or (n9088,s0n9088,s1n9088);
not(notn9088,n22);
and (s0n9088,notn9088,1'b0);
and (s1n9088,n22,n566);
or (n9089,1'b0,n9090,n9091,n9093,n9094);
and (n9090,n5053,n556);
and (n9091,n9092,n567);
and (n9093,n564,n571);
and (n9094,n566,n573);
or (n9095,n9096,n9127);
and (n9096,n9097,n9128);
xor (n9097,n9098,n9109);
xor (n9098,n9099,n9100);
and (n9099,n762,n9087);
and (n9100,n592,n9101);
wire s0n9101,s1n9101,notn9101;
or (n9101,s0n9101,s1n9101);
not(notn9101,n575);
and (s0n9101,notn9101,n9102);
and (s1n9101,n575,n9103);
wire s0n9102,s1n9102,notn9102;
or (n9102,s0n9102,s1n9102);
not(notn9102,n22);
and (s0n9102,notn9102,1'b0);
and (s1n9102,n22,n757);
or (n9103,1'b0,n9104,n9105,n9107,n9108);
and (n9104,n5176,n556);
and (n9105,n9106,n567);
and (n9107,n755,n571);
and (n9108,n757,n573);
or (n9109,n9110,n9127);
and (n9110,n9111,n9124);
xor (n9111,n9112,n9123);
xor (n9112,n9113,n9114);
and (n9113,n765,n9087);
and (n9114,n592,n9115);
wire s0n9115,s1n9115,notn9115;
or (n9115,s0n9115,s1n9115);
not(notn9115,n575);
and (s0n9115,notn9115,n9116);
and (s1n9115,n575,n9117);
wire s0n9116,s1n9116,notn9116;
or (n9116,s0n9116,s1n9116);
not(notn9116,n22);
and (s0n9116,notn9116,1'b0);
and (s1n9116,n22,n781);
or (n9117,1'b0,n9118,n9119,n9121,n9122);
and (n9118,n5299,n556);
and (n9119,n9120,n567);
and (n9121,n779,n571);
and (n9122,n781,n573);
and (n9123,n762,n9101);
and (n9124,n9125,n9126);
and (n9125,n765,n9101);
wire s0n9126,s1n9126,notn9126;
or (n9126,s0n9126,s1n9126);
not(notn9126,n699);
and (s0n9126,notn9126,1'b0);
and (s1n9126,n699,n9087);
and (n9127,n9112,n9123);
or (n9128,n9129,n9258);
and (n9129,n9130,n9151);
xor (n9130,n9131,n9150);
or (n9131,n9132,n9149);
and (n9132,n9133,n9146);
xor (n9133,n9134,n9145);
xor (n9134,n9135,n9136);
xor (n9135,n9125,n9126);
and (n9136,n592,n9137);
wire s0n9137,s1n9137,notn9137;
or (n9137,s0n9137,s1n9137);
not(notn9137,n575);
and (s0n9137,notn9137,n9138);
and (s1n9137,n575,n9139);
wire s0n9138,s1n9138,notn9138;
or (n9138,s0n9138,s1n9138);
not(notn9138,n22);
and (s0n9138,notn9138,1'b0);
and (s1n9138,n22,n797);
or (n9139,1'b0,n9140,n9141,n9143,n9144);
and (n9140,n5422,n556);
and (n9141,n9142,n567);
and (n9143,n795,n571);
and (n9144,n797,n573);
and (n9145,n762,n9115);
and (n9146,n9147,n9148);
wire s0n9147,s1n9147,notn9147;
or (n9147,s0n9147,s1n9147);
not(notn9147,n699);
and (s0n9147,notn9147,1'b0);
and (s1n9147,n699,n9101);
and (n9148,n765,n9115);
and (n9149,n9134,n9145);
xor (n9150,n9111,n9124);
or (n9151,n9152,n9257);
and (n9152,n9153,n9174);
xor (n9153,n9154,n9173);
or (n9154,n9155,n9172);
and (n9155,n9156,n9169);
xor (n9156,n9157,n9158);
and (n9157,n762,n9137);
xor (n9158,n9159,n9160);
xor (n9159,n9147,n9148);
and (n9160,n592,n9161);
wire s0n9161,s1n9161,notn9161;
or (n9161,s0n9161,s1n9161);
not(notn9161,n575);
and (s0n9161,notn9161,n9162);
and (s1n9161,n575,n9163);
wire s0n9162,s1n9162,notn9162;
or (n9162,s0n9162,s1n9162);
not(notn9162,n22);
and (s0n9162,notn9162,1'b0);
and (s1n9162,n22,n813);
or (n9163,1'b0,n9164,n9165,n9167,n9168);
and (n9164,n5545,n556);
and (n9165,n9166,n567);
and (n9167,n811,n571);
and (n9168,n813,n573);
and (n9169,n9170,n9171);
wire s0n9170,s1n9170,notn9170;
or (n9170,s0n9170,s1n9170);
not(notn9170,n699);
and (s0n9170,notn9170,1'b0);
and (s1n9170,n699,n9115);
and (n9171,n765,n9137);
and (n9172,n9157,n9158);
xor (n9173,n9133,n9146);
or (n9174,n9175,n9256);
and (n9175,n9176,n9197);
xor (n9176,n9177,n9196);
or (n9177,n9178,n9195);
and (n9178,n9179,n9192);
xor (n9179,n9180,n9181);
and (n9180,n762,n9161);
xor (n9181,n9182,n9183);
xor (n9182,n9170,n9171);
and (n9183,n592,n9184);
wire s0n9184,s1n9184,notn9184;
or (n9184,s0n9184,s1n9184);
not(notn9184,n575);
and (s0n9184,notn9184,n9185);
and (s1n9184,n575,n9186);
wire s0n9185,s1n9185,notn9185;
or (n9185,s0n9185,s1n9185);
not(notn9185,n22);
and (s0n9185,notn9185,1'b0);
and (s1n9185,n22,n829);
or (n9186,1'b0,n9187,n9188,n9190,n9191);
and (n9187,n5668,n556);
and (n9188,n9189,n567);
and (n9190,n827,n571);
and (n9191,n829,n573);
and (n9192,n9193,n9194);
and (n9193,n765,n9161);
wire s0n9194,s1n9194,notn9194;
or (n9194,s0n9194,s1n9194);
not(notn9194,n699);
and (s0n9194,notn9194,1'b0);
and (s1n9194,n699,n9137);
and (n9195,n9180,n9181);
xor (n9196,n9156,n9169);
or (n9197,n9198,n9255);
and (n9198,n9199,n9220);
xor (n9199,n9200,n9219);
or (n9200,n9201,n9218);
and (n9201,n9202,n9207);
xor (n9202,n9203,n9204);
and (n9203,n762,n9184);
and (n9204,n9205,n9206);
wire s0n9205,s1n9205,notn9205;
or (n9205,s0n9205,s1n9205);
not(notn9205,n699);
and (s0n9205,notn9205,1'b0);
and (s1n9205,n699,n9161);
and (n9206,n765,n9184);
xor (n9207,n9208,n9209);
xor (n9208,n9193,n9194);
and (n9209,n592,n9210);
wire s0n9210,s1n9210,notn9210;
or (n9210,s0n9210,s1n9210);
not(notn9210,n575);
and (s0n9210,notn9210,n9211);
and (s1n9210,n575,n9212);
wire s0n9211,s1n9211,notn9211;
or (n9211,s0n9211,s1n9211);
not(notn9211,n22);
and (s0n9211,notn9211,1'b0);
and (s1n9211,n22,n845);
or (n9212,1'b0,n9213,n9214,n9216,n9217);
and (n9213,n5791,n556);
and (n9214,n9215,n567);
and (n9216,n843,n571);
and (n9217,n845,n573);
and (n9218,n9203,n9204);
xor (n9219,n9179,n9192);
or (n9220,n9221,n9254);
and (n9221,n9222,n9237);
xor (n9222,n9223,n9236);
and (n9223,n9224,n9235);
xor (n9224,n9225,n9234);
and (n9225,n592,n9226);
wire s0n9226,s1n9226,notn9226;
or (n9226,s0n9226,s1n9226);
not(notn9226,n575);
and (s0n9226,notn9226,n9227);
and (s1n9226,n575,n9228);
wire s0n9227,s1n9227,notn9227;
or (n9227,s0n9227,s1n9227);
not(notn9227,n22);
and (s0n9227,notn9227,1'b0);
and (s1n9227,n22,n860);
or (n9228,1'b0,n9229,n9230,n9232,n9233);
and (n9229,n5913,n556);
and (n9230,n9231,n567);
and (n9232,n858,n571);
and (n9233,n860,n573);
and (n9234,n762,n9210);
xor (n9235,n9205,n9206);
xor (n9236,n9202,n9207);
or (n9237,n9238,n9253);
and (n9238,n9239,n9252);
xor (n9239,n9240,n9243);
and (n9240,n9241,n9242);
wire s0n9241,s1n9241,notn9241;
or (n9241,s0n9241,s1n9241);
not(notn9241,n699);
and (s0n9241,notn9241,1'b0);
and (s1n9241,n699,n9184);
and (n9242,n765,n9210);
or (n9243,n9244,n9251);
and (n9244,n9245,n9250);
xor (n9245,n9246,n9249);
and (n9246,n9247,n9248);
and (n9247,n765,n9226);
wire s0n9248,s1n9248,notn9248;
or (n9248,s0n9248,s1n9248);
not(notn9248,n699);
and (s0n9248,notn9248,1'b0);
and (s1n9248,n699,n9210);
xor (n9249,n9241,n9242);
and (n9250,n762,n9226);
and (n9251,n9246,n9249);
xor (n9252,n9224,n9235);
and (n9253,n9240,n9243);
and (n9254,n9223,n9236);
and (n9255,n9200,n9219);
and (n9256,n9177,n9196);
and (n9257,n9154,n9173);
and (n9258,n9131,n9150);
and (n9259,n9260,n9261);
and (n9260,n9084,n979);
or (n9261,n9262,n9266,n9325);
and (n9262,n9263,n9265);
and (n9263,n9264,n979);
xor (n9264,n9097,n9128);
and (n9265,n9084,n1027);
and (n9266,n9265,n9267);
or (n9267,n9268,n9272,n9324);
and (n9268,n9269,n9271);
and (n9269,n9270,n979);
xor (n9270,n9130,n9151);
and (n9271,n9264,n1027);
and (n9272,n9271,n9273);
or (n9273,n9274,n9278,n9323);
and (n9274,n9275,n9277);
and (n9275,n9276,n979);
xor (n9276,n9153,n9174);
and (n9277,n9270,n1027);
and (n9278,n9277,n9279);
or (n9279,n9280,n9284,n9322);
and (n9280,n9281,n9283);
and (n9281,n9282,n979);
xor (n9282,n9176,n9197);
and (n9283,n9276,n1027);
and (n9284,n9283,n9285);
or (n9285,n9286,n9290,n9321);
and (n9286,n9287,n9289);
and (n9287,n9288,n979);
xor (n9288,n9199,n9220);
and (n9289,n9282,n1027);
and (n9290,n9289,n9291);
or (n9291,n9292,n9296,n9320);
and (n9292,n9293,n9295);
and (n9293,n9294,n979);
xor (n9294,n9222,n9237);
and (n9295,n9288,n1027);
and (n9296,n9295,n9297);
or (n9297,n9298,n9302,n9319);
and (n9298,n9299,n9301);
and (n9299,n9300,n979);
xor (n9300,n9239,n9252);
and (n9301,n9294,n1027);
and (n9302,n9301,n9303);
or (n9303,n9304,n9308,n9310);
and (n9304,n9305,n9307);
and (n9305,n9306,n979);
xor (n9306,n9245,n9250);
and (n9307,n9300,n1027);
and (n9308,n9307,n9309);
or (n9309,n9310,n9314,n9315);
and (n9310,n9311,n9313);
and (n9311,n9312,n979);
xor (n9312,n9247,n9248);
and (n9313,n9306,n1027);
and (n9314,n9313,n9315);
and (n9315,n9316,n9318);
wire s0n9316,s1n9316,notn9316;
or (n9316,s0n9316,s1n9316);
not(notn9316,n979);
and (s0n9316,notn9316,1'b0);
and (s1n9316,n979,n9317);
wire s0n9317,s1n9317,notn9317;
or (n9317,s0n9317,s1n9317);
not(notn9317,n699);
and (s0n9317,notn9317,1'b0);
and (s1n9317,n699,n9226);
and (n9318,n9312,n1027);
and (n9319,n9299,n9303);
and (n9320,n9293,n9297);
and (n9321,n9287,n9291);
and (n9322,n9281,n9285);
and (n9323,n9275,n9279);
and (n9324,n9269,n9273);
and (n9325,n9263,n9267);
and (n9326,n9259,n9327);
or (n9327,n9328,n9331,n9392);
and (n9328,n9329,n9330);
and (n9329,n9264,n930);
xor (n9330,n9260,n9261);
and (n9331,n9330,n9332);
or (n9332,n9333,n9337,n9391);
and (n9333,n9334,n9335);
and (n9334,n9270,n930);
xor (n9335,n9336,n9267);
xor (n9336,n9263,n9265);
and (n9337,n9335,n9338);
or (n9338,n9339,n9343,n9390);
and (n9339,n9340,n9341);
and (n9340,n9276,n930);
xor (n9341,n9342,n9273);
xor (n9342,n9269,n9271);
and (n9343,n9341,n9344);
or (n9344,n9345,n9349,n9389);
and (n9345,n9346,n9347);
and (n9346,n9282,n930);
xor (n9347,n9348,n9279);
xor (n9348,n9275,n9277);
and (n9349,n9347,n9350);
or (n9350,n9351,n9355,n9388);
and (n9351,n9352,n9353);
and (n9352,n9288,n930);
xor (n9353,n9354,n9285);
xor (n9354,n9281,n9283);
and (n9355,n9353,n9356);
or (n9356,n9357,n9361,n9387);
and (n9357,n9358,n9359);
and (n9358,n9294,n930);
xor (n9359,n9360,n9291);
xor (n9360,n9287,n9289);
and (n9361,n9359,n9362);
or (n9362,n9363,n9367,n9386);
and (n9363,n9364,n9365);
and (n9364,n9300,n930);
xor (n9365,n9366,n9297);
xor (n9366,n9293,n9295);
and (n9367,n9365,n9368);
or (n9368,n9369,n9373,n9385);
and (n9369,n9370,n9371);
and (n9370,n9306,n930);
xor (n9371,n9372,n9303);
xor (n9372,n9299,n9301);
and (n9373,n9371,n9374);
or (n9374,n9375,n9379,n9384);
and (n9375,n9376,n9377);
and (n9376,n9312,n930);
xor (n9377,n9378,n9309);
xor (n9378,n9305,n9307);
and (n9379,n9377,n9380);
and (n9380,n9381,n9382);
wire s0n9381,s1n9381,notn9381;
or (n9381,s0n9381,s1n9381);
not(notn9381,n930);
and (s0n9381,notn9381,1'b0);
and (s1n9381,n930,n9317);
xor (n9382,n9383,n9315);
xor (n9383,n9311,n9313);
and (n9384,n9376,n9380);
and (n9385,n9370,n9374);
and (n9386,n9364,n9368);
and (n9387,n9358,n9362);
and (n9388,n9352,n9356);
and (n9389,n9346,n9350);
and (n9390,n9340,n9344);
and (n9391,n9334,n9338);
and (n9392,n9329,n9332);
and (n9393,n9083,n9327);
or (n9394,n9395,n9616,n9683);
and (n9395,n9396,n9542);
wire s0n9396,s1n9396,notn9396;
or (n9396,s0n9396,s1n9396);
not(notn9396,n930);
and (s0n9396,notn9396,1'b0);
and (s1n9396,n930,n9397);
or (n9397,n9398,n9495,n9541);
and (n9398,n9399,n9407);
wire s0n9399,s1n9399,notn9399;
or (n9399,s0n9399,s1n9399);
not(notn9399,n594);
and (s0n9399,notn9399,1'b0);
and (s1n9399,n594,n9400);
wire s0n9400,s1n9400,notn9400;
or (n9400,s0n9400,s1n9400);
not(notn9400,n575);
and (s0n9400,notn9400,n9401);
and (s1n9400,n575,n9402);
wire s0n9401,s1n9401,notn9401;
or (n9401,s0n9401,s1n9401);
not(notn9401,n22);
and (s0n9401,notn9401,1'b0);
and (s1n9401,n22,n1253);
or (n9402,1'b0,n9403,n9404,n2750,n9406);
and (n9403,n5050,n556);
and (n9404,n9405,n567);
and (n9406,n1253,n573);
and (n9407,n9408,n9409);
wire s0n9408,s1n9408,notn9408;
or (n9408,s0n9408,s1n9408);
not(notn9408,n651);
and (s0n9408,notn9408,1'b0);
and (s1n9408,n651,n9400);
or (n9409,n9410,n9420,n9494);
and (n9410,n9411,n9419);
wire s0n9411,s1n9411,notn9411;
or (n9411,s0n9411,s1n9411);
not(notn9411,n651);
and (s0n9411,notn9411,1'b0);
and (s1n9411,n651,n9412);
wire s0n9412,s1n9412,notn9412;
or (n9412,s0n9412,s1n9412);
not(notn9412,n575);
and (s0n9412,notn9412,n9413);
and (s1n9412,n575,n9414);
wire s0n9413,s1n9413,notn9413;
or (n9413,s0n9413,s1n9413);
not(notn9413,n22);
and (s0n9413,notn9413,1'b0);
and (s1n9413,n22,n1269);
or (n9414,1'b0,n9415,n9416,n7973,n9418);
and (n9415,n5173,n556);
and (n9416,n9417,n567);
and (n9418,n1269,n573);
wire s0n9419,s1n9419,notn9419;
or (n9419,s0n9419,s1n9419);
not(notn9419,n699);
and (s0n9419,notn9419,1'b0);
and (s1n9419,n699,n9400);
and (n9420,n9419,n9421);
or (n9421,n9422,n9432,n9493);
and (n9422,n9423,n9431);
wire s0n9423,s1n9423,notn9423;
or (n9423,s0n9423,s1n9423);
not(notn9423,n651);
and (s0n9423,notn9423,1'b0);
and (s1n9423,n651,n9424);
wire s0n9424,s1n9424,notn9424;
or (n9424,s0n9424,s1n9424);
not(notn9424,n575);
and (s0n9424,notn9424,n9425);
and (s1n9424,n575,n9426);
wire s0n9425,s1n9425,notn9425;
or (n9425,s0n9425,s1n9425);
not(notn9425,n22);
and (s0n9425,notn9425,1'b0);
and (s1n9425,n22,n1285);
or (n9426,1'b0,n9427,n9428,n8085,n9430);
and (n9427,n5296,n556);
and (n9428,n9429,n567);
and (n9430,n1285,n573);
wire s0n9431,s1n9431,notn9431;
or (n9431,s0n9431,s1n9431);
not(notn9431,n699);
and (s0n9431,notn9431,1'b0);
and (s1n9431,n699,n9412);
and (n9432,n9431,n9433);
or (n9433,n9434,n9444,n9492);
and (n9434,n9435,n9443);
wire s0n9435,s1n9435,notn9435;
or (n9435,s0n9435,s1n9435);
not(notn9435,n651);
and (s0n9435,notn9435,1'b0);
and (s1n9435,n651,n9436);
wire s0n9436,s1n9436,notn9436;
or (n9436,s0n9436,s1n9436);
not(notn9436,n575);
and (s0n9436,notn9436,n9437);
and (s1n9436,n575,n9438);
wire s0n9437,s1n9437,notn9437;
or (n9437,s0n9437,s1n9437);
not(notn9437,n22);
and (s0n9437,notn9437,1'b0);
and (s1n9437,n22,n1301);
or (n9438,1'b0,n9439,n9440,n8197,n9442);
and (n9439,n5419,n556);
and (n9440,n9441,n567);
and (n9442,n1301,n573);
wire s0n9443,s1n9443,notn9443;
or (n9443,s0n9443,s1n9443);
not(notn9443,n699);
and (s0n9443,notn9443,1'b0);
and (s1n9443,n699,n9424);
and (n9444,n9443,n9445);
or (n9445,n9446,n9456,n9491);
and (n9446,n9447,n9455);
wire s0n9447,s1n9447,notn9447;
or (n9447,s0n9447,s1n9447);
not(notn9447,n651);
and (s0n9447,notn9447,1'b0);
and (s1n9447,n651,n9448);
wire s0n9448,s1n9448,notn9448;
or (n9448,s0n9448,s1n9448);
not(notn9448,n575);
and (s0n9448,notn9448,n9449);
and (s1n9448,n575,n9450);
wire s0n9449,s1n9449,notn9449;
or (n9449,s0n9449,s1n9449);
not(notn9449,n22);
and (s0n9449,notn9449,1'b0);
and (s1n9449,n22,n1317);
or (n9450,1'b0,n9451,n9452,n8309,n9454);
and (n9451,n5542,n556);
and (n9452,n9453,n567);
and (n9454,n1317,n573);
wire s0n9455,s1n9455,notn9455;
or (n9455,s0n9455,s1n9455);
not(notn9455,n699);
and (s0n9455,notn9455,1'b0);
and (s1n9455,n699,n9436);
and (n9456,n9455,n9457);
or (n9457,n9458,n9468,n9470);
and (n9458,n9459,n9467);
wire s0n9459,s1n9459,notn9459;
or (n9459,s0n9459,s1n9459);
not(notn9459,n651);
and (s0n9459,notn9459,1'b0);
and (s1n9459,n651,n9460);
wire s0n9460,s1n9460,notn9460;
or (n9460,s0n9460,s1n9460);
not(notn9460,n575);
and (s0n9460,notn9460,n9461);
and (s1n9460,n575,n9462);
wire s0n9461,s1n9461,notn9461;
or (n9461,s0n9461,s1n9461);
not(notn9461,n22);
and (s0n9461,notn9461,1'b0);
and (s1n9461,n22,n1333);
or (n9462,1'b0,n9463,n9464,n8417,n9466);
and (n9463,n5665,n556);
and (n9464,n9465,n567);
and (n9466,n1333,n573);
wire s0n9467,s1n9467,notn9467;
or (n9467,s0n9467,s1n9467);
not(notn9467,n699);
and (s0n9467,notn9467,1'b0);
and (s1n9467,n699,n9448);
and (n9468,n9467,n9469);
or (n9469,n9470,n9480,n9481);
and (n9470,n9471,n9479);
wire s0n9471,s1n9471,notn9471;
or (n9471,s0n9471,s1n9471);
not(notn9471,n651);
and (s0n9471,notn9471,1'b0);
and (s1n9471,n651,n9472);
wire s0n9472,s1n9472,notn9472;
or (n9472,s0n9472,s1n9472);
not(notn9472,n575);
and (s0n9472,notn9472,n9473);
and (s1n9472,n575,n9474);
wire s0n9473,s1n9473,notn9473;
or (n9473,s0n9473,s1n9473);
not(notn9473,n22);
and (s0n9473,notn9473,1'b0);
and (s1n9473,n22,n1349);
or (n9474,1'b0,n9475,n9476,n8525,n9478);
and (n9475,n5788,n556);
and (n9476,n9477,n567);
and (n9478,n1349,n573);
wire s0n9479,s1n9479,notn9479;
or (n9479,s0n9479,s1n9479);
not(notn9479,n699);
and (s0n9479,notn9479,1'b0);
and (s1n9479,n699,n9460);
and (n9480,n9479,n9481);
and (n9481,n9482,n9490);
wire s0n9482,s1n9482,notn9482;
or (n9482,s0n9482,s1n9482);
not(notn9482,n651);
and (s0n9482,notn9482,1'b0);
and (s1n9482,n651,n9483);
wire s0n9483,s1n9483,notn9483;
or (n9483,s0n9483,s1n9483);
not(notn9483,n575);
and (s0n9483,notn9483,n9484);
and (s1n9483,n575,n9485);
wire s0n9484,s1n9484,notn9484;
or (n9484,s0n9484,s1n9484);
not(notn9484,n22);
and (s0n9484,notn9484,1'b0);
and (s1n9484,n22,n1364);
or (n9485,1'b0,n9486,n9487,n8632,n9489);
and (n9486,n5910,n556);
and (n9487,n9488,n567);
and (n9489,n1364,n573);
wire s0n9490,s1n9490,notn9490;
or (n9490,s0n9490,s1n9490);
not(notn9490,n699);
and (s0n9490,notn9490,1'b0);
and (s1n9490,n699,n9472);
and (n9491,n9447,n9457);
and (n9492,n9435,n9445);
and (n9493,n9423,n9433);
and (n9494,n9411,n9421);
and (n9495,n9407,n9496);
or (n9496,n9497,n9500,n9540);
and (n9497,n9498,n9499);
wire s0n9498,s1n9498,notn9498;
or (n9498,s0n9498,s1n9498);
not(notn9498,n594);
and (s0n9498,notn9498,1'b0);
and (s1n9498,n594,n9412);
xor (n9499,n9408,n9409);
and (n9500,n9499,n9501);
or (n9501,n9502,n9506,n9539);
and (n9502,n9503,n9504);
wire s0n9503,s1n9503,notn9503;
or (n9503,s0n9503,s1n9503);
not(notn9503,n594);
and (s0n9503,notn9503,1'b0);
and (s1n9503,n594,n9424);
xor (n9504,n9505,n9421);
xor (n9505,n9411,n9419);
and (n9506,n9504,n9507);
or (n9507,n9508,n9512,n9538);
and (n9508,n9509,n9510);
wire s0n9509,s1n9509,notn9509;
or (n9509,s0n9509,s1n9509);
not(notn9509,n594);
and (s0n9509,notn9509,1'b0);
and (s1n9509,n594,n9436);
xor (n9510,n9511,n9433);
xor (n9511,n9423,n9431);
and (n9512,n9510,n9513);
or (n9513,n9514,n9518,n9537);
and (n9514,n9515,n9516);
wire s0n9515,s1n9515,notn9515;
or (n9515,s0n9515,s1n9515);
not(notn9515,n594);
and (s0n9515,notn9515,1'b0);
and (s1n9515,n594,n9448);
xor (n9516,n9517,n9445);
xor (n9517,n9435,n9443);
and (n9518,n9516,n9519);
or (n9519,n9520,n9524,n9536);
and (n9520,n9521,n9522);
wire s0n9521,s1n9521,notn9521;
or (n9521,s0n9521,s1n9521);
not(notn9521,n594);
and (s0n9521,notn9521,1'b0);
and (s1n9521,n594,n9460);
xor (n9522,n9523,n9457);
xor (n9523,n9447,n9455);
and (n9524,n9522,n9525);
or (n9525,n9526,n9530,n9535);
and (n9526,n9527,n9528);
wire s0n9527,s1n9527,notn9527;
or (n9527,s0n9527,s1n9527);
not(notn9527,n594);
and (s0n9527,notn9527,1'b0);
and (s1n9527,n594,n9472);
xor (n9528,n9529,n9469);
xor (n9529,n9459,n9467);
and (n9530,n9528,n9531);
and (n9531,n9532,n9533);
wire s0n9532,s1n9532,notn9532;
or (n9532,s0n9532,s1n9532);
not(notn9532,n594);
and (s0n9532,notn9532,1'b0);
and (s1n9532,n594,n9483);
xor (n9533,n9534,n9481);
xor (n9534,n9471,n9479);
and (n9535,n9527,n9531);
and (n9536,n9521,n9525);
and (n9537,n9515,n9519);
and (n9538,n9509,n9513);
and (n9539,n9503,n9507);
and (n9540,n9498,n9501);
and (n9541,n9399,n9496);
and (n9542,n9543,n9544);
wire s0n9543,s1n9543,notn9543;
or (n9543,s0n9543,s1n9543);
not(notn9543,n979);
and (s0n9543,notn9543,1'b0);
and (s1n9543,n979,n9397);
or (n9544,n9545,n9550,n9615);
and (n9545,n9546,n9549);
wire s0n9546,s1n9546,notn9546;
or (n9546,s0n9546,s1n9546);
not(notn9546,n979);
and (s0n9546,notn9546,1'b0);
and (s1n9546,n979,n9547);
xor (n9547,n9548,n9496);
xor (n9548,n9399,n9407);
wire s0n9549,s1n9549,notn9549;
or (n9549,s0n9549,s1n9549);
not(notn9549,n1027);
and (s0n9549,notn9549,1'b0);
and (s1n9549,n1027,n9397);
and (n9550,n9549,n9551);
or (n9551,n9552,n9557,n9614);
and (n9552,n9553,n9556);
wire s0n9553,s1n9553,notn9553;
or (n9553,s0n9553,s1n9553);
not(notn9553,n979);
and (s0n9553,notn9553,1'b0);
and (s1n9553,n979,n9554);
xor (n9554,n9555,n9501);
xor (n9555,n9498,n9499);
wire s0n9556,s1n9556,notn9556;
or (n9556,s0n9556,s1n9556);
not(notn9556,n1027);
and (s0n9556,notn9556,1'b0);
and (s1n9556,n1027,n9547);
and (n9557,n9556,n9558);
or (n9558,n9559,n9564,n9613);
and (n9559,n9560,n9563);
wire s0n9560,s1n9560,notn9560;
or (n9560,s0n9560,s1n9560);
not(notn9560,n979);
and (s0n9560,notn9560,1'b0);
and (s1n9560,n979,n9561);
xor (n9561,n9562,n9507);
xor (n9562,n9503,n9504);
wire s0n9563,s1n9563,notn9563;
or (n9563,s0n9563,s1n9563);
not(notn9563,n1027);
and (s0n9563,notn9563,1'b0);
and (s1n9563,n1027,n9554);
and (n9564,n9563,n9565);
or (n9565,n9566,n9571,n9612);
and (n9566,n9567,n9570);
wire s0n9567,s1n9567,notn9567;
or (n9567,s0n9567,s1n9567);
not(notn9567,n979);
and (s0n9567,notn9567,1'b0);
and (s1n9567,n979,n9568);
xor (n9568,n9569,n9513);
xor (n9569,n9509,n9510);
wire s0n9570,s1n9570,notn9570;
or (n9570,s0n9570,s1n9570);
not(notn9570,n1027);
and (s0n9570,notn9570,1'b0);
and (s1n9570,n1027,n9561);
and (n9571,n9570,n9572);
or (n9572,n9573,n9578,n9611);
and (n9573,n9574,n9577);
wire s0n9574,s1n9574,notn9574;
or (n9574,s0n9574,s1n9574);
not(notn9574,n979);
and (s0n9574,notn9574,1'b0);
and (s1n9574,n979,n9575);
xor (n9575,n9576,n9519);
xor (n9576,n9515,n9516);
wire s0n9577,s1n9577,notn9577;
or (n9577,s0n9577,s1n9577);
not(notn9577,n1027);
and (s0n9577,notn9577,1'b0);
and (s1n9577,n1027,n9568);
and (n9578,n9577,n9579);
or (n9579,n9580,n9585,n9610);
and (n9580,n9581,n9584);
wire s0n9581,s1n9581,notn9581;
or (n9581,s0n9581,s1n9581);
not(notn9581,n979);
and (s0n9581,notn9581,1'b0);
and (s1n9581,n979,n9582);
xor (n9582,n9583,n9525);
xor (n9583,n9521,n9522);
wire s0n9584,s1n9584,notn9584;
or (n9584,s0n9584,s1n9584);
not(notn9584,n1027);
and (s0n9584,notn9584,1'b0);
and (s1n9584,n1027,n9575);
and (n9585,n9584,n9586);
or (n9586,n9587,n9592,n9609);
and (n9587,n9588,n9591);
wire s0n9588,s1n9588,notn9588;
or (n9588,s0n9588,s1n9588);
not(notn9588,n979);
and (s0n9588,notn9588,1'b0);
and (s1n9588,n979,n9589);
xor (n9589,n9590,n9531);
xor (n9590,n9527,n9528);
wire s0n9591,s1n9591,notn9591;
or (n9591,s0n9591,s1n9591);
not(notn9591,n1027);
and (s0n9591,notn9591,1'b0);
and (s1n9591,n1027,n9582);
and (n9592,n9591,n9593);
or (n9593,n9594,n9598,n9600);
and (n9594,n9595,n9597);
wire s0n9595,s1n9595,notn9595;
or (n9595,s0n9595,s1n9595);
not(notn9595,n979);
and (s0n9595,notn9595,1'b0);
and (s1n9595,n979,n9596);
xor (n9596,n9532,n9533);
wire s0n9597,s1n9597,notn9597;
or (n9597,s0n9597,s1n9597);
not(notn9597,n1027);
and (s0n9597,notn9597,1'b0);
and (s1n9597,n1027,n9589);
and (n9598,n9597,n9599);
or (n9599,n9600,n9604,n9605);
and (n9600,n9601,n9603);
wire s0n9601,s1n9601,notn9601;
or (n9601,s0n9601,s1n9601);
not(notn9601,n979);
and (s0n9601,notn9601,1'b0);
and (s1n9601,n979,n9602);
xor (n9602,n9482,n9490);
wire s0n9603,s1n9603,notn9603;
or (n9603,s0n9603,s1n9603);
not(notn9603,n1027);
and (s0n9603,notn9603,1'b0);
and (s1n9603,n1027,n9596);
and (n9604,n9603,n9605);
and (n9605,n9606,n9608);
wire s0n9606,s1n9606,notn9606;
or (n9606,s0n9606,s1n9606);
not(notn9606,n979);
and (s0n9606,notn9606,1'b0);
and (s1n9606,n979,n9607);
wire s0n9607,s1n9607,notn9607;
or (n9607,s0n9607,s1n9607);
not(notn9607,n699);
and (s0n9607,notn9607,1'b0);
and (s1n9607,n699,n9483);
wire s0n9608,s1n9608,notn9608;
or (n9608,s0n9608,s1n9608);
not(notn9608,n1027);
and (s0n9608,notn9608,1'b0);
and (s1n9608,n1027,n9602);
and (n9609,n9588,n9593);
and (n9610,n9581,n9586);
and (n9611,n9574,n9579);
and (n9612,n9567,n9572);
and (n9613,n9560,n9565);
and (n9614,n9553,n9558);
and (n9615,n9546,n9551);
and (n9616,n9542,n9617);
or (n9617,n9618,n9621,n9682);
and (n9618,n9619,n9620);
wire s0n9619,s1n9619,notn9619;
or (n9619,s0n9619,s1n9619);
not(notn9619,n930);
and (s0n9619,notn9619,1'b0);
and (s1n9619,n930,n9547);
xor (n9620,n9543,n9544);
and (n9621,n9620,n9622);
or (n9622,n9623,n9627,n9681);
and (n9623,n9624,n9625);
wire s0n9624,s1n9624,notn9624;
or (n9624,s0n9624,s1n9624);
not(notn9624,n930);
and (s0n9624,notn9624,1'b0);
and (s1n9624,n930,n9554);
xor (n9625,n9626,n9551);
xor (n9626,n9546,n9549);
and (n9627,n9625,n9628);
or (n9628,n9629,n9633,n9680);
and (n9629,n9630,n9631);
wire s0n9630,s1n9630,notn9630;
or (n9630,s0n9630,s1n9630);
not(notn9630,n930);
and (s0n9630,notn9630,1'b0);
and (s1n9630,n930,n9561);
xor (n9631,n9632,n9558);
xor (n9632,n9553,n9556);
and (n9633,n9631,n9634);
or (n9634,n9635,n9639,n9679);
and (n9635,n9636,n9637);
wire s0n9636,s1n9636,notn9636;
or (n9636,s0n9636,s1n9636);
not(notn9636,n930);
and (s0n9636,notn9636,1'b0);
and (s1n9636,n930,n9568);
xor (n9637,n9638,n9565);
xor (n9638,n9560,n9563);
and (n9639,n9637,n9640);
or (n9640,n9641,n9645,n9678);
and (n9641,n9642,n9643);
wire s0n9642,s1n9642,notn9642;
or (n9642,s0n9642,s1n9642);
not(notn9642,n930);
and (s0n9642,notn9642,1'b0);
and (s1n9642,n930,n9575);
xor (n9643,n9644,n9572);
xor (n9644,n9567,n9570);
and (n9645,n9643,n9646);
or (n9646,n9647,n9651,n9677);
and (n9647,n9648,n9649);
wire s0n9648,s1n9648,notn9648;
or (n9648,s0n9648,s1n9648);
not(notn9648,n930);
and (s0n9648,notn9648,1'b0);
and (s1n9648,n930,n9582);
xor (n9649,n9650,n9579);
xor (n9650,n9574,n9577);
and (n9651,n9649,n9652);
or (n9652,n9653,n9657,n9676);
and (n9653,n9654,n9655);
wire s0n9654,s1n9654,notn9654;
or (n9654,s0n9654,s1n9654);
not(notn9654,n930);
and (s0n9654,notn9654,1'b0);
and (s1n9654,n930,n9589);
xor (n9655,n9656,n9586);
xor (n9656,n9581,n9584);
and (n9657,n9655,n9658);
or (n9658,n9659,n9663,n9675);
and (n9659,n9660,n9661);
wire s0n9660,s1n9660,notn9660;
or (n9660,s0n9660,s1n9660);
not(notn9660,n930);
and (s0n9660,notn9660,1'b0);
and (s1n9660,n930,n9596);
xor (n9661,n9662,n9593);
xor (n9662,n9588,n9591);
and (n9663,n9661,n9664);
or (n9664,n9665,n9669,n9674);
and (n9665,n9666,n9667);
wire s0n9666,s1n9666,notn9666;
or (n9666,s0n9666,s1n9666);
not(notn9666,n930);
and (s0n9666,notn9666,1'b0);
and (s1n9666,n930,n9602);
xor (n9667,n9668,n9599);
xor (n9668,n9595,n9597);
and (n9669,n9667,n9670);
and (n9670,n9671,n9672);
wire s0n9671,s1n9671,notn9671;
or (n9671,s0n9671,s1n9671);
not(notn9671,n930);
and (s0n9671,notn9671,1'b0);
and (s1n9671,n930,n9607);
xor (n9672,n9673,n9605);
xor (n9673,n9601,n9603);
and (n9674,n9666,n9670);
and (n9675,n9660,n9664);
and (n9676,n9654,n9658);
and (n9677,n9648,n9652);
and (n9678,n9642,n9646);
and (n9679,n9636,n9640);
and (n9680,n9630,n9634);
and (n9681,n9624,n9628);
and (n9682,n9619,n9622);
and (n9683,n9396,n9617);
or (n9684,n9685,n9690,n9778);
and (n9685,n9686,n9688);
xor (n9686,n9687,n9327);
xor (n9687,n9083,n9259);
xor (n9688,n9689,n9617);
xor (n9689,n9396,n9542);
and (n9690,n9688,n9691);
or (n9691,n9692,n9697,n9777);
and (n9692,n9693,n9695);
xor (n9693,n9694,n9332);
xor (n9694,n9329,n9330);
xor (n9695,n9696,n9622);
xor (n9696,n9619,n9620);
and (n9697,n9695,n9698);
or (n9698,n9699,n9704,n9776);
and (n9699,n9700,n9702);
xor (n9700,n9701,n9338);
xor (n9701,n9334,n9335);
xor (n9702,n9703,n9628);
xor (n9703,n9624,n9625);
and (n9704,n9702,n9705);
or (n9705,n9706,n9711,n9775);
and (n9706,n9707,n9709);
xor (n9707,n9708,n9344);
xor (n9708,n9340,n9341);
xor (n9709,n9710,n9634);
xor (n9710,n9630,n9631);
and (n9711,n9709,n9712);
or (n9712,n9713,n9718,n9774);
and (n9713,n9714,n9716);
xor (n9714,n9715,n9350);
xor (n9715,n9346,n9347);
xor (n9716,n9717,n9640);
xor (n9717,n9636,n9637);
and (n9718,n9716,n9719);
or (n9719,n9720,n9725,n9773);
and (n9720,n9721,n9723);
xor (n9721,n9722,n9356);
xor (n9722,n9352,n9353);
xor (n9723,n9724,n9646);
xor (n9724,n9642,n9643);
and (n9725,n9723,n9726);
or (n9726,n9727,n9732,n9772);
and (n9727,n9728,n9730);
xor (n9728,n9729,n9362);
xor (n9729,n9358,n9359);
xor (n9730,n9731,n9652);
xor (n9731,n9648,n9649);
and (n9732,n9730,n9733);
or (n9733,n9734,n9739,n9771);
and (n9734,n9735,n9737);
xor (n9735,n9736,n9368);
xor (n9736,n9364,n9365);
xor (n9737,n9738,n9658);
xor (n9738,n9654,n9655);
and (n9739,n9737,n9740);
or (n9740,n9741,n9746,n9770);
and (n9741,n9742,n9744);
xor (n9742,n9743,n9374);
xor (n9743,n9370,n9371);
xor (n9744,n9745,n9664);
xor (n9745,n9660,n9661);
and (n9746,n9744,n9747);
or (n9747,n9748,n9753,n9769);
and (n9748,n9749,n9751);
xor (n9749,n9750,n9380);
xor (n9750,n9376,n9377);
xor (n9751,n9752,n9670);
xor (n9752,n9666,n9667);
and (n9753,n9751,n9754);
or (n9754,n9755,n9758,n9768);
and (n9755,n9756,n9757);
xor (n9756,n9381,n9382);
xor (n9757,n9671,n9672);
and (n9758,n9757,n9759);
or (n9759,n9760,n9763,n9767);
and (n9760,n9761,n9762);
xor (n9761,n9316,n9318);
xor (n9762,n9606,n9608);
and (n9763,n9762,n9764);
and (n9764,n9765,n9766);
wire s0n9765,s1n9765,notn9765;
or (n9765,s0n9765,s1n9765);
not(notn9765,n1027);
and (s0n9765,notn9765,1'b0);
and (s1n9765,n1027,n9317);
wire s0n9766,s1n9766,notn9766;
or (n9766,s0n9766,s1n9766);
not(notn9766,n1027);
and (s0n9766,notn9766,1'b0);
and (s1n9766,n1027,n9607);
and (n9767,n9761,n9764);
and (n9768,n9756,n9759);
and (n9769,n9749,n9754);
and (n9770,n9742,n9747);
and (n9771,n9735,n9740);
and (n9772,n9728,n9733);
and (n9773,n9721,n9726);
and (n9774,n9714,n9719);
and (n9775,n9707,n9712);
and (n9776,n9700,n9705);
and (n9777,n9693,n9698);
and (n9778,n9686,n9691);
or (n9779,n9780,n9785,n9876);
and (n9780,n9781,n9783);
xor (n9781,n9782,n8994);
xor (n9782,n8989,n8991);
xor (n9783,n9784,n9691);
xor (n9784,n9686,n9688);
and (n9785,n9783,n9786);
or (n9786,n9787,n9792,n9875);
and (n9787,n9788,n9790);
xor (n9788,n9789,n9001);
xor (n9789,n8996,n8998);
xor (n9790,n9791,n9698);
xor (n9791,n9693,n9695);
and (n9792,n9790,n9793);
or (n9793,n9794,n9799,n9874);
and (n9794,n9795,n9797);
xor (n9795,n9796,n9008);
xor (n9796,n9003,n9005);
xor (n9797,n9798,n9705);
xor (n9798,n9700,n9702);
and (n9799,n9797,n9800);
or (n9800,n9801,n9806,n9873);
and (n9801,n9802,n9804);
xor (n9802,n9803,n9015);
xor (n9803,n9010,n9012);
xor (n9804,n9805,n9712);
xor (n9805,n9707,n9709);
and (n9806,n9804,n9807);
or (n9807,n9808,n9813,n9872);
and (n9808,n9809,n9811);
xor (n9809,n9810,n9022);
xor (n9810,n9017,n9019);
xor (n9811,n9812,n9719);
xor (n9812,n9714,n9716);
and (n9813,n9811,n9814);
or (n9814,n9815,n9820,n9871);
and (n9815,n9816,n9818);
xor (n9816,n9817,n9029);
xor (n9817,n9024,n9026);
xor (n9818,n9819,n9726);
xor (n9819,n9721,n9723);
and (n9820,n9818,n9821);
or (n9821,n9822,n9827,n9870);
and (n9822,n9823,n9825);
xor (n9823,n9824,n9036);
xor (n9824,n9031,n9033);
xor (n9825,n9826,n9733);
xor (n9826,n9728,n9730);
and (n9827,n9825,n9828);
or (n9828,n9829,n9834,n9869);
and (n9829,n9830,n9832);
xor (n9830,n9831,n9043);
xor (n9831,n9038,n9040);
xor (n9832,n9833,n9740);
xor (n9833,n9735,n9737);
and (n9834,n9832,n9835);
or (n9835,n9836,n9841,n9868);
and (n9836,n9837,n9839);
xor (n9837,n9838,n9050);
xor (n9838,n9045,n9047);
xor (n9839,n9840,n9747);
xor (n9840,n9742,n9744);
and (n9841,n9839,n9842);
or (n9842,n9843,n9848,n9867);
and (n9843,n9844,n9846);
xor (n9844,n9845,n9057);
xor (n9845,n9052,n9054);
xor (n9846,n9847,n9754);
xor (n9847,n9749,n9751);
and (n9848,n9846,n9849);
or (n9849,n9850,n9855,n9866);
and (n9850,n9851,n9853);
xor (n9851,n9852,n9062);
xor (n9852,n9059,n9060);
xor (n9853,n9854,n9759);
xor (n9854,n9756,n9757);
and (n9855,n9853,n9856);
or (n9856,n9857,n9862,n9865);
and (n9857,n9858,n9860);
xor (n9858,n9859,n2563);
xor (n9859,n9064,n9065);
xor (n9860,n9861,n9764);
xor (n9861,n9761,n9762);
and (n9862,n9860,n9863);
and (n9863,n2664,n9864);
xor (n9864,n9765,n9766);
and (n9865,n9858,n9863);
and (n9866,n9851,n9856);
and (n9867,n9844,n9849);
and (n9868,n9837,n9842);
and (n9869,n9830,n9835);
and (n9870,n9823,n9828);
and (n9871,n9816,n9821);
and (n9872,n9809,n9814);
and (n9873,n9802,n9807);
and (n9874,n9795,n9800);
and (n9875,n9788,n9793);
and (n9876,n9781,n9786);
and (n9877,n9878,n9880);
xor (n9878,n9879,n9786);
xor (n9879,n9781,n9783);
and (n9880,n9881,n9883);
xor (n9881,n9882,n9793);
xor (n9882,n9788,n9790);
and (n9883,n9884,n9886);
xor (n9884,n9885,n9800);
xor (n9885,n9795,n9797);
and (n9886,n9887,n9889);
xor (n9887,n9888,n9807);
xor (n9888,n9802,n9804);
and (n9889,n9890,n9892);
xor (n9890,n9891,n9814);
xor (n9891,n9809,n9811);
and (n9892,n9893,n9895);
xor (n9893,n9894,n9821);
xor (n9894,n9816,n9818);
and (n9895,n9896,n9898);
xor (n9896,n9897,n9828);
xor (n9897,n9823,n9825);
xor (n9898,n9899,n9835);
xor (n9899,n9830,n9832);
wire s0n9900,s1n9900,notn9900;
or (n9900,s0n9900,s1n9900);
not(notn9900,n2755);
and (s0n9900,notn9900,n9901);
and (s1n9900,n2755,n9904);
wire s0n9901,s1n9901,notn9901;
or (n9901,s0n9901,s1n9901);
not(notn9901,n2705);
and (s0n9901,notn9901,1'b0);
and (s1n9901,n2705,n9902);
wire s0n9902,s1n9902,notn9902;
or (n9902,s0n9902,s1n9902);
not(notn9902,n577);
and (s0n9902,notn9902,n1690);
and (s1n9902,n577,n9903);
wire s0n9903,s1n9903,notn9903;
or (n9903,s0n9903,s1n9903);
not(notn9903,n2704);
and (s0n9903,notn9903,1'b0);
and (s1n9903,n2704,n1689);
or (n9904,1'b0,n9905,n9911,n9917,n9923);
and (n9905,n9906,n2718);
or (n9906,1'b0,n9907,n9908,n9909,n9910);
and (n9907,n6831,n556);
and (n9908,n6835,n567);
and (n9909,n6838,n571);
and (n9910,n6841,n573);
and (n9911,n9912,n2730);
or (n9912,1'b0,n9913,n9914,n9915,n9916);
and (n9913,n6846,n556);
and (n9914,n6849,n567);
and (n9915,n6852,n571);
and (n9916,n6855,n573);
and (n9917,n9918,n2742);
or (n9918,1'b0,n9919,n9920,n9921,n9922);
and (n9919,n5012,n556);
and (n9920,n5027,n567);
and (n9921,n5032,n571);
and (n9922,n5037,n573);
and (n9923,n9924,n2752);
or (n9924,1'b0,n9925,n9926,n9927,n9928);
and (n9925,n5044,n556);
and (n9926,n5047,n567);
and (n9927,n5050,n571);
and (n9928,n5053,n573);
or (n9929,n9930,n9933,n9900);
and (n9930,n9931,n8688);
wire s0n9931,s1n9931,notn9931;
or (n9931,s0n9931,s1n9931);
not(notn9931,n4969);
and (s0n9931,notn9931,1'b0);
and (s1n9931,n4969,n9932);
or (n9932,1'b0,n9933,n13857,n13859,n13860,n13861);
and (n9933,n9934,n2907);
wire s0n9934,s1n9934,notn9934;
or (n9934,s0n9934,s1n9934);
not(notn9934,n2902);
and (s0n9934,notn9934,1'b0);
and (s1n9934,n2902,n9935);
xor (n9935,n9936,n13835);
or (n9936,n9937,n13061,n13834);
and (n9937,n9938,n11732);
or (n9938,1'b0,n9939,n9942,n9945,n11671);
and (n9939,n9940,n2893);
wire s0n9940,s1n9940,notn9940;
or (n9940,s0n9940,s1n9940);
not(notn9940,n2891);
and (s0n9940,notn9940,1'b0);
and (s1n9940,n2891,n9941);
and (n9942,n9943,n2907);
wire s0n9943,s1n9943,notn9943;
or (n9943,s0n9943,s1n9943);
not(notn9943,n2902);
and (s0n9943,notn9943,1'b0);
and (s1n9943,n2902,n9944);
and (n9945,n9946,n4883);
wire s0n9946,s1n9946,notn9946;
or (n9946,s0n9946,s1n9946);
not(notn9946,n11666);
and (s0n9946,notn9946,n9947);
and (s1n9946,n11666,1'b0);
wire s0n9947,s1n9947,notn9947;
or (n9947,s0n9947,s1n9947);
not(notn9947,n11661);
and (s0n9947,notn9947,n9948);
and (s1n9947,n11661,1'b1);
wire s0n9948,s1n9948,notn9948;
or (n9948,s0n9948,s1n9948);
not(notn9948,n4861);
and (s0n9948,notn9948,1'b0);
and (s1n9948,n4861,n9949);
xor (n9949,n9950,n11638);
xor (n9950,n9951,n11585);
xor (n9951,n9952,n11147);
xor (n9952,n9953,n11145);
xor (n9953,n9954,n11115);
not (n9954,n9955);
or (n9955,n9956,n10529);
or (n9956,n9957,n10026,n10528);
and (n9957,n9958,n9999);
or (n9958,1'b0,n9959,n9969,n9979,n9989);
and (n9959,n9960,n2718);
or (n9960,1'b0,n9961,n9963,n9965,n9967);
and (n9961,n9962,n2932);
wire s0n9962,s1n9962,notn9962;
or (n9962,s0n9962,s1n9962);
not(notn9962,n2929);
and (s0n9962,notn9962,n6831);
and (s1n9962,n2929,n5088);
and (n9963,n9964,n2955);
wire s0n9964,s1n9964,notn9964;
or (n9964,s0n9964,s1n9964);
not(notn9964,n2929);
and (s0n9964,notn9964,n6835);
and (s1n9964,n2929,n5092);
and (n9965,n9966,n2963);
wire s0n9966,s1n9966,notn9966;
or (n9966,s0n9966,s1n9966);
not(notn9966,n2929);
and (s0n9966,notn9966,n6838);
and (s1n9966,n2929,n5095);
and (n9967,n9968,n2972);
wire s0n9968,s1n9968,notn9968;
or (n9968,s0n9968,s1n9968);
not(notn9968,n2929);
and (s0n9968,notn9968,n6841);
and (s1n9968,n2929,n5098);
and (n9969,n9970,n2730);
or (n9970,1'b0,n9971,n9973,n9975,n9977);
and (n9971,n9972,n2932);
wire s0n9972,s1n9972,notn9972;
or (n9972,s0n9972,s1n9972);
not(notn9972,n2929);
and (s0n9972,notn9972,n6846);
and (s1n9972,n2929,n5103);
and (n9973,n9974,n2955);
wire s0n9974,s1n9974,notn9974;
or (n9974,s0n9974,s1n9974);
not(notn9974,n2929);
and (s0n9974,notn9974,n6849);
and (s1n9974,n2929,n5106);
and (n9975,n9976,n2963);
wire s0n9976,s1n9976,notn9976;
or (n9976,s0n9976,s1n9976);
not(notn9976,n2929);
and (s0n9976,notn9976,n6852);
and (s1n9976,n2929,n5109);
and (n9977,n9978,n2972);
wire s0n9978,s1n9978,notn9978;
or (n9978,s0n9978,s1n9978);
not(notn9978,n2929);
and (s0n9978,notn9978,n6855);
and (s1n9978,n2929,n5112);
and (n9979,n9980,n2742);
or (n9980,1'b0,n9981,n9983,n9985,n9987);
and (n9981,n9982,n2932);
wire s0n9982,s1n9982,notn9982;
or (n9982,s0n9982,s1n9982);
not(notn9982,n2929);
and (s0n9982,notn9982,n5012);
and (s1n9982,n2929,n5117);
and (n9983,n9984,n2955);
wire s0n9984,s1n9984,notn9984;
or (n9984,s0n9984,s1n9984);
not(notn9984,n2929);
and (s0n9984,notn9984,n5027);
and (s1n9984,n2929,n5121);
and (n9985,n9986,n2963);
wire s0n9986,s1n9986,notn9986;
or (n9986,s0n9986,s1n9986);
not(notn9986,n2929);
and (s0n9986,notn9986,n5032);
and (s1n9986,n2929,n5124);
and (n9987,n9988,n2972);
wire s0n9988,s1n9988,notn9988;
or (n9988,s0n9988,s1n9988);
not(notn9988,n2929);
and (s0n9988,notn9988,n5037);
and (s1n9988,n2929,n5127);
and (n9989,n9990,n2752);
or (n9990,1'b0,n9991,n9993,n9995,n9997);
and (n9991,n9992,n2932);
wire s0n9992,s1n9992,notn9992;
or (n9992,s0n9992,s1n9992);
not(notn9992,n2929);
and (s0n9992,notn9992,n5044);
and (s1n9992,n2929,n5132);
and (n9993,n9994,n2955);
wire s0n9994,s1n9994,notn9994;
or (n9994,s0n9994,s1n9994);
not(notn9994,n2929);
and (s0n9994,notn9994,n5047);
and (s1n9994,n2929,n5135);
and (n9995,n9996,n2963);
wire s0n9996,s1n9996,notn9996;
or (n9996,s0n9996,s1n9996);
not(notn9996,n2929);
and (s0n9996,notn9996,n5050);
and (s1n9996,n2929,n5138);
and (n9997,n9998,n2972);
wire s0n9998,s1n9998,notn9998;
or (n9998,s0n9998,s1n9998);
not(notn9998,n2929);
and (s0n9998,notn9998,n5053);
and (s1n9998,n2929,n5141);
or (n9999,1'b0,n10000,n10007,n10013,n10020);
and (n10000,n10001,n2718);
or (n10001,1'b0,n10002,n10004,n10005,n10006);
and (n10002,n10003,n2932);
wire s0n10003,s1n10003,notn10003;
or (n10003,s0n10003,s1n10003);
not(notn10003,n2929);
and (s0n10003,notn10003,n6832);
and (s1n10003,n2929,n5089);
and (n10004,n9962,n2955);
and (n10005,n9964,n2963);
and (n10006,n9966,n2972);
and (n10007,n10008,n2730);
or (n10008,1'b0,n10009,n10010,n10011,n10012);
and (n10009,n9968,n2932);
and (n10010,n9972,n2955);
and (n10011,n9974,n2963);
and (n10012,n9976,n2972);
and (n10013,n10014,n2742);
or (n10014,1'b0,n10015,n10017,n10018,n10019);
and (n10015,n10016,n2932);
wire s0n10016,s1n10016,notn10016;
or (n10016,s0n10016,s1n10016);
not(notn10016,n2929);
and (s0n10016,notn10016,n5013);
and (s1n10016,n2929,n5118);
and (n10017,n9982,n2955);
and (n10018,n9984,n2963);
and (n10019,n9986,n2972);
and (n10020,n10021,n2752);
or (n10021,1'b0,n10022,n10023,n10024,n10025);
and (n10022,n9988,n2932);
and (n10023,n9992,n2955);
and (n10024,n9994,n2963);
and (n10025,n9996,n2972);
and (n10026,n9999,n10027);
or (n10027,n10028,n10097,n10527);
and (n10028,n10029,n10070);
or (n10029,1'b0,n10030,n10040,n10050,n10060);
and (n10030,n10031,n2718);
or (n10031,1'b0,n10032,n10034,n10036,n10038);
and (n10032,n10033,n2932);
wire s0n10033,s1n10033,notn10033;
or (n10033,s0n10033,s1n10033);
not(notn10033,n2929);
and (s0n10033,notn10033,n6900);
and (s1n10033,n2929,n5211);
and (n10034,n10035,n2955);
wire s0n10035,s1n10035,notn10035;
or (n10035,s0n10035,s1n10035);
not(notn10035,n2929);
and (s0n10035,notn10035,n6904);
and (s1n10035,n2929,n5215);
and (n10036,n10037,n2963);
wire s0n10037,s1n10037,notn10037;
or (n10037,s0n10037,s1n10037);
not(notn10037,n2929);
and (s0n10037,notn10037,n6907);
and (s1n10037,n2929,n5218);
and (n10038,n10039,n2972);
wire s0n10039,s1n10039,notn10039;
or (n10039,s0n10039,s1n10039);
not(notn10039,n2929);
and (s0n10039,notn10039,n6910);
and (s1n10039,n2929,n5221);
and (n10040,n10041,n2730);
or (n10041,1'b0,n10042,n10044,n10046,n10048);
and (n10042,n10043,n2932);
wire s0n10043,s1n10043,notn10043;
or (n10043,s0n10043,s1n10043);
not(notn10043,n2929);
and (s0n10043,notn10043,n6915);
and (s1n10043,n2929,n5226);
and (n10044,n10045,n2955);
wire s0n10045,s1n10045,notn10045;
or (n10045,s0n10045,s1n10045);
not(notn10045,n2929);
and (s0n10045,notn10045,n6918);
and (s1n10045,n2929,n5229);
and (n10046,n10047,n2963);
wire s0n10047,s1n10047,notn10047;
or (n10047,s0n10047,s1n10047);
not(notn10047,n2929);
and (s0n10047,notn10047,n6921);
and (s1n10047,n2929,n5232);
and (n10048,n10049,n2972);
wire s0n10049,s1n10049,notn10049;
or (n10049,s0n10049,s1n10049);
not(notn10049,n2929);
and (s0n10049,notn10049,n6924);
and (s1n10049,n2929,n5235);
and (n10050,n10051,n2742);
or (n10051,1'b0,n10052,n10054,n10056,n10058);
and (n10052,n10053,n2932);
wire s0n10053,s1n10053,notn10053;
or (n10053,s0n10053,s1n10053);
not(notn10053,n2929);
and (s0n10053,notn10053,n5152);
and (s1n10053,n2929,n5240);
and (n10054,n10055,n2955);
wire s0n10055,s1n10055,notn10055;
or (n10055,s0n10055,s1n10055);
not(notn10055,n2929);
and (s0n10055,notn10055,n5156);
and (s1n10055,n2929,n5244);
and (n10056,n10057,n2963);
wire s0n10057,s1n10057,notn10057;
or (n10057,s0n10057,s1n10057);
not(notn10057,n2929);
and (s0n10057,notn10057,n5159);
and (s1n10057,n2929,n5247);
and (n10058,n10059,n2972);
wire s0n10059,s1n10059,notn10059;
or (n10059,s0n10059,s1n10059);
not(notn10059,n2929);
and (s0n10059,notn10059,n5162);
and (s1n10059,n2929,n5250);
and (n10060,n10061,n2752);
or (n10061,1'b0,n10062,n10064,n10066,n10068);
and (n10062,n10063,n2932);
wire s0n10063,s1n10063,notn10063;
or (n10063,s0n10063,s1n10063);
not(notn10063,n2929);
and (s0n10063,notn10063,n5167);
and (s1n10063,n2929,n5255);
and (n10064,n10065,n2955);
wire s0n10065,s1n10065,notn10065;
or (n10065,s0n10065,s1n10065);
not(notn10065,n2929);
and (s0n10065,notn10065,n5170);
and (s1n10065,n2929,n5258);
and (n10066,n10067,n2963);
wire s0n10067,s1n10067,notn10067;
or (n10067,s0n10067,s1n10067);
not(notn10067,n2929);
and (s0n10067,notn10067,n5173);
and (s1n10067,n2929,n5261);
and (n10068,n10069,n2972);
wire s0n10069,s1n10069,notn10069;
or (n10069,s0n10069,s1n10069);
not(notn10069,n2929);
and (s0n10069,notn10069,n5176);
and (s1n10069,n2929,n5264);
or (n10070,1'b0,n10071,n10078,n10084,n10091);
and (n10071,n10072,n2718);
or (n10072,1'b0,n10073,n10075,n10076,n10077);
and (n10073,n10074,n2932);
wire s0n10074,s1n10074,notn10074;
or (n10074,s0n10074,s1n10074);
not(notn10074,n2929);
and (s0n10074,notn10074,n6901);
and (s1n10074,n2929,n5212);
and (n10075,n10033,n2955);
and (n10076,n10035,n2963);
and (n10077,n10037,n2972);
and (n10078,n10079,n2730);
or (n10079,1'b0,n10080,n10081,n10082,n10083);
and (n10080,n10039,n2932);
and (n10081,n10043,n2955);
and (n10082,n10045,n2963);
and (n10083,n10047,n2972);
and (n10084,n10085,n2742);
or (n10085,1'b0,n10086,n10088,n10089,n10090);
and (n10086,n10087,n2932);
wire s0n10087,s1n10087,notn10087;
or (n10087,s0n10087,s1n10087);
not(notn10087,n2929);
and (s0n10087,notn10087,n5153);
and (s1n10087,n2929,n5241);
and (n10088,n10053,n2955);
and (n10089,n10055,n2963);
and (n10090,n10057,n2972);
and (n10091,n10092,n2752);
or (n10092,1'b0,n10093,n10094,n10095,n10096);
and (n10093,n10059,n2932);
and (n10094,n10063,n2955);
and (n10095,n10065,n2963);
and (n10096,n10067,n2972);
and (n10097,n10070,n10098);
or (n10098,n10099,n10168,n10526);
and (n10099,n10100,n10141);
or (n10100,1'b0,n10101,n10111,n10121,n10131);
and (n10101,n10102,n2718);
or (n10102,1'b0,n10103,n10105,n10107,n10109);
and (n10103,n10104,n2932);
wire s0n10104,s1n10104,notn10104;
or (n10104,s0n10104,s1n10104);
not(notn10104,n2929);
and (s0n10104,notn10104,n6969);
and (s1n10104,n2929,n5334);
and (n10105,n10106,n2955);
wire s0n10106,s1n10106,notn10106;
or (n10106,s0n10106,s1n10106);
not(notn10106,n2929);
and (s0n10106,notn10106,n6973);
and (s1n10106,n2929,n5338);
and (n10107,n10108,n2963);
wire s0n10108,s1n10108,notn10108;
or (n10108,s0n10108,s1n10108);
not(notn10108,n2929);
and (s0n10108,notn10108,n6976);
and (s1n10108,n2929,n5341);
and (n10109,n10110,n2972);
wire s0n10110,s1n10110,notn10110;
or (n10110,s0n10110,s1n10110);
not(notn10110,n2929);
and (s0n10110,notn10110,n6979);
and (s1n10110,n2929,n5344);
and (n10111,n10112,n2730);
or (n10112,1'b0,n10113,n10115,n10117,n10119);
and (n10113,n10114,n2932);
wire s0n10114,s1n10114,notn10114;
or (n10114,s0n10114,s1n10114);
not(notn10114,n2929);
and (s0n10114,notn10114,n6984);
and (s1n10114,n2929,n5349);
and (n10115,n10116,n2955);
wire s0n10116,s1n10116,notn10116;
or (n10116,s0n10116,s1n10116);
not(notn10116,n2929);
and (s0n10116,notn10116,n6987);
and (s1n10116,n2929,n5352);
and (n10117,n10118,n2963);
wire s0n10118,s1n10118,notn10118;
or (n10118,s0n10118,s1n10118);
not(notn10118,n2929);
and (s0n10118,notn10118,n6990);
and (s1n10118,n2929,n5355);
and (n10119,n10120,n2972);
wire s0n10120,s1n10120,notn10120;
or (n10120,s0n10120,s1n10120);
not(notn10120,n2929);
and (s0n10120,notn10120,n6993);
and (s1n10120,n2929,n5358);
and (n10121,n10122,n2742);
or (n10122,1'b0,n10123,n10125,n10127,n10129);
and (n10123,n10124,n2932);
wire s0n10124,s1n10124,notn10124;
or (n10124,s0n10124,s1n10124);
not(notn10124,n2929);
and (s0n10124,notn10124,n5275);
and (s1n10124,n2929,n5363);
and (n10125,n10126,n2955);
wire s0n10126,s1n10126,notn10126;
or (n10126,s0n10126,s1n10126);
not(notn10126,n2929);
and (s0n10126,notn10126,n5279);
and (s1n10126,n2929,n5367);
and (n10127,n10128,n2963);
wire s0n10128,s1n10128,notn10128;
or (n10128,s0n10128,s1n10128);
not(notn10128,n2929);
and (s0n10128,notn10128,n5282);
and (s1n10128,n2929,n5370);
and (n10129,n10130,n2972);
wire s0n10130,s1n10130,notn10130;
or (n10130,s0n10130,s1n10130);
not(notn10130,n2929);
and (s0n10130,notn10130,n5285);
and (s1n10130,n2929,n5373);
and (n10131,n10132,n2752);
or (n10132,1'b0,n10133,n10135,n10137,n10139);
and (n10133,n10134,n2932);
wire s0n10134,s1n10134,notn10134;
or (n10134,s0n10134,s1n10134);
not(notn10134,n2929);
and (s0n10134,notn10134,n5290);
and (s1n10134,n2929,n5378);
and (n10135,n10136,n2955);
wire s0n10136,s1n10136,notn10136;
or (n10136,s0n10136,s1n10136);
not(notn10136,n2929);
and (s0n10136,notn10136,n5293);
and (s1n10136,n2929,n5381);
and (n10137,n10138,n2963);
wire s0n10138,s1n10138,notn10138;
or (n10138,s0n10138,s1n10138);
not(notn10138,n2929);
and (s0n10138,notn10138,n5296);
and (s1n10138,n2929,n5384);
and (n10139,n10140,n2972);
wire s0n10140,s1n10140,notn10140;
or (n10140,s0n10140,s1n10140);
not(notn10140,n2929);
and (s0n10140,notn10140,n5299);
and (s1n10140,n2929,n5387);
or (n10141,1'b0,n10142,n10149,n10155,n10162);
and (n10142,n10143,n2718);
or (n10143,1'b0,n10144,n10146,n10147,n10148);
and (n10144,n10145,n2932);
wire s0n10145,s1n10145,notn10145;
or (n10145,s0n10145,s1n10145);
not(notn10145,n2929);
and (s0n10145,notn10145,n6970);
and (s1n10145,n2929,n5335);
and (n10146,n10104,n2955);
and (n10147,n10106,n2963);
and (n10148,n10108,n2972);
and (n10149,n10150,n2730);
or (n10150,1'b0,n10151,n10152,n10153,n10154);
and (n10151,n10110,n2932);
and (n10152,n10114,n2955);
and (n10153,n10116,n2963);
and (n10154,n10118,n2972);
and (n10155,n10156,n2742);
or (n10156,1'b0,n10157,n10159,n10160,n10161);
and (n10157,n10158,n2932);
wire s0n10158,s1n10158,notn10158;
or (n10158,s0n10158,s1n10158);
not(notn10158,n2929);
and (s0n10158,notn10158,n5276);
and (s1n10158,n2929,n5364);
and (n10159,n10124,n2955);
and (n10160,n10126,n2963);
and (n10161,n10128,n2972);
and (n10162,n10163,n2752);
or (n10163,1'b0,n10164,n10165,n10166,n10167);
and (n10164,n10130,n2932);
and (n10165,n10134,n2955);
and (n10166,n10136,n2963);
and (n10167,n10138,n2972);
and (n10168,n10141,n10169);
or (n10169,n10170,n10239,n10525);
and (n10170,n10171,n10212);
or (n10171,1'b0,n10172,n10182,n10192,n10202);
and (n10172,n10173,n2718);
or (n10173,1'b0,n10174,n10176,n10178,n10180);
and (n10174,n10175,n2932);
wire s0n10175,s1n10175,notn10175;
or (n10175,s0n10175,s1n10175);
not(notn10175,n2929);
and (s0n10175,notn10175,n7038);
and (s1n10175,n2929,n5457);
and (n10176,n10177,n2955);
wire s0n10177,s1n10177,notn10177;
or (n10177,s0n10177,s1n10177);
not(notn10177,n2929);
and (s0n10177,notn10177,n7042);
and (s1n10177,n2929,n5461);
and (n10178,n10179,n2963);
wire s0n10179,s1n10179,notn10179;
or (n10179,s0n10179,s1n10179);
not(notn10179,n2929);
and (s0n10179,notn10179,n7045);
and (s1n10179,n2929,n5464);
and (n10180,n10181,n2972);
wire s0n10181,s1n10181,notn10181;
or (n10181,s0n10181,s1n10181);
not(notn10181,n2929);
and (s0n10181,notn10181,n7048);
and (s1n10181,n2929,n5467);
and (n10182,n10183,n2730);
or (n10183,1'b0,n10184,n10186,n10188,n10190);
and (n10184,n10185,n2932);
wire s0n10185,s1n10185,notn10185;
or (n10185,s0n10185,s1n10185);
not(notn10185,n2929);
and (s0n10185,notn10185,n7053);
and (s1n10185,n2929,n5472);
and (n10186,n10187,n2955);
wire s0n10187,s1n10187,notn10187;
or (n10187,s0n10187,s1n10187);
not(notn10187,n2929);
and (s0n10187,notn10187,n7056);
and (s1n10187,n2929,n5475);
and (n10188,n10189,n2963);
wire s0n10189,s1n10189,notn10189;
or (n10189,s0n10189,s1n10189);
not(notn10189,n2929);
and (s0n10189,notn10189,n7059);
and (s1n10189,n2929,n5478);
and (n10190,n10191,n2972);
wire s0n10191,s1n10191,notn10191;
or (n10191,s0n10191,s1n10191);
not(notn10191,n2929);
and (s0n10191,notn10191,n7062);
and (s1n10191,n2929,n5481);
and (n10192,n10193,n2742);
or (n10193,1'b0,n10194,n10196,n10198,n10200);
and (n10194,n10195,n2932);
wire s0n10195,s1n10195,notn10195;
or (n10195,s0n10195,s1n10195);
not(notn10195,n2929);
and (s0n10195,notn10195,n5398);
and (s1n10195,n2929,n5486);
and (n10196,n10197,n2955);
wire s0n10197,s1n10197,notn10197;
or (n10197,s0n10197,s1n10197);
not(notn10197,n2929);
and (s0n10197,notn10197,n5402);
and (s1n10197,n2929,n5490);
and (n10198,n10199,n2963);
wire s0n10199,s1n10199,notn10199;
or (n10199,s0n10199,s1n10199);
not(notn10199,n2929);
and (s0n10199,notn10199,n5405);
and (s1n10199,n2929,n5493);
and (n10200,n10201,n2972);
wire s0n10201,s1n10201,notn10201;
or (n10201,s0n10201,s1n10201);
not(notn10201,n2929);
and (s0n10201,notn10201,n5408);
and (s1n10201,n2929,n5496);
and (n10202,n10203,n2752);
or (n10203,1'b0,n10204,n10206,n10208,n10210);
and (n10204,n10205,n2932);
wire s0n10205,s1n10205,notn10205;
or (n10205,s0n10205,s1n10205);
not(notn10205,n2929);
and (s0n10205,notn10205,n5413);
and (s1n10205,n2929,n5501);
and (n10206,n10207,n2955);
wire s0n10207,s1n10207,notn10207;
or (n10207,s0n10207,s1n10207);
not(notn10207,n2929);
and (s0n10207,notn10207,n5416);
and (s1n10207,n2929,n5504);
and (n10208,n10209,n2963);
wire s0n10209,s1n10209,notn10209;
or (n10209,s0n10209,s1n10209);
not(notn10209,n2929);
and (s0n10209,notn10209,n5419);
and (s1n10209,n2929,n5507);
and (n10210,n10211,n2972);
wire s0n10211,s1n10211,notn10211;
or (n10211,s0n10211,s1n10211);
not(notn10211,n2929);
and (s0n10211,notn10211,n5422);
and (s1n10211,n2929,n5510);
or (n10212,1'b0,n10213,n10220,n10226,n10233);
and (n10213,n10214,n2718);
or (n10214,1'b0,n10215,n10217,n10218,n10219);
and (n10215,n10216,n2932);
wire s0n10216,s1n10216,notn10216;
or (n10216,s0n10216,s1n10216);
not(notn10216,n2929);
and (s0n10216,notn10216,n7039);
and (s1n10216,n2929,n5458);
and (n10217,n10175,n2955);
and (n10218,n10177,n2963);
and (n10219,n10179,n2972);
and (n10220,n10221,n2730);
or (n10221,1'b0,n10222,n10223,n10224,n10225);
and (n10222,n10181,n2932);
and (n10223,n10185,n2955);
and (n10224,n10187,n2963);
and (n10225,n10189,n2972);
and (n10226,n10227,n2742);
or (n10227,1'b0,n10228,n10230,n10231,n10232);
and (n10228,n10229,n2932);
wire s0n10229,s1n10229,notn10229;
or (n10229,s0n10229,s1n10229);
not(notn10229,n2929);
and (s0n10229,notn10229,n5399);
and (s1n10229,n2929,n5487);
and (n10230,n10195,n2955);
and (n10231,n10197,n2963);
and (n10232,n10199,n2972);
and (n10233,n10234,n2752);
or (n10234,1'b0,n10235,n10236,n10237,n10238);
and (n10235,n10201,n2932);
and (n10236,n10205,n2955);
and (n10237,n10207,n2963);
and (n10238,n10209,n2972);
and (n10239,n10212,n10240);
or (n10240,n10241,n10310,n10524);
and (n10241,n10242,n10283);
or (n10242,1'b0,n10243,n10253,n10263,n10273);
and (n10243,n10244,n2718);
or (n10244,1'b0,n10245,n10247,n10249,n10251);
and (n10245,n10246,n2932);
wire s0n10246,s1n10246,notn10246;
or (n10246,s0n10246,s1n10246);
not(notn10246,n2929);
and (s0n10246,notn10246,n7107);
and (s1n10246,n2929,n5580);
and (n10247,n10248,n2955);
wire s0n10248,s1n10248,notn10248;
or (n10248,s0n10248,s1n10248);
not(notn10248,n2929);
and (s0n10248,notn10248,n7111);
and (s1n10248,n2929,n5584);
and (n10249,n10250,n2963);
wire s0n10250,s1n10250,notn10250;
or (n10250,s0n10250,s1n10250);
not(notn10250,n2929);
and (s0n10250,notn10250,n7114);
and (s1n10250,n2929,n5587);
and (n10251,n10252,n2972);
wire s0n10252,s1n10252,notn10252;
or (n10252,s0n10252,s1n10252);
not(notn10252,n2929);
and (s0n10252,notn10252,n7117);
and (s1n10252,n2929,n5590);
and (n10253,n10254,n2730);
or (n10254,1'b0,n10255,n10257,n10259,n10261);
and (n10255,n10256,n2932);
wire s0n10256,s1n10256,notn10256;
or (n10256,s0n10256,s1n10256);
not(notn10256,n2929);
and (s0n10256,notn10256,n7122);
and (s1n10256,n2929,n5595);
and (n10257,n10258,n2955);
wire s0n10258,s1n10258,notn10258;
or (n10258,s0n10258,s1n10258);
not(notn10258,n2929);
and (s0n10258,notn10258,n7125);
and (s1n10258,n2929,n5598);
and (n10259,n10260,n2963);
wire s0n10260,s1n10260,notn10260;
or (n10260,s0n10260,s1n10260);
not(notn10260,n2929);
and (s0n10260,notn10260,n7128);
and (s1n10260,n2929,n5601);
and (n10261,n10262,n2972);
wire s0n10262,s1n10262,notn10262;
or (n10262,s0n10262,s1n10262);
not(notn10262,n2929);
and (s0n10262,notn10262,n7131);
and (s1n10262,n2929,n5604);
and (n10263,n10264,n2742);
or (n10264,1'b0,n10265,n10267,n10269,n10271);
and (n10265,n10266,n2932);
wire s0n10266,s1n10266,notn10266;
or (n10266,s0n10266,s1n10266);
not(notn10266,n2929);
and (s0n10266,notn10266,n5521);
and (s1n10266,n2929,n5609);
and (n10267,n10268,n2955);
wire s0n10268,s1n10268,notn10268;
or (n10268,s0n10268,s1n10268);
not(notn10268,n2929);
and (s0n10268,notn10268,n5525);
and (s1n10268,n2929,n5613);
and (n10269,n10270,n2963);
wire s0n10270,s1n10270,notn10270;
or (n10270,s0n10270,s1n10270);
not(notn10270,n2929);
and (s0n10270,notn10270,n5528);
and (s1n10270,n2929,n5616);
and (n10271,n10272,n2972);
wire s0n10272,s1n10272,notn10272;
or (n10272,s0n10272,s1n10272);
not(notn10272,n2929);
and (s0n10272,notn10272,n5531);
and (s1n10272,n2929,n5619);
and (n10273,n10274,n2752);
or (n10274,1'b0,n10275,n10277,n10279,n10281);
and (n10275,n10276,n2932);
wire s0n10276,s1n10276,notn10276;
or (n10276,s0n10276,s1n10276);
not(notn10276,n2929);
and (s0n10276,notn10276,n5536);
and (s1n10276,n2929,n5624);
and (n10277,n10278,n2955);
wire s0n10278,s1n10278,notn10278;
or (n10278,s0n10278,s1n10278);
not(notn10278,n2929);
and (s0n10278,notn10278,n5539);
and (s1n10278,n2929,n5627);
and (n10279,n10280,n2963);
wire s0n10280,s1n10280,notn10280;
or (n10280,s0n10280,s1n10280);
not(notn10280,n2929);
and (s0n10280,notn10280,n5542);
and (s1n10280,n2929,n5630);
and (n10281,n10282,n2972);
wire s0n10282,s1n10282,notn10282;
or (n10282,s0n10282,s1n10282);
not(notn10282,n2929);
and (s0n10282,notn10282,n5545);
and (s1n10282,n2929,n5633);
or (n10283,1'b0,n10284,n10291,n10297,n10304);
and (n10284,n10285,n2718);
or (n10285,1'b0,n10286,n10288,n10289,n10290);
and (n10286,n10287,n2932);
wire s0n10287,s1n10287,notn10287;
or (n10287,s0n10287,s1n10287);
not(notn10287,n2929);
and (s0n10287,notn10287,n7108);
and (s1n10287,n2929,n5581);
and (n10288,n10246,n2955);
and (n10289,n10248,n2963);
and (n10290,n10250,n2972);
and (n10291,n10292,n2730);
or (n10292,1'b0,n10293,n10294,n10295,n10296);
and (n10293,n10252,n2932);
and (n10294,n10256,n2955);
and (n10295,n10258,n2963);
and (n10296,n10260,n2972);
and (n10297,n10298,n2742);
or (n10298,1'b0,n10299,n10301,n10302,n10303);
and (n10299,n10300,n2932);
wire s0n10300,s1n10300,notn10300;
or (n10300,s0n10300,s1n10300);
not(notn10300,n2929);
and (s0n10300,notn10300,n5522);
and (s1n10300,n2929,n5610);
and (n10301,n10266,n2955);
and (n10302,n10268,n2963);
and (n10303,n10270,n2972);
and (n10304,n10305,n2752);
or (n10305,1'b0,n10306,n10307,n10308,n10309);
and (n10306,n10272,n2932);
and (n10307,n10276,n2955);
and (n10308,n10278,n2963);
and (n10309,n10280,n2972);
and (n10310,n10283,n10311);
or (n10311,n10312,n10381,n10523);
and (n10312,n10313,n10354);
or (n10313,1'b0,n10314,n10324,n10334,n10344);
and (n10314,n10315,n2718);
or (n10315,1'b0,n10316,n10318,n10320,n10322);
and (n10316,n10317,n2932);
wire s0n10317,s1n10317,notn10317;
or (n10317,s0n10317,s1n10317);
not(notn10317,n2929);
and (s0n10317,notn10317,n7176);
and (s1n10317,n2929,n5703);
and (n10318,n10319,n2955);
wire s0n10319,s1n10319,notn10319;
or (n10319,s0n10319,s1n10319);
not(notn10319,n2929);
and (s0n10319,notn10319,n7180);
and (s1n10319,n2929,n5707);
and (n10320,n10321,n2963);
wire s0n10321,s1n10321,notn10321;
or (n10321,s0n10321,s1n10321);
not(notn10321,n2929);
and (s0n10321,notn10321,n7183);
and (s1n10321,n2929,n5710);
and (n10322,n10323,n2972);
wire s0n10323,s1n10323,notn10323;
or (n10323,s0n10323,s1n10323);
not(notn10323,n2929);
and (s0n10323,notn10323,n7186);
and (s1n10323,n2929,n5713);
and (n10324,n10325,n2730);
or (n10325,1'b0,n10326,n10328,n10330,n10332);
and (n10326,n10327,n2932);
wire s0n10327,s1n10327,notn10327;
or (n10327,s0n10327,s1n10327);
not(notn10327,n2929);
and (s0n10327,notn10327,n7191);
and (s1n10327,n2929,n5718);
and (n10328,n10329,n2955);
wire s0n10329,s1n10329,notn10329;
or (n10329,s0n10329,s1n10329);
not(notn10329,n2929);
and (s0n10329,notn10329,n7194);
and (s1n10329,n2929,n5721);
and (n10330,n10331,n2963);
wire s0n10331,s1n10331,notn10331;
or (n10331,s0n10331,s1n10331);
not(notn10331,n2929);
and (s0n10331,notn10331,n7197);
and (s1n10331,n2929,n5724);
and (n10332,n10333,n2972);
wire s0n10333,s1n10333,notn10333;
or (n10333,s0n10333,s1n10333);
not(notn10333,n2929);
and (s0n10333,notn10333,n7200);
and (s1n10333,n2929,n5727);
and (n10334,n10335,n2742);
or (n10335,1'b0,n10336,n10338,n10340,n10342);
and (n10336,n10337,n2932);
wire s0n10337,s1n10337,notn10337;
or (n10337,s0n10337,s1n10337);
not(notn10337,n2929);
and (s0n10337,notn10337,n5644);
and (s1n10337,n2929,n5732);
and (n10338,n10339,n2955);
wire s0n10339,s1n10339,notn10339;
or (n10339,s0n10339,s1n10339);
not(notn10339,n2929);
and (s0n10339,notn10339,n5648);
and (s1n10339,n2929,n5736);
and (n10340,n10341,n2963);
wire s0n10341,s1n10341,notn10341;
or (n10341,s0n10341,s1n10341);
not(notn10341,n2929);
and (s0n10341,notn10341,n5651);
and (s1n10341,n2929,n5739);
and (n10342,n10343,n2972);
wire s0n10343,s1n10343,notn10343;
or (n10343,s0n10343,s1n10343);
not(notn10343,n2929);
and (s0n10343,notn10343,n5654);
and (s1n10343,n2929,n5742);
and (n10344,n10345,n2752);
or (n10345,1'b0,n10346,n10348,n10350,n10352);
and (n10346,n10347,n2932);
wire s0n10347,s1n10347,notn10347;
or (n10347,s0n10347,s1n10347);
not(notn10347,n2929);
and (s0n10347,notn10347,n5659);
and (s1n10347,n2929,n5747);
and (n10348,n10349,n2955);
wire s0n10349,s1n10349,notn10349;
or (n10349,s0n10349,s1n10349);
not(notn10349,n2929);
and (s0n10349,notn10349,n5662);
and (s1n10349,n2929,n5750);
and (n10350,n10351,n2963);
wire s0n10351,s1n10351,notn10351;
or (n10351,s0n10351,s1n10351);
not(notn10351,n2929);
and (s0n10351,notn10351,n5665);
and (s1n10351,n2929,n5753);
and (n10352,n10353,n2972);
wire s0n10353,s1n10353,notn10353;
or (n10353,s0n10353,s1n10353);
not(notn10353,n2929);
and (s0n10353,notn10353,n5668);
and (s1n10353,n2929,n5756);
or (n10354,1'b0,n10355,n10362,n10368,n10375);
and (n10355,n10356,n2718);
or (n10356,1'b0,n10357,n10359,n10360,n10361);
and (n10357,n10358,n2932);
wire s0n10358,s1n10358,notn10358;
or (n10358,s0n10358,s1n10358);
not(notn10358,n2929);
and (s0n10358,notn10358,n7177);
and (s1n10358,n2929,n5704);
and (n10359,n10317,n2955);
and (n10360,n10319,n2963);
and (n10361,n10321,n2972);
and (n10362,n10363,n2730);
or (n10363,1'b0,n10364,n10365,n10366,n10367);
and (n10364,n10323,n2932);
and (n10365,n10327,n2955);
and (n10366,n10329,n2963);
and (n10367,n10331,n2972);
and (n10368,n10369,n2742);
or (n10369,1'b0,n10370,n10372,n10373,n10374);
and (n10370,n10371,n2932);
wire s0n10371,s1n10371,notn10371;
or (n10371,s0n10371,s1n10371);
not(notn10371,n2929);
and (s0n10371,notn10371,n5645);
and (s1n10371,n2929,n5733);
and (n10372,n10337,n2955);
and (n10373,n10339,n2963);
and (n10374,n10341,n2972);
and (n10375,n10376,n2752);
or (n10376,1'b0,n10377,n10378,n10379,n10380);
and (n10377,n10343,n2932);
and (n10378,n10347,n2955);
and (n10379,n10349,n2963);
and (n10380,n10351,n2972);
and (n10381,n10354,n10382);
or (n10382,n10383,n10452,n10522);
and (n10383,n10384,n10425);
or (n10384,1'b0,n10385,n10395,n10405,n10415);
and (n10385,n10386,n2718);
or (n10386,1'b0,n10387,n10389,n10391,n10393);
and (n10387,n10388,n2932);
wire s0n10388,s1n10388,notn10388;
or (n10388,s0n10388,s1n10388);
not(notn10388,n2929);
and (s0n10388,notn10388,n7245);
and (s1n10388,n2929,n5826);
and (n10389,n10390,n2955);
wire s0n10390,s1n10390,notn10390;
or (n10390,s0n10390,s1n10390);
not(notn10390,n2929);
and (s0n10390,notn10390,n7249);
and (s1n10390,n2929,n5830);
and (n10391,n10392,n2963);
wire s0n10392,s1n10392,notn10392;
or (n10392,s0n10392,s1n10392);
not(notn10392,n2929);
and (s0n10392,notn10392,n7252);
and (s1n10392,n2929,n5833);
and (n10393,n10394,n2972);
wire s0n10394,s1n10394,notn10394;
or (n10394,s0n10394,s1n10394);
not(notn10394,n2929);
and (s0n10394,notn10394,n7255);
and (s1n10394,n2929,n5836);
and (n10395,n10396,n2730);
or (n10396,1'b0,n10397,n10399,n10401,n10403);
and (n10397,n10398,n2932);
wire s0n10398,s1n10398,notn10398;
or (n10398,s0n10398,s1n10398);
not(notn10398,n2929);
and (s0n10398,notn10398,n7260);
and (s1n10398,n2929,n5841);
and (n10399,n10400,n2955);
wire s0n10400,s1n10400,notn10400;
or (n10400,s0n10400,s1n10400);
not(notn10400,n2929);
and (s0n10400,notn10400,n7263);
and (s1n10400,n2929,n5844);
and (n10401,n10402,n2963);
wire s0n10402,s1n10402,notn10402;
or (n10402,s0n10402,s1n10402);
not(notn10402,n2929);
and (s0n10402,notn10402,n7266);
and (s1n10402,n2929,n5847);
and (n10403,n10404,n2972);
wire s0n10404,s1n10404,notn10404;
or (n10404,s0n10404,s1n10404);
not(notn10404,n2929);
and (s0n10404,notn10404,n7269);
and (s1n10404,n2929,n5850);
and (n10405,n10406,n2742);
or (n10406,1'b0,n10407,n10409,n10411,n10413);
and (n10407,n10408,n2932);
wire s0n10408,s1n10408,notn10408;
or (n10408,s0n10408,s1n10408);
not(notn10408,n2929);
and (s0n10408,notn10408,n5767);
and (s1n10408,n2929,n5855);
and (n10409,n10410,n2955);
wire s0n10410,s1n10410,notn10410;
or (n10410,s0n10410,s1n10410);
not(notn10410,n2929);
and (s0n10410,notn10410,n5771);
and (s1n10410,n2929,n5859);
and (n10411,n10412,n2963);
wire s0n10412,s1n10412,notn10412;
or (n10412,s0n10412,s1n10412);
not(notn10412,n2929);
and (s0n10412,notn10412,n5774);
and (s1n10412,n2929,n5862);
and (n10413,n10414,n2972);
wire s0n10414,s1n10414,notn10414;
or (n10414,s0n10414,s1n10414);
not(notn10414,n2929);
and (s0n10414,notn10414,n5777);
and (s1n10414,n2929,n5865);
and (n10415,n10416,n2752);
or (n10416,1'b0,n10417,n10419,n10421,n10423);
and (n10417,n10418,n2932);
wire s0n10418,s1n10418,notn10418;
or (n10418,s0n10418,s1n10418);
not(notn10418,n2929);
and (s0n10418,notn10418,n5782);
and (s1n10418,n2929,n5870);
and (n10419,n10420,n2955);
wire s0n10420,s1n10420,notn10420;
or (n10420,s0n10420,s1n10420);
not(notn10420,n2929);
and (s0n10420,notn10420,n5785);
and (s1n10420,n2929,n5873);
and (n10421,n10422,n2963);
wire s0n10422,s1n10422,notn10422;
or (n10422,s0n10422,s1n10422);
not(notn10422,n2929);
and (s0n10422,notn10422,n5788);
and (s1n10422,n2929,n5876);
and (n10423,n10424,n2972);
wire s0n10424,s1n10424,notn10424;
or (n10424,s0n10424,s1n10424);
not(notn10424,n2929);
and (s0n10424,notn10424,n5791);
and (s1n10424,n2929,n5879);
or (n10425,1'b0,n10426,n10433,n10439,n10446);
and (n10426,n10427,n2718);
or (n10427,1'b0,n10428,n10430,n10431,n10432);
and (n10428,n10429,n2932);
wire s0n10429,s1n10429,notn10429;
or (n10429,s0n10429,s1n10429);
not(notn10429,n2929);
and (s0n10429,notn10429,n7246);
and (s1n10429,n2929,n5827);
and (n10430,n10388,n2955);
and (n10431,n10390,n2963);
and (n10432,n10392,n2972);
and (n10433,n10434,n2730);
or (n10434,1'b0,n10435,n10436,n10437,n10438);
and (n10435,n10394,n2932);
and (n10436,n10398,n2955);
and (n10437,n10400,n2963);
and (n10438,n10402,n2972);
and (n10439,n10440,n2742);
or (n10440,1'b0,n10441,n10443,n10444,n10445);
and (n10441,n10442,n2932);
wire s0n10442,s1n10442,notn10442;
or (n10442,s0n10442,s1n10442);
not(notn10442,n2929);
and (s0n10442,notn10442,n5768);
and (s1n10442,n2929,n5856);
and (n10443,n10408,n2955);
and (n10444,n10410,n2963);
and (n10445,n10412,n2972);
and (n10446,n10447,n2752);
or (n10447,1'b0,n10448,n10449,n10450,n10451);
and (n10448,n10414,n2932);
and (n10449,n10418,n2955);
and (n10450,n10420,n2963);
and (n10451,n10422,n2972);
and (n10452,n10425,n10453);
and (n10453,n10454,n10495);
or (n10454,1'b0,n10455,n10465,n10475,n10485);
and (n10455,n10456,n2718);
or (n10456,1'b0,n10457,n10459,n10461,n10463);
and (n10457,n10458,n2932);
wire s0n10458,s1n10458,notn10458;
or (n10458,s0n10458,s1n10458);
not(notn10458,n2929);
and (s0n10458,notn10458,n7313);
and (s1n10458,n2929,n5948);
and (n10459,n10460,n2955);
wire s0n10460,s1n10460,notn10460;
or (n10460,s0n10460,s1n10460);
not(notn10460,n2929);
and (s0n10460,notn10460,n7317);
and (s1n10460,n2929,n5952);
and (n10461,n10462,n2963);
wire s0n10462,s1n10462,notn10462;
or (n10462,s0n10462,s1n10462);
not(notn10462,n2929);
and (s0n10462,notn10462,n7320);
and (s1n10462,n2929,n5955);
and (n10463,n10464,n2972);
wire s0n10464,s1n10464,notn10464;
or (n10464,s0n10464,s1n10464);
not(notn10464,n2929);
and (s0n10464,notn10464,n7323);
and (s1n10464,n2929,n5958);
and (n10465,n10466,n2730);
or (n10466,1'b0,n10467,n10469,n10471,n10473);
and (n10467,n10468,n2932);
wire s0n10468,s1n10468,notn10468;
or (n10468,s0n10468,s1n10468);
not(notn10468,n2929);
and (s0n10468,notn10468,n7328);
and (s1n10468,n2929,n5963);
and (n10469,n10470,n2955);
wire s0n10470,s1n10470,notn10470;
or (n10470,s0n10470,s1n10470);
not(notn10470,n2929);
and (s0n10470,notn10470,n7331);
and (s1n10470,n2929,n5966);
and (n10471,n10472,n2963);
wire s0n10472,s1n10472,notn10472;
or (n10472,s0n10472,s1n10472);
not(notn10472,n2929);
and (s0n10472,notn10472,n7334);
and (s1n10472,n2929,n5969);
and (n10473,n10474,n2972);
wire s0n10474,s1n10474,notn10474;
or (n10474,s0n10474,s1n10474);
not(notn10474,n2929);
and (s0n10474,notn10474,n7337);
and (s1n10474,n2929,n5972);
and (n10475,n10476,n2742);
or (n10476,1'b0,n10477,n10479,n10481,n10483);
and (n10477,n10478,n2932);
wire s0n10478,s1n10478,notn10478;
or (n10478,s0n10478,s1n10478);
not(notn10478,n2929);
and (s0n10478,notn10478,n5889);
and (s1n10478,n2929,n5977);
and (n10479,n10480,n2955);
wire s0n10480,s1n10480,notn10480;
or (n10480,s0n10480,s1n10480);
not(notn10480,n2929);
and (s0n10480,notn10480,n5893);
and (s1n10480,n2929,n5981);
and (n10481,n10482,n2963);
wire s0n10482,s1n10482,notn10482;
or (n10482,s0n10482,s1n10482);
not(notn10482,n2929);
and (s0n10482,notn10482,n5896);
and (s1n10482,n2929,n5984);
and (n10483,n10484,n2972);
wire s0n10484,s1n10484,notn10484;
or (n10484,s0n10484,s1n10484);
not(notn10484,n2929);
and (s0n10484,notn10484,n5899);
and (s1n10484,n2929,n5987);
and (n10485,n10486,n2752);
or (n10486,1'b0,n10487,n10489,n10491,n10493);
and (n10487,n10488,n2932);
wire s0n10488,s1n10488,notn10488;
or (n10488,s0n10488,s1n10488);
not(notn10488,n2929);
and (s0n10488,notn10488,n5904);
and (s1n10488,n2929,n5992);
and (n10489,n10490,n2955);
wire s0n10490,s1n10490,notn10490;
or (n10490,s0n10490,s1n10490);
not(notn10490,n2929);
and (s0n10490,notn10490,n5907);
and (s1n10490,n2929,n5995);
and (n10491,n10492,n2963);
wire s0n10492,s1n10492,notn10492;
or (n10492,s0n10492,s1n10492);
not(notn10492,n2929);
and (s0n10492,notn10492,n5910);
and (s1n10492,n2929,n5998);
and (n10493,n10494,n2972);
wire s0n10494,s1n10494,notn10494;
or (n10494,s0n10494,s1n10494);
not(notn10494,n2929);
and (s0n10494,notn10494,n5913);
and (s1n10494,n2929,n6001);
or (n10495,1'b0,n10496,n10503,n10509,n10516);
and (n10496,n10497,n2718);
or (n10497,1'b0,n10498,n10500,n10501,n10502);
and (n10498,n10499,n2932);
wire s0n10499,s1n10499,notn10499;
or (n10499,s0n10499,s1n10499);
not(notn10499,n2929);
and (s0n10499,notn10499,n7314);
and (s1n10499,n2929,n5949);
and (n10500,n10458,n2955);
and (n10501,n10460,n2963);
and (n10502,n10462,n2972);
and (n10503,n10504,n2730);
or (n10504,1'b0,n10505,n10506,n10507,n10508);
and (n10505,n10464,n2932);
and (n10506,n10468,n2955);
and (n10507,n10470,n2963);
and (n10508,n10472,n2972);
and (n10509,n10510,n2742);
or (n10510,1'b0,n10511,n10513,n10514,n10515);
and (n10511,n10512,n2932);
wire s0n10512,s1n10512,notn10512;
or (n10512,s0n10512,s1n10512);
not(notn10512,n2929);
and (s0n10512,notn10512,n5890);
and (s1n10512,n2929,n5978);
and (n10513,n10478,n2955);
and (n10514,n10480,n2963);
and (n10515,n10482,n2972);
and (n10516,n10517,n2752);
or (n10517,1'b0,n10518,n10519,n10520,n10521);
and (n10518,n10484,n2932);
and (n10519,n10488,n2955);
and (n10520,n10490,n2963);
and (n10521,n10492,n2972);
and (n10522,n10384,n10453);
and (n10523,n10313,n10382);
and (n10524,n10242,n10311);
and (n10525,n10171,n10240);
and (n10526,n10100,n10169);
and (n10527,n10029,n10098);
and (n10528,n9958,n10027);
or (n10529,n10530,n10532);
xor (n10530,n10531,n10027);
xor (n10531,n9958,n9999);
or (n10532,n10533,n11063,n11114);
and (n10533,n10534,n10536);
xor (n10534,n10535,n10098);
xor (n10535,n10029,n10070);
not (n10536,n10537);
or (n10537,n10538,n10600,n11062);
and (n10538,n10539,n10569);
or (n10539,1'b0,n10540,n10546,n10555,n10561);
and (n10540,n10541,n2718);
or (n10541,1'b0,n10542,n10543,n10544,n10545);
and (n10542,n9964,n2932);
and (n10543,n9966,n2955);
and (n10544,n9968,n2963);
and (n10545,n9972,n2972);
and (n10546,n10547,n2730);
or (n10547,1'b0,n10548,n10549,n10550,n10551);
and (n10548,n9974,n2932);
and (n10549,n9976,n2955);
and (n10550,n9978,n2963);
and (n10551,n10552,n2972);
wire s0n10552,s1n10552,notn10552;
or (n10552,s0n10552,s1n10552);
not(notn10552,n2929);
and (s0n10552,notn10552,n10553);
and (s1n10552,n2929,n10554);
and (n10555,n10556,n2742);
or (n10556,1'b0,n10557,n10558,n10559,n10560);
and (n10557,n9984,n2932);
and (n10558,n9986,n2955);
and (n10559,n9988,n2963);
and (n10560,n9992,n2972);
and (n10561,n10562,n2752);
or (n10562,1'b0,n10563,n10564,n10565,n10566);
and (n10563,n9994,n2932);
and (n10564,n9996,n2955);
and (n10565,n9998,n2963);
and (n10566,n10567,n2972);
wire s0n10567,s1n10567,notn10567;
or (n10567,s0n10567,s1n10567);
not(notn10567,n2929);
and (s0n10567,notn10567,n9405);
and (s1n10567,n2929,n10568);
or (n10569,1'b0,n10570,n10579,n10585,n10594);
and (n10570,n10571,n2718);
or (n10571,1'b0,n10572,n10576,n10577,n10578);
and (n10572,n10573,n2932);
wire s0n10573,s1n10573,notn10573;
or (n10573,s0n10573,s1n10573);
not(notn10573,n2929);
and (s0n10573,notn10573,n10574);
and (s1n10573,n2929,n10575);
and (n10576,n10003,n2955);
and (n10577,n9962,n2963);
and (n10578,n9964,n2972);
and (n10579,n10580,n2730);
or (n10580,1'b0,n10581,n10582,n10583,n10584);
and (n10581,n9966,n2932);
and (n10582,n9968,n2955);
and (n10583,n9972,n2963);
and (n10584,n9974,n2972);
and (n10585,n10586,n2742);
or (n10586,1'b0,n10587,n10591,n10592,n10593);
and (n10587,n10588,n2932);
wire s0n10588,s1n10588,notn10588;
or (n10588,s0n10588,s1n10588);
not(notn10588,n2929);
and (s0n10588,notn10588,n10589);
and (s1n10588,n2929,n10590);
and (n10591,n10016,n2955);
and (n10592,n9982,n2963);
and (n10593,n9984,n2972);
and (n10594,n10595,n2752);
or (n10595,1'b0,n10596,n10597,n10598,n10599);
and (n10596,n9986,n2932);
and (n10597,n9988,n2955);
and (n10598,n9992,n2963);
and (n10599,n9994,n2972);
and (n10600,n10569,n10601);
or (n10601,n10602,n10664,n11061);
and (n10602,n10603,n10633);
or (n10603,1'b0,n10604,n10610,n10619,n10625);
and (n10604,n10605,n2718);
or (n10605,1'b0,n10606,n10607,n10608,n10609);
and (n10606,n10035,n2932);
and (n10607,n10037,n2955);
and (n10608,n10039,n2963);
and (n10609,n10043,n2972);
and (n10610,n10611,n2730);
or (n10611,1'b0,n10612,n10613,n10614,n10615);
and (n10612,n10045,n2932);
and (n10613,n10047,n2955);
and (n10614,n10049,n2963);
and (n10615,n10616,n2972);
wire s0n10616,s1n10616,notn10616;
or (n10616,s0n10616,s1n10616);
not(notn10616,n2929);
and (s0n10616,notn10616,n10617);
and (s1n10616,n2929,n10618);
and (n10619,n10620,n2742);
or (n10620,1'b0,n10621,n10622,n10623,n10624);
and (n10621,n10055,n2932);
and (n10622,n10057,n2955);
and (n10623,n10059,n2963);
and (n10624,n10063,n2972);
and (n10625,n10626,n2752);
or (n10626,1'b0,n10627,n10628,n10629,n10630);
and (n10627,n10065,n2932);
and (n10628,n10067,n2955);
and (n10629,n10069,n2963);
and (n10630,n10631,n2972);
wire s0n10631,s1n10631,notn10631;
or (n10631,s0n10631,s1n10631);
not(notn10631,n2929);
and (s0n10631,notn10631,n9417);
and (s1n10631,n2929,n10632);
or (n10633,1'b0,n10634,n10643,n10649,n10658);
and (n10634,n10635,n2718);
or (n10635,1'b0,n10636,n10640,n10641,n10642);
and (n10636,n10637,n2932);
wire s0n10637,s1n10637,notn10637;
or (n10637,s0n10637,s1n10637);
not(notn10637,n2929);
and (s0n10637,notn10637,n10638);
and (s1n10637,n2929,n10639);
and (n10640,n10074,n2955);
and (n10641,n10033,n2963);
and (n10642,n10035,n2972);
and (n10643,n10644,n2730);
or (n10644,1'b0,n10645,n10646,n10647,n10648);
and (n10645,n10037,n2932);
and (n10646,n10039,n2955);
and (n10647,n10043,n2963);
and (n10648,n10045,n2972);
and (n10649,n10650,n2742);
or (n10650,1'b0,n10651,n10655,n10656,n10657);
and (n10651,n10652,n2932);
wire s0n10652,s1n10652,notn10652;
or (n10652,s0n10652,s1n10652);
not(notn10652,n2929);
and (s0n10652,notn10652,n10653);
and (s1n10652,n2929,n10654);
and (n10655,n10087,n2955);
and (n10656,n10053,n2963);
and (n10657,n10055,n2972);
and (n10658,n10659,n2752);
or (n10659,1'b0,n10660,n10661,n10662,n10663);
and (n10660,n10057,n2932);
and (n10661,n10059,n2955);
and (n10662,n10063,n2963);
and (n10663,n10065,n2972);
and (n10664,n10633,n10665);
or (n10665,n10666,n10728,n11060);
and (n10666,n10667,n10697);
or (n10667,1'b0,n10668,n10674,n10683,n10689);
and (n10668,n10669,n2718);
or (n10669,1'b0,n10670,n10671,n10672,n10673);
and (n10670,n10106,n2932);
and (n10671,n10108,n2955);
and (n10672,n10110,n2963);
and (n10673,n10114,n2972);
and (n10674,n10675,n2730);
or (n10675,1'b0,n10676,n10677,n10678,n10679);
and (n10676,n10116,n2932);
and (n10677,n10118,n2955);
and (n10678,n10120,n2963);
and (n10679,n10680,n2972);
wire s0n10680,s1n10680,notn10680;
or (n10680,s0n10680,s1n10680);
not(notn10680,n2929);
and (s0n10680,notn10680,n10681);
and (s1n10680,n2929,n10682);
and (n10683,n10684,n2742);
or (n10684,1'b0,n10685,n10686,n10687,n10688);
and (n10685,n10126,n2932);
and (n10686,n10128,n2955);
and (n10687,n10130,n2963);
and (n10688,n10134,n2972);
and (n10689,n10690,n2752);
or (n10690,1'b0,n10691,n10692,n10693,n10694);
and (n10691,n10136,n2932);
and (n10692,n10138,n2955);
and (n10693,n10140,n2963);
and (n10694,n10695,n2972);
wire s0n10695,s1n10695,notn10695;
or (n10695,s0n10695,s1n10695);
not(notn10695,n2929);
and (s0n10695,notn10695,n9429);
and (s1n10695,n2929,n10696);
or (n10697,1'b0,n10698,n10707,n10713,n10722);
and (n10698,n10699,n2718);
or (n10699,1'b0,n10700,n10704,n10705,n10706);
and (n10700,n10701,n2932);
wire s0n10701,s1n10701,notn10701;
or (n10701,s0n10701,s1n10701);
not(notn10701,n2929);
and (s0n10701,notn10701,n10702);
and (s1n10701,n2929,n10703);
and (n10704,n10145,n2955);
and (n10705,n10104,n2963);
and (n10706,n10106,n2972);
and (n10707,n10708,n2730);
or (n10708,1'b0,n10709,n10710,n10711,n10712);
and (n10709,n10108,n2932);
and (n10710,n10110,n2955);
and (n10711,n10114,n2963);
and (n10712,n10116,n2972);
and (n10713,n10714,n2742);
or (n10714,1'b0,n10715,n10719,n10720,n10721);
and (n10715,n10716,n2932);
wire s0n10716,s1n10716,notn10716;
or (n10716,s0n10716,s1n10716);
not(notn10716,n2929);
and (s0n10716,notn10716,n10717);
and (s1n10716,n2929,n10718);
and (n10719,n10158,n2955);
and (n10720,n10124,n2963);
and (n10721,n10126,n2972);
and (n10722,n10723,n2752);
or (n10723,1'b0,n10724,n10725,n10726,n10727);
and (n10724,n10128,n2932);
and (n10725,n10130,n2955);
and (n10726,n10134,n2963);
and (n10727,n10136,n2972);
and (n10728,n10697,n10729);
or (n10729,n10730,n10792,n11059);
and (n10730,n10731,n10761);
or (n10731,1'b0,n10732,n10738,n10747,n10753);
and (n10732,n10733,n2718);
or (n10733,1'b0,n10734,n10735,n10736,n10737);
and (n10734,n10177,n2932);
and (n10735,n10179,n2955);
and (n10736,n10181,n2963);
and (n10737,n10185,n2972);
and (n10738,n10739,n2730);
or (n10739,1'b0,n10740,n10741,n10742,n10743);
and (n10740,n10187,n2932);
and (n10741,n10189,n2955);
and (n10742,n10191,n2963);
and (n10743,n10744,n2972);
wire s0n10744,s1n10744,notn10744;
or (n10744,s0n10744,s1n10744);
not(notn10744,n2929);
and (s0n10744,notn10744,n10745);
and (s1n10744,n2929,n10746);
and (n10747,n10748,n2742);
or (n10748,1'b0,n10749,n10750,n10751,n10752);
and (n10749,n10197,n2932);
and (n10750,n10199,n2955);
and (n10751,n10201,n2963);
and (n10752,n10205,n2972);
and (n10753,n10754,n2752);
or (n10754,1'b0,n10755,n10756,n10757,n10758);
and (n10755,n10207,n2932);
and (n10756,n10209,n2955);
and (n10757,n10211,n2963);
and (n10758,n10759,n2972);
wire s0n10759,s1n10759,notn10759;
or (n10759,s0n10759,s1n10759);
not(notn10759,n2929);
and (s0n10759,notn10759,n9441);
and (s1n10759,n2929,n10760);
or (n10761,1'b0,n10762,n10771,n10777,n10786);
and (n10762,n10763,n2718);
or (n10763,1'b0,n10764,n10768,n10769,n10770);
and (n10764,n10765,n2932);
wire s0n10765,s1n10765,notn10765;
or (n10765,s0n10765,s1n10765);
not(notn10765,n2929);
and (s0n10765,notn10765,n10766);
and (s1n10765,n2929,n10767);
and (n10768,n10216,n2955);
and (n10769,n10175,n2963);
and (n10770,n10177,n2972);
and (n10771,n10772,n2730);
or (n10772,1'b0,n10773,n10774,n10775,n10776);
and (n10773,n10179,n2932);
and (n10774,n10181,n2955);
and (n10775,n10185,n2963);
and (n10776,n10187,n2972);
and (n10777,n10778,n2742);
or (n10778,1'b0,n10779,n10783,n10784,n10785);
and (n10779,n10780,n2932);
wire s0n10780,s1n10780,notn10780;
or (n10780,s0n10780,s1n10780);
not(notn10780,n2929);
and (s0n10780,notn10780,n10781);
and (s1n10780,n2929,n10782);
and (n10783,n10229,n2955);
and (n10784,n10195,n2963);
and (n10785,n10197,n2972);
and (n10786,n10787,n2752);
or (n10787,1'b0,n10788,n10789,n10790,n10791);
and (n10788,n10199,n2932);
and (n10789,n10201,n2955);
and (n10790,n10205,n2963);
and (n10791,n10207,n2972);
and (n10792,n10761,n10793);
or (n10793,n10794,n10859,n11058);
and (n10794,n10795,n10826);
or (n10795,1'b0,n10796,n10803,n10812,n10818);
not (n10796,n10797);
nand (n10797,n10798,n2718);
or (n10798,1'b0,n10799,n10800,n10801,n10802);
and (n10799,n10248,n2932);
and (n10800,n10250,n2955);
and (n10801,n10252,n2963);
and (n10802,n10256,n2972);
and (n10803,n10804,n2730);
or (n10804,1'b0,n10805,n10806,n10807,n10808);
and (n10805,n10258,n2932);
and (n10806,n10260,n2955);
and (n10807,n10262,n2963);
and (n10808,n10809,n2972);
wire s0n10809,s1n10809,notn10809;
or (n10809,s0n10809,s1n10809);
not(notn10809,n2929);
and (s0n10809,notn10809,n10810);
and (s1n10809,n2929,n10811);
and (n10812,n10813,n2742);
or (n10813,1'b0,n10814,n10815,n10816,n10817);
and (n10814,n10268,n2932);
and (n10815,n10270,n2955);
and (n10816,n10272,n2963);
and (n10817,n10276,n2972);
and (n10818,n10819,n2752);
or (n10819,1'b0,n10820,n10821,n10822,n10823);
and (n10820,n10278,n2932);
and (n10821,n10280,n2955);
and (n10822,n10282,n2963);
and (n10823,n10824,n2972);
wire s0n10824,s1n10824,notn10824;
or (n10824,s0n10824,s1n10824);
not(notn10824,n2929);
and (s0n10824,notn10824,n9453);
and (s1n10824,n2929,n10825);
or (n10826,1'b0,n10827,n10836,n10843,n10852);
and (n10827,n10828,n2718);
or (n10828,1'b0,n10829,n10833,n10834,n10835);
and (n10829,n10830,n2932);
wire s0n10830,s1n10830,notn10830;
or (n10830,s0n10830,s1n10830);
not(notn10830,n2929);
and (s0n10830,notn10830,n10831);
and (s1n10830,n2929,n10832);
and (n10833,n10287,n2955);
and (n10834,n10246,n2963);
and (n10835,n10248,n2972);
not (n10836,n10837);
nand (n10837,n10838,n2730);
or (n10838,1'b0,n10839,n10840,n10841,n10842);
and (n10839,n10250,n2932);
and (n10840,n10252,n2955);
and (n10841,n10256,n2963);
and (n10842,n10258,n2972);
and (n10843,n10844,n2742);
or (n10844,1'b0,n10845,n10849,n10850,n10851);
and (n10845,n10846,n2932);
wire s0n10846,s1n10846,notn10846;
or (n10846,s0n10846,s1n10846);
not(notn10846,n2929);
and (s0n10846,notn10846,n10847);
and (s1n10846,n2929,n10848);
and (n10849,n10300,n2955);
and (n10850,n10266,n2963);
and (n10851,n10268,n2972);
not (n10852,n10853);
nand (n10853,n10854,n2752);
or (n10854,1'b0,n10855,n10856,n10857,n10858);
and (n10855,n10270,n2932);
and (n10856,n10272,n2955);
and (n10857,n10276,n2963);
and (n10858,n10278,n2972);
and (n10859,n10826,n10860);
or (n10860,n10861,n10925,n11057);
and (n10861,n10862,n10894);
or (n10862,1'b0,n10863,n10870,n10879,n10886);
not (n10863,n10864);
nand (n10864,n10865,n2718);
or (n10865,1'b0,n10866,n10867,n10868,n10869);
and (n10866,n10319,n2932);
and (n10867,n10321,n2955);
and (n10868,n10323,n2963);
and (n10869,n10327,n2972);
and (n10870,n10871,n2730);
or (n10871,1'b0,n10872,n10873,n10874,n10875);
and (n10872,n10329,n2932);
and (n10873,n10331,n2955);
and (n10874,n10333,n2963);
and (n10875,n10876,n2972);
wire s0n10876,s1n10876,notn10876;
or (n10876,s0n10876,s1n10876);
not(notn10876,n2929);
and (s0n10876,notn10876,n10877);
and (s1n10876,n2929,n10878);
not (n10879,n10880);
nand (n10880,n10881,n2742);
or (n10881,1'b0,n10882,n10883,n10884,n10885);
and (n10882,n10339,n2932);
and (n10883,n10341,n2955);
and (n10884,n10343,n2963);
and (n10885,n10347,n2972);
and (n10886,n10887,n2752);
or (n10887,1'b0,n10888,n10889,n10890,n10891);
and (n10888,n10349,n2932);
and (n10889,n10351,n2955);
and (n10890,n10353,n2963);
and (n10891,n10892,n2972);
wire s0n10892,s1n10892,notn10892;
or (n10892,s0n10892,s1n10892);
not(notn10892,n2929);
and (s0n10892,notn10892,n9465);
and (s1n10892,n2929,n10893);
or (n10894,1'b0,n10895,n10904,n10910,n10919);
and (n10895,n10896,n2718);
or (n10896,1'b0,n10897,n10901,n10902,n10903);
and (n10897,n10898,n2932);
wire s0n10898,s1n10898,notn10898;
or (n10898,s0n10898,s1n10898);
not(notn10898,n2929);
and (s0n10898,notn10898,n10899);
and (s1n10898,n2929,n10900);
and (n10901,n10358,n2955);
and (n10902,n10317,n2963);
and (n10903,n10319,n2972);
and (n10904,n10905,n2730);
or (n10905,1'b0,n10906,n10907,n10908,n10909);
and (n10906,n10321,n2932);
and (n10907,n10323,n2955);
and (n10908,n10327,n2963);
and (n10909,n10329,n2972);
and (n10910,n10911,n2742);
or (n10911,1'b0,n10912,n10916,n10917,n10918);
and (n10912,n10913,n2932);
wire s0n10913,s1n10913,notn10913;
or (n10913,s0n10913,s1n10913);
not(notn10913,n2929);
and (s0n10913,notn10913,n10914);
and (s1n10913,n2929,n10915);
and (n10916,n10371,n2955);
and (n10917,n10337,n2963);
and (n10918,n10339,n2972);
and (n10919,n10920,n2752);
or (n10920,1'b0,n10921,n10922,n10923,n10924);
and (n10921,n10341,n2932);
and (n10922,n10343,n2955);
and (n10923,n10347,n2963);
and (n10924,n10349,n2972);
and (n10925,n10894,n10926);
or (n10926,n10927,n10989,n11056);
and (n10927,n10928,n10958);
or (n10928,1'b0,n10929,n10935,n10944,n10950);
and (n10929,n10930,n2718);
or (n10930,1'b0,n10931,n10932,n10933,n10934);
and (n10931,n10390,n2932);
and (n10932,n10392,n2955);
and (n10933,n10394,n2963);
and (n10934,n10398,n2972);
and (n10935,n10936,n2730);
or (n10936,1'b0,n10937,n10938,n10939,n10940);
and (n10937,n10400,n2932);
and (n10938,n10402,n2955);
and (n10939,n10404,n2963);
and (n10940,n10941,n2972);
wire s0n10941,s1n10941,notn10941;
or (n10941,s0n10941,s1n10941);
not(notn10941,n2929);
and (s0n10941,notn10941,n10942);
and (s1n10941,n2929,n10943);
and (n10944,n10945,n2742);
or (n10945,1'b0,n10946,n10947,n10948,n10949);
and (n10946,n10410,n2932);
and (n10947,n10412,n2955);
and (n10948,n10414,n2963);
and (n10949,n10418,n2972);
and (n10950,n10951,n2752);
or (n10951,1'b0,n10952,n10953,n10954,n10955);
and (n10952,n10420,n2932);
and (n10953,n10422,n2955);
and (n10954,n10424,n2963);
and (n10955,n10956,n2972);
wire s0n10956,s1n10956,notn10956;
or (n10956,s0n10956,s1n10956);
not(notn10956,n2929);
and (s0n10956,notn10956,n9477);
and (s1n10956,n2929,n10957);
or (n10958,1'b0,n10959,n10968,n10974,n10983);
and (n10959,n10960,n2718);
or (n10960,1'b0,n10961,n10965,n10966,n10967);
and (n10961,n10962,n2932);
wire s0n10962,s1n10962,notn10962;
or (n10962,s0n10962,s1n10962);
not(notn10962,n2929);
and (s0n10962,notn10962,n10963);
and (s1n10962,n2929,n10964);
and (n10965,n10429,n2955);
and (n10966,n10388,n2963);
and (n10967,n10390,n2972);
and (n10968,n10969,n2730);
or (n10969,1'b0,n10970,n10971,n10972,n10973);
and (n10970,n10392,n2932);
and (n10971,n10394,n2955);
and (n10972,n10398,n2963);
and (n10973,n10400,n2972);
and (n10974,n10975,n2742);
or (n10975,1'b0,n10976,n10980,n10981,n10982);
and (n10976,n10977,n2932);
wire s0n10977,s1n10977,notn10977;
or (n10977,s0n10977,s1n10977);
not(notn10977,n2929);
and (s0n10977,notn10977,n10978);
and (s1n10977,n2929,n10979);
and (n10980,n10442,n2955);
and (n10981,n10408,n2963);
and (n10982,n10410,n2972);
and (n10983,n10984,n2752);
or (n10984,1'b0,n10985,n10986,n10987,n10988);
and (n10985,n10412,n2932);
and (n10986,n10414,n2955);
and (n10987,n10418,n2963);
and (n10988,n10420,n2972);
and (n10989,n10958,n10990);
and (n10990,n10991,n11023);
or (n10991,1'b0,n10992,n10999,n11008,n11015);
not (n10992,n10993);
nand (n10993,n10994,n2718);
or (n10994,1'b0,n10995,n10996,n10997,n10998);
and (n10995,n10460,n2932);
and (n10996,n10462,n2955);
and (n10997,n10464,n2963);
and (n10998,n10468,n2972);
and (n10999,n11000,n2730);
or (n11000,1'b0,n11001,n11002,n11003,n11004);
and (n11001,n10470,n2932);
and (n11002,n10472,n2955);
and (n11003,n10474,n2963);
and (n11004,n11005,n2972);
wire s0n11005,s1n11005,notn11005;
or (n11005,s0n11005,s1n11005);
not(notn11005,n2929);
and (s0n11005,notn11005,n11006);
and (s1n11005,n2929,n11007);
not (n11008,n11009);
nand (n11009,n11010,n2742);
or (n11010,1'b0,n11011,n11012,n11013,n11014);
and (n11011,n10480,n2932);
and (n11012,n10482,n2955);
and (n11013,n10484,n2963);
and (n11014,n10488,n2972);
and (n11015,n11016,n2752);
or (n11016,1'b0,n11017,n11018,n11019,n11020);
and (n11017,n10490,n2932);
and (n11018,n10492,n2955);
and (n11019,n10494,n2963);
and (n11020,n11021,n2972);
wire s0n11021,s1n11021,notn11021;
or (n11021,s0n11021,s1n11021);
not(notn11021,n2929);
and (s0n11021,notn11021,n9488);
and (s1n11021,n2929,n11022);
or (n11023,1'b0,n11024,n11033,n11040,n11049);
and (n11024,n11025,n2718);
or (n11025,1'b0,n11026,n11030,n11031,n11032);
and (n11026,n11027,n2932);
wire s0n11027,s1n11027,notn11027;
or (n11027,s0n11027,s1n11027);
not(notn11027,n2929);
and (s0n11027,notn11027,n11028);
and (s1n11027,n2929,n11029);
and (n11030,n10499,n2955);
and (n11031,n10458,n2963);
and (n11032,n10460,n2972);
not (n11033,n11034);
nand (n11034,n11035,n2730);
or (n11035,1'b0,n11036,n11037,n11038,n11039);
and (n11036,n10462,n2932);
and (n11037,n10464,n2955);
and (n11038,n10468,n2963);
and (n11039,n10470,n2972);
and (n11040,n11041,n2742);
or (n11041,1'b0,n11042,n11046,n11047,n11048);
and (n11042,n11043,n2932);
wire s0n11043,s1n11043,notn11043;
or (n11043,s0n11043,s1n11043);
not(notn11043,n2929);
and (s0n11043,notn11043,n11044);
and (s1n11043,n2929,n11045);
and (n11046,n10512,n2955);
and (n11047,n10478,n2963);
and (n11048,n10480,n2972);
not (n11049,n11050);
nand (n11050,n11051,n2752);
or (n11051,1'b0,n11052,n11053,n11054,n11055);
and (n11052,n10482,n2932);
and (n11053,n10484,n2955);
and (n11054,n10488,n2963);
and (n11055,n10490,n2972);
and (n11056,n10928,n10990);
and (n11057,n10862,n10926);
and (n11058,n10795,n10860);
and (n11059,n10731,n10793);
and (n11060,n10667,n10729);
and (n11061,n10603,n10665);
and (n11062,n10539,n10601);
and (n11063,n10536,n11064);
or (n11064,n11065,n11071,n11113);
and (n11065,n11066,n11068);
xor (n11066,n11067,n10169);
xor (n11067,n10100,n10141);
not (n11068,n11069);
xor (n11069,n11070,n10601);
xor (n11070,n10539,n10569);
and (n11071,n11068,n11072);
or (n11072,n11073,n11079,n11112);
and (n11073,n11074,n11076);
xor (n11074,n11075,n10240);
xor (n11075,n10171,n10212);
not (n11076,n11077);
xor (n11077,n11078,n10665);
xor (n11078,n10603,n10633);
and (n11079,n11076,n11080);
or (n11080,n11081,n11087,n11111);
and (n11081,n11082,n11084);
xor (n11082,n11083,n10311);
xor (n11083,n10242,n10283);
not (n11084,n11085);
xor (n11085,n11086,n10729);
xor (n11086,n10667,n10697);
and (n11087,n11084,n11088);
or (n11088,n11089,n11095,n11110);
and (n11089,n11090,n11092);
xor (n11090,n11091,n10382);
xor (n11091,n10313,n10354);
not (n11092,n11093);
xor (n11093,n11094,n10793);
xor (n11094,n10731,n10761);
and (n11095,n11092,n11096);
or (n11096,n11097,n11103,n11109);
and (n11097,n11098,n11100);
xor (n11098,n11099,n10453);
xor (n11099,n10384,n10425);
not (n11100,n11101);
xor (n11101,n11102,n10860);
xor (n11102,n10795,n10826);
and (n11103,n11100,n11104);
and (n11104,n11105,n11106);
xor (n11105,n10454,n10495);
not (n11106,n11107);
xor (n11107,n11108,n10926);
xor (n11108,n10862,n10894);
and (n11109,n11098,n11104);
and (n11110,n11090,n11096);
and (n11111,n11082,n11088);
and (n11112,n11074,n11080);
and (n11113,n11066,n11072);
and (n11114,n10534,n11064);
and (n11115,n11116,n11117);
xnor (n11116,n9956,n10529);
and (n11117,n11118,n11119);
xnor (n11118,n10530,n10532);
and (n11119,n11120,n11122);
xor (n11120,n11121,n11064);
xor (n11121,n10534,n10536);
and (n11122,n11123,n11125);
xor (n11123,n11124,n11072);
xor (n11124,n11066,n11068);
and (n11125,n11126,n11128);
xor (n11126,n11127,n11080);
xor (n11127,n11074,n11076);
and (n11128,n11129,n11131);
xor (n11129,n11130,n11088);
xor (n11130,n11082,n11084);
and (n11131,n11132,n11134);
xor (n11132,n11133,n11096);
xor (n11133,n11090,n11092);
and (n11134,n11135,n11137);
xor (n11135,n11136,n11104);
xor (n11136,n11098,n11100);
and (n11137,n11138,n11139);
xor (n11138,n11105,n11106);
and (n11139,n11140,n11143);
not (n11140,n11141);
xor (n11141,n11142,n10990);
xor (n11142,n10928,n10958);
not (n11143,n11144);
xor (n11144,n10991,n11023);
and (n11145,n9953,n11146);
and (n11146,n11147,n11148);
xor (n11147,n11116,n11117);
and (n11148,n11149,n11150);
xor (n11149,n11118,n11119);
or (n11150,n11151,n11532,n11584);
and (n11151,n11152,n11531);
or (n11152,n11153,n11198,n11530);
and (n11153,n11154,n11175);
or (n11154,1'b0,n11155,n11156,n11165,n11167);
and (n11155,n10580,n2718);
and (n11156,n11157,n2730);
or (n11157,1'b0,n11158,n11159,n11160,n11161);
and (n11158,n9976,n2932);
and (n11159,n9978,n2955);
and (n11160,n10552,n2963);
and (n11161,n11162,n2972);
wire s0n11162,s1n11162,notn11162;
or (n11162,s0n11162,s1n11162);
not(notn11162,n2929);
and (s0n11162,notn11162,n11163);
and (s1n11162,n2929,n11164);
not (n11165,n11166);
nand (n11166,n10595,n2742);
and (n11167,n11168,n2752);
or (n11168,1'b0,n11169,n11170,n11171,n11172);
and (n11169,n9996,n2932);
and (n11170,n9998,n2955);
and (n11171,n10567,n2963);
and (n11172,n11173,n2972);
wire s0n11173,s1n11173,notn11173;
or (n11173,s0n11173,s1n11173);
not(notn11173,n2929);
and (s0n11173,notn11173,n9092);
and (s1n11173,n2929,n11174);
or (n11175,1'b0,n11176,n11185,n11187,n11196);
and (n11176,n11177,n2718);
or (n11177,1'b0,n11178,n11182,n11183,n11184);
and (n11178,n11179,n2932);
wire s0n11179,s1n11179,notn11179;
or (n11179,s0n11179,s1n11179);
not(notn11179,n2929);
and (s0n11179,notn11179,n11180);
and (s1n11179,n2929,n11181);
and (n11182,n10573,n2955);
and (n11183,n10003,n2963);
and (n11184,n9962,n2972);
not (n11185,n11186);
nand (n11186,n10541,n2730);
and (n11187,n11188,n2742);
or (n11188,1'b0,n11189,n11193,n11194,n11195);
and (n11189,n11190,n2932);
wire s0n11190,s1n11190,notn11190;
or (n11190,s0n11190,s1n11190);
not(notn11190,n2929);
and (s0n11190,notn11190,n11191);
and (s1n11190,n2929,n11192);
and (n11193,n10588,n2955);
and (n11194,n10016,n2963);
and (n11195,n9982,n2972);
not (n11196,n11197);
nand (n11197,n10556,n2752);
and (n11198,n11175,n11199);
or (n11199,n11200,n11245,n11529);
and (n11200,n11201,n11222);
or (n11201,1'b0,n11202,n11203,n11212,n11214);
and (n11202,n10644,n2718);
and (n11203,n11204,n2730);
or (n11204,1'b0,n11205,n11206,n11207,n11208);
and (n11205,n10047,n2932);
and (n11206,n10049,n2955);
and (n11207,n10616,n2963);
and (n11208,n11209,n2972);
wire s0n11209,s1n11209,notn11209;
or (n11209,s0n11209,s1n11209);
not(notn11209,n2929);
and (s0n11209,notn11209,n11210);
and (s1n11209,n2929,n11211);
not (n11212,n11213);
nand (n11213,n10659,n2742);
and (n11214,n11215,n2752);
or (n11215,1'b0,n11216,n11217,n11218,n11219);
and (n11216,n10067,n2932);
and (n11217,n10069,n2955);
and (n11218,n10631,n2963);
and (n11219,n11220,n2972);
wire s0n11220,s1n11220,notn11220;
or (n11220,s0n11220,s1n11220);
not(notn11220,n2929);
and (s0n11220,notn11220,n9106);
and (s1n11220,n2929,n11221);
or (n11222,1'b0,n11223,n11232,n11234,n11243);
and (n11223,n11224,n2718);
or (n11224,1'b0,n11225,n11229,n11230,n11231);
and (n11225,n11226,n2932);
wire s0n11226,s1n11226,notn11226;
or (n11226,s0n11226,s1n11226);
not(notn11226,n2929);
and (s0n11226,notn11226,n11227);
and (s1n11226,n2929,n11228);
and (n11229,n10637,n2955);
and (n11230,n10074,n2963);
and (n11231,n10033,n2972);
not (n11232,n11233);
nand (n11233,n10605,n2730);
and (n11234,n11235,n2742);
or (n11235,1'b0,n11236,n11240,n11241,n11242);
and (n11236,n11237,n2932);
wire s0n11237,s1n11237,notn11237;
or (n11237,s0n11237,s1n11237);
not(notn11237,n2929);
and (s0n11237,notn11237,n11238);
and (s1n11237,n2929,n11239);
and (n11240,n10652,n2955);
and (n11241,n10087,n2963);
and (n11242,n10053,n2972);
not (n11243,n11244);
nand (n11244,n10620,n2752);
and (n11245,n11222,n11246);
or (n11246,n11247,n11292,n11528);
and (n11247,n11248,n11269);
or (n11248,1'b0,n11249,n11250,n11259,n11261);
and (n11249,n10708,n2718);
and (n11250,n11251,n2730);
or (n11251,1'b0,n11252,n11253,n11254,n11255);
and (n11252,n10118,n2932);
and (n11253,n10120,n2955);
and (n11254,n10680,n2963);
and (n11255,n11256,n2972);
wire s0n11256,s1n11256,notn11256;
or (n11256,s0n11256,s1n11256);
not(notn11256,n2929);
and (s0n11256,notn11256,n11257);
and (s1n11256,n2929,n11258);
not (n11259,n11260);
nand (n11260,n10723,n2742);
and (n11261,n11262,n2752);
or (n11262,1'b0,n11263,n11264,n11265,n11266);
and (n11263,n10138,n2932);
and (n11264,n10140,n2955);
and (n11265,n10695,n2963);
and (n11266,n11267,n2972);
wire s0n11267,s1n11267,notn11267;
or (n11267,s0n11267,s1n11267);
not(notn11267,n2929);
and (s0n11267,notn11267,n9120);
and (s1n11267,n2929,n11268);
or (n11269,1'b0,n11270,n11279,n11281,n11290);
and (n11270,n11271,n2718);
or (n11271,1'b0,n11272,n11276,n11277,n11278);
and (n11272,n11273,n2932);
wire s0n11273,s1n11273,notn11273;
or (n11273,s0n11273,s1n11273);
not(notn11273,n2929);
and (s0n11273,notn11273,n11274);
and (s1n11273,n2929,n11275);
and (n11276,n10701,n2955);
and (n11277,n10145,n2963);
and (n11278,n10104,n2972);
not (n11279,n11280);
nand (n11280,n10669,n2730);
and (n11281,n11282,n2742);
or (n11282,1'b0,n11283,n11287,n11288,n11289);
and (n11283,n11284,n2932);
wire s0n11284,s1n11284,notn11284;
or (n11284,s0n11284,s1n11284);
not(notn11284,n2929);
and (s0n11284,notn11284,n11285);
and (s1n11284,n2929,n11286);
and (n11287,n10716,n2955);
and (n11288,n10158,n2963);
and (n11289,n10124,n2972);
not (n11290,n11291);
nand (n11291,n10684,n2752);
and (n11292,n11269,n11293);
or (n11293,n11294,n11339,n11527);
and (n11294,n11295,n11316);
or (n11295,1'b0,n11296,n11297,n11306,n11308);
and (n11296,n10772,n2718);
and (n11297,n11298,n2730);
or (n11298,1'b0,n11299,n11300,n11301,n11302);
and (n11299,n10189,n2932);
and (n11300,n10191,n2955);
and (n11301,n10744,n2963);
and (n11302,n11303,n2972);
wire s0n11303,s1n11303,notn11303;
or (n11303,s0n11303,s1n11303);
not(notn11303,n2929);
and (s0n11303,notn11303,n11304);
and (s1n11303,n2929,n11305);
not (n11306,n11307);
nand (n11307,n10787,n2742);
and (n11308,n11309,n2752);
or (n11309,1'b0,n11310,n11311,n11312,n11313);
and (n11310,n10209,n2932);
and (n11311,n10211,n2955);
and (n11312,n10759,n2963);
and (n11313,n11314,n2972);
wire s0n11314,s1n11314,notn11314;
or (n11314,s0n11314,s1n11314);
not(notn11314,n2929);
and (s0n11314,notn11314,n9142);
and (s1n11314,n2929,n11315);
or (n11316,1'b0,n11317,n11326,n11328,n11337);
and (n11317,n11318,n2718);
or (n11318,1'b0,n11319,n11323,n11324,n11325);
and (n11319,n11320,n2932);
wire s0n11320,s1n11320,notn11320;
or (n11320,s0n11320,s1n11320);
not(notn11320,n2929);
and (s0n11320,notn11320,n11321);
and (s1n11320,n2929,n11322);
and (n11323,n10765,n2955);
and (n11324,n10216,n2963);
and (n11325,n10175,n2972);
not (n11326,n11327);
nand (n11327,n10733,n2730);
and (n11328,n11329,n2742);
or (n11329,1'b0,n11330,n11334,n11335,n11336);
and (n11330,n11331,n2932);
wire s0n11331,s1n11331,notn11331;
or (n11331,s0n11331,s1n11331);
not(notn11331,n2929);
and (s0n11331,notn11331,n11332);
and (s1n11331,n2929,n11333);
and (n11334,n10780,n2955);
and (n11335,n10229,n2963);
and (n11336,n10195,n2972);
not (n11337,n11338);
nand (n11338,n10748,n2752);
and (n11339,n11316,n11340);
or (n11340,n11341,n11384,n11526);
and (n11341,n11342,n11363);
or (n11342,1'b0,n11343,n11344,n11353,n11355);
and (n11343,n10838,n2718);
and (n11344,n11345,n2730);
or (n11345,1'b0,n11346,n11347,n11348,n11349);
and (n11346,n10260,n2932);
and (n11347,n10262,n2955);
and (n11348,n10809,n2963);
and (n11349,n11350,n2972);
wire s0n11350,s1n11350,notn11350;
or (n11350,s0n11350,s1n11350);
not(notn11350,n2929);
and (s0n11350,notn11350,n11351);
and (s1n11350,n2929,n11352);
not (n11353,n11354);
nand (n11354,n10854,n2742);
and (n11355,n11356,n2752);
or (n11356,1'b0,n11357,n11358,n11359,n11360);
and (n11357,n10280,n2932);
and (n11358,n10282,n2955);
and (n11359,n10824,n2963);
and (n11360,n11361,n2972);
wire s0n11361,s1n11361,notn11361;
or (n11361,s0n11361,s1n11361);
not(notn11361,n2929);
and (s0n11361,notn11361,n9166);
and (s1n11361,n2929,n11362);
or (n11363,1'b0,n11364,n11373,n11374,n11383);
and (n11364,n11365,n2718);
or (n11365,1'b0,n11366,n11370,n11371,n11372);
and (n11366,n11367,n2932);
wire s0n11367,s1n11367,notn11367;
or (n11367,s0n11367,s1n11367);
not(notn11367,n2929);
and (s0n11367,notn11367,n11368);
and (s1n11367,n2929,n11369);
and (n11370,n10830,n2955);
and (n11371,n10287,n2963);
and (n11372,n10246,n2972);
and (n11373,n10798,n2730);
and (n11374,n11375,n2742);
or (n11375,1'b0,n11376,n11380,n11381,n11382);
and (n11376,n11377,n2932);
wire s0n11377,s1n11377,notn11377;
or (n11377,s0n11377,s1n11377);
not(notn11377,n2929);
and (s0n11377,notn11377,n11378);
and (s1n11377,n2929,n11379);
and (n11380,n10846,n2955);
and (n11381,n10300,n2963);
and (n11382,n10266,n2972);
and (n11383,n10813,n2752);
and (n11384,n11363,n11385);
or (n11385,n11386,n11431,n11525);
and (n11386,n11387,n11408);
or (n11387,1'b0,n11388,n11389,n11398,n11400);
and (n11388,n10905,n2718);
and (n11389,n11390,n2730);
or (n11390,1'b0,n11391,n11392,n11393,n11394);
and (n11391,n10331,n2932);
and (n11392,n10333,n2955);
and (n11393,n10876,n2963);
and (n11394,n11395,n2972);
wire s0n11395,s1n11395,notn11395;
or (n11395,s0n11395,s1n11395);
not(notn11395,n2929);
and (s0n11395,notn11395,n11396);
and (s1n11395,n2929,n11397);
not (n11398,n11399);
nand (n11399,n10920,n2742);
and (n11400,n11401,n2752);
or (n11401,1'b0,n11402,n11403,n11404,n11405);
and (n11402,n10351,n2932);
and (n11403,n10353,n2955);
and (n11404,n10892,n2963);
and (n11405,n11406,n2972);
wire s0n11406,s1n11406,notn11406;
or (n11406,s0n11406,s1n11406);
not(notn11406,n2929);
and (s0n11406,notn11406,n9189);
and (s1n11406,n2929,n11407);
or (n11408,1'b0,n11409,n11418,n11420,n11429);
and (n11409,n11410,n2718);
or (n11410,1'b0,n11411,n11415,n11416,n11417);
and (n11411,n11412,n2932);
wire s0n11412,s1n11412,notn11412;
or (n11412,s0n11412,s1n11412);
not(notn11412,n2929);
and (s0n11412,notn11412,n11413);
and (s1n11412,n2929,n11414);
and (n11415,n10898,n2955);
and (n11416,n10358,n2963);
and (n11417,n10317,n2972);
not (n11418,n11419);
nand (n11419,n10865,n2730);
and (n11420,n11421,n2742);
or (n11421,1'b0,n11422,n11426,n11427,n11428);
and (n11422,n11423,n2932);
wire s0n11423,s1n11423,notn11423;
or (n11423,s0n11423,s1n11423);
not(notn11423,n2929);
and (s0n11423,notn11423,n11424);
and (s1n11423,n2929,n11425);
and (n11426,n10913,n2955);
and (n11427,n10371,n2963);
and (n11428,n10337,n2972);
not (n11429,n11430);
nand (n11430,n10881,n2752);
and (n11431,n11408,n11432);
or (n11432,n11433,n11478,n11524);
and (n11433,n11434,n11455);
or (n11434,1'b0,n11435,n11436,n11445,n11447);
and (n11435,n10969,n2718);
and (n11436,n11437,n2730);
or (n11437,1'b0,n11438,n11439,n11440,n11441);
and (n11438,n10402,n2932);
and (n11439,n10404,n2955);
and (n11440,n10941,n2963);
and (n11441,n11442,n2972);
wire s0n11442,s1n11442,notn11442;
or (n11442,s0n11442,s1n11442);
not(notn11442,n2929);
and (s0n11442,notn11442,n11443);
and (s1n11442,n2929,n11444);
not (n11445,n11446);
nand (n11446,n10984,n2742);
and (n11447,n11448,n2752);
or (n11448,1'b0,n11449,n11450,n11451,n11452);
and (n11449,n10422,n2932);
and (n11450,n10424,n2955);
and (n11451,n10956,n2963);
and (n11452,n11453,n2972);
wire s0n11453,s1n11453,notn11453;
or (n11453,s0n11453,s1n11453);
not(notn11453,n2929);
and (s0n11453,notn11453,n9215);
and (s1n11453,n2929,n11454);
or (n11455,1'b0,n11456,n11465,n11467,n11476);
and (n11456,n11457,n2718);
or (n11457,1'b0,n11458,n11462,n11463,n11464);
and (n11458,n11459,n2932);
wire s0n11459,s1n11459,notn11459;
or (n11459,s0n11459,s1n11459);
not(notn11459,n2929);
and (s0n11459,notn11459,n11460);
and (s1n11459,n2929,n11461);
and (n11462,n10962,n2955);
and (n11463,n10429,n2963);
and (n11464,n10388,n2972);
not (n11465,n11466);
nand (n11466,n10930,n2730);
and (n11467,n11468,n2742);
or (n11468,1'b0,n11469,n11473,n11474,n11475);
and (n11469,n11470,n2932);
wire s0n11470,s1n11470,notn11470;
or (n11470,s0n11470,s1n11470);
not(notn11470,n2929);
and (s0n11470,notn11470,n11471);
and (s1n11470,n2929,n11472);
and (n11473,n10977,n2955);
and (n11474,n10442,n2963);
and (n11475,n10408,n2972);
not (n11476,n11477);
nand (n11477,n10945,n2752);
and (n11478,n11455,n11479);
and (n11479,n11480,n11501);
or (n11480,1'b0,n11481,n11482,n11491,n11493);
and (n11481,n11035,n2718);
and (n11482,n11483,n2730);
or (n11483,1'b0,n11484,n11485,n11486,n11487);
and (n11484,n10472,n2932);
and (n11485,n10474,n2955);
and (n11486,n11005,n2963);
and (n11487,n11488,n2972);
wire s0n11488,s1n11488,notn11488;
or (n11488,s0n11488,s1n11488);
not(notn11488,n2929);
and (s0n11488,notn11488,n11489);
and (s1n11488,n2929,n11490);
not (n11491,n11492);
nand (n11492,n11051,n2742);
and (n11493,n11494,n2752);
or (n11494,1'b0,n11495,n11496,n11497,n11498);
and (n11495,n10492,n2932);
and (n11496,n10494,n2955);
and (n11497,n11021,n2963);
and (n11498,n11499,n2972);
wire s0n11499,s1n11499,notn11499;
or (n11499,s0n11499,s1n11499);
not(notn11499,n2929);
and (s0n11499,notn11499,n9231);
and (s1n11499,n2929,n11500);
or (n11501,1'b0,n11502,n11511,n11513,n11522);
and (n11502,n11503,n2718);
or (n11503,1'b0,n11504,n11508,n11509,n11510);
and (n11504,n11505,n2932);
wire s0n11505,s1n11505,notn11505;
or (n11505,s0n11505,s1n11505);
not(notn11505,n2929);
and (s0n11505,notn11505,n11506);
and (s1n11505,n2929,n11507);
and (n11508,n11027,n2955);
and (n11509,n10499,n2963);
and (n11510,n10458,n2972);
not (n11511,n11512);
nand (n11512,n10994,n2730);
and (n11513,n11514,n2742);
or (n11514,1'b0,n11515,n11519,n11520,n11521);
and (n11515,n11516,n2932);
wire s0n11516,s1n11516,notn11516;
or (n11516,s0n11516,s1n11516);
not(notn11516,n2929);
and (s0n11516,notn11516,n11517);
and (s1n11516,n2929,n11518);
and (n11519,n11043,n2955);
and (n11520,n10512,n2963);
and (n11521,n10478,n2972);
not (n11522,n11523);
nand (n11523,n11010,n2752);
and (n11524,n11434,n11479);
and (n11525,n11387,n11432);
and (n11526,n11342,n11385);
and (n11527,n11295,n11340);
and (n11528,n11248,n11293);
and (n11529,n11201,n11246);
and (n11530,n11154,n11199);
xor (n11531,n11120,n11122);
and (n11532,n11531,n11533);
or (n11533,n11534,n11538,n11583);
and (n11534,n11535,n11537);
xor (n11535,n11536,n11199);
xor (n11536,n11154,n11175);
xor (n11537,n11123,n11125);
and (n11538,n11537,n11539);
or (n11539,n11540,n11544,n11582);
and (n11540,n11541,n11543);
xor (n11541,n11542,n11246);
xor (n11542,n11201,n11222);
xor (n11543,n11126,n11128);
and (n11544,n11543,n11545);
or (n11545,n11546,n11550,n11581);
and (n11546,n11547,n11549);
xor (n11547,n11548,n11293);
xor (n11548,n11248,n11269);
xor (n11549,n11129,n11131);
and (n11550,n11549,n11551);
or (n11551,n11552,n11556,n11580);
and (n11552,n11553,n11555);
xor (n11553,n11554,n11340);
xor (n11554,n11295,n11316);
xor (n11555,n11132,n11134);
and (n11556,n11555,n11557);
or (n11557,n11558,n11562,n11579);
and (n11558,n11559,n11561);
xor (n11559,n11560,n11385);
xor (n11560,n11342,n11363);
xor (n11561,n11135,n11137);
and (n11562,n11561,n11563);
or (n11563,n11564,n11568,n11578);
and (n11564,n11565,n11567);
xor (n11565,n11566,n11432);
xor (n11566,n11387,n11408);
xor (n11567,n11138,n11139);
and (n11568,n11567,n11569);
or (n11569,n11570,n11574,n11577);
and (n11570,n11571,n11573);
xor (n11571,n11572,n11479);
xor (n11572,n11434,n11455);
xor (n11573,n11140,n11143);
and (n11574,n11573,n11575);
and (n11575,n11576,n11144);
xor (n11576,n11480,n11501);
and (n11577,n11571,n11575);
and (n11578,n11565,n11569);
and (n11579,n11559,n11563);
and (n11580,n11553,n11557);
and (n11581,n11547,n11551);
and (n11582,n11541,n11545);
and (n11583,n11535,n11539);
and (n11584,n11152,n11533);
or (n11585,n11586,n11587,n11637);
xor (n11586,n9953,n11146);
and (n11587,n11149,n11588);
or (n11588,n11589,n11591,n11636);
and (n11589,n11590,n11531);
xor (n11590,n11147,n11148);
and (n11591,n11531,n11592);
or (n11592,n11593,n11595,n11635);
and (n11593,n11594,n11537);
xor (n11594,n11149,n11150);
and (n11595,n11537,n11596);
or (n11596,n11597,n11600,n11634);
and (n11597,n11598,n11543);
xor (n11598,n11599,n11533);
xor (n11599,n11152,n11531);
and (n11600,n11543,n11601);
or (n11601,n11602,n11605,n11633);
and (n11602,n11603,n11549);
xor (n11603,n11604,n11539);
xor (n11604,n11535,n11537);
and (n11605,n11549,n11606);
or (n11606,n11607,n11610,n11632);
and (n11607,n11608,n11555);
xor (n11608,n11609,n11545);
xor (n11609,n11541,n11543);
and (n11610,n11555,n11611);
or (n11611,n11612,n11615,n11631);
and (n11612,n11613,n11561);
xor (n11613,n11614,n11551);
xor (n11614,n11547,n11549);
and (n11615,n11561,n11616);
or (n11616,n11617,n11620,n11630);
and (n11617,n11618,n11567);
xor (n11618,n11619,n11557);
xor (n11619,n11553,n11555);
and (n11620,n11567,n11621);
or (n11621,n11622,n11625,n11629);
and (n11622,n11623,n11573);
xor (n11623,n11624,n11563);
xor (n11624,n11559,n11561);
and (n11625,n11573,n11626);
and (n11626,n11627,n11144);
xor (n11627,n11628,n11569);
xor (n11628,n11565,n11567);
and (n11629,n11623,n11626);
and (n11630,n11618,n11621);
and (n11631,n11613,n11616);
and (n11632,n11608,n11611);
and (n11633,n11603,n11606);
and (n11634,n11598,n11601);
and (n11635,n11594,n11596);
and (n11636,n11590,n11592);
and (n11637,n11586,n11588);
and (n11638,n11639,n11641);
xor (n11639,n11640,n11588);
xor (n11640,n11586,n11149);
and (n11641,n11642,n11644);
xor (n11642,n11643,n11592);
xor (n11643,n11590,n11531);
and (n11644,n11645,n11647);
xor (n11645,n11646,n11596);
xor (n11646,n11594,n11537);
and (n11647,n11648,n11650);
xor (n11648,n11649,n11601);
xor (n11649,n11598,n11543);
and (n11650,n11651,n11653);
xor (n11651,n11652,n11606);
xor (n11652,n11603,n11549);
and (n11653,n11654,n11656);
xor (n11654,n11655,n11611);
xor (n11655,n11608,n11555);
and (n11656,n11657,n11659);
xor (n11657,n11658,n11616);
xor (n11658,n11613,n11561);
xor (n11659,n11660,n11621);
xor (n11660,n11618,n11567);
wire s0n11661,s1n11661,notn11661;
or (n11661,s0n11661,s1n11661);
not(notn11661,n4861);
and (s0n11661,notn11661,1'b0);
and (s1n11661,n4861,n11662);
xor (n11662,n11663,n11665);
xor (n11663,n11145,n11664);
and (n11664,n11147,n11585);
and (n11665,n9950,n11638);
wire s0n11666,s1n11666,notn11666;
or (n11666,s0n11666,s1n11666);
not(notn11666,n4861);
and (s0n11666,notn11666,1'b0);
and (s1n11666,n4861,n11667);
xor (n11667,n11668,n11670);
xor (n11668,n11145,n11669);
and (n11669,n9953,n11664);
and (n11670,n11663,n11665);
or (n11671,1'b0,n11672,n11687,n11702,n11717);
and (n11672,n11673,n2718);
or (n11673,1'b0,n11674,n11680,n11686);
and (n11674,n11675,n4895);
or (n11675,1'b0,n11676,n11677,n11678,n11679);
and (n11676,n5088,n556);
and (n11677,n5092,n567);
and (n11678,n5095,n571);
and (n11679,n5098,n573);
and (n11680,n11681,n2944);
or (n11681,1'b0,n11682,n11683,n11684,n11685);
and (n11682,n6832,n556);
and (n11683,n6831,n567);
and (n11684,n6835,n571);
and (n11685,n6838,n573);
and (n11686,n9906,n4903);
and (n11687,n11688,n2730);
or (n11688,1'b0,n11689,n11695,n11701);
and (n11689,n11690,n4895);
or (n11690,1'b0,n11691,n11692,n11693,n11694);
and (n11691,n5103,n556);
and (n11692,n5106,n567);
and (n11693,n5109,n571);
and (n11694,n5112,n573);
and (n11695,n11696,n2944);
or (n11696,1'b0,n11697,n11698,n11699,n11700);
and (n11697,n6841,n556);
and (n11698,n6846,n567);
and (n11699,n6849,n571);
and (n11700,n6852,n573);
and (n11701,n9912,n4903);
and (n11702,n11703,n2742);
or (n11703,1'b0,n11704,n11710,n11716);
and (n11704,n11705,n4895);
or (n11705,1'b0,n11706,n11707,n11708,n11709);
and (n11706,n5117,n556);
and (n11707,n5121,n567);
and (n11708,n5124,n571);
and (n11709,n5127,n573);
and (n11710,n11711,n2944);
or (n11711,1'b0,n11712,n11713,n11714,n11715);
and (n11712,n5013,n556);
and (n11713,n5012,n567);
and (n11714,n5027,n571);
and (n11715,n5032,n573);
and (n11716,n9918,n4903);
and (n11717,n11718,n2752);
or (n11718,1'b0,n11719,n11725,n11731);
and (n11719,n11720,n4895);
or (n11720,1'b0,n11721,n11722,n11723,n11724);
and (n11721,n5132,n556);
and (n11722,n5135,n567);
and (n11723,n5138,n571);
and (n11724,n5141,n573);
and (n11725,n11726,n2944);
or (n11726,1'b0,n11727,n11728,n11729,n11730);
and (n11727,n5037,n556);
and (n11728,n5044,n567);
and (n11729,n5047,n571);
and (n11730,n5050,n573);
and (n11731,n9924,n4903);
or (n11732,1'b0,n11733,n13057,n13059,n13060);
and (n11733,n11734,n2893);
wire s0n11734,s1n11734,notn11734;
or (n11734,s0n11734,s1n11734);
not(notn11734,n2891);
and (s0n11734,notn11734,1'b0);
and (s1n11734,n2891,n11735);
wire s0n11735,s1n11735,notn11735;
or (n11735,s0n11735,s1n11735);
not(notn11735,n13046);
and (s0n11735,notn11735,n11736);
and (s1n11735,n13046,1'b0);
wire s0n11736,s1n11736,notn11736;
or (n11736,s0n11736,s1n11736);
not(notn11736,n13031);
and (s0n11736,notn11736,n11737);
and (s1n11736,n13031,1'b1);
wire s0n11737,s1n11737,notn11737;
or (n11737,s0n11737,s1n11737);
not(notn11737,n4966);
and (s0n11737,notn11737,n11738);
and (s1n11737,n4966,n12815);
wire s0n11738,s1n11738,notn11738;
or (n11738,s0n11738,s1n11738);
not(notn11738,n4966);
and (s0n11738,notn11738,n11739);
and (s1n11738,n4966,n12812);
xor (n11739,n11740,n12789);
xor (n11740,n11741,n12732);
xor (n11741,n11742,n12663);
xor (n11742,n11743,n12653);
xor (n11743,n11744,n12073);
xor (n11744,n11745,n11748);
xor (n11745,n7684,n11746);
wire s0n11746,s1n11746,notn11746;
or (n11746,s0n11746,s1n11746);
not(notn11746,n4966);
and (s0n11746,notn11746,1'b0);
and (s1n11746,n4966,n11747);
or (n11748,n11749,n11752,n12072);
and (n11749,n7691,n11750);
wire s0n11750,s1n11750,notn11750;
or (n11750,s0n11750,s1n11750);
not(notn11750,n4966);
and (s0n11750,notn11750,1'b0);
and (s1n11750,n4966,n11751);
and (n11752,n11750,n11753);
or (n11753,n11754,n11757,n12071);
and (n11754,n6019,n11755);
wire s0n11755,s1n11755,notn11755;
or (n11755,s0n11755,s1n11755);
not(notn11755,n4966);
and (s0n11755,notn11755,1'b0);
and (s1n11755,n4966,n11756);
and (n11757,n11755,n11758);
or (n11758,n11759,n11762,n12070);
and (n11759,n6025,n11760);
wire s0n11760,s1n11760,notn11760;
or (n11760,s0n11760,s1n11760);
not(notn11760,n4966);
and (s0n11760,notn11760,1'b0);
and (s1n11760,n4966,n11761);
and (n11762,n11760,n11763);
or (n11763,n11764,n11767,n12069);
and (n11764,n6032,n11765);
wire s0n11765,s1n11765,notn11765;
or (n11765,s0n11765,s1n11765);
not(notn11765,n4966);
and (s0n11765,notn11765,1'b0);
and (s1n11765,n4966,n11766);
and (n11767,n11765,n11768);
or (n11768,n11769,n11804,n12068);
and (n11769,n6039,n11770);
wire s0n11770,s1n11770,notn11770;
or (n11770,s0n11770,s1n11770);
not(notn11770,n4966);
and (s0n11770,notn11770,n11771);
and (s1n11770,n4966,n11803);
or (n11771,1'b0,n11772,n11787,n11801,n11802);
and (n11772,n11773,n2718);
or (n11773,1'b0,n11774,n11778,n11781,n11784);
and (n11774,n11775,n5016);
wire s0n11775,s1n11775,notn11775;
or (n11775,s0n11775,s1n11775);
not(notn11775,n5014);
and (s0n11775,notn11775,n11776);
and (s1n11775,n5014,n11777);
and (n11778,n11779,n5028);
wire s0n11779,s1n11779,notn11779;
or (n11779,s0n11779,s1n11779);
not(notn11779,n5014);
and (s0n11779,notn11779,n11780);
and (s1n11779,n5014,n11776);
and (n11781,n11782,n5033);
wire s0n11782,s1n11782,notn11782;
or (n11782,s0n11782,s1n11782);
not(notn11782,n5014);
and (s0n11782,notn11782,n11783);
and (s1n11782,n5014,n11780);
and (n11784,n11785,n5038);
wire s0n11785,s1n11785,notn11785;
or (n11785,s0n11785,s1n11785);
not(notn11785,n5014);
and (s0n11785,notn11785,n11786);
and (s1n11785,n5014,n11783);
and (n11787,n11788,n2730);
or (n11788,1'b0,n11789,n11792,n11795,n11798);
and (n11789,n11790,n5016);
wire s0n11790,s1n11790,notn11790;
or (n11790,s0n11790,s1n11790);
not(notn11790,n5014);
and (s0n11790,notn11790,n11791);
and (s1n11790,n5014,n11786);
and (n11792,n11793,n5028);
wire s0n11793,s1n11793,notn11793;
or (n11793,s0n11793,s1n11793);
not(notn11793,n5014);
and (s0n11793,notn11793,n11794);
and (s1n11793,n5014,n11791);
and (n11795,n11796,n5033);
wire s0n11796,s1n11796,notn11796;
or (n11796,s0n11796,s1n11796);
not(notn11796,n5014);
and (s0n11796,notn11796,n11797);
and (s1n11796,n5014,n11794);
and (n11798,n11799,n5038);
wire s0n11799,s1n11799,notn11799;
or (n11799,s0n11799,s1n11799);
not(notn11799,n5014);
and (s0n11799,notn11799,n11800);
and (s1n11799,n5014,n11797);
and (n11801,n6085,n2742);
and (n11802,n6095,n2752);
and (n11804,n11770,n11805);
or (n11805,n11806,n11841,n12067);
and (n11806,n6128,n11807);
wire s0n11807,s1n11807,notn11807;
or (n11807,s0n11807,s1n11807);
not(notn11807,n4966);
and (s0n11807,notn11807,n11808);
and (s1n11807,n4966,n11840);
or (n11808,1'b0,n11809,n11824,n11838,n11839);
and (n11809,n11810,n2718);
or (n11810,1'b0,n11811,n11815,n11818,n11821);
and (n11811,n11812,n5016);
wire s0n11812,s1n11812,notn11812;
or (n11812,s0n11812,s1n11812);
not(notn11812,n5014);
and (s0n11812,notn11812,n11813);
and (s1n11812,n5014,n11814);
and (n11815,n11816,n5028);
wire s0n11816,s1n11816,notn11816;
or (n11816,s0n11816,s1n11816);
not(notn11816,n5014);
and (s0n11816,notn11816,n11817);
and (s1n11816,n5014,n11813);
and (n11818,n11819,n5033);
wire s0n11819,s1n11819,notn11819;
or (n11819,s0n11819,s1n11819);
not(notn11819,n5014);
and (s0n11819,notn11819,n11820);
and (s1n11819,n5014,n11817);
and (n11821,n11822,n5038);
wire s0n11822,s1n11822,notn11822;
or (n11822,s0n11822,s1n11822);
not(notn11822,n5014);
and (s0n11822,notn11822,n11823);
and (s1n11822,n5014,n11820);
and (n11824,n11825,n2730);
or (n11825,1'b0,n11826,n11829,n11832,n11835);
and (n11826,n11827,n5016);
wire s0n11827,s1n11827,notn11827;
or (n11827,s0n11827,s1n11827);
not(notn11827,n5014);
and (s0n11827,notn11827,n11828);
and (s1n11827,n5014,n11823);
and (n11829,n11830,n5028);
wire s0n11830,s1n11830,notn11830;
or (n11830,s0n11830,s1n11830);
not(notn11830,n5014);
and (s0n11830,notn11830,n11831);
and (s1n11830,n5014,n11828);
and (n11832,n11833,n5033);
wire s0n11833,s1n11833,notn11833;
or (n11833,s0n11833,s1n11833);
not(notn11833,n5014);
and (s0n11833,notn11833,n11834);
and (s1n11833,n5014,n11831);
and (n11835,n11836,n5038);
wire s0n11836,s1n11836,notn11836;
or (n11836,s0n11836,s1n11836);
not(notn11836,n5014);
and (s0n11836,notn11836,n11837);
and (s1n11836,n5014,n11834);
and (n11838,n6174,n2742);
and (n11839,n6184,n2752);
and (n11841,n11807,n11842);
or (n11842,n11843,n11878,n12066);
and (n11843,n6217,n11844);
wire s0n11844,s1n11844,notn11844;
or (n11844,s0n11844,s1n11844);
not(notn11844,n4966);
and (s0n11844,notn11844,n11845);
and (s1n11844,n4966,n11877);
or (n11845,1'b0,n11846,n11861,n11875,n11876);
and (n11846,n11847,n2718);
or (n11847,1'b0,n11848,n11852,n11855,n11858);
and (n11848,n11849,n5016);
wire s0n11849,s1n11849,notn11849;
or (n11849,s0n11849,s1n11849);
not(notn11849,n5014);
and (s0n11849,notn11849,n11850);
and (s1n11849,n5014,n11851);
and (n11852,n11853,n5028);
wire s0n11853,s1n11853,notn11853;
or (n11853,s0n11853,s1n11853);
not(notn11853,n5014);
and (s0n11853,notn11853,n11854);
and (s1n11853,n5014,n11850);
and (n11855,n11856,n5033);
wire s0n11856,s1n11856,notn11856;
or (n11856,s0n11856,s1n11856);
not(notn11856,n5014);
and (s0n11856,notn11856,n11857);
and (s1n11856,n5014,n11854);
and (n11858,n11859,n5038);
wire s0n11859,s1n11859,notn11859;
or (n11859,s0n11859,s1n11859);
not(notn11859,n5014);
and (s0n11859,notn11859,n11860);
and (s1n11859,n5014,n11857);
and (n11861,n11862,n2730);
or (n11862,1'b0,n11863,n11866,n11869,n11872);
and (n11863,n11864,n5016);
wire s0n11864,s1n11864,notn11864;
or (n11864,s0n11864,s1n11864);
not(notn11864,n5014);
and (s0n11864,notn11864,n11865);
and (s1n11864,n5014,n11860);
and (n11866,n11867,n5028);
wire s0n11867,s1n11867,notn11867;
or (n11867,s0n11867,s1n11867);
not(notn11867,n5014);
and (s0n11867,notn11867,n11868);
and (s1n11867,n5014,n11865);
and (n11869,n11870,n5033);
wire s0n11870,s1n11870,notn11870;
or (n11870,s0n11870,s1n11870);
not(notn11870,n5014);
and (s0n11870,notn11870,n11871);
and (s1n11870,n5014,n11868);
and (n11872,n11873,n5038);
wire s0n11873,s1n11873,notn11873;
or (n11873,s0n11873,s1n11873);
not(notn11873,n5014);
and (s0n11873,notn11873,n11874);
and (s1n11873,n5014,n11871);
and (n11875,n6263,n2742);
and (n11876,n6273,n2752);
and (n11878,n11844,n11879);
or (n11879,n11880,n11915,n12065);
and (n11880,n6306,n11881);
wire s0n11881,s1n11881,notn11881;
or (n11881,s0n11881,s1n11881);
not(notn11881,n4966);
and (s0n11881,notn11881,n11882);
and (s1n11881,n4966,n11914);
or (n11882,1'b0,n11883,n11898,n11912,n11913);
and (n11883,n11884,n2718);
or (n11884,1'b0,n11885,n11889,n11892,n11895);
and (n11885,n11886,n5016);
wire s0n11886,s1n11886,notn11886;
or (n11886,s0n11886,s1n11886);
not(notn11886,n5014);
and (s0n11886,notn11886,n11887);
and (s1n11886,n5014,n11888);
and (n11889,n11890,n5028);
wire s0n11890,s1n11890,notn11890;
or (n11890,s0n11890,s1n11890);
not(notn11890,n5014);
and (s0n11890,notn11890,n11891);
and (s1n11890,n5014,n11887);
and (n11892,n11893,n5033);
wire s0n11893,s1n11893,notn11893;
or (n11893,s0n11893,s1n11893);
not(notn11893,n5014);
and (s0n11893,notn11893,n11894);
and (s1n11893,n5014,n11891);
and (n11895,n11896,n5038);
wire s0n11896,s1n11896,notn11896;
or (n11896,s0n11896,s1n11896);
not(notn11896,n5014);
and (s0n11896,notn11896,n11897);
and (s1n11896,n5014,n11894);
and (n11898,n11899,n2730);
or (n11899,1'b0,n11900,n11903,n11906,n11909);
and (n11900,n11901,n5016);
wire s0n11901,s1n11901,notn11901;
or (n11901,s0n11901,s1n11901);
not(notn11901,n5014);
and (s0n11901,notn11901,n11902);
and (s1n11901,n5014,n11897);
and (n11903,n11904,n5028);
wire s0n11904,s1n11904,notn11904;
or (n11904,s0n11904,s1n11904);
not(notn11904,n5014);
and (s0n11904,notn11904,n11905);
and (s1n11904,n5014,n11902);
and (n11906,n11907,n5033);
wire s0n11907,s1n11907,notn11907;
or (n11907,s0n11907,s1n11907);
not(notn11907,n5014);
and (s0n11907,notn11907,n11908);
and (s1n11907,n5014,n11905);
and (n11909,n11910,n5038);
wire s0n11910,s1n11910,notn11910;
or (n11910,s0n11910,s1n11910);
not(notn11910,n5014);
and (s0n11910,notn11910,n11911);
and (s1n11910,n5014,n11908);
and (n11912,n6352,n2742);
and (n11913,n6362,n2752);
and (n11915,n11881,n11916);
or (n11916,n11917,n11952,n12064);
and (n11917,n6395,n11918);
wire s0n11918,s1n11918,notn11918;
or (n11918,s0n11918,s1n11918);
not(notn11918,n4966);
and (s0n11918,notn11918,n11919);
and (s1n11918,n4966,n11951);
or (n11919,1'b0,n11920,n11935,n11949,n11950);
and (n11920,n11921,n2718);
or (n11921,1'b0,n11922,n11926,n11929,n11932);
and (n11922,n11923,n5016);
wire s0n11923,s1n11923,notn11923;
or (n11923,s0n11923,s1n11923);
not(notn11923,n5014);
and (s0n11923,notn11923,n11924);
and (s1n11923,n5014,n11925);
and (n11926,n11927,n5028);
wire s0n11927,s1n11927,notn11927;
or (n11927,s0n11927,s1n11927);
not(notn11927,n5014);
and (s0n11927,notn11927,n11928);
and (s1n11927,n5014,n11924);
and (n11929,n11930,n5033);
wire s0n11930,s1n11930,notn11930;
or (n11930,s0n11930,s1n11930);
not(notn11930,n5014);
and (s0n11930,notn11930,n11931);
and (s1n11930,n5014,n11928);
and (n11932,n11933,n5038);
wire s0n11933,s1n11933,notn11933;
or (n11933,s0n11933,s1n11933);
not(notn11933,n5014);
and (s0n11933,notn11933,n11934);
and (s1n11933,n5014,n11931);
and (n11935,n11936,n2730);
or (n11936,1'b0,n11937,n11940,n11943,n11946);
and (n11937,n11938,n5016);
wire s0n11938,s1n11938,notn11938;
or (n11938,s0n11938,s1n11938);
not(notn11938,n5014);
and (s0n11938,notn11938,n11939);
and (s1n11938,n5014,n11934);
and (n11940,n11941,n5028);
wire s0n11941,s1n11941,notn11941;
or (n11941,s0n11941,s1n11941);
not(notn11941,n5014);
and (s0n11941,notn11941,n11942);
and (s1n11941,n5014,n11939);
and (n11943,n11944,n5033);
wire s0n11944,s1n11944,notn11944;
or (n11944,s0n11944,s1n11944);
not(notn11944,n5014);
and (s0n11944,notn11944,n11945);
and (s1n11944,n5014,n11942);
and (n11946,n11947,n5038);
wire s0n11947,s1n11947,notn11947;
or (n11947,s0n11947,s1n11947);
not(notn11947,n5014);
and (s0n11947,notn11947,n11948);
and (s1n11947,n5014,n11945);
and (n11949,n6441,n2742);
and (n11950,n6451,n2752);
and (n11952,n11918,n11953);
or (n11953,n11954,n11989,n12063);
and (n11954,n6484,n11955);
wire s0n11955,s1n11955,notn11955;
or (n11955,s0n11955,s1n11955);
not(notn11955,n4966);
and (s0n11955,notn11955,n11956);
and (s1n11955,n4966,n11988);
or (n11956,1'b0,n11957,n11972,n11986,n11987);
and (n11957,n11958,n2718);
or (n11958,1'b0,n11959,n11963,n11966,n11969);
and (n11959,n11960,n5016);
wire s0n11960,s1n11960,notn11960;
or (n11960,s0n11960,s1n11960);
not(notn11960,n5014);
and (s0n11960,notn11960,n11961);
and (s1n11960,n5014,n11962);
and (n11963,n11964,n5028);
wire s0n11964,s1n11964,notn11964;
or (n11964,s0n11964,s1n11964);
not(notn11964,n5014);
and (s0n11964,notn11964,n11965);
and (s1n11964,n5014,n11961);
and (n11966,n11967,n5033);
wire s0n11967,s1n11967,notn11967;
or (n11967,s0n11967,s1n11967);
not(notn11967,n5014);
and (s0n11967,notn11967,n11968);
and (s1n11967,n5014,n11965);
and (n11969,n11970,n5038);
wire s0n11970,s1n11970,notn11970;
or (n11970,s0n11970,s1n11970);
not(notn11970,n5014);
and (s0n11970,notn11970,n11971);
and (s1n11970,n5014,n11968);
and (n11972,n11973,n2730);
or (n11973,1'b0,n11974,n11977,n11980,n11983);
and (n11974,n11975,n5016);
wire s0n11975,s1n11975,notn11975;
or (n11975,s0n11975,s1n11975);
not(notn11975,n5014);
and (s0n11975,notn11975,n11976);
and (s1n11975,n5014,n11971);
and (n11977,n11978,n5028);
wire s0n11978,s1n11978,notn11978;
or (n11978,s0n11978,s1n11978);
not(notn11978,n5014);
and (s0n11978,notn11978,n11979);
and (s1n11978,n5014,n11976);
and (n11980,n11981,n5033);
wire s0n11981,s1n11981,notn11981;
or (n11981,s0n11981,s1n11981);
not(notn11981,n5014);
and (s0n11981,notn11981,n11982);
and (s1n11981,n5014,n11979);
and (n11983,n11984,n5038);
wire s0n11984,s1n11984,notn11984;
or (n11984,s0n11984,s1n11984);
not(notn11984,n5014);
and (s0n11984,notn11984,n11985);
and (s1n11984,n5014,n11982);
and (n11986,n6530,n2742);
and (n11987,n6540,n2752);
and (n11989,n11955,n11990);
or (n11990,n11991,n12026,n12062);
and (n11991,n6573,n11992);
wire s0n11992,s1n11992,notn11992;
or (n11992,s0n11992,s1n11992);
not(notn11992,n4966);
and (s0n11992,notn11992,n11993);
and (s1n11992,n4966,n12025);
or (n11993,1'b0,n11994,n12009,n12023,n12024);
and (n11994,n11995,n2718);
or (n11995,1'b0,n11996,n12000,n12003,n12006);
and (n11996,n11997,n5016);
wire s0n11997,s1n11997,notn11997;
or (n11997,s0n11997,s1n11997);
not(notn11997,n5014);
and (s0n11997,notn11997,n11998);
and (s1n11997,n5014,n11999);
and (n12000,n12001,n5028);
wire s0n12001,s1n12001,notn12001;
or (n12001,s0n12001,s1n12001);
not(notn12001,n5014);
and (s0n12001,notn12001,n12002);
and (s1n12001,n5014,n11998);
and (n12003,n12004,n5033);
wire s0n12004,s1n12004,notn12004;
or (n12004,s0n12004,s1n12004);
not(notn12004,n5014);
and (s0n12004,notn12004,n12005);
and (s1n12004,n5014,n12002);
and (n12006,n12007,n5038);
wire s0n12007,s1n12007,notn12007;
or (n12007,s0n12007,s1n12007);
not(notn12007,n5014);
and (s0n12007,notn12007,n12008);
and (s1n12007,n5014,n12005);
and (n12009,n12010,n2730);
or (n12010,1'b0,n12011,n12014,n12017,n12020);
and (n12011,n12012,n5016);
wire s0n12012,s1n12012,notn12012;
or (n12012,s0n12012,s1n12012);
not(notn12012,n5014);
and (s0n12012,notn12012,n12013);
and (s1n12012,n5014,n12008);
and (n12014,n12015,n5028);
wire s0n12015,s1n12015,notn12015;
or (n12015,s0n12015,s1n12015);
not(notn12015,n5014);
and (s0n12015,notn12015,n12016);
and (s1n12015,n5014,n12013);
and (n12017,n12018,n5033);
wire s0n12018,s1n12018,notn12018;
or (n12018,s0n12018,s1n12018);
not(notn12018,n5014);
and (s0n12018,notn12018,n12019);
and (s1n12018,n5014,n12016);
and (n12020,n12021,n5038);
wire s0n12021,s1n12021,notn12021;
or (n12021,s0n12021,s1n12021);
not(notn12021,n5014);
and (s0n12021,notn12021,n12022);
and (s1n12021,n5014,n12019);
and (n12023,n6619,n2742);
and (n12024,n6629,n2752);
and (n12026,n11992,n12027);
and (n12027,n6661,n12028);
wire s0n12028,s1n12028,notn12028;
or (n12028,s0n12028,s1n12028);
not(notn12028,n4966);
and (s0n12028,notn12028,n12029);
and (s1n12028,n4966,n12061);
or (n12029,1'b0,n12030,n12045,n12059,n12060);
and (n12030,n12031,n2718);
or (n12031,1'b0,n12032,n12036,n12039,n12042);
and (n12032,n12033,n5016);
wire s0n12033,s1n12033,notn12033;
or (n12033,s0n12033,s1n12033);
not(notn12033,n5014);
and (s0n12033,notn12033,n12034);
and (s1n12033,n5014,n12035);
and (n12036,n12037,n5028);
wire s0n12037,s1n12037,notn12037;
or (n12037,s0n12037,s1n12037);
not(notn12037,n5014);
and (s0n12037,notn12037,n12038);
and (s1n12037,n5014,n12034);
and (n12039,n12040,n5033);
wire s0n12040,s1n12040,notn12040;
or (n12040,s0n12040,s1n12040);
not(notn12040,n5014);
and (s0n12040,notn12040,n12041);
and (s1n12040,n5014,n12038);
and (n12042,n12043,n5038);
wire s0n12043,s1n12043,notn12043;
or (n12043,s0n12043,s1n12043);
not(notn12043,n5014);
and (s0n12043,notn12043,n12044);
and (s1n12043,n5014,n12041);
and (n12045,n12046,n2730);
or (n12046,1'b0,n12047,n12050,n12053,n12056);
and (n12047,n12048,n5016);
wire s0n12048,s1n12048,notn12048;
or (n12048,s0n12048,s1n12048);
not(notn12048,n5014);
and (s0n12048,notn12048,n12049);
and (s1n12048,n5014,n12044);
and (n12050,n12051,n5028);
wire s0n12051,s1n12051,notn12051;
or (n12051,s0n12051,s1n12051);
not(notn12051,n5014);
and (s0n12051,notn12051,n12052);
and (s1n12051,n5014,n12049);
and (n12053,n12054,n5033);
wire s0n12054,s1n12054,notn12054;
or (n12054,s0n12054,s1n12054);
not(notn12054,n5014);
and (s0n12054,notn12054,n12055);
and (s1n12054,n5014,n12052);
and (n12056,n12057,n5038);
wire s0n12057,s1n12057,notn12057;
or (n12057,s0n12057,s1n12057);
not(notn12057,n5014);
and (s0n12057,notn12057,n12058);
and (s1n12057,n5014,n12055);
and (n12059,n6707,n2742);
and (n12060,n6717,n2752);
and (n12062,n6573,n12027);
and (n12063,n6484,n11990);
and (n12064,n6395,n11953);
and (n12065,n6306,n11916);
and (n12066,n6217,n11879);
and (n12067,n6128,n11842);
and (n12068,n6039,n11805);
and (n12069,n6032,n11768);
and (n12070,n6025,n11763);
and (n12071,n6019,n11758);
and (n12072,n7691,n11753);
xor (n12073,n12074,n12618);
xor (n12074,n12075,n12459);
xor (n12075,n12076,n12115);
xor (n12076,n12077,n12078);
xor (n12077,n6774,n4987);
or (n12078,n12079,n12080,n12114);
and (n12079,n6781,n4994);
and (n12080,n4994,n12081);
or (n12081,n12082,n12083,n12113);
and (n12082,n6788,n5001);
and (n12083,n5001,n12084);
or (n12084,n12085,n12086,n12112);
and (n12085,n6825,n5082);
and (n12086,n5082,n12087);
or (n12087,n12088,n12089,n12111);
and (n12088,n6894,n5205);
and (n12089,n5205,n12090);
or (n12090,n12091,n12092,n12110);
and (n12091,n6963,n5328);
and (n12092,n5328,n12093);
or (n12093,n12094,n12095,n12109);
and (n12094,n7032,n5451);
and (n12095,n5451,n12096);
or (n12096,n12097,n12098,n12108);
and (n12097,n7101,n5574);
and (n12098,n5574,n12099);
or (n12099,n12100,n12101,n12107);
and (n12100,n7170,n5697);
and (n12101,n5697,n12102);
or (n12102,n12103,n12104,n12106);
and (n12103,n7239,n5820);
and (n12104,n5820,n12105);
and (n12105,n7307,n5942);
and (n12106,n7239,n12105);
and (n12107,n7170,n12102);
and (n12108,n7101,n12099);
and (n12109,n7032,n12096);
and (n12110,n6963,n12093);
and (n12111,n6894,n12090);
and (n12112,n6825,n12087);
and (n12113,n6788,n12084);
and (n12114,n6781,n12081);
not (n12115,n12116);
nor (n12116,n12117,n12456);
and (n12117,n12118,n12453);
nand (n12118,n12119,n12437);
or (n12119,n12120,n12135);
nand (n12120,n12121,n12128);
and (n12121,n12122,n12125);
or (n12122,n6034,n12123);
wire s0n12123,s1n12123,notn12123;
or (n12123,s0n12123,s1n12123);
not(notn12123,n4966);
and (s0n12123,notn12123,1'b0);
and (s1n12123,n4966,n12124);
or (n12125,n6027,n12126);
wire s0n12126,s1n12126,notn12126;
or (n12126,s0n12126,s1n12126);
not(notn12126,n4966);
and (s0n12126,notn12126,1'b0);
and (s1n12126,n4966,n12127);
nor (n12128,n12129,n12132);
nor (n12129,n7693,n12130);
wire s0n12130,s1n12130,notn12130;
or (n12130,s0n12130,s1n12130);
not(notn12130,n4966);
and (s0n12130,notn12130,1'b0);
and (s1n12130,n4966,n12131);
nor (n12132,n6021,n12133);
wire s0n12133,s1n12133,notn12133;
or (n12133,s0n12133,s1n12133);
not(notn12133,n4966);
and (s0n12133,notn12133,1'b0);
and (s1n12133,n4966,n12134);
not (n12135,n12136);
or (n12136,n12137,n12172,n12436);
and (n12137,n6082,n12138);
wire s0n12138,s1n12138,notn12138;
or (n12138,s0n12138,s1n12138);
not(notn12138,n4966);
and (s0n12138,notn12138,n12139);
and (s1n12138,n4966,n12171);
or (n12139,1'b0,n12140,n12155,n12169,n12170);
and (n12140,n12141,n2718);
or (n12141,1'b0,n12142,n12146,n12149,n12152);
and (n12142,n12143,n5016);
wire s0n12143,s1n12143,notn12143;
or (n12143,s0n12143,s1n12143);
not(notn12143,n5014);
and (s0n12143,notn12143,n12144);
and (s1n12143,n5014,n12145);
and (n12146,n12147,n5028);
wire s0n12147,s1n12147,notn12147;
or (n12147,s0n12147,s1n12147);
not(notn12147,n5014);
and (s0n12147,notn12147,n12148);
and (s1n12147,n5014,n12144);
and (n12149,n12150,n5033);
wire s0n12150,s1n12150,notn12150;
or (n12150,s0n12150,s1n12150);
not(notn12150,n5014);
and (s0n12150,notn12150,n12151);
and (s1n12150,n5014,n12148);
and (n12152,n12153,n5038);
wire s0n12153,s1n12153,notn12153;
or (n12153,s0n12153,s1n12153);
not(notn12153,n5014);
and (s0n12153,notn12153,n12154);
and (s1n12153,n5014,n12151);
and (n12155,n12156,n2730);
or (n12156,1'b0,n12157,n12160,n12163,n12166);
and (n12157,n12158,n5016);
wire s0n12158,s1n12158,notn12158;
or (n12158,s0n12158,s1n12158);
not(notn12158,n5014);
and (s0n12158,notn12158,n12159);
and (s1n12158,n5014,n12154);
and (n12160,n12161,n5028);
wire s0n12161,s1n12161,notn12161;
or (n12161,s0n12161,s1n12161);
not(notn12161,n5014);
and (s0n12161,notn12161,n12162);
and (s1n12161,n5014,n12159);
and (n12163,n12164,n5033);
wire s0n12164,s1n12164,notn12164;
or (n12164,s0n12164,s1n12164);
not(notn12164,n5014);
and (s0n12164,notn12164,n12165);
and (s1n12164,n5014,n12162);
and (n12166,n12167,n5038);
wire s0n12167,s1n12167,notn12167;
or (n12167,s0n12167,s1n12167);
not(notn12167,n5014);
and (s0n12167,notn12167,n12168);
and (s1n12167,n5014,n12165);
and (n12169,n6042,n2742);
and (n12170,n6052,n2752);
and (n12172,n12138,n12173);
or (n12173,n12174,n12209,n12435);
and (n12174,n6171,n12175);
wire s0n12175,s1n12175,notn12175;
or (n12175,s0n12175,s1n12175);
not(notn12175,n4966);
and (s0n12175,notn12175,n12176);
and (s1n12175,n4966,n12208);
or (n12176,1'b0,n12177,n12192,n12206,n12207);
and (n12177,n12178,n2718);
or (n12178,1'b0,n12179,n12183,n12186,n12189);
and (n12179,n12180,n5016);
wire s0n12180,s1n12180,notn12180;
or (n12180,s0n12180,s1n12180);
not(notn12180,n5014);
and (s0n12180,notn12180,n12181);
and (s1n12180,n5014,n12182);
and (n12183,n12184,n5028);
wire s0n12184,s1n12184,notn12184;
or (n12184,s0n12184,s1n12184);
not(notn12184,n5014);
and (s0n12184,notn12184,n12185);
and (s1n12184,n5014,n12181);
and (n12186,n12187,n5033);
wire s0n12187,s1n12187,notn12187;
or (n12187,s0n12187,s1n12187);
not(notn12187,n5014);
and (s0n12187,notn12187,n12188);
and (s1n12187,n5014,n12185);
and (n12189,n12190,n5038);
wire s0n12190,s1n12190,notn12190;
or (n12190,s0n12190,s1n12190);
not(notn12190,n5014);
and (s0n12190,notn12190,n12191);
and (s1n12190,n5014,n12188);
and (n12192,n12193,n2730);
or (n12193,1'b0,n12194,n12197,n12200,n12203);
and (n12194,n12195,n5016);
wire s0n12195,s1n12195,notn12195;
or (n12195,s0n12195,s1n12195);
not(notn12195,n5014);
and (s0n12195,notn12195,n12196);
and (s1n12195,n5014,n12191);
and (n12197,n12198,n5028);
wire s0n12198,s1n12198,notn12198;
or (n12198,s0n12198,s1n12198);
not(notn12198,n5014);
and (s0n12198,notn12198,n12199);
and (s1n12198,n5014,n12196);
and (n12200,n12201,n5033);
wire s0n12201,s1n12201,notn12201;
or (n12201,s0n12201,s1n12201);
not(notn12201,n5014);
and (s0n12201,notn12201,n12202);
and (s1n12201,n5014,n12199);
and (n12203,n12204,n5038);
wire s0n12204,s1n12204,notn12204;
or (n12204,s0n12204,s1n12204);
not(notn12204,n5014);
and (s0n12204,notn12204,n12205);
and (s1n12204,n5014,n12202);
and (n12206,n6131,n2742);
and (n12207,n6141,n2752);
and (n12209,n12175,n12210);
or (n12210,n12211,n12246,n12434);
and (n12211,n6260,n12212);
wire s0n12212,s1n12212,notn12212;
or (n12212,s0n12212,s1n12212);
not(notn12212,n4966);
and (s0n12212,notn12212,n12213);
and (s1n12212,n4966,n12245);
or (n12213,1'b0,n12214,n12229,n12243,n12244);
and (n12214,n12215,n2718);
or (n12215,1'b0,n12216,n12220,n12223,n12226);
and (n12216,n12217,n5016);
wire s0n12217,s1n12217,notn12217;
or (n12217,s0n12217,s1n12217);
not(notn12217,n5014);
and (s0n12217,notn12217,n12218);
and (s1n12217,n5014,n12219);
and (n12220,n12221,n5028);
wire s0n12221,s1n12221,notn12221;
or (n12221,s0n12221,s1n12221);
not(notn12221,n5014);
and (s0n12221,notn12221,n12222);
and (s1n12221,n5014,n12218);
and (n12223,n12224,n5033);
wire s0n12224,s1n12224,notn12224;
or (n12224,s0n12224,s1n12224);
not(notn12224,n5014);
and (s0n12224,notn12224,n12225);
and (s1n12224,n5014,n12222);
and (n12226,n12227,n5038);
wire s0n12227,s1n12227,notn12227;
or (n12227,s0n12227,s1n12227);
not(notn12227,n5014);
and (s0n12227,notn12227,n12228);
and (s1n12227,n5014,n12225);
and (n12229,n12230,n2730);
or (n12230,1'b0,n12231,n12234,n12237,n12240);
and (n12231,n12232,n5016);
wire s0n12232,s1n12232,notn12232;
or (n12232,s0n12232,s1n12232);
not(notn12232,n5014);
and (s0n12232,notn12232,n12233);
and (s1n12232,n5014,n12228);
and (n12234,n12235,n5028);
wire s0n12235,s1n12235,notn12235;
or (n12235,s0n12235,s1n12235);
not(notn12235,n5014);
and (s0n12235,notn12235,n12236);
and (s1n12235,n5014,n12233);
and (n12237,n12238,n5033);
wire s0n12238,s1n12238,notn12238;
or (n12238,s0n12238,s1n12238);
not(notn12238,n5014);
and (s0n12238,notn12238,n12239);
and (s1n12238,n5014,n12236);
and (n12240,n12241,n5038);
wire s0n12241,s1n12241,notn12241;
or (n12241,s0n12241,s1n12241);
not(notn12241,n5014);
and (s0n12241,notn12241,n12242);
and (s1n12241,n5014,n12239);
and (n12243,n6220,n2742);
and (n12244,n6230,n2752);
and (n12246,n12212,n12247);
or (n12247,n12248,n12283,n12433);
and (n12248,n6349,n12249);
wire s0n12249,s1n12249,notn12249;
or (n12249,s0n12249,s1n12249);
not(notn12249,n4966);
and (s0n12249,notn12249,n12250);
and (s1n12249,n4966,n12282);
or (n12250,1'b0,n12251,n12266,n12280,n12281);
and (n12251,n12252,n2718);
or (n12252,1'b0,n12253,n12257,n12260,n12263);
and (n12253,n12254,n5016);
wire s0n12254,s1n12254,notn12254;
or (n12254,s0n12254,s1n12254);
not(notn12254,n5014);
and (s0n12254,notn12254,n12255);
and (s1n12254,n5014,n12256);
and (n12257,n12258,n5028);
wire s0n12258,s1n12258,notn12258;
or (n12258,s0n12258,s1n12258);
not(notn12258,n5014);
and (s0n12258,notn12258,n12259);
and (s1n12258,n5014,n12255);
and (n12260,n12261,n5033);
wire s0n12261,s1n12261,notn12261;
or (n12261,s0n12261,s1n12261);
not(notn12261,n5014);
and (s0n12261,notn12261,n12262);
and (s1n12261,n5014,n12259);
and (n12263,n12264,n5038);
wire s0n12264,s1n12264,notn12264;
or (n12264,s0n12264,s1n12264);
not(notn12264,n5014);
and (s0n12264,notn12264,n12265);
and (s1n12264,n5014,n12262);
and (n12266,n12267,n2730);
or (n12267,1'b0,n12268,n12271,n12274,n12277);
and (n12268,n12269,n5016);
wire s0n12269,s1n12269,notn12269;
or (n12269,s0n12269,s1n12269);
not(notn12269,n5014);
and (s0n12269,notn12269,n12270);
and (s1n12269,n5014,n12265);
and (n12271,n12272,n5028);
wire s0n12272,s1n12272,notn12272;
or (n12272,s0n12272,s1n12272);
not(notn12272,n5014);
and (s0n12272,notn12272,n12273);
and (s1n12272,n5014,n12270);
and (n12274,n12275,n5033);
wire s0n12275,s1n12275,notn12275;
or (n12275,s0n12275,s1n12275);
not(notn12275,n5014);
and (s0n12275,notn12275,n12276);
and (s1n12275,n5014,n12273);
and (n12277,n12278,n5038);
wire s0n12278,s1n12278,notn12278;
or (n12278,s0n12278,s1n12278);
not(notn12278,n5014);
and (s0n12278,notn12278,n12279);
and (s1n12278,n5014,n12276);
and (n12280,n6309,n2742);
and (n12281,n6319,n2752);
and (n12283,n12249,n12284);
or (n12284,n12285,n12320,n12432);
and (n12285,n6438,n12286);
wire s0n12286,s1n12286,notn12286;
or (n12286,s0n12286,s1n12286);
not(notn12286,n4966);
and (s0n12286,notn12286,n12287);
and (s1n12286,n4966,n12319);
or (n12287,1'b0,n12288,n12303,n12317,n12318);
and (n12288,n12289,n2718);
or (n12289,1'b0,n12290,n12294,n12297,n12300);
and (n12290,n12291,n5016);
wire s0n12291,s1n12291,notn12291;
or (n12291,s0n12291,s1n12291);
not(notn12291,n5014);
and (s0n12291,notn12291,n12292);
and (s1n12291,n5014,n12293);
and (n12294,n12295,n5028);
wire s0n12295,s1n12295,notn12295;
or (n12295,s0n12295,s1n12295);
not(notn12295,n5014);
and (s0n12295,notn12295,n12296);
and (s1n12295,n5014,n12292);
and (n12297,n12298,n5033);
wire s0n12298,s1n12298,notn12298;
or (n12298,s0n12298,s1n12298);
not(notn12298,n5014);
and (s0n12298,notn12298,n12299);
and (s1n12298,n5014,n12296);
and (n12300,n12301,n5038);
wire s0n12301,s1n12301,notn12301;
or (n12301,s0n12301,s1n12301);
not(notn12301,n5014);
and (s0n12301,notn12301,n12302);
and (s1n12301,n5014,n12299);
and (n12303,n12304,n2730);
or (n12304,1'b0,n12305,n12308,n12311,n12314);
and (n12305,n12306,n5016);
wire s0n12306,s1n12306,notn12306;
or (n12306,s0n12306,s1n12306);
not(notn12306,n5014);
and (s0n12306,notn12306,n12307);
and (s1n12306,n5014,n12302);
and (n12308,n12309,n5028);
wire s0n12309,s1n12309,notn12309;
or (n12309,s0n12309,s1n12309);
not(notn12309,n5014);
and (s0n12309,notn12309,n12310);
and (s1n12309,n5014,n12307);
and (n12311,n12312,n5033);
wire s0n12312,s1n12312,notn12312;
or (n12312,s0n12312,s1n12312);
not(notn12312,n5014);
and (s0n12312,notn12312,n12313);
and (s1n12312,n5014,n12310);
and (n12314,n12315,n5038);
wire s0n12315,s1n12315,notn12315;
or (n12315,s0n12315,s1n12315);
not(notn12315,n5014);
and (s0n12315,notn12315,n12316);
and (s1n12315,n5014,n12313);
and (n12317,n6398,n2742);
and (n12318,n6408,n2752);
and (n12320,n12286,n12321);
or (n12321,n12322,n12357,n12431);
and (n12322,n6527,n12323);
wire s0n12323,s1n12323,notn12323;
or (n12323,s0n12323,s1n12323);
not(notn12323,n4966);
and (s0n12323,notn12323,n12324);
and (s1n12323,n4966,n12356);
or (n12324,1'b0,n12325,n12340,n12354,n12355);
and (n12325,n12326,n2718);
or (n12326,1'b0,n12327,n12331,n12334,n12337);
and (n12327,n12328,n5016);
wire s0n12328,s1n12328,notn12328;
or (n12328,s0n12328,s1n12328);
not(notn12328,n5014);
and (s0n12328,notn12328,n12329);
and (s1n12328,n5014,n12330);
and (n12331,n12332,n5028);
wire s0n12332,s1n12332,notn12332;
or (n12332,s0n12332,s1n12332);
not(notn12332,n5014);
and (s0n12332,notn12332,n12333);
and (s1n12332,n5014,n12329);
and (n12334,n12335,n5033);
wire s0n12335,s1n12335,notn12335;
or (n12335,s0n12335,s1n12335);
not(notn12335,n5014);
and (s0n12335,notn12335,n12336);
and (s1n12335,n5014,n12333);
and (n12337,n12338,n5038);
wire s0n12338,s1n12338,notn12338;
or (n12338,s0n12338,s1n12338);
not(notn12338,n5014);
and (s0n12338,notn12338,n12339);
and (s1n12338,n5014,n12336);
and (n12340,n12341,n2730);
or (n12341,1'b0,n12342,n12345,n12348,n12351);
and (n12342,n12343,n5016);
wire s0n12343,s1n12343,notn12343;
or (n12343,s0n12343,s1n12343);
not(notn12343,n5014);
and (s0n12343,notn12343,n12344);
and (s1n12343,n5014,n12339);
and (n12345,n12346,n5028);
wire s0n12346,s1n12346,notn12346;
or (n12346,s0n12346,s1n12346);
not(notn12346,n5014);
and (s0n12346,notn12346,n12347);
and (s1n12346,n5014,n12344);
and (n12348,n12349,n5033);
wire s0n12349,s1n12349,notn12349;
or (n12349,s0n12349,s1n12349);
not(notn12349,n5014);
and (s0n12349,notn12349,n12350);
and (s1n12349,n5014,n12347);
and (n12351,n12352,n5038);
wire s0n12352,s1n12352,notn12352;
or (n12352,s0n12352,s1n12352);
not(notn12352,n5014);
and (s0n12352,notn12352,n12353);
and (s1n12352,n5014,n12350);
and (n12354,n6487,n2742);
and (n12355,n6497,n2752);
and (n12357,n12323,n12358);
or (n12358,n12359,n12394,n12430);
and (n12359,n6616,n12360);
wire s0n12360,s1n12360,notn12360;
or (n12360,s0n12360,s1n12360);
not(notn12360,n4966);
and (s0n12360,notn12360,n12361);
and (s1n12360,n4966,n12393);
or (n12361,1'b0,n12362,n12377,n12391,n12392);
and (n12362,n12363,n2718);
or (n12363,1'b0,n12364,n12368,n12371,n12374);
and (n12364,n12365,n5016);
wire s0n12365,s1n12365,notn12365;
or (n12365,s0n12365,s1n12365);
not(notn12365,n5014);
and (s0n12365,notn12365,n12366);
and (s1n12365,n5014,n12367);
and (n12368,n12369,n5028);
wire s0n12369,s1n12369,notn12369;
or (n12369,s0n12369,s1n12369);
not(notn12369,n5014);
and (s0n12369,notn12369,n12370);
and (s1n12369,n5014,n12366);
and (n12371,n12372,n5033);
wire s0n12372,s1n12372,notn12372;
or (n12372,s0n12372,s1n12372);
not(notn12372,n5014);
and (s0n12372,notn12372,n12373);
and (s1n12372,n5014,n12370);
and (n12374,n12375,n5038);
wire s0n12375,s1n12375,notn12375;
or (n12375,s0n12375,s1n12375);
not(notn12375,n5014);
and (s0n12375,notn12375,n12376);
and (s1n12375,n5014,n12373);
and (n12377,n12378,n2730);
or (n12378,1'b0,n12379,n12382,n12385,n12388);
and (n12379,n12380,n5016);
wire s0n12380,s1n12380,notn12380;
or (n12380,s0n12380,s1n12380);
not(notn12380,n5014);
and (s0n12380,notn12380,n12381);
and (s1n12380,n5014,n12376);
and (n12382,n12383,n5028);
wire s0n12383,s1n12383,notn12383;
or (n12383,s0n12383,s1n12383);
not(notn12383,n5014);
and (s0n12383,notn12383,n12384);
and (s1n12383,n5014,n12381);
and (n12385,n12386,n5033);
wire s0n12386,s1n12386,notn12386;
or (n12386,s0n12386,s1n12386);
not(notn12386,n5014);
and (s0n12386,notn12386,n12387);
and (s1n12386,n5014,n12384);
and (n12388,n12389,n5038);
wire s0n12389,s1n12389,notn12389;
or (n12389,s0n12389,s1n12389);
not(notn12389,n5014);
and (s0n12389,notn12389,n12390);
and (s1n12389,n5014,n12387);
and (n12391,n6576,n2742);
and (n12392,n6586,n2752);
and (n12394,n12360,n12395);
and (n12395,n6704,n12396);
wire s0n12396,s1n12396,notn12396;
or (n12396,s0n12396,s1n12396);
not(notn12396,n4966);
and (s0n12396,notn12396,n12397);
and (s1n12396,n4966,n12429);
or (n12397,1'b0,n12398,n12413,n12427,n12428);
and (n12398,n12399,n2718);
or (n12399,1'b0,n12400,n12404,n12407,n12410);
and (n12400,n12401,n5016);
wire s0n12401,s1n12401,notn12401;
or (n12401,s0n12401,s1n12401);
not(notn12401,n5014);
and (s0n12401,notn12401,n12402);
and (s1n12401,n5014,n12403);
and (n12404,n12405,n5028);
wire s0n12405,s1n12405,notn12405;
or (n12405,s0n12405,s1n12405);
not(notn12405,n5014);
and (s0n12405,notn12405,n12406);
and (s1n12405,n5014,n12402);
and (n12407,n12408,n5033);
wire s0n12408,s1n12408,notn12408;
or (n12408,s0n12408,s1n12408);
not(notn12408,n5014);
and (s0n12408,notn12408,n12409);
and (s1n12408,n5014,n12406);
and (n12410,n12411,n5038);
wire s0n12411,s1n12411,notn12411;
or (n12411,s0n12411,s1n12411);
not(notn12411,n5014);
and (s0n12411,notn12411,n12412);
and (s1n12411,n5014,n12409);
and (n12413,n12414,n2730);
or (n12414,1'b0,n12415,n12418,n12421,n12424);
and (n12415,n12416,n5016);
wire s0n12416,s1n12416,notn12416;
or (n12416,s0n12416,s1n12416);
not(notn12416,n5014);
and (s0n12416,notn12416,n12417);
and (s1n12416,n5014,n12412);
and (n12418,n12419,n5028);
wire s0n12419,s1n12419,notn12419;
or (n12419,s0n12419,s1n12419);
not(notn12419,n5014);
and (s0n12419,notn12419,n12420);
and (s1n12419,n5014,n12417);
and (n12421,n12422,n5033);
wire s0n12422,s1n12422,notn12422;
or (n12422,s0n12422,s1n12422);
not(notn12422,n5014);
and (s0n12422,notn12422,n12423);
and (s1n12422,n5014,n12420);
and (n12424,n12425,n5038);
wire s0n12425,s1n12425,notn12425;
or (n12425,s0n12425,s1n12425);
not(notn12425,n5014);
and (s0n12425,notn12425,n12426);
and (s1n12425,n5014,n12423);
and (n12427,n6664,n2742);
and (n12428,n6674,n2752);
and (n12430,n6616,n12395);
and (n12431,n6527,n12358);
and (n12432,n6438,n12321);
and (n12433,n6349,n12284);
and (n12434,n6260,n12247);
and (n12435,n6171,n12210);
and (n12436,n6082,n12173);
not (n12437,n12438);
nand (n12438,n12439,n12448);
or (n12439,n12440,n12441);
not (n12440,n12128);
not (n12441,n12442);
nand (n12442,n12443,n12447);
or (n12443,n12444,n12445);
not (n12444,n12125);
not (n12445,n12446);
and (n12446,n6034,n12123);
nand (n12447,n6027,n12126);
nor (n12448,n12449,n12452);
and (n12449,n12450,n12451);
not (n12450,n12129);
and (n12451,n6021,n12133);
and (n12452,n7693,n12130);
xor (n12453,n7686,n12454);
wire s0n12454,s1n12454,notn12454;
or (n12454,s0n12454,s1n12454);
not(notn12454,n4966);
and (s0n12454,notn12454,1'b0);
and (s1n12454,n4966,n12455);
and (n12456,n12457,n12458);
not (n12457,n12118);
not (n12458,n12453);
or (n12459,n12460,n12477,n12617);
and (n12460,n12461,n12463);
xor (n12461,n12462,n12081);
xor (n12462,n6781,n4994);
not (n12463,n12464);
nand (n12464,n12465,n12476);
or (n12465,n12466,n12468);
not (n12466,n12467);
xor (n12467,n7693,n12130);
nand (n12468,n12469,n12473);
or (n12469,n12470,n12135);
not (n12470,n12471);
nor (n12471,n12472,n12132);
not (n12472,n12121);
nor (n12473,n12474,n12451);
and (n12474,n12442,n12475);
not (n12475,n12132);
nand (n12476,n12468,n12466);
and (n12477,n12463,n12478);
or (n12478,n12479,n12544,n12616);
and (n12479,n12480,n12482);
xor (n12480,n12481,n12084);
xor (n12481,n6788,n5001);
not (n12482,n12483);
xor (n12483,n12484,n12485);
xor (n12484,n6021,n12133);
nand (n12485,n12486,n12529);
or (n12486,n12487,n12508);
not (n12487,n12488);
and (n12488,n12489,n12501);
nor (n12489,n12490,n12497);
nand (n12490,n12491,n12494);
nand (n12491,n12492,n12493);
not (n12492,n6349);
not (n12493,n12249);
nand (n12494,n12495,n12496);
not (n12495,n6438);
not (n12496,n12286);
not (n12497,n12498);
nand (n12498,n12499,n12500);
not (n12499,n6082);
not (n12500,n12138);
not (n12501,n12502);
nor (n12502,n12503,n12505);
not (n12503,n12504);
not (n12504,n12285);
nand (n12505,n12506,n12507);
not (n12506,n12323);
not (n12507,n6527);
not (n12508,n12509);
nor (n12509,n12510,n12519);
nand (n12510,n12511,n12121);
not (n12511,n12512);
nand (n12512,n12513,n12516);
nand (n12513,n12514,n12515);
not (n12514,n6260);
not (n12515,n12212);
nand (n12516,n12517,n12518);
not (n12517,n6171);
not (n12518,n12175);
not (n12519,n12520);
nand (n12520,n12521,n12523,n12528);
and (n12521,n12522,n12504);
not (n12522,n12359);
nand (n12523,n12524,n12526);
not (n12524,n12525);
nor (n12525,n6616,n12360);
not (n12526,n12527);
not (n12527,n12395);
not (n12528,n12322);
nor (n12529,n12530,n12537);
and (n12530,n12531,n12532,n12121);
and (n12531,n12498,n12516);
not (n12532,n12533);
nand (n12533,n12534,n12513);
nand (n12534,n12535,n12536);
not (n12535,n12248);
not (n12536,n12211);
nand (n12537,n12538,n12441);
or (n12538,n12472,n12539);
not (n12539,n12540);
nand (n12540,n12541,n12543);
or (n12541,n12542,n12497);
not (n12542,n12174);
not (n12543,n12137);
and (n12544,n12482,n12545);
or (n12545,n12546,n12555,n12615);
and (n12546,n12547,n12549);
xor (n12547,n12548,n12087);
xor (n12548,n6825,n5082);
not (n12549,n12550);
xor (n12550,n12551,n12552);
xor (n12551,n6027,n12126);
or (n12552,n12446,n12553,n12554);
and (n12553,n12123,n12136);
and (n12554,n6034,n12136);
and (n12555,n12549,n12556);
or (n12556,n12557,n12563,n12614);
and (n12557,n12558,n12560);
xor (n12558,n12559,n12090);
xor (n12559,n6894,n5205);
not (n12560,n12561);
xor (n12561,n12562,n12136);
xor (n12562,n6034,n12123);
and (n12563,n12560,n12564);
or (n12564,n12565,n12571,n12613);
and (n12565,n12566,n12568);
xor (n12566,n12567,n12093);
xor (n12567,n6963,n5328);
not (n12568,n12569);
xor (n12569,n12570,n12173);
xor (n12570,n6082,n12138);
and (n12571,n12568,n12572);
or (n12572,n12573,n12579,n12612);
and (n12573,n12574,n12576);
xor (n12574,n12575,n12096);
xor (n12575,n7032,n5451);
not (n12576,n12577);
xor (n12577,n12578,n12210);
xor (n12578,n6171,n12175);
and (n12579,n12576,n12580);
or (n12580,n12581,n12587,n12611);
and (n12581,n12582,n12584);
xor (n12582,n12583,n12099);
xor (n12583,n7101,n5574);
not (n12584,n12585);
xor (n12585,n12586,n12247);
xor (n12586,n6260,n12212);
and (n12587,n12584,n12588);
or (n12588,n12589,n12595,n12610);
and (n12589,n12590,n12592);
xor (n12590,n12591,n12102);
xor (n12591,n7170,n5697);
not (n12592,n12593);
xor (n12593,n12594,n12284);
xor (n12594,n6349,n12249);
and (n12595,n12592,n12596);
or (n12596,n12597,n12603,n12609);
and (n12597,n12598,n12600);
xor (n12598,n12599,n12105);
xor (n12599,n7239,n5820);
not (n12600,n12601);
xor (n12601,n12602,n12321);
xor (n12602,n6438,n12286);
and (n12603,n12600,n12604);
and (n12604,n12605,n12606);
xor (n12605,n7307,n5942);
not (n12606,n12607);
xor (n12607,n12608,n12358);
xor (n12608,n6527,n12323);
and (n12609,n12598,n12604);
and (n12610,n12590,n12596);
and (n12611,n12582,n12588);
and (n12612,n12574,n12580);
and (n12613,n12566,n12572);
and (n12614,n12558,n12564);
and (n12615,n12547,n12556);
and (n12616,n12480,n12545);
and (n12617,n12461,n12478);
and (n12618,n12619,n12621);
xor (n12619,n12620,n12478);
xor (n12620,n12461,n12463);
and (n12621,n12622,n12624);
xor (n12622,n12623,n12545);
xor (n12623,n12480,n12482);
and (n12624,n12625,n12627);
xor (n12625,n12626,n12556);
xor (n12626,n12547,n12549);
and (n12627,n12628,n12630);
xor (n12628,n12629,n12564);
xor (n12629,n12558,n12560);
and (n12630,n12631,n12633);
xor (n12631,n12632,n12572);
xor (n12632,n12566,n12568);
and (n12633,n12634,n12636);
xor (n12634,n12635,n12580);
xor (n12635,n12574,n12576);
and (n12636,n12637,n12639);
xor (n12637,n12638,n12588);
xor (n12638,n12582,n12584);
and (n12639,n12640,n12642);
xor (n12640,n12641,n12596);
xor (n12641,n12590,n12592);
and (n12642,n12643,n12645);
xor (n12643,n12644,n12604);
xor (n12644,n12598,n12600);
and (n12645,n12646,n12647);
xor (n12646,n12605,n12606);
and (n12647,n12648,n12651);
not (n12648,n12649);
xor (n12649,n12650,n12395);
xor (n12650,n6616,n12360);
not (n12651,n12652);
xor (n12652,n6704,n12396);
or (n12653,n12654,n12658,n12731);
and (n12654,n12655,n12657);
xor (n12655,n12656,n11753);
xor (n12656,n7691,n11750);
xor (n12657,n12619,n12621);
and (n12658,n12657,n12659);
or (n12659,n12660,n12664,n12730);
and (n12660,n12661,n12663);
xor (n12661,n12662,n11758);
xor (n12662,n6019,n11755);
xor (n12663,n12622,n12624);
and (n12664,n12663,n12665);
or (n12665,n12666,n12670,n12729);
and (n12666,n12667,n12669);
xor (n12667,n12668,n11763);
xor (n12668,n6025,n11760);
xor (n12669,n12625,n12627);
and (n12670,n12669,n12671);
or (n12671,n12672,n12676,n12728);
and (n12672,n12673,n12675);
xor (n12673,n12674,n11768);
xor (n12674,n6032,n11765);
xor (n12675,n12628,n12630);
and (n12676,n12675,n12677);
or (n12677,n12678,n12682,n12727);
and (n12678,n12679,n12681);
xor (n12679,n12680,n11805);
xor (n12680,n6039,n11770);
xor (n12681,n12631,n12633);
and (n12682,n12681,n12683);
or (n12683,n12684,n12688,n12726);
and (n12684,n12685,n12687);
xor (n12685,n12686,n11842);
xor (n12686,n6128,n11807);
xor (n12687,n12634,n12636);
and (n12688,n12687,n12689);
or (n12689,n12690,n12694,n12725);
and (n12690,n12691,n12693);
xor (n12691,n12692,n11879);
xor (n12692,n6217,n11844);
xor (n12693,n12637,n12639);
and (n12694,n12693,n12695);
or (n12695,n12696,n12700,n12724);
and (n12696,n12697,n12699);
xor (n12697,n12698,n11916);
xor (n12698,n6306,n11881);
xor (n12699,n12640,n12642);
and (n12700,n12699,n12701);
or (n12701,n12702,n12706,n12723);
and (n12702,n12703,n12705);
xor (n12703,n12704,n11953);
xor (n12704,n6395,n11918);
xor (n12705,n12643,n12645);
and (n12706,n12705,n12707);
or (n12707,n12708,n12712,n12722);
and (n12708,n12709,n12711);
xor (n12709,n12710,n11990);
xor (n12710,n6484,n11955);
xor (n12711,n12646,n12647);
and (n12712,n12711,n12713);
or (n12713,n12714,n12718,n12721);
and (n12714,n12715,n12717);
xor (n12715,n12716,n12027);
xor (n12716,n6573,n11992);
xor (n12717,n12648,n12651);
and (n12718,n12717,n12719);
and (n12719,n12720,n12652);
xor (n12720,n6661,n12028);
and (n12721,n12715,n12719);
and (n12722,n12709,n12713);
and (n12723,n12703,n12707);
and (n12724,n12697,n12701);
and (n12725,n12691,n12695);
and (n12726,n12685,n12689);
and (n12727,n12679,n12683);
and (n12728,n12673,n12677);
and (n12729,n12667,n12671);
and (n12730,n12661,n12665);
and (n12731,n12655,n12659);
or (n12732,n12733,n12736,n12788);
and (n12733,n12734,n12669);
xor (n12734,n12735,n12659);
xor (n12735,n12655,n12657);
and (n12736,n12669,n12737);
or (n12737,n12738,n12741,n12787);
and (n12738,n12739,n12675);
xor (n12739,n12740,n12665);
xor (n12740,n12661,n12663);
and (n12741,n12675,n12742);
or (n12742,n12743,n12746,n12786);
and (n12743,n12744,n12681);
xor (n12744,n12745,n12671);
xor (n12745,n12667,n12669);
and (n12746,n12681,n12747);
or (n12747,n12748,n12751,n12785);
and (n12748,n12749,n12687);
xor (n12749,n12750,n12677);
xor (n12750,n12673,n12675);
and (n12751,n12687,n12752);
or (n12752,n12753,n12756,n12784);
and (n12753,n12754,n12693);
xor (n12754,n12755,n12683);
xor (n12755,n12679,n12681);
and (n12756,n12693,n12757);
or (n12757,n12758,n12761,n12783);
and (n12758,n12759,n12699);
xor (n12759,n12760,n12689);
xor (n12760,n12685,n12687);
and (n12761,n12699,n12762);
or (n12762,n12763,n12766,n12782);
and (n12763,n12764,n12705);
xor (n12764,n12765,n12695);
xor (n12765,n12691,n12693);
and (n12766,n12705,n12767);
or (n12767,n12768,n12771,n12781);
and (n12768,n12769,n12711);
xor (n12769,n12770,n12701);
xor (n12770,n12697,n12699);
and (n12771,n12711,n12772);
or (n12772,n12773,n12776,n12780);
and (n12773,n12774,n12717);
xor (n12774,n12775,n12707);
xor (n12775,n12703,n12705);
and (n12776,n12717,n12777);
and (n12777,n12778,n12652);
xor (n12778,n12779,n12713);
xor (n12779,n12709,n12711);
and (n12780,n12774,n12777);
and (n12781,n12769,n12772);
and (n12782,n12764,n12767);
and (n12783,n12759,n12762);
and (n12784,n12754,n12757);
and (n12785,n12749,n12752);
and (n12786,n12744,n12747);
and (n12787,n12739,n12742);
and (n12788,n12734,n12737);
and (n12789,n12790,n12792);
xor (n12790,n12791,n12737);
xor (n12791,n12734,n12669);
and (n12792,n12793,n12795);
xor (n12793,n12794,n12742);
xor (n12794,n12739,n12675);
and (n12795,n12796,n12798);
xor (n12796,n12797,n12747);
xor (n12797,n12744,n12681);
and (n12798,n12799,n12801);
xor (n12799,n12800,n12752);
xor (n12800,n12749,n12687);
and (n12801,n12802,n12804);
xor (n12802,n12803,n12757);
xor (n12803,n12754,n12693);
and (n12804,n12805,n12807);
xor (n12805,n12806,n12762);
xor (n12806,n12759,n12699);
and (n12807,n12808,n12810);
xor (n12808,n12809,n12767);
xor (n12809,n12764,n12705);
xor (n12810,n12811,n12772);
xor (n12811,n12769,n12711);
xor (n12812,n11740,n12813);
and (n12813,n12790,n12814);
and (n12814,n12793,n12796);
wire s0n12815,s1n12815,notn12815;
or (n12815,s0n12815,s1n12815);
not(notn12815,n4966);
and (s0n12815,notn12815,n12816);
and (s1n12815,n4966,n13025);
xor (n12816,n12817,n13012);
xor (n12817,n12818,n12984);
xor (n12818,n12819,n12963);
xor (n12819,n12820,n12957);
xor (n12820,n12821,n12839);
xor (n12821,n12822,n12825);
xor (n12822,n7668,n12823);
wire s0n12823,s1n12823,notn12823;
or (n12823,s0n12823,s1n12823);
not(notn12823,n4966);
and (s0n12823,notn12823,1'b0);
and (s1n12823,n4966,n12824);
or (n12825,n12826,n12827,n12838);
and (n12826,n7668,n12823);
and (n12827,n12823,n12828);
or (n12828,n12829,n12832,n12837);
and (n12829,n7677,n12830);
wire s0n12830,s1n12830,notn12830;
or (n12830,s0n12830,s1n12830);
not(notn12830,n4966);
and (s0n12830,notn12830,1'b0);
and (s1n12830,n4966,n12831);
and (n12832,n12830,n12833);
or (n12833,n12834,n12835,n12836);
and (n12834,n7684,n11746);
and (n12835,n11746,n11748);
and (n12836,n7684,n11748);
and (n12837,n7677,n12833);
and (n12838,n7668,n12828);
xor (n12839,n12840,n12944);
xor (n12840,n12841,n12889);
xor (n12841,n12842,n12864);
xor (n12842,n12843,n12844);
xor (n12843,n7709,n7645);
or (n12844,n12845,n12846,n12863);
and (n12845,n7709,n7645);
and (n12846,n7645,n12847);
or (n12847,n12848,n12849,n12862);
and (n12848,n7718,n7654);
and (n12849,n7654,n12850);
or (n12850,n12851,n12852,n12861);
and (n12851,n6761,n4974);
and (n12852,n4974,n12853);
or (n12853,n12854,n12855,n12860);
and (n12854,n6767,n4980);
and (n12855,n4980,n12856);
or (n12856,n12857,n12858,n12859);
and (n12857,n6774,n4987);
and (n12858,n4987,n12078);
and (n12859,n6774,n12078);
and (n12860,n6767,n12856);
and (n12861,n6761,n12853);
and (n12862,n7718,n12850);
and (n12863,n7709,n12847);
not (n12864,n12865);
nor (n12865,n12866,n12878);
and (n12866,n12136,n12867);
nor (n12867,n12868,n12120);
not (n12868,n12869);
nor (n12869,n12870,n12875);
nand (n12870,n12871,n12872);
or (n12871,n7686,n12454);
or (n12872,n7679,n12873);
wire s0n12873,s1n12873,notn12873;
or (n12873,s0n12873,s1n12873);
not(notn12873,n4966);
and (s0n12873,notn12873,1'b0);
and (s1n12873,n4966,n12874);
and (n12875,n7670,n12876);
wire s0n12876,s1n12876,notn12876;
or (n12876,s0n12876,s1n12876);
not(notn12876,n4966);
and (s0n12876,notn12876,1'b0);
and (s1n12876,n4966,n12877);
nand (n12878,n12879,n12880);
or (n12879,n12437,n12868);
nor (n12880,n12881,n12888);
and (n12881,n12882,n12887);
nand (n12882,n12883,n12886);
or (n12883,n12884,n12885);
nand (n12884,n7686,n12454);
not (n12885,n12872);
nand (n12886,n7679,n12873);
not (n12887,n12875);
nor (n12888,n7670,n12876);
or (n12889,n12890,n12892,n12943);
and (n12890,n12891,n12864);
xor (n12891,n12843,n12847);
and (n12892,n12864,n12893);
or (n12893,n12894,n12897,n12942);
and (n12894,n12895,n12864);
xor (n12895,n12896,n12850);
xor (n12896,n7718,n7654);
and (n12897,n12864,n12898);
or (n12898,n12899,n12915,n12941);
and (n12899,n12900,n12902);
xor (n12900,n12901,n12853);
xor (n12901,n6761,n4974);
not (n12902,n12903);
nand (n12903,n12904,n12914);
or (n12904,n12905,n12907);
not (n12905,n12906);
xor (n12906,n7670,n12876);
nand (n12907,n12908,n12911);
or (n12908,n12909,n12135);
not (n12909,n12910);
nor (n12910,n12120,n12870);
nor (n12911,n12912,n12882);
and (n12912,n12438,n12913);
not (n12913,n12870);
nand (n12914,n12907,n12905);
and (n12915,n12902,n12916);
or (n12916,n12917,n12935,n12940);
and (n12917,n12918,n12920);
xor (n12918,n12919,n12856);
xor (n12919,n6767,n4980);
not (n12920,n12921);
nor (n12921,n12922,n12932);
and (n12922,n12923,n12931);
nand (n12923,n12924,n12928);
or (n12924,n12925,n12135);
not (n12925,n12926);
nor (n12926,n12927,n12120);
not (n12927,n12871);
nor (n12928,n12929,n12930);
and (n12929,n12438,n12871);
not (n12930,n12884);
xor (n12931,n7679,n12873);
and (n12932,n12933,n12934);
not (n12933,n12923);
not (n12934,n12931);
and (n12935,n12920,n12936);
or (n12936,n12937,n12938,n12939);
and (n12937,n12076,n12115);
and (n12938,n12115,n12459);
and (n12939,n12076,n12459);
and (n12940,n12918,n12936);
and (n12941,n12900,n12916);
and (n12942,n12895,n12898);
and (n12943,n12891,n12893);
and (n12944,n12945,n12947);
xor (n12945,n12946,n12893);
xor (n12946,n12891,n12864);
and (n12947,n12948,n12950);
xor (n12948,n12949,n12898);
xor (n12949,n12895,n12864);
and (n12950,n12951,n12953);
xor (n12951,n12952,n12916);
xor (n12952,n12900,n12902);
and (n12953,n12954,n12956);
xor (n12954,n12955,n12936);
xor (n12955,n12918,n12920);
and (n12956,n12074,n12618);
or (n12957,n12958,n12960,n12983);
and (n12958,n12821,n12959);
xor (n12959,n12945,n12947);
and (n12960,n12959,n12961);
or (n12961,n12962,n12964,n12982);
and (n12962,n12821,n12963);
xor (n12963,n12948,n12950);
and (n12964,n12963,n12965);
or (n12965,n12966,n12969,n12981);
and (n12966,n12967,n12968);
xor (n12967,n12822,n12828);
xor (n12968,n12951,n12953);
and (n12969,n12968,n12970);
or (n12970,n12971,n12975,n12980);
and (n12971,n12972,n12974);
xor (n12972,n12973,n12833);
xor (n12973,n7677,n12830);
xor (n12974,n12954,n12956);
and (n12975,n12974,n12976);
or (n12976,n12977,n12978,n12979);
and (n12977,n11744,n12073);
and (n12978,n12073,n12653);
and (n12979,n11744,n12653);
and (n12980,n12972,n12976);
and (n12981,n12967,n12970);
and (n12982,n12821,n12965);
and (n12983,n12821,n12961);
or (n12984,n12985,n12988,n13011);
and (n12985,n12986,n12968);
xor (n12986,n12987,n12961);
xor (n12987,n12821,n12959);
and (n12988,n12968,n12989);
or (n12989,n12990,n12993,n13010);
and (n12990,n12991,n12974);
xor (n12991,n12992,n12965);
xor (n12992,n12821,n12963);
and (n12993,n12974,n12994);
or (n12994,n12995,n12998,n13009);
and (n12995,n12996,n12073);
xor (n12996,n12997,n12970);
xor (n12997,n12967,n12968);
and (n12998,n12073,n12999);
or (n12999,n13000,n13003,n13008);
and (n13000,n13001,n12657);
xor (n13001,n13002,n12976);
xor (n13002,n12972,n12974);
and (n13003,n12657,n13004);
or (n13004,n13005,n13006,n13007);
and (n13005,n11742,n12663);
and (n13006,n12663,n12732);
and (n13007,n11742,n12732);
and (n13008,n13001,n13004);
and (n13009,n12996,n12999);
and (n13010,n12991,n12994);
and (n13011,n12986,n12989);
and (n13012,n13013,n13015);
xor (n13013,n13014,n12989);
xor (n13014,n12986,n12968);
and (n13015,n13016,n13018);
xor (n13016,n13017,n12994);
xor (n13017,n12991,n12974);
and (n13018,n13019,n13021);
xor (n13019,n13020,n12999);
xor (n13020,n12996,n12073);
and (n13021,n13022,n13024);
xor (n13022,n13023,n13004);
xor (n13023,n13001,n12657);
and (n13024,n11740,n12789);
xor (n13025,n12817,n13026);
and (n13026,n13013,n13027);
and (n13027,n13016,n13028);
and (n13028,n13019,n13029);
and (n13029,n13022,n13030);
and (n13030,n11740,n12813);
wire s0n13031,s1n13031,notn13031;
or (n13031,s0n13031,s1n13031);
not(notn13031,n4966);
and (s0n13031,notn13031,n13032);
and (s1n13031,n4966,n13035);
wire s0n13032,s1n13032,notn13032;
or (n13032,s0n13032,s1n13032);
not(notn13032,n4966);
and (s0n13032,notn13032,n13033);
and (s1n13032,n4966,n13034);
xor (n13033,n13022,n13024);
xor (n13034,n13022,n13030);
wire s0n13035,s1n13035,notn13035;
or (n13035,s0n13035,s1n13035);
not(notn13035,n4966);
and (s0n13035,notn13035,n13036);
and (s1n13035,n4966,n13044);
xor (n13036,n13037,n13043);
xor (n13037,n13038,n13039);
xor (n13038,n12819,n12959);
or (n13039,n13040,n13041,n13042);
and (n13040,n12819,n12963);
and (n13041,n12963,n12984);
and (n13042,n12819,n12984);
and (n13043,n12817,n13012);
xor (n13044,n13037,n13045);
and (n13045,n12817,n13026);
wire s0n13046,s1n13046,notn13046;
or (n13046,s0n13046,s1n13046);
not(notn13046,n4966);
and (s0n13046,notn13046,n13047);
and (s1n13046,n4966,n13055);
xor (n13047,n13048,n13054);
xor (n13048,n13049,n13050);
xor (n13049,n12819,n12839);
or (n13050,n13051,n13052,n13053);
and (n13051,n12819,n12959);
and (n13052,n12959,n13039);
and (n13053,n12819,n13039);
and (n13054,n13037,n13043);
xor (n13055,n13048,n13056);
and (n13056,n13037,n13045);
and (n13057,n13058,n2907);
wire s0n13058,s1n13058,notn13058;
or (n13058,s0n13058,s1n13058);
not(notn13058,n2902);
and (s0n13058,notn13058,1'b0);
and (s1n13058,n2902,n11735);
and (n13059,n11735,n7875);
and (n13060,n9946,n7878);
and (n13061,n11732,n13062);
or (n13062,n13063,n13173,n13833);
and (n13063,n13064,n13157);
or (n13064,1'b0,n13065,n13068,n13071,n13076);
and (n13065,n13066,n2893);
wire s0n13066,s1n13066,notn13066;
or (n13066,s0n13066,s1n13066);
not(notn13066,n2891);
and (s0n13066,notn13066,1'b0);
and (s1n13066,n2891,n13067);
and (n13068,n13069,n2907);
wire s0n13069,s1n13069,notn13069;
or (n13069,s0n13069,s1n13069);
not(notn13069,n2902);
and (s0n13069,notn13069,1'b0);
and (s1n13069,n2902,n13070);
and (n13071,n13072,n4883);
wire s0n13072,s1n13072,notn13072;
or (n13072,s0n13072,s1n13072);
not(notn13072,n11666);
and (s0n13072,notn13072,n13073);
and (s1n13072,n11666,1'b0);
wire s0n13073,s1n13073,notn13073;
or (n13073,s0n13073,s1n13073);
not(notn13073,n11661);
and (s0n13073,notn13073,n13074);
and (s1n13073,n11661,1'b1);
wire s0n13074,s1n13074,notn13074;
or (n13074,s0n13074,s1n13074);
not(notn13074,n4861);
and (s0n13074,notn13074,1'b0);
and (s1n13074,n4861,n13075);
xor (n13075,n11639,n11641);
or (n13076,1'b0,n13077,n13097,n13117,n13137);
and (n13077,n13078,n2718);
or (n13078,1'b0,n13079,n13085,n13091);
and (n13079,n13080,n4895);
or (n13080,1'b0,n13081,n13082,n13083,n13084);
and (n13081,n5211,n556);
and (n13082,n5215,n567);
and (n13083,n5218,n571);
and (n13084,n5221,n573);
and (n13085,n13086,n2944);
or (n13086,1'b0,n13087,n13088,n13089,n13090);
and (n13087,n6901,n556);
and (n13088,n6900,n567);
and (n13089,n6904,n571);
and (n13090,n6907,n573);
and (n13091,n13092,n4903);
or (n13092,1'b0,n13093,n13094,n13095,n13096);
and (n13093,n6900,n556);
and (n13094,n6904,n567);
and (n13095,n6907,n571);
and (n13096,n6910,n573);
and (n13097,n13098,n2730);
or (n13098,1'b0,n13099,n13105,n13111);
and (n13099,n13100,n4895);
or (n13100,1'b0,n13101,n13102,n13103,n13104);
and (n13101,n5226,n556);
and (n13102,n5229,n567);
and (n13103,n5232,n571);
and (n13104,n5235,n573);
and (n13105,n13106,n2944);
or (n13106,1'b0,n13107,n13108,n13109,n13110);
and (n13107,n6910,n556);
and (n13108,n6915,n567);
and (n13109,n6918,n571);
and (n13110,n6921,n573);
and (n13111,n13112,n4903);
or (n13112,1'b0,n13113,n13114,n13115,n13116);
and (n13113,n6915,n556);
and (n13114,n6918,n567);
and (n13115,n6921,n571);
and (n13116,n6924,n573);
and (n13117,n13118,n2742);
or (n13118,1'b0,n13119,n13125,n13131);
and (n13119,n13120,n4895);
or (n13120,1'b0,n13121,n13122,n13123,n13124);
and (n13121,n5240,n556);
and (n13122,n5244,n567);
and (n13123,n5247,n571);
and (n13124,n5250,n573);
and (n13125,n13126,n2944);
or (n13126,1'b0,n13127,n13128,n13129,n13130);
and (n13127,n5153,n556);
and (n13128,n5152,n567);
and (n13129,n5156,n571);
and (n13130,n5159,n573);
and (n13131,n13132,n4903);
or (n13132,1'b0,n13133,n13134,n13135,n13136);
and (n13133,n5152,n556);
and (n13134,n5156,n567);
and (n13135,n5159,n571);
and (n13136,n5162,n573);
and (n13137,n13138,n2752);
or (n13138,1'b0,n13139,n13145,n13151);
and (n13139,n13140,n4895);
or (n13140,1'b0,n13141,n13142,n13143,n13144);
and (n13141,n5255,n556);
and (n13142,n5258,n567);
and (n13143,n5261,n571);
and (n13144,n5264,n573);
and (n13145,n13146,n2944);
or (n13146,1'b0,n13147,n13148,n13149,n13150);
and (n13147,n5162,n556);
and (n13148,n5167,n567);
and (n13149,n5170,n571);
and (n13150,n5173,n573);
and (n13151,n13152,n4903);
or (n13152,1'b0,n13153,n13154,n13155,n13156);
and (n13153,n5167,n556);
and (n13154,n5170,n567);
and (n13155,n5173,n571);
and (n13156,n5176,n573);
or (n13157,1'b0,n13158,n13169,n13171,n13172);
and (n13158,n13159,n2893);
wire s0n13159,s1n13159,notn13159;
or (n13159,s0n13159,s1n13159);
not(notn13159,n2891);
and (s0n13159,notn13159,1'b0);
and (s1n13159,n2891,n13160);
wire s0n13160,s1n13160,notn13160;
or (n13160,s0n13160,s1n13160);
not(notn13160,n13046);
and (s0n13160,notn13160,n13161);
and (s1n13160,n13046,1'b0);
wire s0n13161,s1n13161,notn13161;
or (n13161,s0n13161,s1n13161);
not(notn13161,n13031);
and (s0n13161,notn13161,n13162);
and (s1n13161,n13031,1'b1);
wire s0n13162,s1n13162,notn13162;
or (n13162,s0n13162,s1n13162);
not(notn13162,n4966);
and (s0n13162,notn13162,n13163);
and (s1n13162,n4966,n13166);
wire s0n13163,s1n13163,notn13163;
or (n13163,s0n13163,s1n13163);
not(notn13163,n4966);
and (s0n13163,notn13163,n13164);
and (s1n13163,n4966,n13165);
xor (n13164,n12790,n12792);
xor (n13165,n12790,n12814);
wire s0n13166,s1n13166,notn13166;
or (n13166,s0n13166,s1n13166);
not(notn13166,n4966);
and (s0n13166,notn13166,n13167);
and (s1n13166,n4966,n13168);
xor (n13167,n13013,n13015);
xor (n13168,n13013,n13027);
and (n13169,n13170,n2907);
wire s0n13170,s1n13170,notn13170;
or (n13170,s0n13170,s1n13170);
not(notn13170,n2902);
and (s0n13170,notn13170,1'b0);
and (s1n13170,n2902,n13160);
and (n13171,n13160,n7875);
and (n13172,n13072,n7878);
and (n13173,n13157,n13174);
or (n13174,n13175,n13285,n13832);
and (n13175,n13176,n13269);
or (n13176,1'b0,n13177,n13180,n13183,n13188);
and (n13177,n13178,n2893);
wire s0n13178,s1n13178,notn13178;
or (n13178,s0n13178,s1n13178);
not(notn13178,n2891);
and (s0n13178,notn13178,1'b0);
and (s1n13178,n2891,n13179);
and (n13180,n13181,n2907);
wire s0n13181,s1n13181,notn13181;
or (n13181,s0n13181,s1n13181);
not(notn13181,n2902);
and (s0n13181,notn13181,1'b0);
and (s1n13181,n2902,n13182);
and (n13183,n13184,n4883);
wire s0n13184,s1n13184,notn13184;
or (n13184,s0n13184,s1n13184);
not(notn13184,n11666);
and (s0n13184,notn13184,n13185);
and (s1n13184,n11666,1'b0);
wire s0n13185,s1n13185,notn13185;
or (n13185,s0n13185,s1n13185);
not(notn13185,n11661);
and (s0n13185,notn13185,n13186);
and (s1n13185,n11661,1'b1);
wire s0n13186,s1n13186,notn13186;
or (n13186,s0n13186,s1n13186);
not(notn13186,n4861);
and (s0n13186,notn13186,1'b0);
and (s1n13186,n4861,n13187);
xor (n13187,n11642,n11644);
or (n13188,1'b0,n13189,n13209,n13229,n13249);
and (n13189,n13190,n2718);
or (n13190,1'b0,n13191,n13197,n13203);
and (n13191,n13192,n4895);
or (n13192,1'b0,n13193,n13194,n13195,n13196);
and (n13193,n5334,n556);
and (n13194,n5338,n567);
and (n13195,n5341,n571);
and (n13196,n5344,n573);
and (n13197,n13198,n2944);
or (n13198,1'b0,n13199,n13200,n13201,n13202);
and (n13199,n6970,n556);
and (n13200,n6969,n567);
and (n13201,n6973,n571);
and (n13202,n6976,n573);
and (n13203,n13204,n4903);
or (n13204,1'b0,n13205,n13206,n13207,n13208);
and (n13205,n6969,n556);
and (n13206,n6973,n567);
and (n13207,n6976,n571);
and (n13208,n6979,n573);
and (n13209,n13210,n2730);
or (n13210,1'b0,n13211,n13217,n13223);
and (n13211,n13212,n4895);
or (n13212,1'b0,n13213,n13214,n13215,n13216);
and (n13213,n5349,n556);
and (n13214,n5352,n567);
and (n13215,n5355,n571);
and (n13216,n5358,n573);
and (n13217,n13218,n2944);
or (n13218,1'b0,n13219,n13220,n13221,n13222);
and (n13219,n6979,n556);
and (n13220,n6984,n567);
and (n13221,n6987,n571);
and (n13222,n6990,n573);
and (n13223,n13224,n4903);
or (n13224,1'b0,n13225,n13226,n13227,n13228);
and (n13225,n6984,n556);
and (n13226,n6987,n567);
and (n13227,n6990,n571);
and (n13228,n6993,n573);
and (n13229,n13230,n2742);
or (n13230,1'b0,n13231,n13237,n13243);
and (n13231,n13232,n4895);
or (n13232,1'b0,n13233,n13234,n13235,n13236);
and (n13233,n5363,n556);
and (n13234,n5367,n567);
and (n13235,n5370,n571);
and (n13236,n5373,n573);
and (n13237,n13238,n2944);
or (n13238,1'b0,n13239,n13240,n13241,n13242);
and (n13239,n5276,n556);
and (n13240,n5275,n567);
and (n13241,n5279,n571);
and (n13242,n5282,n573);
and (n13243,n13244,n4903);
or (n13244,1'b0,n13245,n13246,n13247,n13248);
and (n13245,n5275,n556);
and (n13246,n5279,n567);
and (n13247,n5282,n571);
and (n13248,n5285,n573);
and (n13249,n13250,n2752);
or (n13250,1'b0,n13251,n13257,n13263);
and (n13251,n13252,n4895);
or (n13252,1'b0,n13253,n13254,n13255,n13256);
and (n13253,n5378,n556);
and (n13254,n5381,n567);
and (n13255,n5384,n571);
and (n13256,n5387,n573);
and (n13257,n13258,n2944);
or (n13258,1'b0,n13259,n13260,n13261,n13262);
and (n13259,n5285,n556);
and (n13260,n5290,n567);
and (n13261,n5293,n571);
and (n13262,n5296,n573);
and (n13263,n13264,n4903);
or (n13264,1'b0,n13265,n13266,n13267,n13268);
and (n13265,n5290,n556);
and (n13266,n5293,n567);
and (n13267,n5296,n571);
and (n13268,n5299,n573);
or (n13269,1'b0,n13270,n13281,n13283,n13284);
and (n13270,n13271,n2893);
wire s0n13271,s1n13271,notn13271;
or (n13271,s0n13271,s1n13271);
not(notn13271,n2891);
and (s0n13271,notn13271,1'b0);
and (s1n13271,n2891,n13272);
wire s0n13272,s1n13272,notn13272;
or (n13272,s0n13272,s1n13272);
not(notn13272,n13046);
and (s0n13272,notn13272,n13273);
and (s1n13272,n13046,1'b0);
wire s0n13273,s1n13273,notn13273;
or (n13273,s0n13273,s1n13273);
not(notn13273,n13031);
and (s0n13273,notn13273,n13274);
and (s1n13273,n13031,1'b1);
wire s0n13274,s1n13274,notn13274;
or (n13274,s0n13274,s1n13274);
not(notn13274,n4966);
and (s0n13274,notn13274,n13275);
and (s1n13274,n4966,n13278);
wire s0n13275,s1n13275,notn13275;
or (n13275,s0n13275,s1n13275);
not(notn13275,n4966);
and (s0n13275,notn13275,n13276);
and (s1n13275,n4966,n13277);
xor (n13276,n12793,n12795);
xor (n13277,n12793,n12796);
wire s0n13278,s1n13278,notn13278;
or (n13278,s0n13278,s1n13278);
not(notn13278,n4966);
and (s0n13278,notn13278,n13279);
and (s1n13278,n4966,n13280);
xor (n13279,n13016,n13018);
xor (n13280,n13016,n13028);
and (n13281,n13282,n2907);
wire s0n13282,s1n13282,notn13282;
or (n13282,s0n13282,s1n13282);
not(notn13282,n2902);
and (s0n13282,notn13282,1'b0);
and (s1n13282,n2902,n13272);
and (n13283,n13272,n7875);
and (n13284,n13184,n7878);
and (n13285,n13269,n13286);
or (n13286,n13287,n13397,n13831);
and (n13287,n13288,n13381);
or (n13288,1'b0,n13289,n13292,n13295,n13300);
and (n13289,n13290,n2893);
wire s0n13290,s1n13290,notn13290;
or (n13290,s0n13290,s1n13290);
not(notn13290,n2891);
and (s0n13290,notn13290,1'b0);
and (s1n13290,n2891,n13291);
and (n13292,n13293,n2907);
wire s0n13293,s1n13293,notn13293;
or (n13293,s0n13293,s1n13293);
not(notn13293,n2902);
and (s0n13293,notn13293,1'b0);
and (s1n13293,n2902,n13294);
and (n13295,n13296,n4883);
wire s0n13296,s1n13296,notn13296;
or (n13296,s0n13296,s1n13296);
not(notn13296,n11666);
and (s0n13296,notn13296,n13297);
and (s1n13296,n11666,1'b0);
wire s0n13297,s1n13297,notn13297;
or (n13297,s0n13297,s1n13297);
not(notn13297,n11661);
and (s0n13297,notn13297,n13298);
and (s1n13297,n11661,1'b1);
wire s0n13298,s1n13298,notn13298;
or (n13298,s0n13298,s1n13298);
not(notn13298,n4861);
and (s0n13298,notn13298,1'b0);
and (s1n13298,n4861,n13299);
xor (n13299,n11645,n11647);
or (n13300,1'b0,n13301,n13321,n13341,n13361);
and (n13301,n13302,n2718);
or (n13302,1'b0,n13303,n13309,n13315);
and (n13303,n13304,n4895);
or (n13304,1'b0,n13305,n13306,n13307,n13308);
and (n13305,n5457,n556);
and (n13306,n5461,n567);
and (n13307,n5464,n571);
and (n13308,n5467,n573);
and (n13309,n13310,n2944);
or (n13310,1'b0,n13311,n13312,n13313,n13314);
and (n13311,n7039,n556);
and (n13312,n7038,n567);
and (n13313,n7042,n571);
and (n13314,n7045,n573);
and (n13315,n13316,n4903);
or (n13316,1'b0,n13317,n13318,n13319,n13320);
and (n13317,n7038,n556);
and (n13318,n7042,n567);
and (n13319,n7045,n571);
and (n13320,n7048,n573);
and (n13321,n13322,n2730);
or (n13322,1'b0,n13323,n13329,n13335);
and (n13323,n13324,n4895);
or (n13324,1'b0,n13325,n13326,n13327,n13328);
and (n13325,n5472,n556);
and (n13326,n5475,n567);
and (n13327,n5478,n571);
and (n13328,n5481,n573);
and (n13329,n13330,n2944);
or (n13330,1'b0,n13331,n13332,n13333,n13334);
and (n13331,n7048,n556);
and (n13332,n7053,n567);
and (n13333,n7056,n571);
and (n13334,n7059,n573);
and (n13335,n13336,n4903);
or (n13336,1'b0,n13337,n13338,n13339,n13340);
and (n13337,n7053,n556);
and (n13338,n7056,n567);
and (n13339,n7059,n571);
and (n13340,n7062,n573);
and (n13341,n13342,n2742);
or (n13342,1'b0,n13343,n13349,n13355);
and (n13343,n13344,n4895);
or (n13344,1'b0,n13345,n13346,n13347,n13348);
and (n13345,n5486,n556);
and (n13346,n5490,n567);
and (n13347,n5493,n571);
and (n13348,n5496,n573);
and (n13349,n13350,n2944);
or (n13350,1'b0,n13351,n13352,n13353,n13354);
and (n13351,n5399,n556);
and (n13352,n5398,n567);
and (n13353,n5402,n571);
and (n13354,n5405,n573);
and (n13355,n13356,n4903);
or (n13356,1'b0,n13357,n13358,n13359,n13360);
and (n13357,n5398,n556);
and (n13358,n5402,n567);
and (n13359,n5405,n571);
and (n13360,n5408,n573);
and (n13361,n13362,n2752);
or (n13362,1'b0,n13363,n13369,n13375);
and (n13363,n13364,n4895);
or (n13364,1'b0,n13365,n13366,n13367,n13368);
and (n13365,n5501,n556);
and (n13366,n5504,n567);
and (n13367,n5507,n571);
and (n13368,n5510,n573);
and (n13369,n13370,n2944);
or (n13370,1'b0,n13371,n13372,n13373,n13374);
and (n13371,n5408,n556);
and (n13372,n5413,n567);
and (n13373,n5416,n571);
and (n13374,n5419,n573);
and (n13375,n13376,n4903);
or (n13376,1'b0,n13377,n13378,n13379,n13380);
and (n13377,n5413,n556);
and (n13378,n5416,n567);
and (n13379,n5419,n571);
and (n13380,n5422,n573);
or (n13381,1'b0,n13382,n13393,n13395,n13396);
and (n13382,n13383,n2893);
wire s0n13383,s1n13383,notn13383;
or (n13383,s0n13383,s1n13383);
not(notn13383,n2891);
and (s0n13383,notn13383,1'b0);
and (s1n13383,n2891,n13384);
wire s0n13384,s1n13384,notn13384;
or (n13384,s0n13384,s1n13384);
not(notn13384,n13046);
and (s0n13384,notn13384,n13385);
and (s1n13384,n13046,1'b0);
wire s0n13385,s1n13385,notn13385;
or (n13385,s0n13385,s1n13385);
not(notn13385,n13031);
and (s0n13385,notn13385,n13386);
and (s1n13385,n13031,1'b1);
wire s0n13386,s1n13386,notn13386;
or (n13386,s0n13386,s1n13386);
not(notn13386,n4966);
and (s0n13386,notn13386,n13387);
and (s1n13386,n4966,n13390);
wire s0n13387,s1n13387,notn13387;
or (n13387,s0n13387,s1n13387);
not(notn13387,n4966);
and (s0n13387,notn13387,n13388);
and (s1n13387,n4966,n13389);
xor (n13388,n12796,n12798);
not (n13389,n12796);
wire s0n13390,s1n13390,notn13390;
or (n13390,s0n13390,s1n13390);
not(notn13390,n4966);
and (s0n13390,notn13390,n13391);
and (s1n13390,n4966,n13392);
xor (n13391,n13019,n13021);
xor (n13392,n13019,n13029);
and (n13393,n13394,n2907);
wire s0n13394,s1n13394,notn13394;
or (n13394,s0n13394,s1n13394);
not(notn13394,n2902);
and (s0n13394,notn13394,1'b0);
and (s1n13394,n2902,n13384);
and (n13395,n13384,n7875);
and (n13396,n13296,n7878);
and (n13397,n13381,n13398);
or (n13398,n13399,n13505,n13830);
and (n13399,n13400,n13493);
or (n13400,1'b0,n13401,n13404,n13407,n13412);
and (n13401,n13402,n2893);
wire s0n13402,s1n13402,notn13402;
or (n13402,s0n13402,s1n13402);
not(notn13402,n2891);
and (s0n13402,notn13402,1'b0);
and (s1n13402,n2891,n13403);
and (n13404,n13405,n2907);
wire s0n13405,s1n13405,notn13405;
or (n13405,s0n13405,s1n13405);
not(notn13405,n2902);
and (s0n13405,notn13405,1'b0);
and (s1n13405,n2902,n13406);
and (n13407,n13408,n4883);
wire s0n13408,s1n13408,notn13408;
or (n13408,s0n13408,s1n13408);
not(notn13408,n11666);
and (s0n13408,notn13408,n13409);
and (s1n13408,n11666,1'b0);
wire s0n13409,s1n13409,notn13409;
or (n13409,s0n13409,s1n13409);
not(notn13409,n11661);
and (s0n13409,notn13409,n13410);
and (s1n13409,n11661,1'b1);
wire s0n13410,s1n13410,notn13410;
or (n13410,s0n13410,s1n13410);
not(notn13410,n4861);
and (s0n13410,notn13410,1'b0);
and (s1n13410,n4861,n13411);
xor (n13411,n11648,n11650);
or (n13412,1'b0,n13413,n13433,n13453,n13473);
and (n13413,n13414,n2718);
or (n13414,1'b0,n13415,n13421,n13427);
and (n13415,n13416,n4895);
or (n13416,1'b0,n13417,n13418,n13419,n13420);
and (n13417,n5580,n556);
and (n13418,n5584,n567);
and (n13419,n5587,n571);
and (n13420,n5590,n573);
and (n13421,n13422,n2944);
or (n13422,1'b0,n13423,n13424,n13425,n13426);
and (n13423,n7108,n556);
and (n13424,n7107,n567);
and (n13425,n7111,n571);
and (n13426,n7114,n573);
and (n13427,n13428,n4903);
or (n13428,1'b0,n13429,n13430,n13431,n13432);
and (n13429,n7107,n556);
and (n13430,n7111,n567);
and (n13431,n7114,n571);
and (n13432,n7117,n573);
and (n13433,n13434,n2730);
or (n13434,1'b0,n13435,n13441,n13447);
and (n13435,n13436,n4895);
or (n13436,1'b0,n13437,n13438,n13439,n13440);
and (n13437,n5595,n556);
and (n13438,n5598,n567);
and (n13439,n5601,n571);
and (n13440,n5604,n573);
and (n13441,n13442,n2944);
or (n13442,1'b0,n13443,n13444,n13445,n13446);
and (n13443,n7117,n556);
and (n13444,n7122,n567);
and (n13445,n7125,n571);
and (n13446,n7128,n573);
and (n13447,n13448,n4903);
or (n13448,1'b0,n13449,n13450,n13451,n13452);
and (n13449,n7122,n556);
and (n13450,n7125,n567);
and (n13451,n7128,n571);
and (n13452,n7131,n573);
and (n13453,n13454,n2742);
or (n13454,1'b0,n13455,n13461,n13467);
and (n13455,n13456,n4895);
or (n13456,1'b0,n13457,n13458,n13459,n13460);
and (n13457,n5609,n556);
and (n13458,n5613,n567);
and (n13459,n5616,n571);
and (n13460,n5619,n573);
and (n13461,n13462,n2944);
or (n13462,1'b0,n13463,n13464,n13465,n13466);
and (n13463,n5522,n556);
and (n13464,n5521,n567);
and (n13465,n5525,n571);
and (n13466,n5528,n573);
and (n13467,n13468,n4903);
or (n13468,1'b0,n13469,n13470,n13471,n13472);
and (n13469,n5521,n556);
and (n13470,n5525,n567);
and (n13471,n5528,n571);
and (n13472,n5531,n573);
and (n13473,n13474,n2752);
or (n13474,1'b0,n13475,n13481,n13487);
and (n13475,n13476,n4895);
or (n13476,1'b0,n13477,n13478,n13479,n13480);
and (n13477,n5624,n556);
and (n13478,n5627,n567);
and (n13479,n5630,n571);
and (n13480,n5633,n573);
and (n13481,n13482,n2944);
or (n13482,1'b0,n13483,n13484,n13485,n13486);
and (n13483,n5531,n556);
and (n13484,n5536,n567);
and (n13485,n5539,n571);
and (n13486,n5542,n573);
and (n13487,n13488,n4903);
or (n13488,1'b0,n13489,n13490,n13491,n13492);
and (n13489,n5536,n556);
and (n13490,n5539,n567);
and (n13491,n5542,n571);
and (n13492,n5545,n573);
or (n13493,1'b0,n13494,n13501,n13503,n13504);
and (n13494,n13495,n2893);
wire s0n13495,s1n13495,notn13495;
or (n13495,s0n13495,s1n13495);
not(notn13495,n2891);
and (s0n13495,notn13495,1'b0);
and (s1n13495,n2891,n13496);
wire s0n13496,s1n13496,notn13496;
or (n13496,s0n13496,s1n13496);
not(notn13496,n13046);
and (s0n13496,notn13496,n13497);
and (s1n13496,n13046,1'b0);
wire s0n13497,s1n13497,notn13497;
or (n13497,s0n13497,s1n13497);
not(notn13497,n13031);
and (s0n13497,notn13497,n13498);
and (s1n13497,n13031,1'b1);
wire s0n13498,s1n13498,notn13498;
or (n13498,s0n13498,s1n13498);
not(notn13498,n4966);
and (s0n13498,notn13498,n13499);
and (s1n13498,n4966,n13032);
wire s0n13499,s1n13499,notn13499;
or (n13499,s0n13499,s1n13499);
not(notn13499,n4966);
and (s0n13499,notn13499,n13500);
and (s1n13499,n4966,n12799);
xor (n13500,n12799,n12801);
and (n13501,n13502,n2907);
wire s0n13502,s1n13502,notn13502;
or (n13502,s0n13502,s1n13502);
not(notn13502,n2902);
and (s0n13502,notn13502,1'b0);
and (s1n13502,n2902,n13496);
and (n13503,n13496,n7875);
and (n13504,n13408,n7878);
and (n13505,n13493,n13506);
or (n13506,n13507,n13613,n13829);
and (n13507,n13508,n13601);
or (n13508,1'b0,n13509,n13512,n13515,n13520);
and (n13509,n13510,n2893);
wire s0n13510,s1n13510,notn13510;
or (n13510,s0n13510,s1n13510);
not(notn13510,n2891);
and (s0n13510,notn13510,1'b0);
and (s1n13510,n2891,n13511);
and (n13512,n13513,n2907);
wire s0n13513,s1n13513,notn13513;
or (n13513,s0n13513,s1n13513);
not(notn13513,n2902);
and (s0n13513,notn13513,1'b0);
and (s1n13513,n2902,n13514);
and (n13515,n13516,n4883);
wire s0n13516,s1n13516,notn13516;
or (n13516,s0n13516,s1n13516);
not(notn13516,n11666);
and (s0n13516,notn13516,n13517);
and (s1n13516,n11666,1'b0);
wire s0n13517,s1n13517,notn13517;
or (n13517,s0n13517,s1n13517);
not(notn13517,n11661);
and (s0n13517,notn13517,n13518);
and (s1n13517,n11661,1'b1);
wire s0n13518,s1n13518,notn13518;
or (n13518,s0n13518,s1n13518);
not(notn13518,n4861);
and (s0n13518,notn13518,1'b0);
and (s1n13518,n4861,n13519);
xor (n13519,n11651,n11653);
or (n13520,1'b0,n13521,n13541,n13561,n13581);
and (n13521,n13522,n2718);
or (n13522,1'b0,n13523,n13529,n13535);
and (n13523,n13524,n4895);
or (n13524,1'b0,n13525,n13526,n13527,n13528);
and (n13525,n5703,n556);
and (n13526,n5707,n567);
and (n13527,n5710,n571);
and (n13528,n5713,n573);
and (n13529,n13530,n2944);
or (n13530,1'b0,n13531,n13532,n13533,n13534);
and (n13531,n7177,n556);
and (n13532,n7176,n567);
and (n13533,n7180,n571);
and (n13534,n7183,n573);
and (n13535,n13536,n4903);
or (n13536,1'b0,n13537,n13538,n13539,n13540);
and (n13537,n7176,n556);
and (n13538,n7180,n567);
and (n13539,n7183,n571);
and (n13540,n7186,n573);
and (n13541,n13542,n2730);
or (n13542,1'b0,n13543,n13549,n13555);
and (n13543,n13544,n4895);
or (n13544,1'b0,n13545,n13546,n13547,n13548);
and (n13545,n5718,n556);
and (n13546,n5721,n567);
and (n13547,n5724,n571);
and (n13548,n5727,n573);
and (n13549,n13550,n2944);
or (n13550,1'b0,n13551,n13552,n13553,n13554);
and (n13551,n7186,n556);
and (n13552,n7191,n567);
and (n13553,n7194,n571);
and (n13554,n7197,n573);
and (n13555,n13556,n4903);
or (n13556,1'b0,n13557,n13558,n13559,n13560);
and (n13557,n7191,n556);
and (n13558,n7194,n567);
and (n13559,n7197,n571);
and (n13560,n7200,n573);
and (n13561,n13562,n2742);
or (n13562,1'b0,n13563,n13569,n13575);
and (n13563,n13564,n4895);
or (n13564,1'b0,n13565,n13566,n13567,n13568);
and (n13565,n5732,n556);
and (n13566,n5736,n567);
and (n13567,n5739,n571);
and (n13568,n5742,n573);
and (n13569,n13570,n2944);
or (n13570,1'b0,n13571,n13572,n13573,n13574);
and (n13571,n5645,n556);
and (n13572,n5644,n567);
and (n13573,n5648,n571);
and (n13574,n5651,n573);
and (n13575,n13576,n4903);
or (n13576,1'b0,n13577,n13578,n13579,n13580);
and (n13577,n5644,n556);
and (n13578,n5648,n567);
and (n13579,n5651,n571);
and (n13580,n5654,n573);
and (n13581,n13582,n2752);
or (n13582,1'b0,n13583,n13589,n13595);
and (n13583,n13584,n4895);
or (n13584,1'b0,n13585,n13586,n13587,n13588);
and (n13585,n5747,n556);
and (n13586,n5750,n567);
and (n13587,n5753,n571);
and (n13588,n5756,n573);
and (n13589,n13590,n2944);
or (n13590,1'b0,n13591,n13592,n13593,n13594);
and (n13591,n5654,n556);
and (n13592,n5659,n567);
and (n13593,n5662,n571);
and (n13594,n5665,n573);
and (n13595,n13596,n4903);
or (n13596,1'b0,n13597,n13598,n13599,n13600);
and (n13597,n5659,n556);
and (n13598,n5662,n567);
and (n13599,n5665,n571);
and (n13600,n5668,n573);
or (n13601,1'b0,n13602,n13609,n13611,n13612);
and (n13602,n13603,n2893);
wire s0n13603,s1n13603,notn13603;
or (n13603,s0n13603,s1n13603);
not(notn13603,n2891);
and (s0n13603,notn13603,1'b0);
and (s1n13603,n2891,n13604);
wire s0n13604,s1n13604,notn13604;
or (n13604,s0n13604,s1n13604);
not(notn13604,n13046);
and (s0n13604,notn13604,n13605);
and (s1n13604,n13046,1'b0);
wire s0n13605,s1n13605,notn13605;
or (n13605,s0n13605,s1n13605);
not(notn13605,n13031);
and (s0n13605,notn13605,n13606);
and (s1n13605,n13031,1'b1);
wire s0n13606,s1n13606,notn13606;
or (n13606,s0n13606,s1n13606);
not(notn13606,n4966);
and (s0n13606,notn13606,n13607);
and (s1n13606,n4966,n11738);
wire s0n13607,s1n13607,notn13607;
or (n13607,s0n13607,s1n13607);
not(notn13607,n4966);
and (s0n13607,notn13607,n13608);
and (s1n13607,n4966,n12802);
xor (n13608,n12802,n12804);
and (n13609,n13610,n2907);
wire s0n13610,s1n13610,notn13610;
or (n13610,s0n13610,s1n13610);
not(notn13610,n2902);
and (s0n13610,notn13610,1'b0);
and (s1n13610,n2902,n13604);
and (n13611,n13604,n7875);
and (n13612,n13516,n7878);
and (n13613,n13601,n13614);
or (n13614,n13615,n13721,n13828);
and (n13615,n13616,n13709);
or (n13616,1'b0,n13617,n13620,n13623,n13628);
and (n13617,n13618,n2893);
wire s0n13618,s1n13618,notn13618;
or (n13618,s0n13618,s1n13618);
not(notn13618,n2891);
and (s0n13618,notn13618,1'b0);
and (s1n13618,n2891,n13619);
and (n13620,n13621,n2907);
wire s0n13621,s1n13621,notn13621;
or (n13621,s0n13621,s1n13621);
not(notn13621,n2902);
and (s0n13621,notn13621,1'b0);
and (s1n13621,n2902,n13622);
and (n13623,n13624,n4883);
wire s0n13624,s1n13624,notn13624;
or (n13624,s0n13624,s1n13624);
not(notn13624,n11666);
and (s0n13624,notn13624,n13625);
and (s1n13624,n11666,1'b0);
wire s0n13625,s1n13625,notn13625;
or (n13625,s0n13625,s1n13625);
not(notn13625,n11661);
and (s0n13625,notn13625,n13626);
and (s1n13625,n11661,1'b1);
wire s0n13626,s1n13626,notn13626;
or (n13626,s0n13626,s1n13626);
not(notn13626,n4861);
and (s0n13626,notn13626,1'b0);
and (s1n13626,n4861,n13627);
xor (n13627,n11654,n11656);
or (n13628,1'b0,n13629,n13649,n13669,n13689);
and (n13629,n13630,n2718);
or (n13630,1'b0,n13631,n13637,n13643);
and (n13631,n13632,n4895);
or (n13632,1'b0,n13633,n13634,n13635,n13636);
and (n13633,n5826,n556);
and (n13634,n5830,n567);
and (n13635,n5833,n571);
and (n13636,n5836,n573);
and (n13637,n13638,n2944);
or (n13638,1'b0,n13639,n13640,n13641,n13642);
and (n13639,n7246,n556);
and (n13640,n7245,n567);
and (n13641,n7249,n571);
and (n13642,n7252,n573);
and (n13643,n13644,n4903);
or (n13644,1'b0,n13645,n13646,n13647,n13648);
and (n13645,n7245,n556);
and (n13646,n7249,n567);
and (n13647,n7252,n571);
and (n13648,n7255,n573);
and (n13649,n13650,n2730);
or (n13650,1'b0,n13651,n13657,n13663);
and (n13651,n13652,n4895);
or (n13652,1'b0,n13653,n13654,n13655,n13656);
and (n13653,n5841,n556);
and (n13654,n5844,n567);
and (n13655,n5847,n571);
and (n13656,n5850,n573);
and (n13657,n13658,n2944);
or (n13658,1'b0,n13659,n13660,n13661,n13662);
and (n13659,n7255,n556);
and (n13660,n7260,n567);
and (n13661,n7263,n571);
and (n13662,n7266,n573);
and (n13663,n13664,n4903);
or (n13664,1'b0,n13665,n13666,n13667,n13668);
and (n13665,n7260,n556);
and (n13666,n7263,n567);
and (n13667,n7266,n571);
and (n13668,n7269,n573);
and (n13669,n13670,n2742);
or (n13670,1'b0,n13671,n13677,n13683);
and (n13671,n13672,n4895);
or (n13672,1'b0,n13673,n13674,n13675,n13676);
and (n13673,n5855,n556);
and (n13674,n5859,n567);
and (n13675,n5862,n571);
and (n13676,n5865,n573);
and (n13677,n13678,n2944);
or (n13678,1'b0,n13679,n13680,n13681,n13682);
and (n13679,n5768,n556);
and (n13680,n5767,n567);
and (n13681,n5771,n571);
and (n13682,n5774,n573);
and (n13683,n13684,n4903);
or (n13684,1'b0,n13685,n13686,n13687,n13688);
and (n13685,n5767,n556);
and (n13686,n5771,n567);
and (n13687,n5774,n571);
and (n13688,n5777,n573);
and (n13689,n13690,n2752);
or (n13690,1'b0,n13691,n13697,n13703);
and (n13691,n13692,n4895);
or (n13692,1'b0,n13693,n13694,n13695,n13696);
and (n13693,n5870,n556);
and (n13694,n5873,n567);
and (n13695,n5876,n571);
and (n13696,n5879,n573);
and (n13697,n13698,n2944);
or (n13698,1'b0,n13699,n13700,n13701,n13702);
and (n13699,n5777,n556);
and (n13700,n5782,n567);
and (n13701,n5785,n571);
and (n13702,n5788,n573);
and (n13703,n13704,n4903);
or (n13704,1'b0,n13705,n13706,n13707,n13708);
and (n13705,n5782,n556);
and (n13706,n5785,n567);
and (n13707,n5788,n571);
and (n13708,n5791,n573);
or (n13709,1'b0,n13710,n13717,n13719,n13720);
and (n13710,n13711,n2893);
wire s0n13711,s1n13711,notn13711;
or (n13711,s0n13711,s1n13711);
not(notn13711,n2891);
and (s0n13711,notn13711,1'b0);
and (s1n13711,n2891,n13712);
wire s0n13712,s1n13712,notn13712;
or (n13712,s0n13712,s1n13712);
not(notn13712,n13046);
and (s0n13712,notn13712,n13713);
and (s1n13712,n13046,1'b0);
wire s0n13713,s1n13713,notn13713;
or (n13713,s0n13713,s1n13713);
not(notn13713,n13031);
and (s0n13713,notn13713,n13714);
and (s1n13713,n13031,1'b1);
wire s0n13714,s1n13714,notn13714;
or (n13714,s0n13714,s1n13714);
not(notn13714,n4966);
and (s0n13714,notn13714,n13715);
and (s1n13714,n4966,n13163);
wire s0n13715,s1n13715,notn13715;
or (n13715,s0n13715,s1n13715);
not(notn13715,n4966);
and (s0n13715,notn13715,n13716);
and (s1n13715,n4966,n12805);
xor (n13716,n12805,n12807);
and (n13717,n13718,n2907);
wire s0n13718,s1n13718,notn13718;
or (n13718,s0n13718,s1n13718);
not(notn13718,n2902);
and (s0n13718,notn13718,1'b0);
and (s1n13718,n2902,n13712);
and (n13719,n13712,n7875);
and (n13720,n13624,n7878);
and (n13721,n13709,n13722);
and (n13722,n13723,n13816);
or (n13723,1'b0,n13724,n13727,n13730,n13735);
and (n13724,n13725,n2893);
wire s0n13725,s1n13725,notn13725;
or (n13725,s0n13725,s1n13725);
not(notn13725,n2891);
and (s0n13725,notn13725,1'b0);
and (s1n13725,n2891,n13726);
and (n13727,n13728,n2907);
wire s0n13728,s1n13728,notn13728;
or (n13728,s0n13728,s1n13728);
not(notn13728,n2902);
and (s0n13728,notn13728,1'b0);
and (s1n13728,n2902,n13729);
and (n13730,n13731,n4883);
wire s0n13731,s1n13731,notn13731;
or (n13731,s0n13731,s1n13731);
not(notn13731,n11666);
and (s0n13731,notn13731,n13732);
and (s1n13731,n11666,1'b0);
wire s0n13732,s1n13732,notn13732;
or (n13732,s0n13732,s1n13732);
not(notn13732,n11661);
and (s0n13732,notn13732,n13733);
and (s1n13732,n11661,1'b1);
wire s0n13733,s1n13733,notn13733;
or (n13733,s0n13733,s1n13733);
not(notn13733,n4861);
and (s0n13733,notn13733,1'b0);
and (s1n13733,n4861,n13734);
xor (n13734,n11657,n11659);
or (n13735,1'b0,n13736,n13756,n13776,n13796);
and (n13736,n13737,n2718);
or (n13737,1'b0,n13738,n13744,n13750);
and (n13738,n13739,n4895);
or (n13739,1'b0,n13740,n13741,n13742,n13743);
and (n13740,n5948,n556);
and (n13741,n5952,n567);
and (n13742,n5955,n571);
and (n13743,n5958,n573);
and (n13744,n13745,n2944);
or (n13745,1'b0,n13746,n13747,n13748,n13749);
and (n13746,n7314,n556);
and (n13747,n7313,n567);
and (n13748,n7317,n571);
and (n13749,n7320,n573);
and (n13750,n13751,n4903);
or (n13751,1'b0,n13752,n13753,n13754,n13755);
and (n13752,n7313,n556);
and (n13753,n7317,n567);
and (n13754,n7320,n571);
and (n13755,n7323,n573);
and (n13756,n13757,n2730);
or (n13757,1'b0,n13758,n13764,n13770);
and (n13758,n13759,n4895);
or (n13759,1'b0,n13760,n13761,n13762,n13763);
and (n13760,n5963,n556);
and (n13761,n5966,n567);
and (n13762,n5969,n571);
and (n13763,n5972,n573);
and (n13764,n13765,n2944);
or (n13765,1'b0,n13766,n13767,n13768,n13769);
and (n13766,n7323,n556);
and (n13767,n7328,n567);
and (n13768,n7331,n571);
and (n13769,n7334,n573);
and (n13770,n13771,n4903);
or (n13771,1'b0,n13772,n13773,n13774,n13775);
and (n13772,n7328,n556);
and (n13773,n7331,n567);
and (n13774,n7334,n571);
and (n13775,n7337,n573);
and (n13776,n13777,n2742);
or (n13777,1'b0,n13778,n13784,n13790);
and (n13778,n13779,n4895);
or (n13779,1'b0,n13780,n13781,n13782,n13783);
and (n13780,n5977,n556);
and (n13781,n5981,n567);
and (n13782,n5984,n571);
and (n13783,n5987,n573);
and (n13784,n13785,n2944);
or (n13785,1'b0,n13786,n13787,n13788,n13789);
and (n13786,n5890,n556);
and (n13787,n5889,n567);
and (n13788,n5893,n571);
and (n13789,n5896,n573);
and (n13790,n13791,n4903);
or (n13791,1'b0,n13792,n13793,n13794,n13795);
and (n13792,n5889,n556);
and (n13793,n5893,n567);
and (n13794,n5896,n571);
and (n13795,n5899,n573);
and (n13796,n13797,n2752);
or (n13797,1'b0,n13798,n13804,n13810);
and (n13798,n13799,n4895);
or (n13799,1'b0,n13800,n13801,n13802,n13803);
and (n13800,n5992,n556);
and (n13801,n5995,n567);
and (n13802,n5998,n571);
and (n13803,n6001,n573);
and (n13804,n13805,n2944);
or (n13805,1'b0,n13806,n13807,n13808,n13809);
and (n13806,n5899,n556);
and (n13807,n5904,n567);
and (n13808,n5907,n571);
and (n13809,n5910,n573);
and (n13810,n13811,n4903);
or (n13811,1'b0,n13812,n13813,n13814,n13815);
and (n13812,n5904,n556);
and (n13813,n5907,n567);
and (n13814,n5910,n571);
and (n13815,n5913,n573);
or (n13816,1'b0,n13817,n13824,n13826,n13827);
and (n13817,n13818,n2893);
wire s0n13818,s1n13818,notn13818;
or (n13818,s0n13818,s1n13818);
not(notn13818,n2891);
and (s0n13818,notn13818,1'b0);
and (s1n13818,n2891,n13819);
wire s0n13819,s1n13819,notn13819;
or (n13819,s0n13819,s1n13819);
not(notn13819,n13046);
and (s0n13819,notn13819,n13820);
and (s1n13819,n13046,1'b0);
wire s0n13820,s1n13820,notn13820;
or (n13820,s0n13820,s1n13820);
not(notn13820,n13031);
and (s0n13820,notn13820,n13821);
and (s1n13820,n13031,1'b1);
wire s0n13821,s1n13821,notn13821;
or (n13821,s0n13821,s1n13821);
not(notn13821,n4966);
and (s0n13821,notn13821,n13822);
and (s1n13821,n4966,n13275);
wire s0n13822,s1n13822,notn13822;
or (n13822,s0n13822,s1n13822);
not(notn13822,n4966);
and (s0n13822,notn13822,n13823);
and (s1n13822,n4966,n12808);
xor (n13823,n12808,n12810);
and (n13824,n13825,n2907);
wire s0n13825,s1n13825,notn13825;
or (n13825,s0n13825,s1n13825);
not(notn13825,n2902);
and (s0n13825,notn13825,1'b0);
and (s1n13825,n2902,n13819);
and (n13826,n13819,n7875);
and (n13827,n13731,n7878);
and (n13828,n13616,n13722);
and (n13829,n13508,n13614);
and (n13830,n13400,n13506);
and (n13831,n13288,n13398);
and (n13832,n13176,n13286);
and (n13833,n13064,n13174);
and (n13834,n9938,n13062);
and (n13835,n13836,n13838);
xor (n13836,n13837,n13062);
xor (n13837,n9938,n11732);
and (n13838,n13839,n13841);
xor (n13839,n13840,n13174);
xor (n13840,n13064,n13157);
and (n13841,n13842,n13844);
xor (n13842,n13843,n13286);
xor (n13843,n13176,n13269);
and (n13844,n13845,n13847);
xor (n13845,n13846,n13398);
xor (n13846,n13288,n13381);
and (n13847,n13848,n13850);
xor (n13848,n13849,n13506);
xor (n13849,n13400,n13493);
and (n13850,n13851,n13853);
xor (n13851,n13852,n13614);
xor (n13852,n13508,n13601);
and (n13853,n13854,n13856);
xor (n13854,n13855,n13722);
xor (n13855,n13616,n13709);
xor (n13856,n13723,n13816);
and (n13857,n13858,n8677);
wire s0n13858,s1n13858,notn13858;
or (n13858,s0n13858,s1n13858);
not(notn13858,n4969);
and (s0n13858,notn13858,1'b0);
and (s1n13858,n4969,n9935);
and (n13859,n11734,n2950);
and (n13860,n11735,n5024);
and (n13861,n9946,n2941);
and (n13862,n3,n13863);
not (n13863,n573);
or (n13864,n13865,n13866);
and (n13865,n8700,n2905);
and (n13866,n3,n13867);
not (n13867,n2905);
wire s0n13868,s1n13868,notn13868;
or (n13868,s0n13868,s1n13868);
not(notn13868,n19815);
and (s0n13868,notn13868,n13869);
and (s1n13868,n19815,n19814);
wire s0n13869,s1n13869,notn13869;
or (n13869,s0n13869,s1n13869);
not(notn13869,n19813);
and (s0n13869,notn13869,n13870);
and (s1n13869,n19813,n17724);
or (n13870,n13871,n17723);
and (n13871,n13872,n14131);
wire s0n13872,s1n13872,notn13872;
or (n13872,s0n13872,s1n13872);
not(notn13872,n17028);
and (s0n13872,notn13872,n13873);
and (s1n13872,n17028,n13883);
wire s0n13873,s1n13873,notn13873;
or (n13873,s0n13873,s1n13873);
not(notn13873,n14503);
and (s0n13873,notn13873,n13874);
and (s1n13873,n14503,n17618);
wire s0n13874,s1n13874,notn13874;
or (n13874,s0n13874,s1n13874);
not(notn13874,n14503);
and (s0n13874,notn13874,n13875);
and (s1n13874,n14503,n17537);
wire s0n13875,s1n13875,notn13875;
or (n13875,s0n13875,s1n13875);
not(notn13875,n17294);
and (s0n13875,notn13875,n13876);
and (s1n13875,n17294,n17444);
wire s0n13876,s1n13876,notn13876;
or (n13876,s0n13876,s1n13876);
not(notn13876,n17443);
and (s0n13876,notn13876,n13877);
and (s1n13876,n17443,n17392);
xor (n13877,n13878,n17363);
xor (n13878,n13879,n17298);
xor (n13879,n13880,n17040);
wire s0n13880,s1n13880,notn13880;
or (n13880,s0n13880,s1n13880);
not(notn13880,n17028);
and (s0n13880,notn13880,n13881);
and (s1n13880,n17028,1'b0);
xor (n13881,n13882,n14633);
xor (n13882,n13883,n14550);
nand (n13883,n13884,n14334,n14514);
nor (n13884,n13885,n14132);
and (n13885,n13886,n14108);
or (n13886,1'b0,n13887,n13895,n13898,n13901);
and (n13887,n13888,n13889);
and (n13889,n13890,n13891,n13893);
not (n13891,n13892);
not (n13893,n13894);
and (n13895,n13896,n13897);
nor (n13897,n13890,n13891,n13894);
and (n13898,n13899,n13900);
and (n13900,n13890,n13892,n13893);
and (n13901,n13902,n14131);
wire s0n13902,s1n13902,notn13902;
or (n13902,s0n13902,s1n13902);
not(notn13902,n14123);
and (s0n13902,notn13902,1'b0);
and (s1n13902,n14123,n13903);
wire s0n13903,s1n13903,notn13903;
or (n13903,s0n13903,s1n13903);
not(notn13903,n555);
and (s0n13903,notn13903,n13904);
and (s1n13903,n555,n14112);
wire s0n13904,s1n13904,notn13904;
or (n13904,s0n13904,s1n13904);
not(notn13904,n13948);
and (s0n13904,notn13904,n13905);
and (s1n13904,n13948,n13910);
wire s0n13905,s1n13905,notn13905;
or (n13905,s0n13905,s1n13905);
not(notn13905,n13907);
and (s0n13905,notn13905,1'b0);
and (s1n13905,n13907,n13906);
and (n13907,n13908,n13909);
or (n13910,n13911,n13918,n13921,n13926,n13933,n13940);
and (n13911,n13912,n13913);
or (n13913,n13914,n13917);
or (n13914,n13915,n13916);
nor (n13915,n28,n29,n585,n582);
nor (n13916,n33,n2773,n585,n582);
and (n13917,n33,n29,n581,n582);
and (n13918,n13919,n13920);
and (n13920,n33,n2773,n581,n582);
and (n13921,n13922,n13923);
or (n13923,n13924,n13925);
and (n13924,n28,n2773,n585,n582);
and (n13925,n28,n29,n581,n582);
and (n13926,n13927,n13928);
or (n13928,n13929,n13932);
or (n13929,n13930,n13931);
nor (n13930,n33,n29,n581,n582);
nor (n13931,n28,n2773,n585,n582);
and (n13932,n28,n29,n585,n582);
and (n13933,n13934,n13935);
or (n13935,n13936,n13939);
or (n13936,n13937,n13938);
nor (n13937,n33,n2773,n581,n582);
nor (n13938,n33,n29,n585,n582);
and (n13939,n28,n2773,n581,n582);
and (n13940,n13906,n13941);
or (n13941,n13942,n13947);
or (n13942,n13943,n13946);
or (n13943,n13944,n13945);
nor (n13944,n28,n29,n581,n582);
nor (n13945,n28,n2773,n581,n582);
and (n13946,n33,n2773,n585,n582);
and (n13947,n33,n29,n585,n582);
or (n13948,n13949,n14111);
or (n13949,n13950,n14108);
nor (n13950,n13951,n14005,n14039,n14074);
wire s0n13951,s1n13951,notn13951;
or (n13951,s0n13951,s1n13951);
not(notn13951,n13985);
and (s0n13951,notn13951,1'b1);
and (s1n13951,n13985,n13952);
or (n13952,n555,n13953,n13955,n13957,n13959,n13961,n13963,n13965,n13967,n13969,n13971,n13973,n13975,n13977,n13979,n13981,n13983);
and (n13953,n13954,n2768);
and (n13955,n13956,n2770);
and (n13957,n13958,n2772);
and (n13959,n13960,n2775);
and (n13961,n13962,n2777);
and (n13963,n13964,n2779);
and (n13965,n13966,n2781);
and (n13967,n13968,n2783);
and (n13969,n13970,n2785);
and (n13971,n13972,n2787);
and (n13973,n13974,n2789);
and (n13975,n13976,n2791);
and (n13977,n13978,n2793);
and (n13979,n13980,n2795);
and (n13981,n13982,n2797);
and (n13983,n13984,n2799);
and (n13985,n13986,n13994,n14000,n42);
not (n13986,n13987);
wire s0n13987,s1n13987,notn13987;
or (n13987,s0n13987,s1n13987);
not(notn13987,n554);
and (s0n13987,notn13987,n13988);
and (s1n13987,n554,1'b1);
wire s0n13988,s1n13988,notn13988;
or (n13988,s0n13988,s1n13988);
not(notn13988,n184);
and (s0n13988,notn13988,n13989);
and (s1n13988,n184,n13990);
wire s0n13990,s1n13990,notn13990;
or (n13990,s0n13990,s1n13990);
not(notn13990,n547);
and (s0n13990,notn13990,n13991);
and (s1n13990,n547,n529);
or (n13991,n47,1'b0,1'b0,1'b0,n545,1'b0,n13992,1'b0);
or (n13992,n543,n13993);
nor (n13993,n297,n543,n544,n545,n546,n520,n497,n498,n499,n500,n501,n502,n503,n504,n54,n479,n481,n483,n484,n486,n487,n488,n512,n513,n514,n515,n516,n517,n518,n519);
not (n13994,n13995);
wire s0n13995,s1n13995,notn13995;
or (n13995,s0n13995,s1n13995);
not(notn13995,n554);
and (s0n13995,notn13995,n13996);
and (s1n13995,n554,1'b0);
wire s0n13996,s1n13996,notn13996;
or (n13996,s0n13996,s1n13996);
not(notn13996,n184);
and (s0n13996,notn13996,n13997);
and (s1n13996,n184,n13998);
wire s0n13998,s1n13998,notn13998;
or (n13998,s0n13998,s1n13998);
not(notn13998,n547);
and (s0n13998,notn13998,n13999);
and (s1n13998,n547,n522);
or (n13999,1'b0,1'b0,1'b0,1'b0,n545,n544,1'b0,1'b0);
wire s0n14000,s1n14000,notn14000;
or (n14000,s0n14000,s1n14000);
not(notn14000,n554);
and (s0n14000,notn14000,n14001);
and (s1n14000,n554,1'b1);
wire s0n14001,s1n14001,notn14001;
or (n14001,s0n14001,s1n14001);
not(notn14001,n184);
and (s0n14001,notn14001,n14002);
and (s1n14001,n184,n14003);
wire s0n14003,s1n14003,notn14003;
or (n14003,s0n14003,s1n14003);
not(notn14003,n547);
and (s0n14003,notn14003,n14004);
and (s1n14003,n547,n297);
or (n14004,1'b0,1'b0,n520,n546,1'b0,1'b0,1'b0,1'b0);
wire s0n14005,s1n14005,notn14005;
or (n14005,s0n14005,s1n14005);
not(notn14005,n13985);
and (s0n14005,notn14005,1'b1);
and (s1n14005,n13985,n14006);
or (n14006,n555,n14007,n14009,n14011,n14013,n14015,n14017,n14019,n14021,n14023,n14025,n14027,n14029,n14031,n14033,n14035,n14037);
and (n14007,n14008,n2768);
and (n14009,n14010,n2770);
and (n14011,n14012,n2772);
and (n14013,n14014,n2775);
and (n14015,n14016,n2777);
and (n14017,n14018,n2779);
and (n14019,n14020,n2781);
and (n14021,n14022,n2783);
and (n14023,n14024,n2785);
and (n14025,n14026,n2787);
and (n14027,n14028,n2789);
and (n14029,n14030,n2791);
and (n14031,n14032,n2793);
and (n14033,n14034,n2795);
and (n14035,n14036,n2797);
and (n14037,n14038,n2799);
not (n14039,n14040);
wire s0n14040,s1n14040,notn14040;
or (n14040,s0n14040,s1n14040);
not(notn14040,n13985);
and (s0n14040,notn14040,1'b1);
and (s1n14040,n13985,n14041);
or (n14041,n555,n14042,n14044,n14046,n14048,n14050,n14052,n14054,n14056,n14058,n14060,n14062,n14064,n14066,n14068,n14070,n14072);
and (n14042,n14043,n2768);
and (n14044,n14045,n2770);
and (n14046,n14047,n2772);
and (n14048,n14049,n2775);
and (n14050,n14051,n2777);
and (n14052,n14053,n2779);
and (n14054,n14055,n2781);
and (n14056,n14057,n2783);
and (n14058,n14059,n2785);
and (n14060,n14061,n2787);
and (n14062,n14063,n2789);
and (n14064,n14065,n2791);
and (n14066,n14067,n2793);
and (n14068,n14069,n2795);
and (n14070,n14071,n2797);
and (n14072,n14073,n2799);
wire s0n14074,s1n14074,notn14074;
or (n14074,s0n14074,s1n14074);
not(notn14074,n13985);
and (s0n14074,notn14074,1'b1);
and (s1n14074,n13985,n14075);
or (n14075,n555,n14076,n14078,n14080,n14082,n14084,n14086,n14088,n14090,n14092,n14094,n14096,n14098,n14100,n14102,n14104,n14106);
and (n14076,n14077,n2768);
and (n14078,n14079,n2770);
and (n14080,n14081,n2772);
and (n14082,n14083,n2775);
and (n14084,n14085,n2777);
and (n14086,n14087,n2779);
and (n14088,n14089,n2781);
and (n14090,n14091,n2783);
and (n14092,n14093,n2785);
and (n14094,n14095,n2787);
and (n14096,n14097,n2789);
and (n14098,n14099,n2791);
and (n14100,n14101,n2793);
and (n14102,n14103,n2795);
and (n14104,n14105,n2797);
and (n14106,n14107,n2799);
and (n14108,n13951,n14109,n14040,n14110);
not (n14109,n14005);
not (n14110,n14074);
nor (n14111,n13951,n14109,n14039,n14074);
wire s0n14112,s1n14112,notn14112;
or (n14112,s0n14112,s1n14112);
not(notn14112,n14119);
and (s0n14112,notn14112,1'b0);
and (s1n14112,n14119,n14113);
wire s0n14113,s1n14113,notn14113;
or (n14113,s0n14113,s1n14113);
not(notn14113,n14116);
and (s0n14113,notn14113,n14114);
and (s1n14113,n14116,n14115);
not (n14116,n14117);
and (n14117,n555,n14118);
not (n14118,n589);
and (n14119,n555,n14120);
and (n14120,n14121,n14122);
and (n14123,n42,n14124);
or (n14124,n14125,n14126);
or (n14125,n13890,n13892,n13894);
or (n14126,n14127,n14128,n14129,n14130);
nor (n14131,n13890,n13892,n13893);
nand (n14132,n14133,n14244,n14259);
nor (n14133,n14134,n14231,n14241);
and (n14134,n14135,n14138);
not (n14135,n14136);
nand (n14136,n14137,n13889);
and (n14137,n13951,n14005,n14040,n14110);
wire s0n14138,s1n14138,notn14138;
or (n14138,s0n14138,s1n14138);
not(notn14138,n14227);
and (s0n14138,notn14138,1'b0);
and (s1n14138,n14227,n14139);
or (n14139,1'b0,n14140,n14197,n14201,n14203,n14207,n14224);
and (n14140,n14141,n14193);
wire s0n14141,s1n14141,notn14141;
or (n14141,s0n14141,s1n14141);
not(notn14141,n42);
and (s0n14141,notn14141,1'b0);
and (s1n14141,n42,n14142);
wire s0n14142,s1n14142,notn14142;
or (n14142,s0n14142,s1n14142);
not(notn14142,n14187);
and (s0n14142,notn14142,n14143);
and (s1n14142,n14187,n14168);
wire s0n14143,s1n14143,notn14143;
or (n14143,s0n14143,s1n14143);
not(notn14143,n14163);
and (s0n14143,notn14143,1'b0);
and (s1n14143,n14163,n14144);
or (n14144,1'b0,n14145,n14154);
and (n14145,n14146,n14147);
or (n14147,n14148,n14153);
or (n14148,n14149,n14152);
or (n14149,n14150,n14151);
nor (n14150,n33,n29,n581,n582,n591);
nor (n14151,n33,n2773,n581,n582,n591);
nor (n14152,n33,n29,n585,n582,n591);
nor (n14153,n33,n2773,n585,n582,n591);
and (n14154,n14155,n14156);
or (n14156,n14157,n14162);
or (n14157,n14158,n14161);
or (n14158,n14159,n14160);
nor (n14159,n28,n29,n581,n582,n591);
nor (n14160,n28,n2773,n581,n582,n591);
nor (n14161,n28,n29,n585,n582,n591);
nor (n14162,n28,n2773,n585,n582,n591);
and (n14163,n14164,n14125);
and (n14164,n14165,n14167);
and (n14165,n555,n14166);
nand (n14166,n582,n555);
not (n14167,n14121);
or (n14168,1'b0,n14169,n14174,n14179,n14183);
and (n14169,n14170,n14171);
or (n14171,n14172,n2768);
or (n14172,n14173,n2772);
or (n14173,n2789,n2785);
and (n14174,n14175,n14176);
or (n14176,n14177,n2770);
or (n14177,n14178,n2775);
or (n14178,n2791,n2787);
and (n14179,n14146,n14180);
or (n14180,n14181,n2777);
or (n14181,n14182,n2781);
or (n14182,n2797,n2793);
and (n14183,n14155,n14184);
or (n14184,n14185,n2779);
or (n14185,n14186,n2783);
or (n14186,n2799,n2795);
and (n14187,n14188,n14189);
and (n14188,n591,n14125);
or (n14189,n14000,n14190);
and (n14190,n14191,n14192);
not (n14191,n14000);
nor (n14192,n13908,n13909);
or (n14193,n14194,n2768);
or (n14194,n14195,n2772);
or (n14195,n14196,n2785);
or (n14196,n2793,n2777);
and (n14197,n14198,n14199);
or (n14199,n14200,n2770);
or (n14200,n2787,n2775);
and (n14201,n14202,n2781);
and (n14203,n14204,n14205);
or (n14205,n14206,n2779);
or (n14206,n2795,n2783);
and (n14207,n14208,n2789);
wire s0n14208,s1n14208,notn14208;
or (n14208,s0n14208,s1n14208);
not(notn14208,n14210);
and (s0n14208,notn14208,n14170);
and (s1n14208,n14210,n14209);
and (n14210,n14211,n14217);
and (n14211,n42,n14212);
or (n14212,n14213,n14214,n14215,n14216);
nand (n14217,n14218,n14220,n14221,n14223);
not (n14218,n14219);
not (n14221,n14222);
and (n14224,n14209,n14225);
or (n14225,n14226,n2791);
or (n14226,n2799,n2797);
nor (n14227,n14074,n14228);
nand (n14228,n14005,n13951,n14229);
nor (n14229,n14191,n14230);
nand (n14230,n42,n14125,n591);
and (n14231,n14232,n14240);
nand (n14232,n14233,n14238);
or (n14233,n14234,n14236);
not (n14234,n14235);
or (n14235,n13897,n13889);
not (n14236,n14237);
nor (n14237,n13951,n14005,n14040,n14110);
nand (n14238,n14239,n13900);
and (n14239,n13951,n14005,n14039,n14110);
and (n14241,n14242,n14141);
and (n14242,n14137,n14243);
or (n14243,n13900,n13897);
not (n14244,n14245);
and (n14245,n14246,n14137);
and (n14246,n14247,n14131);
wire s0n14247,s1n14247,notn14247;
or (n14247,s0n14247,s1n14247);
not(notn14247,n42);
and (s0n14247,notn14247,1'b0);
and (s1n14247,n42,n14248);
wire s0n14248,s1n14248,notn14248;
or (n14248,s0n14248,s1n14248);
not(notn14248,n14187);
and (s0n14248,notn14248,n14249);
and (s1n14248,n14187,n14254);
wire s0n14249,s1n14249,notn14249;
or (n14249,s0n14249,s1n14249);
not(notn14249,n14163);
and (s0n14249,notn14249,1'b0);
and (s1n14249,n14163,n14250);
or (n14250,1'b0,n14251,n14252);
and (n14251,n14204,n14147);
and (n14252,n14253,n14156);
or (n14254,1'b0,n14255,n14256,n14257,n14258);
and (n14255,n14198,n14171);
and (n14256,n14202,n14176);
and (n14257,n14204,n14180);
and (n14258,n14253,n14184);
not (n14259,n14260);
nand (n14260,n14261,n14329);
nor (n14261,n14262,n14295,n14312);
and (n14262,n14263,n14280);
and (n14263,n14264,n13897);
nand (n14264,n14265,n14267);
not (n14265,n14266);
nor (n14266,n13951,n14005,n14040,n14074);
nor (n14267,n14268,n14274);
and (n14268,n14269,n14273);
nor (n14269,n14270,n13909);
not (n14270,n14271);
and (n14271,n14272,n591);
and (n14272,n14191,n42);
not (n14273,n13908);
nor (n14274,n14275,n14121);
not (n14275,n14276);
nor (n14276,n14277,n14278);
not (n14277,n14122);
not (n14278,n14279);
and (n14279,n42,n555);
wire s0n14280,s1n14280,notn14280;
or (n14280,s0n14280,s1n14280);
not(notn14280,n42);
and (s0n14280,notn14280,1'b0);
and (s1n14280,n42,n14281);
wire s0n14281,s1n14281,notn14281;
or (n14281,s0n14281,s1n14281);
not(notn14281,n14187);
and (s0n14281,notn14281,n14282);
and (s1n14281,n14187,n14288);
wire s0n14282,s1n14282,notn14282;
or (n14282,s0n14282,s1n14282);
not(notn14282,n14163);
and (s0n14282,notn14282,1'b0);
and (s1n14282,n14163,n14283);
or (n14283,1'b0,n14284,n14286);
and (n14284,n14285,n14147);
and (n14286,n14287,n14156);
or (n14288,1'b0,n14289,n14291,n14293,n14294);
and (n14289,n14290,n14171);
and (n14291,n14292,n14176);
and (n14293,n14285,n14180);
and (n14294,n14287,n14184);
and (n14295,n14296,n14297);
and (n14296,n14264,n14131);
wire s0n14297,s1n14297,notn14297;
or (n14297,s0n14297,s1n14297);
not(notn14297,n42);
and (s0n14297,notn14297,1'b0);
and (s1n14297,n42,n14298);
wire s0n14298,s1n14298,notn14298;
or (n14298,s0n14298,s1n14298);
not(notn14298,n14187);
and (s0n14298,notn14298,n14299);
and (s1n14298,n14187,n14305);
wire s0n14299,s1n14299,notn14299;
or (n14299,s0n14299,s1n14299);
not(notn14299,n14163);
and (s0n14299,notn14299,1'b0);
and (s1n14299,n14163,n14300);
or (n14300,1'b0,n14301,n14303);
and (n14301,n14302,n14147);
and (n14303,n14304,n14156);
or (n14305,1'b0,n14306,n14308,n14310,n14311);
and (n14306,n14307,n14171);
and (n14308,n14309,n14176);
and (n14310,n14302,n14180);
and (n14311,n14304,n14184);
wire s0n14312,s1n14312,notn14312;
or (n14312,s0n14312,s1n14312);
not(notn14312,n14326);
and (s0n14312,notn14312,n14313);
and (s1n14312,n14326,n14318);
wire s0n14313,s1n14313,notn14313;
or (n14313,s0n14313,s1n14313);
not(notn14313,n14315);
and (s0n14313,notn14313,1'b0);
and (s1n14313,n14315,n14314);
and (n14315,n14316,n14279);
and (n14316,n14317,n14120);
and (n14317,n14131,n33);
or (n14318,1'b0,n14319,n14322,n14325);
and (n14319,n14320,n14321);
or (n14321,n2787,n2770);
and (n14322,n14323,n14324);
or (n14324,n2791,n2775);
and (n14325,n14314,n14184);
and (n14326,n14327,n591);
and (n14327,n14328,n14131);
and (n14328,n14272,n13907);
nor (n14329,n14330,n14332);
and (n14330,n14331,n14141);
and (n14331,n14264,n13889);
and (n14332,n14333,n14247);
and (n14333,n14264,n13900);
nor (n14334,n14335,n14342);
and (n14335,n14336,n14341);
nand (n14336,n14337,n14340);
or (n14337,n14338,n14339);
not (n14338,n13900);
not (n14339,n13950);
nand (n14340,n14111,n13897);
nand (n14342,n14343,n14432,n14442,n14487);
nor (n14343,n14344,n14425,n14429);
and (n14344,n14345,n14346);
and (n14345,n14131,n14111);
wire s0n14346,s1n14346,notn14346;
or (n14346,s0n14346,s1n14346);
not(notn14346,n42);
and (s0n14346,notn14346,1'b0);
and (s1n14346,n42,n14347);
wire s0n14347,s1n14347,notn14347;
or (n14347,s0n14347,s1n14347);
not(notn14347,n14422);
and (s0n14347,notn14347,n14348);
and (s1n14347,n14422,n14370);
wire s0n14348,s1n14348,notn14348;
or (n14348,s0n14348,s1n14348);
not(notn14348,n14362);
and (s0n14348,notn14348,1'b0);
and (s1n14348,n14362,n14349);
or (n14349,1'b0,n14350,n14353,n14356,n14359);
and (n14350,n14351,n14352);
or (n14352,n14162,n14153);
and (n14353,n14354,n14355);
or (n14355,n14161,n14152);
and (n14356,n14357,n14358);
or (n14358,n14160,n14151);
and (n14359,n14360,n14361);
or (n14361,n14159,n14150);
and (n14362,n14363,n14364);
and (n14363,n555,n14125);
or (n14364,n14365,n14366);
and (n14365,n14121,n14277);
and (n14366,n14367,n14368);
nor (n14367,n14121,n14122);
and (n14368,n42,n14369);
or (n14369,n14219,n14220,n14222,n14223);
or (n14370,1'b0,n14371,n14390,n14396,n14415);
and (n14371,n14372,n14387);
wire s0n14372,s1n14372,notn14372;
or (n14372,s0n14372,s1n14372);
not(notn14372,n14374);
and (s0n14372,notn14372,1'b0);
and (s1n14372,n14374,n14373);
and (n14374,n42,n14375);
and (n14375,n591,n14376);
or (n14376,n14000,n14377);
and (n14377,n14191,n14378);
or (n14378,n14379,n14386);
or (n14379,n14380,n14383);
and (n14380,n14381,n14125);
and (n14381,n13908,n14382);
not (n14382,n13909);
and (n14383,n14384,n14368);
and (n14384,n14385,n14125);
nor (n14385,n13908,n14382);
and (n14386,n13907,n14126);
or (n14387,n14388,n2768);
or (n14388,n14389,n2770);
or (n14389,n2779,n2777);
and (n14390,n14391,n14393);
wire s0n14391,s1n14391,notn14391;
or (n14391,s0n14391,s1n14391);
not(notn14391,n14374);
and (s0n14391,notn14391,1'b0);
and (s1n14391,n14374,n14392);
or (n14393,n14394,n2772);
or (n14394,n14395,n2775);
or (n14395,n2783,n2781);
and (n14396,n14397,n14412);
wire s0n14397,s1n14397,notn14397;
or (n14397,s0n14397,s1n14397);
not(notn14397,n42);
and (s0n14397,notn14397,1'b0);
and (s1n14397,n42,n14398);
wire s0n14398,s1n14398,notn14398;
or (n14398,s0n14398,s1n14398);
not(notn14398,n14375);
and (s0n14398,notn14398,n14399);
and (s1n14398,n14375,n14411);
wire s0n14399,s1n14399,notn14399;
or (n14399,s0n14399,s1n14399);
not(notn14399,n14409);
and (s0n14399,notn14399,n14400);
and (s1n14399,n14409,n14357);
wire s0n14400,s1n14400,notn14400;
or (n14400,s0n14400,s1n14400);
not(notn14400,n14401);
and (s0n14400,notn14400,1'b0);
and (s1n14400,n14401,n14351);
and (n14401,n14402,n14403);
and (n14402,n14117,n14166);
or (n14403,n14404,n14408);
or (n14404,n14405,n14406);
and (n14405,n14365,n14125);
and (n14406,n14407,n14368);
and (n14407,n14367,n14125);
and (n14408,n14120,n14126);
and (n14409,n14410,n14403);
and (n14410,n555,n14116);
or (n14412,n14413,n2785);
or (n14413,n14414,n2787);
or (n14414,n2795,n2793);
and (n14415,n14416,n14421);
wire s0n14416,s1n14416,notn14416;
or (n14416,s0n14416,s1n14416);
not(notn14416,n42);
and (s0n14416,notn14416,1'b0);
and (s1n14416,n42,n14417);
wire s0n14417,s1n14417,notn14417;
or (n14417,s0n14417,s1n14417);
not(notn14417,n14375);
and (s0n14417,notn14417,n14418);
and (s1n14417,n14375,n14420);
wire s0n14418,s1n14418,notn14418;
or (n14418,s0n14418,s1n14418);
not(notn14418,n14409);
and (s0n14418,notn14418,n14419);
and (s1n14418,n14409,n14360);
wire s0n14419,s1n14419,notn14419;
or (n14419,s0n14419,s1n14419);
not(notn14419,n14401);
and (s0n14419,notn14419,1'b0);
and (s1n14419,n14401,n14354);
or (n14421,n14225,n2789);
and (n14422,n14188,n14423);
or (n14423,n14000,n14424);
and (n14424,n14191,n14381);
and (n14425,n14426,n14428);
not (n14426,n14427);
nand (n14427,n14239,n13897);
and (n14429,n14430,n13899);
not (n14430,n14431);
nand (n14431,n13950,n13897);
nor (n14432,n14433,n14437);
and (n14433,n14434,n14436);
not (n14434,n14435);
nand (n14435,n14111,n13889);
and (n14437,n14438,n14441);
nor (n14438,n14439,n14440);
not (n14439,n14239);
not (n14440,n13889);
nand (n14442,n14443,n14456);
not (n14443,n14444);
nor (n14444,n14445,n14453);
and (n14445,n14446,n14125);
nand (n14446,n14447,n14450);
not (n14447,n14448);
nor (n14448,n14449,n14005,n14040,n14074);
not (n14449,n13951);
nor (n14450,n14451,n14452);
and (n14451,n14269,n13908);
nor (n14452,n14167,n14278,n14122);
nor (n14453,n14236,n14454);
not (n14454,n14455);
or (n14455,n14131,n13900);
wire s0n14456,s1n14456,notn14456;
or (n14456,s0n14456,s1n14456);
not(notn14456,n42);
and (s0n14456,notn14456,1'b0);
and (s1n14456,n42,n14457);
wire s0n14457,s1n14457,notn14457;
or (n14457,s0n14457,s1n14457);
not(notn14457,n14422);
and (s0n14457,notn14457,n14458);
and (s1n14457,n14422,n14468);
wire s0n14458,s1n14458,notn14458;
or (n14458,s0n14458,s1n14458);
not(notn14458,n14362);
and (s0n14458,notn14458,1'b0);
and (s1n14458,n14362,n14459);
or (n14459,1'b0,n14460,n14462,n14464,n14466);
and (n14460,n14461,n14352);
and (n14462,n14463,n14355);
and (n14464,n14465,n14358);
and (n14466,n14467,n14361);
or (n14468,1'b0,n14469,n14472,n14475,n14481);
and (n14469,n14470,n14387);
wire s0n14470,s1n14470,notn14470;
or (n14470,s0n14470,s1n14470);
not(notn14470,n14374);
and (s0n14470,notn14470,1'b0);
and (s1n14470,n14374,n14471);
and (n14472,n14473,n14393);
wire s0n14473,s1n14473,notn14473;
or (n14473,s0n14473,s1n14473);
not(notn14473,n14374);
and (s0n14473,notn14473,1'b0);
and (s1n14473,n14374,n14474);
and (n14475,n14476,n14412);
wire s0n14476,s1n14476,notn14476;
or (n14476,s0n14476,s1n14476);
not(notn14476,n42);
and (s0n14476,notn14476,1'b0);
and (s1n14476,n42,n14477);
wire s0n14477,s1n14477,notn14477;
or (n14477,s0n14477,s1n14477);
not(notn14477,n14375);
and (s0n14477,notn14477,n14478);
and (s1n14477,n14375,n14480);
wire s0n14478,s1n14478,notn14478;
or (n14478,s0n14478,s1n14478);
not(notn14478,n14409);
and (s0n14478,notn14478,n14479);
and (s1n14478,n14409,n14465);
wire s0n14479,s1n14479,notn14479;
or (n14479,s0n14479,s1n14479);
not(notn14479,n14401);
and (s0n14479,notn14479,1'b0);
and (s1n14479,n14401,n14461);
and (n14481,n14482,n14421);
wire s0n14482,s1n14482,notn14482;
or (n14482,s0n14482,s1n14482);
not(notn14482,n42);
and (s0n14482,notn14482,1'b0);
and (s1n14482,n42,n14483);
wire s0n14483,s1n14483,notn14483;
or (n14483,s0n14483,s1n14483);
not(notn14483,n14375);
and (s0n14483,notn14483,n14484);
and (s1n14483,n14375,n14486);
wire s0n14484,s1n14484,notn14484;
or (n14484,s0n14484,s1n14484);
not(notn14484,n14409);
and (s0n14484,notn14484,n14485);
and (s1n14484,n14409,n14467);
wire s0n14485,s1n14485,notn14485;
or (n14485,s0n14485,s1n14485);
not(notn14485,n14401);
and (s0n14485,notn14485,1'b0);
and (s1n14485,n14401,n14463);
nor (n14487,n14488,n14492,n14508);
and (n14488,n14489,n13896);
not (n14489,n14490);
nand (n14490,n13949,n14491);
nor (n14491,n13951,n14440);
and (n14492,n14493,n14507);
not (n14493,n14494);
nor (n14494,n14495,n14501);
not (n14495,n14496);
nand (n14496,n14497,n13900);
nor (n14497,n14270,n14498);
nand (n14498,n14499,n14500,n585,n13909);
nor (n14499,n582,n29);
nor (n14500,n28,n13908);
nor (n14501,n14502,n14317);
not (n14502,n14503);
wire s0n14503,s1n14503,notn14503;
or (n14503,s0n14503,s1n14503);
not(notn14503,n14271);
and (s0n14503,notn14503,n14504);
and (s1n14503,n14271,n14506);
and (n14504,n14505,n14279);
and (n14505,n14125,n14120);
and (n14506,n14125,n13907);
and (n14508,n14509,n14511);
wire s0n14509,s1n14509,notn14509;
or (n14509,s0n14509,s1n14509);
not(notn14509,n14374);
and (s0n14509,notn14509,1'b0);
and (s1n14509,n14374,n14510);
nor (n14511,n14512,n14513);
not (n14512,n14497);
nand (n14513,n14368,n14131);
nor (n14514,n14515,n14548);
and (n14515,n14516,n14519);
nand (n14516,n14517,n14518);
nand (n14517,n14111,n13900);
nand (n14518,n13950,n14131);
wire s0n14519,s1n14519,notn14519;
or (n14519,s0n14519,s1n14519);
not(notn14519,n42);
and (s0n14519,notn14519,1'b0);
and (s1n14519,n42,n14520);
wire s0n14520,s1n14520,notn14520;
or (n14520,s0n14520,s1n14520);
not(notn14520,n14422);
and (s0n14520,notn14520,n14521);
and (s1n14520,n14422,n14531);
wire s0n14521,s1n14521,notn14521;
or (n14521,s0n14521,s1n14521);
not(notn14521,n14362);
and (s0n14521,notn14521,1'b0);
and (s1n14521,n14362,n14522);
or (n14522,1'b0,n14523,n14525,n14527,n14529);
and (n14523,n14524,n14352);
and (n14525,n14526,n14355);
and (n14527,n14528,n14358);
and (n14529,n14530,n14361);
or (n14531,1'b0,n14532,n14535,n14536,n14542);
and (n14532,n14533,n14387);
wire s0n14533,s1n14533,notn14533;
or (n14533,s0n14533,s1n14533);
not(notn14533,n14374);
and (s0n14533,notn14533,1'b0);
and (s1n14533,n14374,n14534);
and (n14535,n14509,n14393);
and (n14536,n14537,n14412);
wire s0n14537,s1n14537,notn14537;
or (n14537,s0n14537,s1n14537);
not(notn14537,n42);
and (s0n14537,notn14537,1'b0);
and (s1n14537,n42,n14538);
wire s0n14538,s1n14538,notn14538;
or (n14538,s0n14538,s1n14538);
not(notn14538,n14375);
and (s0n14538,notn14538,n14539);
and (s1n14538,n14375,n14541);
wire s0n14539,s1n14539,notn14539;
or (n14539,s0n14539,s1n14539);
not(notn14539,n14409);
and (s0n14539,notn14539,n14540);
and (s1n14539,n14409,n14528);
wire s0n14540,s1n14540,notn14540;
or (n14540,s0n14540,s1n14540);
not(notn14540,n14401);
and (s0n14540,notn14540,1'b0);
and (s1n14540,n14401,n14524);
and (n14542,n14543,n14421);
wire s0n14543,s1n14543,notn14543;
or (n14543,s0n14543,s1n14543);
not(notn14543,n42);
and (s0n14543,notn14543,1'b0);
and (s1n14543,n42,n14544);
wire s0n14544,s1n14544,notn14544;
or (n14544,s0n14544,s1n14544);
not(notn14544,n14375);
and (s0n14544,notn14544,n14545);
and (s1n14544,n14375,n14547);
wire s0n14545,s1n14545,notn14545;
or (n14545,s0n14545,s1n14545);
not(notn14545,n14409);
and (s0n14545,notn14545,n14546);
and (s1n14545,n14409,n14530);
wire s0n14546,s1n14546,notn14546;
or (n14546,s0n14546,s1n14546);
not(notn14546,n14401);
and (s0n14546,notn14546,1'b0);
and (s1n14546,n14401,n14526);
and (n14548,n14549,n14239);
and (n14549,n14280,n14131);
wire s0n14550,s1n14550,notn14550;
or (n14550,s0n14550,s1n14550);
not(notn14550,n14631);
and (s0n14550,notn14550,n14551);
and (s1n14550,n14631,n14574);
wire s0n14551,s1n14551,notn14551;
or (n14551,s0n14551,s1n14551);
not(notn14551,n14271);
and (s0n14551,notn14551,n14552);
and (s1n14551,n14271,n14558);
wire s0n14552,s1n14552,notn14552;
or (n14552,s0n14552,s1n14552);
not(notn14552,n14279);
and (s0n14552,notn14552,1'b0);
and (s1n14552,n14279,n14553);
and (n14553,n14554,n14120);
wire s0n14554,s1n14554,notn14554;
or (n14554,s0n14554,s1n14554);
not(notn14554,n14125);
and (s0n14554,notn14554,1'b0);
and (s1n14554,n14125,n14555);
wire s0n14555,s1n14555,notn14555;
or (n14555,s0n14555,s1n14555);
not(notn14555,n14317);
and (s0n14555,notn14555,n14556);
and (s1n14555,n14317,n14557);
or (n14558,n14559,n14565,1'b0);
and (n14559,n14560,n13907);
wire s0n14560,s1n14560,notn14560;
or (n14560,s0n14560,s1n14560);
not(notn14560,n14125);
and (s0n14560,notn14560,1'b0);
and (s1n14560,n14125,n14561);
wire s0n14561,s1n14561,notn14561;
or (n14561,s0n14561,s1n14561);
not(notn14561,n14563);
and (s0n14561,notn14561,n14556);
and (s1n14561,n14563,n14562);
and (n14563,n14564,n33);
and (n14564,n14131,n585);
and (n14565,n14566,n14385);
wire s0n14566,s1n14566,notn14566;
or (n14566,s0n14566,s1n14566);
not(notn14566,n2799);
and (s0n14566,notn14566,1'b0);
and (s1n14566,n2799,n14567);
or (n14567,1'b0,n14568,n14571);
and (n14568,n14569,n13900);
wire s0n14569,s1n14569,notn14569;
or (n14569,s0n14569,s1n14569);
not(notn14569,n14570);
and (s0n14569,notn14569,n14202);
and (s1n14569,n14570,1'b0);
not (n14570,n14211);
and (n14571,n14572,n14131);
wire s0n14572,s1n14572,notn14572;
or (n14572,s0n14572,s1n14572);
not(notn14572,n14573);
and (s0n14572,notn14572,n14391);
and (s1n14572,n14573,1'b0);
not (n14573,n14368);
or (n14574,n14575,n14608,n14621,n14623,n14627,n14629,1'b0);
and (n14575,n14576,n14237);
wire s0n14576,s1n14576,notn14576;
or (n14576,s0n14576,s1n14576);
not(notn14576,n14455);
and (s0n14576,notn14576,1'b0);
and (s1n14576,n14455,n14577);
wire s0n14577,s1n14577,notn14577;
or (n14577,s0n14577,s1n14577);
not(notn14577,n42);
and (s0n14577,notn14577,1'b0);
and (s1n14577,n42,n14578);
wire s0n14578,s1n14578,notn14578;
or (n14578,s0n14578,s1n14578);
not(notn14578,n14422);
and (s0n14578,notn14578,n14579);
and (s1n14578,n14422,n14589);
wire s0n14579,s1n14579,notn14579;
or (n14579,s0n14579,s1n14579);
not(notn14579,n14362);
and (s0n14579,notn14579,1'b0);
and (s1n14579,n14362,n14580);
or (n14580,1'b0,n14581,n14583,n14585,n14587);
and (n14581,n14582,n14352);
and (n14583,n14584,n14355);
and (n14585,n14586,n14358);
and (n14587,n14588,n14361);
or (n14589,1'b0,n14590,n14593,n14596,n14602);
and (n14590,n14591,n14387);
wire s0n14591,s1n14591,notn14591;
or (n14591,s0n14591,s1n14591);
not(notn14591,n14374);
and (s0n14591,notn14591,1'b0);
and (s1n14591,n14374,n14592);
and (n14593,n14594,n14393);
wire s0n14594,s1n14594,notn14594;
or (n14594,s0n14594,s1n14594);
not(notn14594,n14374);
and (s0n14594,notn14594,1'b0);
and (s1n14594,n14374,n14595);
and (n14596,n14597,n14412);
wire s0n14597,s1n14597,notn14597;
or (n14597,s0n14597,s1n14597);
not(notn14597,n42);
and (s0n14597,notn14597,1'b0);
and (s1n14597,n42,n14598);
wire s0n14598,s1n14598,notn14598;
or (n14598,s0n14598,s1n14598);
not(notn14598,n14375);
and (s0n14598,notn14598,n14599);
and (s1n14598,n14375,n14601);
wire s0n14599,s1n14599,notn14599;
or (n14599,s0n14599,s1n14599);
not(notn14599,n14409);
and (s0n14599,notn14599,n14600);
and (s1n14599,n14409,n14586);
wire s0n14600,s1n14600,notn14600;
or (n14600,s0n14600,s1n14600);
not(notn14600,n14401);
and (s0n14600,notn14600,1'b0);
and (s1n14600,n14401,n14582);
and (n14602,n14603,n14421);
wire s0n14603,s1n14603,notn14603;
or (n14603,s0n14603,s1n14603);
not(notn14603,n42);
and (s0n14603,notn14603,1'b0);
and (s1n14603,n42,n14604);
wire s0n14604,s1n14604,notn14604;
or (n14604,s0n14604,s1n14604);
not(notn14604,n14375);
and (s0n14604,notn14604,n14605);
and (s1n14604,n14375,n14607);
wire s0n14605,s1n14605,notn14605;
or (n14605,s0n14605,s1n14605);
not(notn14605,n14409);
and (s0n14605,notn14605,n14606);
and (s1n14605,n14409,n14588);
wire s0n14606,s1n14606,notn14606;
or (n14606,s0n14606,s1n14606);
not(notn14606,n14401);
and (s0n14606,notn14606,1'b0);
and (s1n14606,n14401,n14584);
and (n14608,n14609,n14137);
or (n14609,1'b0,n14610,n14620);
and (n14610,n14611,n14235);
wire s0n14611,s1n14611,notn14611;
or (n14611,s0n14611,s1n14611);
not(notn14611,n14227);
and (s0n14611,notn14611,1'b0);
and (s1n14611,n14227,n14612);
or (n14612,1'b0,n14140,n14613,n14614,n14615,n14616,n14619);
and (n14613,n14307,n14199);
and (n14614,n14309,n2781);
and (n14615,n14302,n14205);
and (n14616,n14617,n2789);
wire s0n14617,s1n14617,notn14617;
or (n14617,s0n14617,s1n14617);
not(notn14617,n14210);
and (s0n14617,notn14617,n14170);
and (s1n14617,n14210,n14618);
and (n14619,n14618,n14225);
and (n14620,n14280,n14455);
and (n14621,n14622,n14111);
wire s0n14622,s1n14622,notn14622;
or (n14622,s0n14622,s1n14622);
not(notn14622,n14455);
and (s0n14622,notn14622,1'b0);
and (s1n14622,n14455,n14456);
not (n14623,n14624);
nand (n14624,n14625,n14346);
not (n14625,n14626);
nand (n14626,n14108,n14131);
and (n14627,n14628,n13950);
wire s0n14628,s1n14628,notn14628;
or (n14628,s0n14628,s1n14628);
not(notn14628,n14131);
and (s0n14628,notn14628,1'b0);
and (s1n14628,n14131,n14456);
and (n14629,n14630,n14239);
wire s0n14630,s1n14630,notn14630;
or (n14630,s0n14630,s1n14630);
not(notn14630,n14131);
and (s0n14630,notn14630,1'b0);
and (s1n14630,n14131,n14611);
and (n14631,n14632,n591);
and (n14632,n14000,n42);
or (n14633,n14634,n14970,n17027);
and (n14634,n14635,n14898);
wire s0n14635,s1n14635,notn14635;
or (n14635,s0n14635,s1n14635);
not(notn14635,n14631);
and (s0n14635,notn14635,n14636);
and (s1n14635,n14631,n14763);
wire s0n14636,s1n14636,notn14636;
or (n14636,s0n14636,s1n14636);
not(notn14636,n14271);
and (s0n14636,notn14636,n14637);
and (s1n14636,n14271,n14751);
wire s0n14637,s1n14637,notn14637;
or (n14637,s0n14637,s1n14637);
not(notn14637,n14279);
and (s0n14637,notn14637,1'b0);
and (s1n14637,n14279,n14638);
or (n14638,1'b0,n14639,n14652,n14719);
and (n14639,n14640,n14120);
wire s0n14640,s1n14640,notn14640;
or (n14640,s0n14640,s1n14640);
not(notn14640,n14125);
and (s0n14640,notn14640,1'b0);
and (s1n14640,n14125,n14641);
wire s0n14641,s1n14641,notn14641;
or (n14641,s0n14641,s1n14641);
not(notn14641,n14317);
and (s0n14641,notn14641,n14642);
and (s1n14641,n14317,n14643);
wire s0n14643,s1n14643,notn14643;
or (n14643,s0n14643,s1n14643);
not(notn14643,n14326);
and (s0n14643,notn14643,n14644);
and (s1n14643,n14326,n14646);
wire s0n14644,s1n14644,notn14644;
or (n14644,s0n14644,s1n14644);
not(notn14644,n14315);
and (s0n14644,notn14644,1'b0);
and (s1n14644,n14315,n14645);
or (n14646,1'b0,n14647,n14649,n14651);
and (n14647,n14648,n14321);
and (n14649,n14650,n14324);
and (n14651,n14645,n14184);
and (n14652,n14653,n14718);
or (n14653,1'b0,n14654,n14670,n14686,n14702);
and (n14654,n14655,n13889);
wire s0n14655,s1n14655,notn14655;
or (n14655,s0n14655,s1n14655);
not(notn14655,n42);
and (s0n14655,notn14655,1'b0);
and (s1n14655,n42,n14656);
wire s0n14656,s1n14656,notn14656;
or (n14656,s0n14656,s1n14656);
not(notn14656,n14187);
and (s0n14656,notn14656,n14657);
and (s1n14656,n14187,n14663);
wire s0n14657,s1n14657,notn14657;
or (n14657,s0n14657,s1n14657);
not(notn14657,n14163);
and (s0n14657,notn14657,1'b0);
and (s1n14657,n14163,n14658);
or (n14658,1'b0,n14659,n14661);
and (n14659,n14660,n14147);
and (n14661,n14662,n14156);
or (n14663,1'b0,n14664,n14666,n14668,n14669);
and (n14664,n14665,n14171);
and (n14666,n14667,n14176);
and (n14668,n14660,n14180);
and (n14669,n14662,n14184);
and (n14670,n14671,n13897);
wire s0n14671,s1n14671,notn14671;
or (n14671,s0n14671,s1n14671);
not(notn14671,n42);
and (s0n14671,notn14671,1'b0);
and (s1n14671,n42,n14672);
wire s0n14672,s1n14672,notn14672;
or (n14672,s0n14672,s1n14672);
not(notn14672,n14187);
and (s0n14672,notn14672,n14673);
and (s1n14672,n14187,n14679);
wire s0n14673,s1n14673,notn14673;
or (n14673,s0n14673,s1n14673);
not(notn14673,n14163);
and (s0n14673,notn14673,1'b0);
and (s1n14673,n14163,n14674);
or (n14674,1'b0,n14675,n14677);
and (n14675,n14676,n14147);
and (n14677,n14678,n14156);
or (n14679,1'b0,n14680,n14682,n14684,n14685);
and (n14680,n14681,n14171);
and (n14682,n14683,n14176);
and (n14684,n14676,n14180);
and (n14685,n14678,n14184);
and (n14686,n14687,n13900);
wire s0n14687,s1n14687,notn14687;
or (n14687,s0n14687,s1n14687);
not(notn14687,n42);
and (s0n14687,notn14687,1'b0);
and (s1n14687,n42,n14688);
wire s0n14688,s1n14688,notn14688;
or (n14688,s0n14688,s1n14688);
not(notn14688,n14187);
and (s0n14688,notn14688,n14689);
and (s1n14688,n14187,n14695);
wire s0n14689,s1n14689,notn14689;
or (n14689,s0n14689,s1n14689);
not(notn14689,n14163);
and (s0n14689,notn14689,1'b0);
and (s1n14689,n14163,n14690);
or (n14690,1'b0,n14691,n14693);
and (n14691,n14692,n14147);
and (n14693,n14694,n14156);
or (n14695,1'b0,n14696,n14698,n14700,n14701);
and (n14696,n14697,n14171);
and (n14698,n14699,n14176);
and (n14700,n14692,n14180);
and (n14701,n14694,n14184);
and (n14702,n14703,n14131);
wire s0n14703,s1n14703,notn14703;
or (n14703,s0n14703,s1n14703);
not(notn14703,n42);
and (s0n14703,notn14703,1'b0);
and (s1n14703,n42,n14704);
wire s0n14704,s1n14704,notn14704;
or (n14704,s0n14704,s1n14704);
not(notn14704,n14187);
and (s0n14704,notn14704,n14705);
and (s1n14704,n14187,n14711);
wire s0n14705,s1n14705,notn14705;
or (n14705,s0n14705,s1n14705);
not(notn14705,n14163);
and (s0n14705,notn14705,1'b0);
and (s1n14705,n14163,n14706);
or (n14706,1'b0,n14707,n14709);
and (n14707,n14708,n14147);
and (n14709,n14710,n14156);
or (n14711,1'b0,n14712,n14714,n14716,n14717);
and (n14712,n14713,n14171);
and (n14714,n14715,n14176);
and (n14716,n14708,n14180);
and (n14717,n14710,n14184);
nor (n14718,n14121,n14277);
and (n14719,n14720,n14365);
wire s0n14720,s1n14720,notn14720;
or (n14720,s0n14720,s1n14720);
not(notn14720,n42);
and (s0n14720,notn14720,1'b0);
and (s1n14720,n42,n14721);
wire s0n14721,s1n14721,notn14721;
or (n14721,s0n14721,s1n14721);
not(notn14721,n14422);
and (s0n14721,notn14721,n14722);
and (s1n14721,n14422,n14732);
wire s0n14722,s1n14722,notn14722;
or (n14722,s0n14722,s1n14722);
not(notn14722,n14362);
and (s0n14722,notn14722,1'b0);
and (s1n14722,n14362,n14723);
or (n14723,1'b0,n14724,n14726,n14728,n14730);
and (n14724,n14725,n14352);
and (n14726,n14727,n14355);
and (n14728,n14729,n14358);
and (n14730,n14731,n14361);
or (n14732,1'b0,n14733,n14736,n14739,n14745);
and (n14733,n14734,n14387);
wire s0n14734,s1n14734,notn14734;
or (n14734,s0n14734,s1n14734);
not(notn14734,n14374);
and (s0n14734,notn14734,1'b0);
and (s1n14734,n14374,n14735);
and (n14736,n14737,n14393);
wire s0n14737,s1n14737,notn14737;
or (n14737,s0n14737,s1n14737);
not(notn14737,n14374);
and (s0n14737,notn14737,1'b0);
and (s1n14737,n14374,n14738);
and (n14739,n14740,n14412);
wire s0n14740,s1n14740,notn14740;
or (n14740,s0n14740,s1n14740);
not(notn14740,n42);
and (s0n14740,notn14740,1'b0);
and (s1n14740,n42,n14741);
wire s0n14741,s1n14741,notn14741;
or (n14741,s0n14741,s1n14741);
not(notn14741,n14375);
and (s0n14741,notn14741,n14742);
and (s1n14741,n14375,n14744);
wire s0n14742,s1n14742,notn14742;
or (n14742,s0n14742,s1n14742);
not(notn14742,n14409);
and (s0n14742,notn14742,n14743);
and (s1n14742,n14409,n14729);
wire s0n14743,s1n14743,notn14743;
or (n14743,s0n14743,s1n14743);
not(notn14743,n14401);
and (s0n14743,notn14743,1'b0);
and (s1n14743,n14401,n14725);
and (n14745,n14746,n14421);
wire s0n14746,s1n14746,notn14746;
or (n14746,s0n14746,s1n14746);
not(notn14746,n42);
and (s0n14746,notn14746,1'b0);
and (s1n14746,n42,n14747);
wire s0n14747,s1n14747,notn14747;
or (n14747,s0n14747,s1n14747);
not(notn14747,n14375);
and (s0n14747,notn14747,n14748);
and (s1n14747,n14375,n14750);
wire s0n14748,s1n14748,notn14748;
or (n14748,s0n14748,s1n14748);
not(notn14748,n14409);
and (s0n14748,notn14748,n14749);
and (s1n14748,n14409,n14731);
wire s0n14749,s1n14749,notn14749;
or (n14749,s0n14749,s1n14749);
not(notn14749,n14401);
and (s0n14749,notn14749,1'b0);
and (s1n14749,n14401,n14727);
or (n14751,n14752,n14753,n14761,n14762);
and (n14752,n14640,n13907);
and (n14753,n14754,n14385);
wire s0n14754,s1n14754,notn14754;
or (n14754,s0n14754,s1n14754);
not(notn14754,n2799);
and (s0n14754,notn14754,1'b0);
and (s1n14754,n2799,n14755);
or (n14755,1'b0,n14756,n14757);
and (n14756,n14642,n13900);
and (n14757,n14758,n14131);
wire s0n14758,s1n14758,notn14758;
or (n14758,s0n14758,s1n14758);
not(notn14758,n14573);
and (s0n14758,notn14758,n14759);
and (s1n14758,n14573,1'b0);
wire s0n14759,s1n14759,notn14759;
or (n14759,s0n14759,s1n14759);
not(notn14759,n14374);
and (s0n14759,notn14759,1'b0);
and (s1n14759,n14374,n14760);
and (n14761,n14720,n14381);
and (n14762,n14653,n14192);
or (n14763,1'b0,n14764,n14769,n14784,n14852,n14882,n14888,n14896,n14897);
and (n14764,n14765,n14237);
or (n14765,1'b0,n14766,n14768);
and (n14766,n14767,n14235);
wire s0n14768,s1n14768,notn14768;
or (n14768,s0n14768,s1n14768);
not(notn14768,n14455);
and (s0n14768,notn14768,1'b0);
and (s1n14768,n14455,n14720);
and (n14769,n14770,n14137);
or (n14770,1'b0,n14771,n14782,n14783);
and (n14771,n14772,n13889);
wire s0n14772,s1n14772,notn14772;
or (n14772,s0n14772,s1n14772);
not(notn14772,n14227);
and (s0n14772,notn14772,1'b0);
and (s1n14772,n14227,n14773);
or (n14773,1'b0,n14774,n14775,n14776,n14777,n14778,n14781);
and (n14774,n14655,n14193);
and (n14775,n14697,n14199);
and (n14776,n14699,n2781);
and (n14777,n14692,n14205);
and (n14778,n14779,n2789);
wire s0n14779,s1n14779,notn14779;
or (n14779,s0n14779,s1n14779);
not(notn14779,n14210);
and (s0n14779,notn14779,n14665);
and (s1n14779,n14210,n14780);
and (n14781,n14780,n14225);
and (n14782,n14655,n14243);
and (n14783,n14687,n14131);
and (n14784,n14785,n14111);
or (n14785,1'b0,n14786,n14788,n14790,n14820);
and (n14786,n14787,n13889);
and (n14788,n14789,n13897);
and (n14790,n14791,n13900);
wire s0n14791,s1n14791,notn14791;
or (n14791,s0n14791,s1n14791);
not(notn14791,n42);
and (s0n14791,notn14791,1'b0);
and (s1n14791,n42,n14792);
wire s0n14792,s1n14792,notn14792;
or (n14792,s0n14792,s1n14792);
not(notn14792,n14422);
and (s0n14792,notn14792,n14793);
and (s1n14792,n14422,n14803);
wire s0n14793,s1n14793,notn14793;
or (n14793,s0n14793,s1n14793);
not(notn14793,n14362);
and (s0n14793,notn14793,1'b0);
and (s1n14793,n14362,n14794);
or (n14794,1'b0,n14795,n14797,n14799,n14801);
and (n14795,n14796,n14352);
and (n14797,n14798,n14355);
and (n14799,n14800,n14358);
and (n14801,n14802,n14361);
or (n14803,1'b0,n14804,n14807,n14808,n14814);
and (n14804,n14805,n14387);
wire s0n14805,s1n14805,notn14805;
or (n14805,s0n14805,s1n14805);
not(notn14805,n14374);
and (s0n14805,notn14805,1'b0);
and (s1n14805,n14374,n14806);
and (n14807,n14759,n14393);
and (n14808,n14809,n14412);
wire s0n14809,s1n14809,notn14809;
or (n14809,s0n14809,s1n14809);
not(notn14809,n42);
and (s0n14809,notn14809,1'b0);
and (s1n14809,n42,n14810);
wire s0n14810,s1n14810,notn14810;
or (n14810,s0n14810,s1n14810);
not(notn14810,n14375);
and (s0n14810,notn14810,n14811);
and (s1n14810,n14375,n14813);
wire s0n14811,s1n14811,notn14811;
or (n14811,s0n14811,s1n14811);
not(notn14811,n14409);
and (s0n14811,notn14811,n14812);
and (s1n14811,n14409,n14800);
wire s0n14812,s1n14812,notn14812;
or (n14812,s0n14812,s1n14812);
not(notn14812,n14401);
and (s0n14812,notn14812,1'b0);
and (s1n14812,n14401,n14796);
and (n14814,n14815,n14421);
wire s0n14815,s1n14815,notn14815;
or (n14815,s0n14815,s1n14815);
not(notn14815,n42);
and (s0n14815,notn14815,1'b0);
and (s1n14815,n42,n14816);
wire s0n14816,s1n14816,notn14816;
or (n14816,s0n14816,s1n14816);
not(notn14816,n14375);
and (s0n14816,notn14816,n14817);
and (s1n14816,n14375,n14819);
wire s0n14817,s1n14817,notn14817;
or (n14817,s0n14817,s1n14817);
not(notn14817,n14409);
and (s0n14817,notn14817,n14818);
and (s1n14817,n14409,n14802);
wire s0n14818,s1n14818,notn14818;
or (n14818,s0n14818,s1n14818);
not(notn14818,n14401);
and (s0n14818,notn14818,1'b0);
and (s1n14818,n14401,n14798);
wire s0n14820,s1n14820,notn14820;
or (n14820,s0n14820,s1n14820);
not(notn14820,n14131);
and (s0n14820,notn14820,1'b0);
and (s1n14820,n14131,n14821);
wire s0n14821,s1n14821,notn14821;
or (n14821,s0n14821,s1n14821);
not(notn14821,n42);
and (s0n14821,notn14821,1'b0);
and (s1n14821,n42,n14822);
wire s0n14822,s1n14822,notn14822;
or (n14822,s0n14822,s1n14822);
not(notn14822,n14422);
and (s0n14822,notn14822,n14823);
and (s1n14822,n14422,n14833);
wire s0n14823,s1n14823,notn14823;
or (n14823,s0n14823,s1n14823);
not(notn14823,n14362);
and (s0n14823,notn14823,1'b0);
and (s1n14823,n14362,n14824);
or (n14824,1'b0,n14825,n14827,n14829,n14831);
and (n14825,n14826,n14352);
and (n14827,n14828,n14355);
and (n14829,n14830,n14358);
and (n14831,n14832,n14361);
or (n14833,1'b0,n14834,n14837,n14840,n14846);
and (n14834,n14835,n14387);
wire s0n14835,s1n14835,notn14835;
or (n14835,s0n14835,s1n14835);
not(notn14835,n14374);
and (s0n14835,notn14835,1'b0);
and (s1n14835,n14374,n14836);
and (n14837,n14838,n14393);
wire s0n14838,s1n14838,notn14838;
or (n14838,s0n14838,s1n14838);
not(notn14838,n14374);
and (s0n14838,notn14838,1'b0);
and (s1n14838,n14374,n14839);
and (n14840,n14841,n14412);
wire s0n14841,s1n14841,notn14841;
or (n14841,s0n14841,s1n14841);
not(notn14841,n42);
and (s0n14841,notn14841,1'b0);
and (s1n14841,n42,n14842);
wire s0n14842,s1n14842,notn14842;
or (n14842,s0n14842,s1n14842);
not(notn14842,n14375);
and (s0n14842,notn14842,n14843);
and (s1n14842,n14375,n14845);
wire s0n14843,s1n14843,notn14843;
or (n14843,s0n14843,s1n14843);
not(notn14843,n14409);
and (s0n14843,notn14843,n14844);
and (s1n14843,n14409,n14830);
wire s0n14844,s1n14844,notn14844;
or (n14844,s0n14844,s1n14844);
not(notn14844,n14401);
and (s0n14844,notn14844,1'b0);
and (s1n14844,n14401,n14826);
and (n14846,n14847,n14421);
wire s0n14847,s1n14847,notn14847;
or (n14847,s0n14847,s1n14847);
not(notn14847,n42);
and (s0n14847,notn14847,1'b0);
and (s1n14847,n42,n14848);
wire s0n14848,s1n14848,notn14848;
or (n14848,s0n14848,s1n14848);
not(notn14848,n14375);
and (s0n14848,notn14848,n14849);
and (s1n14848,n14375,n14851);
wire s0n14849,s1n14849,notn14849;
or (n14849,s0n14849,s1n14849);
not(notn14849,n14409);
and (s0n14849,notn14849,n14850);
and (s1n14849,n14409,n14832);
wire s0n14850,s1n14850,notn14850;
or (n14850,s0n14850,s1n14850);
not(notn14850,n14401);
and (s0n14850,notn14850,1'b0);
and (s1n14850,n14401,n14828);
and (n14852,n14853,n14108);
or (n14853,1'b0,n14854,n14856,n14858,n14860);
and (n14854,n14855,n13889);
and (n14856,n14857,n13897);
and (n14858,n14859,n13900);
and (n14860,n14861,n14131);
wire s0n14861,s1n14861,notn14861;
or (n14861,s0n14861,s1n14861);
not(notn14861,n14123);
and (s0n14861,notn14861,1'b0);
and (s1n14861,n14123,n14862);
wire s0n14862,s1n14862,notn14862;
or (n14862,s0n14862,s1n14862);
not(notn14862,n555);
and (s0n14862,notn14862,n14863);
and (s1n14862,n555,n14878);
wire s0n14863,s1n14863,notn14863;
or (n14863,s0n14863,s1n14863);
not(notn14863,n13948);
and (s0n14863,notn14863,n14864);
and (s1n14863,n13948,n14866);
wire s0n14864,s1n14864,notn14864;
or (n14864,s0n14864,s1n14864);
not(notn14864,n13907);
and (s0n14864,notn14864,1'b0);
and (s1n14864,n13907,n14865);
or (n14866,n14867,n14869,n14871,n14873,n14875,n14877);
and (n14867,n14868,n13913);
and (n14869,n14870,n13920);
and (n14871,n14872,n13923);
and (n14873,n14874,n13928);
and (n14875,n14876,n13935);
and (n14877,n14865,n13941);
wire s0n14878,s1n14878,notn14878;
or (n14878,s0n14878,s1n14878);
not(notn14878,n14119);
and (s0n14878,notn14878,1'b0);
and (s1n14878,n14119,n14879);
wire s0n14879,s1n14879,notn14879;
or (n14879,s0n14879,s1n14879);
not(notn14879,n14116);
and (s0n14879,notn14879,n14880);
and (s1n14879,n14116,n14881);
and (n14882,n14883,n13950);
or (n14883,1'b0,n14884,n14885,n14886,n14887);
and (n14884,n14857,n13889);
and (n14885,n14859,n13897);
and (n14886,n14789,n13900);
wire s0n14887,s1n14887,notn14887;
or (n14887,s0n14887,s1n14887);
not(notn14887,n14131);
and (s0n14887,notn14887,1'b0);
and (s1n14887,n14131,n14791);
and (n14888,n14889,n14239);
or (n14889,1'b0,n14890,n14892,n14894,n14895);
and (n14890,n14891,n13889);
and (n14892,n14893,n13897);
and (n14894,n14767,n13900);
and (n14895,n14671,n14131);
and (n14896,n14720,n14448);
and (n14897,n14653,n14266);
wire s0n14898,s1n14898,notn14898;
or (n14898,s0n14898,s1n14898);
not(notn14898,n14631);
and (s0n14898,notn14898,n14899);
and (s1n14898,n14631,n14917);
wire s0n14899,s1n14899,notn14899;
or (n14899,s0n14899,s1n14899);
not(notn14899,n14271);
and (s0n14899,notn14899,n14900);
and (s1n14899,n14271,n14905);
wire s0n14900,s1n14900,notn14900;
or (n14900,s0n14900,s1n14900);
not(notn14900,n14279);
and (s0n14900,notn14900,1'b0);
and (s1n14900,n14279,n14901);
and (n14901,n14902,n14120);
wire s0n14902,s1n14902,notn14902;
or (n14902,s0n14902,s1n14902);
not(notn14902,n14125);
and (s0n14902,notn14902,1'b0);
and (s1n14902,n14125,n14903);
wire s0n14903,s1n14903,notn14903;
or (n14903,s0n14903,s1n14903);
not(notn14903,n14317);
and (s0n14903,notn14903,n14904);
and (s1n14903,n14317,n14562);
or (n14905,n14906,n14910,1'b0);
and (n14906,n14907,n13907);
wire s0n14907,s1n14907,notn14907;
or (n14907,s0n14907,s1n14907);
not(notn14907,n14125);
and (s0n14907,notn14907,1'b0);
and (s1n14907,n14125,n14908);
wire s0n14908,s1n14908,notn14908;
or (n14908,s0n14908,s1n14908);
not(notn14908,n14563);
and (s0n14908,notn14908,n14904);
and (s1n14908,n14563,n14909);
and (n14910,n14911,n14385);
wire s0n14911,s1n14911,notn14911;
or (n14911,s0n14911,s1n14911);
not(notn14911,n2799);
and (s0n14911,notn14911,1'b0);
and (s1n14911,n2799,n14912);
or (n14912,1'b0,n14913,n14915);
and (n14913,n14914,n13900);
wire s0n14914,s1n14914,notn14914;
or (n14914,s0n14914,s1n14914);
not(notn14914,n14570);
and (s0n14914,notn14914,n14699);
and (s1n14914,n14570,1'b0);
and (n14915,n14916,n14131);
wire s0n14916,s1n14916,notn14916;
or (n14916,s0n14916,s1n14916);
not(notn14916,n14573);
and (s0n14916,notn14916,n14838);
and (s1n14916,n14573,1'b0);
or (n14917,n14918,n14951,n14964,n14965,n14966,n14968,1'b0);
and (n14918,n14919,n14237);
wire s0n14919,s1n14919,notn14919;
or (n14919,s0n14919,s1n14919);
not(notn14919,n14455);
and (s0n14919,notn14919,1'b0);
and (s1n14919,n14455,n14920);
wire s0n14920,s1n14920,notn14920;
or (n14920,s0n14920,s1n14920);
not(notn14920,n42);
and (s0n14920,notn14920,1'b0);
and (s1n14920,n42,n14921);
wire s0n14921,s1n14921,notn14921;
or (n14921,s0n14921,s1n14921);
not(notn14921,n14422);
and (s0n14921,notn14921,n14922);
and (s1n14921,n14422,n14932);
wire s0n14922,s1n14922,notn14922;
or (n14922,s0n14922,s1n14922);
not(notn14922,n14362);
and (s0n14922,notn14922,1'b0);
and (s1n14922,n14362,n14923);
or (n14923,1'b0,n14924,n14926,n14928,n14930);
and (n14924,n14925,n14352);
and (n14926,n14927,n14355);
and (n14928,n14929,n14358);
and (n14930,n14931,n14361);
or (n14932,1'b0,n14933,n14936,n14939,n14945);
and (n14933,n14934,n14387);
wire s0n14934,s1n14934,notn14934;
or (n14934,s0n14934,s1n14934);
not(notn14934,n14374);
and (s0n14934,notn14934,1'b0);
and (s1n14934,n14374,n14935);
and (n14936,n14937,n14393);
wire s0n14937,s1n14937,notn14937;
or (n14937,s0n14937,s1n14937);
not(notn14937,n14374);
and (s0n14937,notn14937,1'b0);
and (s1n14937,n14374,n14938);
and (n14939,n14940,n14412);
wire s0n14940,s1n14940,notn14940;
or (n14940,s0n14940,s1n14940);
not(notn14940,n42);
and (s0n14940,notn14940,1'b0);
and (s1n14940,n42,n14941);
wire s0n14941,s1n14941,notn14941;
or (n14941,s0n14941,s1n14941);
not(notn14941,n14375);
and (s0n14941,notn14941,n14942);
and (s1n14941,n14375,n14944);
wire s0n14942,s1n14942,notn14942;
or (n14942,s0n14942,s1n14942);
not(notn14942,n14409);
and (s0n14942,notn14942,n14943);
and (s1n14942,n14409,n14929);
wire s0n14943,s1n14943,notn14943;
or (n14943,s0n14943,s1n14943);
not(notn14943,n14401);
and (s0n14943,notn14943,1'b0);
and (s1n14943,n14401,n14925);
and (n14945,n14946,n14421);
wire s0n14946,s1n14946,notn14946;
or (n14946,s0n14946,s1n14946);
not(notn14946,n42);
and (s0n14946,notn14946,1'b0);
and (s1n14946,n42,n14947);
wire s0n14947,s1n14947,notn14947;
or (n14947,s0n14947,s1n14947);
not(notn14947,n14375);
and (s0n14947,notn14947,n14948);
and (s1n14947,n14375,n14950);
wire s0n14948,s1n14948,notn14948;
or (n14948,s0n14948,s1n14948);
not(notn14948,n14409);
and (s0n14948,notn14948,n14949);
and (s1n14948,n14409,n14931);
wire s0n14949,s1n14949,notn14949;
or (n14949,s0n14949,s1n14949);
not(notn14949,n14401);
and (s0n14949,notn14949,1'b0);
and (s1n14949,n14401,n14927);
and (n14951,n14952,n14137);
or (n14952,1'b0,n14953,n14963);
and (n14953,n14954,n14235);
wire s0n14954,s1n14954,notn14954;
or (n14954,s0n14954,s1n14954);
not(notn14954,n14227);
and (s0n14954,notn14954,1'b0);
and (s1n14954,n14227,n14955);
or (n14955,1'b0,n14774,n14956,n14957,n14958,n14959,n14962);
and (n14956,n14713,n14199);
and (n14957,n14715,n2781);
and (n14958,n14708,n14205);
and (n14959,n14960,n2789);
wire s0n14960,s1n14960,notn14960;
or (n14960,s0n14960,s1n14960);
not(notn14960,n14210);
and (s0n14960,notn14960,n14665);
and (s1n14960,n14210,n14961);
and (n14962,n14961,n14225);
and (n14963,n14671,n14455);
and (n14964,n14768,n14111);
and (n14965,n14820,n14108);
and (n14966,n14967,n13950);
wire s0n14967,s1n14967,notn14967;
or (n14967,s0n14967,s1n14967);
not(notn14967,n14131);
and (s0n14967,notn14967,1'b0);
and (s1n14967,n14131,n14720);
and (n14968,n14969,n14239);
wire s0n14969,s1n14969,notn14969;
or (n14969,s0n14969,s1n14969);
not(notn14969,n14131);
and (s0n14969,notn14969,1'b0);
and (s1n14969,n14131,n14954);
and (n14970,n14898,n14971);
or (n14971,n14972,n15296,n17026);
and (n14972,n14973,n15222);
nand (n14973,n14974,n15105,n15189);
nor (n14974,n14975,n15005);
and (n14975,n14976,n14108);
or (n14976,1'b0,n14977,n14979,n14981,n14983);
and (n14977,n14978,n13889);
and (n14979,n14980,n13897);
and (n14981,n14982,n13900);
and (n14983,n14984,n14131);
wire s0n14984,s1n14984,notn14984;
or (n14984,s0n14984,s1n14984);
not(notn14984,n14123);
and (s0n14984,notn14984,1'b0);
and (s1n14984,n14123,n14985);
wire s0n14985,s1n14985,notn14985;
or (n14985,s0n14985,s1n14985);
not(notn14985,n555);
and (s0n14985,notn14985,n14986);
and (s1n14985,n555,n15001);
wire s0n14986,s1n14986,notn14986;
or (n14986,s0n14986,s1n14986);
not(notn14986,n13948);
and (s0n14986,notn14986,n14987);
and (s1n14986,n13948,n14989);
wire s0n14987,s1n14987,notn14987;
or (n14987,s0n14987,s1n14987);
not(notn14987,n13907);
and (s0n14987,notn14987,1'b0);
and (s1n14987,n13907,n14988);
or (n14989,n14990,n14992,n14994,n14996,n14998,n15000);
and (n14990,n14991,n13913);
and (n14992,n14993,n13920);
and (n14994,n14995,n13923);
and (n14996,n14997,n13928);
and (n14998,n14999,n13935);
and (n15000,n14988,n13941);
wire s0n15001,s1n15001,notn15001;
or (n15001,s0n15001,s1n15001);
not(notn15001,n14119);
and (s0n15001,notn15001,1'b0);
and (s1n15001,n14119,n15002);
wire s0n15002,s1n15002,notn15002;
or (n15002,s0n15002,s1n15002);
not(notn15002,n14116);
and (s0n15002,notn15002,n15003);
and (s1n15002,n14116,n15004);
nand (n15005,n15006,n15087,n15102);
not (n15006,n15007);
nand (n15007,n15008,n15054);
nor (n15008,n15009,n15038);
nand (n15009,n15010,n15028);
or (n15010,n15011,n15027);
not (n15011,n15012);
wire s0n15012,s1n15012,notn15012;
or (n15012,s0n15012,s1n15012);
not(notn15012,n42);
and (s0n15012,notn15012,1'b0);
and (s1n15012,n42,n15013);
wire s0n15013,s1n15013,notn15013;
or (n15013,s0n15013,s1n15013);
not(notn15013,n14187);
and (s0n15013,notn15013,n15014);
and (s1n15013,n14187,n15020);
wire s0n15014,s1n15014,notn15014;
or (n15014,s0n15014,s1n15014);
not(notn15014,n14163);
and (s0n15014,notn15014,1'b0);
and (s1n15014,n14163,n15015);
or (n15015,1'b0,n15016,n15018);
and (n15016,n15017,n14147);
and (n15018,n15019,n14156);
or (n15020,1'b0,n15021,n15023,n15025,n15026);
and (n15021,n15022,n14171);
and (n15023,n15024,n14176);
and (n15025,n15017,n14180);
and (n15026,n15019,n14184);
not (n15027,n14296);
not (n15028,n15029);
wire s0n15029,s1n15029,notn15029;
or (n15029,s0n15029,s1n15029);
not(notn15029,n14326);
and (s0n15029,notn15029,n15030);
and (s1n15029,n14326,n15032);
wire s0n15030,s1n15030,notn15030;
or (n15030,s0n15030,s1n15030);
not(notn15030,n14315);
and (s0n15030,notn15030,1'b0);
and (s1n15030,n14315,n15031);
or (n15032,1'b0,n15033,n15035,n15037);
and (n15033,n15034,n14321);
and (n15035,n15036,n14324);
and (n15037,n15031,n14184);
and (n15038,n14263,n15039);
wire s0n15039,s1n15039,notn15039;
or (n15039,s0n15039,s1n15039);
not(notn15039,n42);
and (s0n15039,notn15039,1'b0);
and (s1n15039,n42,n15040);
wire s0n15040,s1n15040,notn15040;
or (n15040,s0n15040,s1n15040);
not(notn15040,n14187);
and (s0n15040,notn15040,n15041);
and (s1n15040,n14187,n15047);
wire s0n15041,s1n15041,notn15041;
or (n15041,s0n15041,s1n15041);
not(notn15041,n14163);
and (s0n15041,notn15041,1'b0);
and (s1n15041,n14163,n15042);
or (n15042,1'b0,n15043,n15045);
and (n15043,n15044,n14147);
and (n15045,n15046,n14156);
or (n15047,1'b0,n15048,n15050,n15052,n15053);
and (n15048,n15049,n14171);
and (n15050,n15051,n14176);
and (n15052,n15044,n14180);
and (n15053,n15046,n14184);
nor (n15054,n15055,n15071);
and (n15055,n14331,n15056);
wire s0n15056,s1n15056,notn15056;
or (n15056,s0n15056,s1n15056);
not(notn15056,n42);
and (s0n15056,notn15056,1'b0);
and (s1n15056,n42,n15057);
wire s0n15057,s1n15057,notn15057;
or (n15057,s0n15057,s1n15057);
not(notn15057,n14187);
and (s0n15057,notn15057,n15058);
and (s1n15057,n14187,n15064);
wire s0n15058,s1n15058,notn15058;
or (n15058,s0n15058,s1n15058);
not(notn15058,n14163);
and (s0n15058,notn15058,1'b0);
and (s1n15058,n14163,n15059);
or (n15059,1'b0,n15060,n15062);
and (n15060,n15061,n14147);
and (n15062,n15063,n14156);
or (n15064,1'b0,n15065,n15067,n15069,n15070);
and (n15065,n15066,n14171);
and (n15067,n15068,n14176);
and (n15069,n15061,n14180);
and (n15070,n15063,n14184);
and (n15071,n14333,n15072);
wire s0n15072,s1n15072,notn15072;
or (n15072,s0n15072,s1n15072);
not(notn15072,n42);
and (s0n15072,notn15072,1'b0);
and (s1n15072,n42,n15073);
wire s0n15073,s1n15073,notn15073;
or (n15073,s0n15073,s1n15073);
not(notn15073,n14187);
and (s0n15073,notn15073,n15074);
and (s1n15073,n14187,n15080);
wire s0n15074,s1n15074,notn15074;
or (n15074,s0n15074,s1n15074);
not(notn15074,n14163);
and (s0n15074,notn15074,1'b0);
and (s1n15074,n14163,n15075);
or (n15075,1'b0,n15076,n15078);
and (n15076,n15077,n14147);
and (n15078,n15079,n14156);
or (n15080,1'b0,n15081,n15083,n15085,n15086);
and (n15081,n15082,n14171);
and (n15083,n15084,n14176);
and (n15085,n15077,n14180);
and (n15086,n15079,n14184);
nor (n15087,n15088,n15099,n15101);
and (n15088,n14135,n15089);
wire s0n15089,s1n15089,notn15089;
or (n15089,s0n15089,s1n15089);
not(notn15089,n14227);
and (s0n15089,notn15089,1'b0);
and (s1n15089,n14227,n15090);
or (n15090,1'b0,n15091,n15092,n15093,n15094,n15095,n15098);
and (n15091,n15056,n14193);
and (n15092,n15082,n14199);
and (n15093,n15084,n2781);
and (n15094,n15077,n14205);
and (n15095,n15096,n2789);
wire s0n15096,s1n15096,notn15096;
or (n15096,s0n15096,s1n15096);
not(notn15096,n14210);
and (s0n15096,notn15096,n15066);
and (s1n15096,n14210,n15097);
and (n15098,n15097,n14225);
and (n15099,n14232,n15100);
and (n15101,n14242,n15056);
not (n15102,n15103);
and (n15103,n15104,n14137);
and (n15104,n15072,n14131);
nor (n15105,n15106,n15108);
and (n15106,n14336,n15107);
nand (n15108,n15109,n15115,n15150,n15182);
nor (n15109,n15110,n15112,n15114);
and (n15110,n14438,n15111);
and (n15112,n14426,n15113);
and (n15114,n14430,n14982);
nor (n15115,n15116,n15118);
and (n15116,n14434,n15117);
and (n15118,n14345,n15119);
wire s0n15119,s1n15119,notn15119;
or (n15119,s0n15119,s1n15119);
not(notn15119,n42);
and (s0n15119,notn15119,1'b0);
and (s1n15119,n42,n15120);
wire s0n15120,s1n15120,notn15120;
or (n15120,s0n15120,s1n15120);
not(notn15120,n14422);
and (s0n15120,notn15120,n15121);
and (s1n15120,n14422,n15131);
wire s0n15121,s1n15121,notn15121;
or (n15121,s0n15121,s1n15121);
not(notn15121,n14362);
and (s0n15121,notn15121,1'b0);
and (s1n15121,n14362,n15122);
or (n15122,1'b0,n15123,n15125,n15127,n15129);
and (n15123,n15124,n14352);
and (n15125,n15126,n14355);
and (n15127,n15128,n14358);
and (n15129,n15130,n14361);
or (n15131,1'b0,n15132,n15135,n15138,n15144);
and (n15132,n15133,n14387);
wire s0n15133,s1n15133,notn15133;
or (n15133,s0n15133,s1n15133);
not(notn15133,n14374);
and (s0n15133,notn15133,1'b0);
and (s1n15133,n14374,n15134);
and (n15135,n15136,n14393);
wire s0n15136,s1n15136,notn15136;
or (n15136,s0n15136,s1n15136);
not(notn15136,n14374);
and (s0n15136,notn15136,1'b0);
and (s1n15136,n14374,n15137);
and (n15138,n15139,n14412);
wire s0n15139,s1n15139,notn15139;
or (n15139,s0n15139,s1n15139);
not(notn15139,n42);
and (s0n15139,notn15139,1'b0);
and (s1n15139,n42,n15140);
wire s0n15140,s1n15140,notn15140;
or (n15140,s0n15140,s1n15140);
not(notn15140,n14375);
and (s0n15140,notn15140,n15141);
and (s1n15140,n14375,n15143);
wire s0n15141,s1n15141,notn15141;
or (n15141,s0n15141,s1n15141);
not(notn15141,n14409);
and (s0n15141,notn15141,n15142);
and (s1n15141,n14409,n15128);
wire s0n15142,s1n15142,notn15142;
or (n15142,s0n15142,s1n15142);
not(notn15142,n14401);
and (s0n15142,notn15142,1'b0);
and (s1n15142,n14401,n15124);
and (n15144,n15145,n14421);
wire s0n15145,s1n15145,notn15145;
or (n15145,s0n15145,s1n15145);
not(notn15145,n42);
and (s0n15145,notn15145,1'b0);
and (s1n15145,n42,n15146);
wire s0n15146,s1n15146,notn15146;
or (n15146,s0n15146,s1n15146);
not(notn15146,n14375);
and (s0n15146,notn15146,n15147);
and (s1n15146,n14375,n15149);
wire s0n15147,s1n15147,notn15147;
or (n15147,s0n15147,s1n15147);
not(notn15147,n14409);
and (s0n15147,notn15147,n15148);
and (s1n15147,n14409,n15130);
wire s0n15148,s1n15148,notn15148;
or (n15148,s0n15148,s1n15148);
not(notn15148,n14401);
and (s0n15148,notn15148,1'b0);
and (s1n15148,n14401,n15126);
nand (n15150,n14443,n15151);
wire s0n15151,s1n15151,notn15151;
or (n15151,s0n15151,s1n15151);
not(notn15151,n42);
and (s0n15151,notn15151,1'b0);
and (s1n15151,n42,n15152);
wire s0n15152,s1n15152,notn15152;
or (n15152,s0n15152,s1n15152);
not(notn15152,n14422);
and (s0n15152,notn15152,n15153);
and (s1n15152,n14422,n15163);
wire s0n15153,s1n15153,notn15153;
or (n15153,s0n15153,s1n15153);
not(notn15153,n14362);
and (s0n15153,notn15153,1'b0);
and (s1n15153,n14362,n15154);
or (n15154,1'b0,n15155,n15157,n15159,n15161);
and (n15155,n15156,n14352);
and (n15157,n15158,n14355);
and (n15159,n15160,n14358);
and (n15161,n15162,n14361);
or (n15163,1'b0,n15164,n15167,n15170,n15176);
and (n15164,n15165,n14387);
wire s0n15165,s1n15165,notn15165;
or (n15165,s0n15165,s1n15165);
not(notn15165,n14374);
and (s0n15165,notn15165,1'b0);
and (s1n15165,n14374,n15166);
and (n15167,n15168,n14393);
wire s0n15168,s1n15168,notn15168;
or (n15168,s0n15168,s1n15168);
not(notn15168,n14374);
and (s0n15168,notn15168,1'b0);
and (s1n15168,n14374,n15169);
and (n15170,n15171,n14412);
wire s0n15171,s1n15171,notn15171;
or (n15171,s0n15171,s1n15171);
not(notn15171,n42);
and (s0n15171,notn15171,1'b0);
and (s1n15171,n42,n15172);
wire s0n15172,s1n15172,notn15172;
or (n15172,s0n15172,s1n15172);
not(notn15172,n14375);
and (s0n15172,notn15172,n15173);
and (s1n15172,n14375,n15175);
wire s0n15173,s1n15173,notn15173;
or (n15173,s0n15173,s1n15173);
not(notn15173,n14409);
and (s0n15173,notn15173,n15174);
and (s1n15173,n14409,n15160);
wire s0n15174,s1n15174,notn15174;
or (n15174,s0n15174,s1n15174);
not(notn15174,n14401);
and (s0n15174,notn15174,1'b0);
and (s1n15174,n14401,n15156);
and (n15176,n15177,n14421);
wire s0n15177,s1n15177,notn15177;
or (n15177,s0n15177,s1n15177);
not(notn15177,n42);
and (s0n15177,notn15177,1'b0);
and (s1n15177,n42,n15178);
wire s0n15178,s1n15178,notn15178;
or (n15178,s0n15178,s1n15178);
not(notn15178,n14375);
and (s0n15178,notn15178,n15179);
and (s1n15178,n14375,n15181);
wire s0n15179,s1n15179,notn15179;
or (n15179,s0n15179,s1n15179);
not(notn15179,n14409);
and (s0n15179,notn15179,n15180);
and (s1n15179,n14409,n15162);
wire s0n15180,s1n15180,notn15180;
or (n15180,s0n15180,s1n15180);
not(notn15180,n14401);
and (s0n15180,notn15180,1'b0);
and (s1n15180,n14401,n15158);
nor (n15182,n15183,n15184,n15186);
and (n15183,n14489,n14980);
and (n15184,n14493,n15185);
and (n15186,n15187,n14511);
wire s0n15187,s1n15187,notn15187;
or (n15187,s0n15187,s1n15187);
not(notn15187,n14374);
and (s0n15187,notn15187,1'b0);
and (s1n15187,n14374,n15188);
nor (n15189,n15190,n15220);
and (n15190,n14516,n15191);
wire s0n15191,s1n15191,notn15191;
or (n15191,s0n15191,s1n15191);
not(notn15191,n42);
and (s0n15191,notn15191,1'b0);
and (s1n15191,n42,n15192);
wire s0n15192,s1n15192,notn15192;
or (n15192,s0n15192,s1n15192);
not(notn15192,n14422);
and (s0n15192,notn15192,n15193);
and (s1n15192,n14422,n15203);
wire s0n15193,s1n15193,notn15193;
or (n15193,s0n15193,s1n15193);
not(notn15193,n14362);
and (s0n15193,notn15193,1'b0);
and (s1n15193,n14362,n15194);
or (n15194,1'b0,n15195,n15197,n15199,n15201);
and (n15195,n15196,n14352);
and (n15197,n15198,n14355);
and (n15199,n15200,n14358);
and (n15201,n15202,n14361);
or (n15203,1'b0,n15204,n15207,n15208,n15214);
and (n15204,n15205,n14387);
wire s0n15205,s1n15205,notn15205;
or (n15205,s0n15205,s1n15205);
not(notn15205,n14374);
and (s0n15205,notn15205,1'b0);
and (s1n15205,n14374,n15206);
and (n15207,n15187,n14393);
and (n15208,n15209,n14412);
wire s0n15209,s1n15209,notn15209;
or (n15209,s0n15209,s1n15209);
not(notn15209,n42);
and (s0n15209,notn15209,1'b0);
and (s1n15209,n42,n15210);
wire s0n15210,s1n15210,notn15210;
or (n15210,s0n15210,s1n15210);
not(notn15210,n14375);
and (s0n15210,notn15210,n15211);
and (s1n15210,n14375,n15213);
wire s0n15211,s1n15211,notn15211;
or (n15211,s0n15211,s1n15211);
not(notn15211,n14409);
and (s0n15211,notn15211,n15212);
and (s1n15211,n14409,n15200);
wire s0n15212,s1n15212,notn15212;
or (n15212,s0n15212,s1n15212);
not(notn15212,n14401);
and (s0n15212,notn15212,1'b0);
and (s1n15212,n14401,n15196);
and (n15214,n15215,n14421);
wire s0n15215,s1n15215,notn15215;
or (n15215,s0n15215,s1n15215);
not(notn15215,n42);
and (s0n15215,notn15215,1'b0);
and (s1n15215,n42,n15216);
wire s0n15216,s1n15216,notn15216;
or (n15216,s0n15216,s1n15216);
not(notn15216,n14375);
and (s0n15216,notn15216,n15217);
and (s1n15216,n14375,n15219);
wire s0n15217,s1n15217,notn15217;
or (n15217,s0n15217,s1n15217);
not(notn15217,n14409);
and (s0n15217,notn15217,n15218);
and (s1n15217,n14409,n15202);
wire s0n15218,s1n15218,notn15218;
or (n15218,s0n15218,s1n15218);
not(notn15218,n14401);
and (s0n15218,notn15218,1'b0);
and (s1n15218,n14401,n15198);
and (n15220,n15221,n14239);
and (n15221,n15039,n14131);
wire s0n15222,s1n15222,notn15222;
or (n15222,s0n15222,s1n15222);
not(notn15222,n14631);
and (s0n15222,notn15222,n15223);
and (s1n15222,n14631,n15241);
wire s0n15223,s1n15223,notn15223;
or (n15223,s0n15223,s1n15223);
not(notn15223,n14271);
and (s0n15223,notn15223,n15224);
and (s1n15223,n14271,n15229);
wire s0n15224,s1n15224,notn15224;
or (n15224,s0n15224,s1n15224);
not(notn15224,n14279);
and (s0n15224,notn15224,1'b0);
and (s1n15224,n14279,n15225);
and (n15225,n15226,n14120);
wire s0n15226,s1n15226,notn15226;
or (n15226,s0n15226,s1n15226);
not(notn15226,n14125);
and (s0n15226,notn15226,1'b0);
and (s1n15226,n14125,n15227);
wire s0n15227,s1n15227,notn15227;
or (n15227,s0n15227,s1n15227);
not(notn15227,n14317);
and (s0n15227,notn15227,n15228);
and (s1n15227,n14317,n14909);
or (n15229,n15230,n15234,1'b0);
and (n15230,n15231,n13907);
wire s0n15231,s1n15231,notn15231;
or (n15231,s0n15231,s1n15231);
not(notn15231,n14125);
and (s0n15231,notn15231,1'b0);
and (s1n15231,n14125,n15232);
wire s0n15232,s1n15232,notn15232;
or (n15232,s0n15232,s1n15232);
not(notn15232,n14563);
and (s0n15232,notn15232,n15228);
and (s1n15232,n14563,n15233);
and (n15234,n15235,n14385);
wire s0n15235,s1n15235,notn15235;
or (n15235,s0n15235,s1n15235);
not(notn15235,n2799);
and (s0n15235,notn15235,1'b0);
and (s1n15235,n2799,n15236);
or (n15236,1'b0,n15237,n15239);
and (n15237,n15238,n13900);
wire s0n15238,s1n15238,notn15238;
or (n15238,s0n15238,s1n15238);
not(notn15238,n14570);
and (s0n15238,notn15238,n15084);
and (s1n15238,n14570,1'b0);
and (n15239,n15240,n14131);
wire s0n15240,s1n15240,notn15240;
or (n15240,s0n15240,s1n15240);
not(notn15240,n14573);
and (s0n15240,notn15240,n15136);
and (s1n15240,n14573,1'b0);
or (n15241,n15242,n15275,n15288,n15290,n15292,n15294,1'b0);
and (n15242,n15243,n14237);
wire s0n15243,s1n15243,notn15243;
or (n15243,s0n15243,s1n15243);
not(notn15243,n14455);
and (s0n15243,notn15243,1'b0);
and (s1n15243,n14455,n15244);
wire s0n15244,s1n15244,notn15244;
or (n15244,s0n15244,s1n15244);
not(notn15244,n42);
and (s0n15244,notn15244,1'b0);
and (s1n15244,n42,n15245);
wire s0n15245,s1n15245,notn15245;
or (n15245,s0n15245,s1n15245);
not(notn15245,n14422);
and (s0n15245,notn15245,n15246);
and (s1n15245,n14422,n15256);
wire s0n15246,s1n15246,notn15246;
or (n15246,s0n15246,s1n15246);
not(notn15246,n14362);
and (s0n15246,notn15246,1'b0);
and (s1n15246,n14362,n15247);
or (n15247,1'b0,n15248,n15250,n15252,n15254);
and (n15248,n15249,n14352);
and (n15250,n15251,n14355);
and (n15252,n15253,n14358);
and (n15254,n15255,n14361);
or (n15256,1'b0,n15257,n15260,n15263,n15269);
and (n15257,n15258,n14387);
wire s0n15258,s1n15258,notn15258;
or (n15258,s0n15258,s1n15258);
not(notn15258,n14374);
and (s0n15258,notn15258,1'b0);
and (s1n15258,n14374,n15259);
and (n15260,n15261,n14393);
wire s0n15261,s1n15261,notn15261;
or (n15261,s0n15261,s1n15261);
not(notn15261,n14374);
and (s0n15261,notn15261,1'b0);
and (s1n15261,n14374,n15262);
and (n15263,n15264,n14412);
wire s0n15264,s1n15264,notn15264;
or (n15264,s0n15264,s1n15264);
not(notn15264,n42);
and (s0n15264,notn15264,1'b0);
and (s1n15264,n42,n15265);
wire s0n15265,s1n15265,notn15265;
or (n15265,s0n15265,s1n15265);
not(notn15265,n14375);
and (s0n15265,notn15265,n15266);
and (s1n15265,n14375,n15268);
wire s0n15266,s1n15266,notn15266;
or (n15266,s0n15266,s1n15266);
not(notn15266,n14409);
and (s0n15266,notn15266,n15267);
and (s1n15266,n14409,n15253);
wire s0n15267,s1n15267,notn15267;
or (n15267,s0n15267,s1n15267);
not(notn15267,n14401);
and (s0n15267,notn15267,1'b0);
and (s1n15267,n14401,n15249);
and (n15269,n15270,n14421);
wire s0n15270,s1n15270,notn15270;
or (n15270,s0n15270,s1n15270);
not(notn15270,n42);
and (s0n15270,notn15270,1'b0);
and (s1n15270,n42,n15271);
wire s0n15271,s1n15271,notn15271;
or (n15271,s0n15271,s1n15271);
not(notn15271,n14375);
and (s0n15271,notn15271,n15272);
and (s1n15271,n14375,n15274);
wire s0n15272,s1n15272,notn15272;
or (n15272,s0n15272,s1n15272);
not(notn15272,n14409);
and (s0n15272,notn15272,n15273);
and (s1n15272,n14409,n15255);
wire s0n15273,s1n15273,notn15273;
or (n15273,s0n15273,s1n15273);
not(notn15273,n14401);
and (s0n15273,notn15273,1'b0);
and (s1n15273,n14401,n15251);
and (n15275,n15276,n14137);
or (n15276,1'b0,n15277,n15287);
and (n15277,n15278,n14235);
wire s0n15278,s1n15278,notn15278;
or (n15278,s0n15278,s1n15278);
not(notn15278,n14227);
and (s0n15278,notn15278,1'b0);
and (s1n15278,n14227,n15279);
or (n15279,1'b0,n15091,n15280,n15281,n15282,n15283,n15286);
and (n15280,n15022,n14199);
and (n15281,n15024,n2781);
and (n15282,n15017,n14205);
and (n15283,n15284,n2789);
wire s0n15284,s1n15284,notn15284;
or (n15284,s0n15284,s1n15284);
not(notn15284,n14210);
and (s0n15284,notn15284,n15066);
and (s1n15284,n14210,n15285);
and (n15286,n15285,n14225);
and (n15287,n15039,n14455);
and (n15288,n15289,n14111);
wire s0n15289,s1n15289,notn15289;
or (n15289,s0n15289,s1n15289);
not(notn15289,n14455);
and (s0n15289,notn15289,1'b0);
and (s1n15289,n14455,n15151);
and (n15290,n15291,n14108);
wire s0n15291,s1n15291,notn15291;
or (n15291,s0n15291,s1n15291);
not(notn15291,n14131);
and (s0n15291,notn15291,1'b0);
and (s1n15291,n14131,n15119);
and (n15292,n15293,n13950);
wire s0n15293,s1n15293,notn15293;
or (n15293,s0n15293,s1n15293);
not(notn15293,n14131);
and (s0n15293,notn15293,1'b0);
and (s1n15293,n14131,n15151);
and (n15294,n15295,n14239);
wire s0n15295,s1n15295,notn15295;
or (n15295,s0n15295,s1n15295);
not(notn15295,n14131);
and (s0n15295,notn15295,1'b0);
and (s1n15295,n14131,n15278);
and (n15296,n15222,n15297);
or (n15297,n15298,n15635,n17025);
and (n15298,n15299,n15562);
wire s0n15299,s1n15299,notn15299;
or (n15299,s0n15299,s1n15299);
not(notn15299,n14631);
and (s0n15299,notn15299,n15300);
and (s1n15299,n14631,n15426);
wire s0n15300,s1n15300,notn15300;
or (n15300,s0n15300,s1n15300);
not(notn15300,n14271);
and (s0n15300,notn15300,n15301);
and (s1n15300,n14271,n15414);
wire s0n15301,s1n15301,notn15301;
or (n15301,s0n15301,s1n15301);
not(notn15301,n14279);
and (s0n15301,notn15301,1'b0);
and (s1n15301,n14279,n15302);
or (n15302,1'b0,n15303,n15316,n15382);
and (n15303,n15304,n14120);
wire s0n15304,s1n15304,notn15304;
or (n15304,s0n15304,s1n15304);
not(notn15304,n14125);
and (s0n15304,notn15304,1'b0);
and (s1n15304,n14125,n15305);
wire s0n15305,s1n15305,notn15305;
or (n15305,s0n15305,s1n15305);
not(notn15305,n14317);
and (s0n15305,notn15305,n15306);
and (s1n15305,n14317,n15307);
wire s0n15307,s1n15307,notn15307;
or (n15307,s0n15307,s1n15307);
not(notn15307,n14326);
and (s0n15307,notn15307,n15308);
and (s1n15307,n14326,n15310);
wire s0n15308,s1n15308,notn15308;
or (n15308,s0n15308,s1n15308);
not(notn15308,n14315);
and (s0n15308,notn15308,1'b0);
and (s1n15308,n14315,n15309);
or (n15310,1'b0,n15311,n15313,n15315);
and (n15311,n15312,n14321);
and (n15313,n15314,n14324);
and (n15315,n15309,n14184);
and (n15316,n15317,n14718);
or (n15317,1'b0,n15318,n15334,n15350,n15366);
and (n15318,n15319,n13889);
wire s0n15319,s1n15319,notn15319;
or (n15319,s0n15319,s1n15319);
not(notn15319,n42);
and (s0n15319,notn15319,1'b0);
and (s1n15319,n42,n15320);
wire s0n15320,s1n15320,notn15320;
or (n15320,s0n15320,s1n15320);
not(notn15320,n14187);
and (s0n15320,notn15320,n15321);
and (s1n15320,n14187,n15327);
wire s0n15321,s1n15321,notn15321;
or (n15321,s0n15321,s1n15321);
not(notn15321,n14163);
and (s0n15321,notn15321,1'b0);
and (s1n15321,n14163,n15322);
or (n15322,1'b0,n15323,n15325);
and (n15323,n15324,n14147);
and (n15325,n15326,n14156);
or (n15327,1'b0,n15328,n15330,n15332,n15333);
and (n15328,n15329,n14171);
and (n15330,n15331,n14176);
and (n15332,n15324,n14180);
and (n15333,n15326,n14184);
and (n15334,n15335,n13897);
wire s0n15335,s1n15335,notn15335;
or (n15335,s0n15335,s1n15335);
not(notn15335,n42);
and (s0n15335,notn15335,1'b0);
and (s1n15335,n42,n15336);
wire s0n15336,s1n15336,notn15336;
or (n15336,s0n15336,s1n15336);
not(notn15336,n14187);
and (s0n15336,notn15336,n15337);
and (s1n15336,n14187,n15343);
wire s0n15337,s1n15337,notn15337;
or (n15337,s0n15337,s1n15337);
not(notn15337,n14163);
and (s0n15337,notn15337,1'b0);
and (s1n15337,n14163,n15338);
or (n15338,1'b0,n15339,n15341);
and (n15339,n15340,n14147);
and (n15341,n15342,n14156);
or (n15343,1'b0,n15344,n15346,n15348,n15349);
and (n15344,n15345,n14171);
and (n15346,n15347,n14176);
and (n15348,n15340,n14180);
and (n15349,n15342,n14184);
and (n15350,n15351,n13900);
wire s0n15351,s1n15351,notn15351;
or (n15351,s0n15351,s1n15351);
not(notn15351,n42);
and (s0n15351,notn15351,1'b0);
and (s1n15351,n42,n15352);
wire s0n15352,s1n15352,notn15352;
or (n15352,s0n15352,s1n15352);
not(notn15352,n14187);
and (s0n15352,notn15352,n15353);
and (s1n15352,n14187,n15359);
wire s0n15353,s1n15353,notn15353;
or (n15353,s0n15353,s1n15353);
not(notn15353,n14163);
and (s0n15353,notn15353,1'b0);
and (s1n15353,n14163,n15354);
or (n15354,1'b0,n15355,n15357);
and (n15355,n15356,n14147);
and (n15357,n15358,n14156);
or (n15359,1'b0,n15360,n15362,n15364,n15365);
and (n15360,n15361,n14171);
and (n15362,n15363,n14176);
and (n15364,n15356,n14180);
and (n15365,n15358,n14184);
and (n15366,n15367,n14131);
wire s0n15367,s1n15367,notn15367;
or (n15367,s0n15367,s1n15367);
not(notn15367,n42);
and (s0n15367,notn15367,1'b0);
and (s1n15367,n42,n15368);
wire s0n15368,s1n15368,notn15368;
or (n15368,s0n15368,s1n15368);
not(notn15368,n14187);
and (s0n15368,notn15368,n15369);
and (s1n15368,n14187,n15375);
wire s0n15369,s1n15369,notn15369;
or (n15369,s0n15369,s1n15369);
not(notn15369,n14163);
and (s0n15369,notn15369,1'b0);
and (s1n15369,n14163,n15370);
or (n15370,1'b0,n15371,n15373);
and (n15371,n15372,n14147);
and (n15373,n15374,n14156);
or (n15375,1'b0,n15376,n15378,n15380,n15381);
and (n15376,n15377,n14171);
and (n15378,n15379,n14176);
and (n15380,n15372,n14180);
and (n15381,n15374,n14184);
and (n15382,n15383,n14365);
wire s0n15383,s1n15383,notn15383;
or (n15383,s0n15383,s1n15383);
not(notn15383,n42);
and (s0n15383,notn15383,1'b0);
and (s1n15383,n42,n15384);
wire s0n15384,s1n15384,notn15384;
or (n15384,s0n15384,s1n15384);
not(notn15384,n14422);
and (s0n15384,notn15384,n15385);
and (s1n15384,n14422,n15395);
wire s0n15385,s1n15385,notn15385;
or (n15385,s0n15385,s1n15385);
not(notn15385,n14362);
and (s0n15385,notn15385,1'b0);
and (s1n15385,n14362,n15386);
or (n15386,1'b0,n15387,n15389,n15391,n15393);
and (n15387,n15388,n14352);
and (n15389,n15390,n14355);
and (n15391,n15392,n14358);
and (n15393,n15394,n14361);
or (n15395,1'b0,n15396,n15399,n15402,n15408);
and (n15396,n15397,n14387);
wire s0n15397,s1n15397,notn15397;
or (n15397,s0n15397,s1n15397);
not(notn15397,n14374);
and (s0n15397,notn15397,1'b0);
and (s1n15397,n14374,n15398);
and (n15399,n15400,n14393);
wire s0n15400,s1n15400,notn15400;
or (n15400,s0n15400,s1n15400);
not(notn15400,n14374);
and (s0n15400,notn15400,1'b0);
and (s1n15400,n14374,n15401);
and (n15402,n15403,n14412);
wire s0n15403,s1n15403,notn15403;
or (n15403,s0n15403,s1n15403);
not(notn15403,n42);
and (s0n15403,notn15403,1'b0);
and (s1n15403,n42,n15404);
wire s0n15404,s1n15404,notn15404;
or (n15404,s0n15404,s1n15404);
not(notn15404,n14375);
and (s0n15404,notn15404,n15405);
and (s1n15404,n14375,n15407);
wire s0n15405,s1n15405,notn15405;
or (n15405,s0n15405,s1n15405);
not(notn15405,n14409);
and (s0n15405,notn15405,n15406);
and (s1n15405,n14409,n15392);
wire s0n15406,s1n15406,notn15406;
or (n15406,s0n15406,s1n15406);
not(notn15406,n14401);
and (s0n15406,notn15406,1'b0);
and (s1n15406,n14401,n15388);
and (n15408,n15409,n14421);
wire s0n15409,s1n15409,notn15409;
or (n15409,s0n15409,s1n15409);
not(notn15409,n42);
and (s0n15409,notn15409,1'b0);
and (s1n15409,n42,n15410);
wire s0n15410,s1n15410,notn15410;
or (n15410,s0n15410,s1n15410);
not(notn15410,n14375);
and (s0n15410,notn15410,n15411);
and (s1n15410,n14375,n15413);
wire s0n15411,s1n15411,notn15411;
or (n15411,s0n15411,s1n15411);
not(notn15411,n14409);
and (s0n15411,notn15411,n15412);
and (s1n15411,n14409,n15394);
wire s0n15412,s1n15412,notn15412;
or (n15412,s0n15412,s1n15412);
not(notn15412,n14401);
and (s0n15412,notn15412,1'b0);
and (s1n15412,n14401,n15390);
or (n15414,n15415,n15416,n15424,n15425);
and (n15415,n15304,n13907);
and (n15416,n15417,n14385);
wire s0n15417,s1n15417,notn15417;
or (n15417,s0n15417,s1n15417);
not(notn15417,n2799);
and (s0n15417,notn15417,1'b0);
and (s1n15417,n2799,n15418);
or (n15418,1'b0,n15419,n15420);
and (n15419,n15306,n13900);
and (n15420,n15421,n14131);
wire s0n15421,s1n15421,notn15421;
or (n15421,s0n15421,s1n15421);
not(notn15421,n14573);
and (s0n15421,notn15421,n15422);
and (s1n15421,n14573,1'b0);
wire s0n15422,s1n15422,notn15422;
or (n15422,s0n15422,s1n15422);
not(notn15422,n14374);
and (s0n15422,notn15422,1'b0);
and (s1n15422,n14374,n15423);
and (n15424,n15383,n14381);
and (n15425,n15317,n14192);
or (n15426,1'b0,n15427,n15432,n15447,n15515,n15546,n15552,n15560,n15561);
and (n15427,n15428,n14237);
or (n15428,1'b0,n15429,n15431);
and (n15429,n15430,n14235);
wire s0n15431,s1n15431,notn15431;
or (n15431,s0n15431,s1n15431);
not(notn15431,n14455);
and (s0n15431,notn15431,1'b0);
and (s1n15431,n14455,n15383);
and (n15432,n15433,n14137);
or (n15433,1'b0,n15434,n15445,n15446);
and (n15434,n15435,n13889);
wire s0n15435,s1n15435,notn15435;
or (n15435,s0n15435,s1n15435);
not(notn15435,n14227);
and (s0n15435,notn15435,1'b0);
and (s1n15435,n14227,n15436);
or (n15436,1'b0,n15437,n15438,n15439,n15440,n15441,n15444);
and (n15437,n15319,n14193);
and (n15438,n15361,n14199);
and (n15439,n15363,n2781);
and (n15440,n15356,n14205);
and (n15441,n15442,n2789);
wire s0n15442,s1n15442,notn15442;
or (n15442,s0n15442,s1n15442);
not(notn15442,n14210);
and (s0n15442,notn15442,n15329);
and (s1n15442,n14210,n15443);
and (n15444,n15443,n14225);
and (n15445,n15319,n14243);
and (n15446,n15351,n14131);
and (n15447,n15448,n14111);
or (n15448,1'b0,n15449,n15451,n15453,n15483);
and (n15449,n15450,n13889);
and (n15451,n15452,n13897);
and (n15453,n15454,n13900);
wire s0n15454,s1n15454,notn15454;
or (n15454,s0n15454,s1n15454);
not(notn15454,n42);
and (s0n15454,notn15454,1'b0);
and (s1n15454,n42,n15455);
wire s0n15455,s1n15455,notn15455;
or (n15455,s0n15455,s1n15455);
not(notn15455,n14422);
and (s0n15455,notn15455,n15456);
and (s1n15455,n14422,n15466);
wire s0n15456,s1n15456,notn15456;
or (n15456,s0n15456,s1n15456);
not(notn15456,n14362);
and (s0n15456,notn15456,1'b0);
and (s1n15456,n14362,n15457);
or (n15457,1'b0,n15458,n15460,n15462,n15464);
and (n15458,n15459,n14352);
and (n15460,n15461,n14355);
and (n15462,n15463,n14358);
and (n15464,n15465,n14361);
or (n15466,1'b0,n15467,n15470,n15471,n15477);
and (n15467,n15468,n14387);
wire s0n15468,s1n15468,notn15468;
or (n15468,s0n15468,s1n15468);
not(notn15468,n14374);
and (s0n15468,notn15468,1'b0);
and (s1n15468,n14374,n15469);
and (n15470,n15422,n14393);
and (n15471,n15472,n14412);
wire s0n15472,s1n15472,notn15472;
or (n15472,s0n15472,s1n15472);
not(notn15472,n42);
and (s0n15472,notn15472,1'b0);
and (s1n15472,n42,n15473);
wire s0n15473,s1n15473,notn15473;
or (n15473,s0n15473,s1n15473);
not(notn15473,n14375);
and (s0n15473,notn15473,n15474);
and (s1n15473,n14375,n15476);
wire s0n15474,s1n15474,notn15474;
or (n15474,s0n15474,s1n15474);
not(notn15474,n14409);
and (s0n15474,notn15474,n15475);
and (s1n15474,n14409,n15463);
wire s0n15475,s1n15475,notn15475;
or (n15475,s0n15475,s1n15475);
not(notn15475,n14401);
and (s0n15475,notn15475,1'b0);
and (s1n15475,n14401,n15459);
and (n15477,n15478,n14421);
wire s0n15478,s1n15478,notn15478;
or (n15478,s0n15478,s1n15478);
not(notn15478,n42);
and (s0n15478,notn15478,1'b0);
and (s1n15478,n42,n15479);
wire s0n15479,s1n15479,notn15479;
or (n15479,s0n15479,s1n15479);
not(notn15479,n14375);
and (s0n15479,notn15479,n15480);
and (s1n15479,n14375,n15482);
wire s0n15480,s1n15480,notn15480;
or (n15480,s0n15480,s1n15480);
not(notn15480,n14409);
and (s0n15480,notn15480,n15481);
and (s1n15480,n14409,n15465);
wire s0n15481,s1n15481,notn15481;
or (n15481,s0n15481,s1n15481);
not(notn15481,n14401);
and (s0n15481,notn15481,1'b0);
and (s1n15481,n14401,n15461);
wire s0n15483,s1n15483,notn15483;
or (n15483,s0n15483,s1n15483);
not(notn15483,n14131);
and (s0n15483,notn15483,1'b0);
and (s1n15483,n14131,n15484);
wire s0n15484,s1n15484,notn15484;
or (n15484,s0n15484,s1n15484);
not(notn15484,n42);
and (s0n15484,notn15484,1'b0);
and (s1n15484,n42,n15485);
wire s0n15485,s1n15485,notn15485;
or (n15485,s0n15485,s1n15485);
not(notn15485,n14422);
and (s0n15485,notn15485,n15486);
and (s1n15485,n14422,n15496);
wire s0n15486,s1n15486,notn15486;
or (n15486,s0n15486,s1n15486);
not(notn15486,n14362);
and (s0n15486,notn15486,1'b0);
and (s1n15486,n14362,n15487);
or (n15487,1'b0,n15488,n15490,n15492,n15494);
and (n15488,n15489,n14352);
and (n15490,n15491,n14355);
and (n15492,n15493,n14358);
and (n15494,n15495,n14361);
or (n15496,1'b0,n15497,n15500,n15503,n15509);
and (n15497,n15498,n14387);
wire s0n15498,s1n15498,notn15498;
or (n15498,s0n15498,s1n15498);
not(notn15498,n14374);
and (s0n15498,notn15498,1'b0);
and (s1n15498,n14374,n15499);
and (n15500,n15501,n14393);
wire s0n15501,s1n15501,notn15501;
or (n15501,s0n15501,s1n15501);
not(notn15501,n14374);
and (s0n15501,notn15501,1'b0);
and (s1n15501,n14374,n15502);
and (n15503,n15504,n14412);
wire s0n15504,s1n15504,notn15504;
or (n15504,s0n15504,s1n15504);
not(notn15504,n42);
and (s0n15504,notn15504,1'b0);
and (s1n15504,n42,n15505);
wire s0n15505,s1n15505,notn15505;
or (n15505,s0n15505,s1n15505);
not(notn15505,n14375);
and (s0n15505,notn15505,n15506);
and (s1n15505,n14375,n15508);
wire s0n15506,s1n15506,notn15506;
or (n15506,s0n15506,s1n15506);
not(notn15506,n14409);
and (s0n15506,notn15506,n15507);
and (s1n15506,n14409,n15493);
wire s0n15507,s1n15507,notn15507;
or (n15507,s0n15507,s1n15507);
not(notn15507,n14401);
and (s0n15507,notn15507,1'b0);
and (s1n15507,n14401,n15489);
and (n15509,n15510,n14421);
wire s0n15510,s1n15510,notn15510;
or (n15510,s0n15510,s1n15510);
not(notn15510,n42);
and (s0n15510,notn15510,1'b0);
and (s1n15510,n42,n15511);
wire s0n15511,s1n15511,notn15511;
or (n15511,s0n15511,s1n15511);
not(notn15511,n14375);
and (s0n15511,notn15511,n15512);
and (s1n15511,n14375,n15514);
wire s0n15512,s1n15512,notn15512;
or (n15512,s0n15512,s1n15512);
not(notn15512,n14409);
and (s0n15512,notn15512,n15513);
and (s1n15512,n14409,n15495);
wire s0n15513,s1n15513,notn15513;
or (n15513,s0n15513,s1n15513);
not(notn15513,n14401);
and (s0n15513,notn15513,1'b0);
and (s1n15513,n14401,n15491);
not (n15515,n15516);
nand (n15516,n15517,n14108);
or (n15517,1'b0,n15518,n15520,n15522,n15524);
and (n15518,n15519,n13889);
and (n15520,n15521,n13897);
and (n15522,n15523,n13900);
and (n15524,n15525,n14131);
wire s0n15525,s1n15525,notn15525;
or (n15525,s0n15525,s1n15525);
not(notn15525,n14123);
and (s0n15525,notn15525,1'b0);
and (s1n15525,n14123,n15526);
wire s0n15526,s1n15526,notn15526;
or (n15526,s0n15526,s1n15526);
not(notn15526,n555);
and (s0n15526,notn15526,n15527);
and (s1n15526,n555,n15542);
wire s0n15527,s1n15527,notn15527;
or (n15527,s0n15527,s1n15527);
not(notn15527,n13948);
and (s0n15527,notn15527,n15528);
and (s1n15527,n13948,n15530);
wire s0n15528,s1n15528,notn15528;
or (n15528,s0n15528,s1n15528);
not(notn15528,n13907);
and (s0n15528,notn15528,1'b0);
and (s1n15528,n13907,n15529);
or (n15530,n15531,n15533,n15535,n15537,n15539,n15541);
and (n15531,n15532,n13913);
and (n15533,n15534,n13920);
and (n15535,n15536,n13923);
and (n15537,n15538,n13928);
and (n15539,n15540,n13935);
and (n15541,n15529,n13941);
wire s0n15542,s1n15542,notn15542;
or (n15542,s0n15542,s1n15542);
not(notn15542,n14119);
and (s0n15542,notn15542,1'b0);
and (s1n15542,n14119,n15543);
wire s0n15543,s1n15543,notn15543;
or (n15543,s0n15543,s1n15543);
not(notn15543,n14116);
and (s0n15543,notn15543,n15544);
and (s1n15543,n14116,n15545);
and (n15546,n15547,n13950);
or (n15547,1'b0,n15548,n15549,n15550,n15551);
and (n15548,n15521,n13889);
and (n15549,n15523,n13897);
and (n15550,n15452,n13900);
wire s0n15551,s1n15551,notn15551;
or (n15551,s0n15551,s1n15551);
not(notn15551,n14131);
and (s0n15551,notn15551,1'b0);
and (s1n15551,n14131,n15454);
and (n15552,n15553,n14239);
or (n15553,1'b0,n15554,n15556,n15558,n15559);
and (n15554,n15555,n13889);
and (n15556,n15557,n13897);
and (n15558,n15430,n13900);
and (n15559,n15335,n14131);
and (n15560,n15383,n14448);
and (n15561,n15317,n14266);
wire s0n15562,s1n15562,notn15562;
or (n15562,s0n15562,s1n15562);
not(notn15562,n14631);
and (s0n15562,notn15562,n15563);
and (s1n15562,n14631,n15581);
wire s0n15563,s1n15563,notn15563;
or (n15563,s0n15563,s1n15563);
not(notn15563,n14271);
and (s0n15563,notn15563,n15564);
and (s1n15563,n14271,n15569);
wire s0n15564,s1n15564,notn15564;
or (n15564,s0n15564,s1n15564);
not(notn15564,n14279);
and (s0n15564,notn15564,1'b0);
and (s1n15564,n14279,n15565);
and (n15565,n15566,n14120);
wire s0n15566,s1n15566,notn15566;
or (n15566,s0n15566,s1n15566);
not(notn15566,n14125);
and (s0n15566,notn15566,1'b0);
and (s1n15566,n14125,n15567);
wire s0n15567,s1n15567,notn15567;
or (n15567,s0n15567,s1n15567);
not(notn15567,n14317);
and (s0n15567,notn15567,n15568);
and (s1n15567,n14317,n15233);
or (n15569,n15570,n15574,1'b0);
and (n15570,n15571,n13907);
wire s0n15571,s1n15571,notn15571;
or (n15571,s0n15571,s1n15571);
not(notn15571,n14125);
and (s0n15571,notn15571,1'b0);
and (s1n15571,n14125,n15572);
wire s0n15572,s1n15572,notn15572;
or (n15572,s0n15572,s1n15572);
not(notn15572,n14563);
and (s0n15572,notn15572,n15568);
and (s1n15572,n14563,n15573);
and (n15574,n15575,n14385);
wire s0n15575,s1n15575,notn15575;
or (n15575,s0n15575,s1n15575);
not(notn15575,n2799);
and (s0n15575,notn15575,1'b0);
and (s1n15575,n2799,n15576);
or (n15576,1'b0,n15577,n15579);
and (n15577,n15578,n13900);
wire s0n15578,s1n15578,notn15578;
or (n15578,s0n15578,s1n15578);
not(notn15578,n14570);
and (s0n15578,notn15578,n15363);
and (s1n15578,n14570,1'b0);
and (n15579,n15580,n14131);
wire s0n15580,s1n15580,notn15580;
or (n15580,s0n15580,s1n15580);
not(notn15580,n14573);
and (s0n15580,notn15580,n15501);
and (s1n15580,n14573,1'b0);
or (n15581,n15582,n15615,n15628,n15629,n15631,n15633,1'b0);
and (n15582,n15583,n14237);
wire s0n15583,s1n15583,notn15583;
or (n15583,s0n15583,s1n15583);
not(notn15583,n14455);
and (s0n15583,notn15583,1'b0);
and (s1n15583,n14455,n15584);
wire s0n15584,s1n15584,notn15584;
or (n15584,s0n15584,s1n15584);
not(notn15584,n42);
and (s0n15584,notn15584,1'b0);
and (s1n15584,n42,n15585);
wire s0n15585,s1n15585,notn15585;
or (n15585,s0n15585,s1n15585);
not(notn15585,n14422);
and (s0n15585,notn15585,n15586);
and (s1n15585,n14422,n15596);
wire s0n15586,s1n15586,notn15586;
or (n15586,s0n15586,s1n15586);
not(notn15586,n14362);
and (s0n15586,notn15586,1'b0);
and (s1n15586,n14362,n15587);
or (n15587,1'b0,n15588,n15590,n15592,n15594);
and (n15588,n15589,n14352);
and (n15590,n15591,n14355);
and (n15592,n15593,n14358);
and (n15594,n15595,n14361);
or (n15596,1'b0,n15597,n15600,n15603,n15609);
and (n15597,n15598,n14387);
wire s0n15598,s1n15598,notn15598;
or (n15598,s0n15598,s1n15598);
not(notn15598,n14374);
and (s0n15598,notn15598,1'b0);
and (s1n15598,n14374,n15599);
and (n15600,n15601,n14393);
wire s0n15601,s1n15601,notn15601;
or (n15601,s0n15601,s1n15601);
not(notn15601,n14374);
and (s0n15601,notn15601,1'b0);
and (s1n15601,n14374,n15602);
and (n15603,n15604,n14412);
wire s0n15604,s1n15604,notn15604;
or (n15604,s0n15604,s1n15604);
not(notn15604,n42);
and (s0n15604,notn15604,1'b0);
and (s1n15604,n42,n15605);
wire s0n15605,s1n15605,notn15605;
or (n15605,s0n15605,s1n15605);
not(notn15605,n14375);
and (s0n15605,notn15605,n15606);
and (s1n15605,n14375,n15608);
wire s0n15606,s1n15606,notn15606;
or (n15606,s0n15606,s1n15606);
not(notn15606,n14409);
and (s0n15606,notn15606,n15607);
and (s1n15606,n14409,n15593);
wire s0n15607,s1n15607,notn15607;
or (n15607,s0n15607,s1n15607);
not(notn15607,n14401);
and (s0n15607,notn15607,1'b0);
and (s1n15607,n14401,n15589);
and (n15609,n15610,n14421);
wire s0n15610,s1n15610,notn15610;
or (n15610,s0n15610,s1n15610);
not(notn15610,n42);
and (s0n15610,notn15610,1'b0);
and (s1n15610,n42,n15611);
wire s0n15611,s1n15611,notn15611;
or (n15611,s0n15611,s1n15611);
not(notn15611,n14375);
and (s0n15611,notn15611,n15612);
and (s1n15611,n14375,n15614);
wire s0n15612,s1n15612,notn15612;
or (n15612,s0n15612,s1n15612);
not(notn15612,n14409);
and (s0n15612,notn15612,n15613);
and (s1n15612,n14409,n15595);
wire s0n15613,s1n15613,notn15613;
or (n15613,s0n15613,s1n15613);
not(notn15613,n14401);
and (s0n15613,notn15613,1'b0);
and (s1n15613,n14401,n15591);
and (n15615,n15616,n14137);
or (n15616,1'b0,n15617,n15627);
and (n15617,n15618,n14235);
wire s0n15618,s1n15618,notn15618;
or (n15618,s0n15618,s1n15618);
not(notn15618,n14227);
and (s0n15618,notn15618,1'b0);
and (s1n15618,n14227,n15619);
or (n15619,1'b0,n15437,n15620,n15621,n15622,n15623,n15626);
and (n15620,n15377,n14199);
and (n15621,n15379,n2781);
and (n15622,n15372,n14205);
and (n15623,n15624,n2789);
wire s0n15624,s1n15624,notn15624;
or (n15624,s0n15624,s1n15624);
not(notn15624,n14210);
and (s0n15624,notn15624,n15329);
and (s1n15624,n14210,n15625);
and (n15626,n15625,n14225);
and (n15627,n15335,n14455);
and (n15628,n15431,n14111);
not (n15629,n15630);
nand (n15630,n14625,n15484);
and (n15631,n15632,n13950);
wire s0n15632,s1n15632,notn15632;
or (n15632,s0n15632,s1n15632);
not(notn15632,n14131);
and (s0n15632,notn15632,1'b0);
and (s1n15632,n14131,n15383);
and (n15633,n15634,n14239);
wire s0n15634,s1n15634,notn15634;
or (n15634,s0n15634,s1n15634);
not(notn15634,n14131);
and (s0n15634,notn15634,1'b0);
and (s1n15634,n14131,n15618);
and (n15635,n15562,n15636);
or (n15636,n15637,n15975,n17024);
and (n15637,n15638,n15901);
wire s0n15638,s1n15638,notn15638;
or (n15638,s0n15638,s1n15638);
not(notn15638,n14631);
and (s0n15638,notn15638,n15639);
and (s1n15638,n14631,n15765);
wire s0n15639,s1n15639,notn15639;
or (n15639,s0n15639,s1n15639);
not(notn15639,n14271);
and (s0n15639,notn15639,n15640);
and (s1n15639,n14271,n15753);
wire s0n15640,s1n15640,notn15640;
or (n15640,s0n15640,s1n15640);
not(notn15640,n14279);
and (s0n15640,notn15640,1'b0);
and (s1n15640,n14279,n15641);
or (n15641,1'b0,n15642,n15655,n15721);
and (n15642,n15643,n14120);
wire s0n15643,s1n15643,notn15643;
or (n15643,s0n15643,s1n15643);
not(notn15643,n14125);
and (s0n15643,notn15643,1'b0);
and (s1n15643,n14125,n15644);
wire s0n15644,s1n15644,notn15644;
or (n15644,s0n15644,s1n15644);
not(notn15644,n14317);
and (s0n15644,notn15644,n15645);
and (s1n15644,n14317,n15646);
wire s0n15646,s1n15646,notn15646;
or (n15646,s0n15646,s1n15646);
not(notn15646,n14326);
and (s0n15646,notn15646,n15647);
and (s1n15646,n14326,n15649);
wire s0n15647,s1n15647,notn15647;
or (n15647,s0n15647,s1n15647);
not(notn15647,n14315);
and (s0n15647,notn15647,1'b0);
and (s1n15647,n14315,n15648);
or (n15649,1'b0,n15650,n15652,n15654);
and (n15650,n15651,n14321);
and (n15652,n15653,n14324);
and (n15654,n15648,n14184);
and (n15655,n15656,n14718);
or (n15656,1'b0,n15657,n15673,n15689,n15705);
and (n15657,n15658,n13889);
wire s0n15658,s1n15658,notn15658;
or (n15658,s0n15658,s1n15658);
not(notn15658,n42);
and (s0n15658,notn15658,1'b0);
and (s1n15658,n42,n15659);
wire s0n15659,s1n15659,notn15659;
or (n15659,s0n15659,s1n15659);
not(notn15659,n14187);
and (s0n15659,notn15659,n15660);
and (s1n15659,n14187,n15666);
wire s0n15660,s1n15660,notn15660;
or (n15660,s0n15660,s1n15660);
not(notn15660,n14163);
and (s0n15660,notn15660,1'b0);
and (s1n15660,n14163,n15661);
or (n15661,1'b0,n15662,n15664);
and (n15662,n15663,n14147);
and (n15664,n15665,n14156);
or (n15666,1'b0,n15667,n15669,n15671,n15672);
and (n15667,n15668,n14171);
and (n15669,n15670,n14176);
and (n15671,n15663,n14180);
and (n15672,n15665,n14184);
and (n15673,n15674,n13897);
wire s0n15674,s1n15674,notn15674;
or (n15674,s0n15674,s1n15674);
not(notn15674,n42);
and (s0n15674,notn15674,1'b0);
and (s1n15674,n42,n15675);
wire s0n15675,s1n15675,notn15675;
or (n15675,s0n15675,s1n15675);
not(notn15675,n14187);
and (s0n15675,notn15675,n15676);
and (s1n15675,n14187,n15682);
wire s0n15676,s1n15676,notn15676;
or (n15676,s0n15676,s1n15676);
not(notn15676,n14163);
and (s0n15676,notn15676,1'b0);
and (s1n15676,n14163,n15677);
or (n15677,1'b0,n15678,n15680);
and (n15678,n15679,n14147);
and (n15680,n15681,n14156);
or (n15682,1'b0,n15683,n15685,n15687,n15688);
and (n15683,n15684,n14171);
and (n15685,n15686,n14176);
and (n15687,n15679,n14180);
and (n15688,n15681,n14184);
and (n15689,n15690,n13900);
wire s0n15690,s1n15690,notn15690;
or (n15690,s0n15690,s1n15690);
not(notn15690,n42);
and (s0n15690,notn15690,1'b0);
and (s1n15690,n42,n15691);
wire s0n15691,s1n15691,notn15691;
or (n15691,s0n15691,s1n15691);
not(notn15691,n14187);
and (s0n15691,notn15691,n15692);
and (s1n15691,n14187,n15698);
wire s0n15692,s1n15692,notn15692;
or (n15692,s0n15692,s1n15692);
not(notn15692,n14163);
and (s0n15692,notn15692,1'b0);
and (s1n15692,n14163,n15693);
or (n15693,1'b0,n15694,n15696);
and (n15694,n15695,n14147);
and (n15696,n15697,n14156);
or (n15698,1'b0,n15699,n15701,n15703,n15704);
and (n15699,n15700,n14171);
and (n15701,n15702,n14176);
and (n15703,n15695,n14180);
and (n15704,n15697,n14184);
and (n15705,n15706,n14131);
wire s0n15706,s1n15706,notn15706;
or (n15706,s0n15706,s1n15706);
not(notn15706,n42);
and (s0n15706,notn15706,1'b0);
and (s1n15706,n42,n15707);
wire s0n15707,s1n15707,notn15707;
or (n15707,s0n15707,s1n15707);
not(notn15707,n14187);
and (s0n15707,notn15707,n15708);
and (s1n15707,n14187,n15714);
wire s0n15708,s1n15708,notn15708;
or (n15708,s0n15708,s1n15708);
not(notn15708,n14163);
and (s0n15708,notn15708,1'b0);
and (s1n15708,n14163,n15709);
or (n15709,1'b0,n15710,n15712);
and (n15710,n15711,n14147);
and (n15712,n15713,n14156);
or (n15714,1'b0,n15715,n15717,n15719,n15720);
and (n15715,n15716,n14171);
and (n15717,n15718,n14176);
and (n15719,n15711,n14180);
and (n15720,n15713,n14184);
and (n15721,n15722,n14365);
wire s0n15722,s1n15722,notn15722;
or (n15722,s0n15722,s1n15722);
not(notn15722,n42);
and (s0n15722,notn15722,1'b0);
and (s1n15722,n42,n15723);
wire s0n15723,s1n15723,notn15723;
or (n15723,s0n15723,s1n15723);
not(notn15723,n14422);
and (s0n15723,notn15723,n15724);
and (s1n15723,n14422,n15734);
wire s0n15724,s1n15724,notn15724;
or (n15724,s0n15724,s1n15724);
not(notn15724,n14362);
and (s0n15724,notn15724,1'b0);
and (s1n15724,n14362,n15725);
or (n15725,1'b0,n15726,n15728,n15730,n15732);
and (n15726,n15727,n14352);
and (n15728,n15729,n14355);
and (n15730,n15731,n14358);
and (n15732,n15733,n14361);
or (n15734,1'b0,n15735,n15738,n15741,n15747);
and (n15735,n15736,n14387);
wire s0n15736,s1n15736,notn15736;
or (n15736,s0n15736,s1n15736);
not(notn15736,n14374);
and (s0n15736,notn15736,1'b0);
and (s1n15736,n14374,n15737);
and (n15738,n15739,n14393);
wire s0n15739,s1n15739,notn15739;
or (n15739,s0n15739,s1n15739);
not(notn15739,n14374);
and (s0n15739,notn15739,1'b0);
and (s1n15739,n14374,n15740);
and (n15741,n15742,n14412);
wire s0n15742,s1n15742,notn15742;
or (n15742,s0n15742,s1n15742);
not(notn15742,n42);
and (s0n15742,notn15742,1'b0);
and (s1n15742,n42,n15743);
wire s0n15743,s1n15743,notn15743;
or (n15743,s0n15743,s1n15743);
not(notn15743,n14375);
and (s0n15743,notn15743,n15744);
and (s1n15743,n14375,n15746);
wire s0n15744,s1n15744,notn15744;
or (n15744,s0n15744,s1n15744);
not(notn15744,n14409);
and (s0n15744,notn15744,n15745);
and (s1n15744,n14409,n15731);
wire s0n15745,s1n15745,notn15745;
or (n15745,s0n15745,s1n15745);
not(notn15745,n14401);
and (s0n15745,notn15745,1'b0);
and (s1n15745,n14401,n15727);
and (n15747,n15748,n14421);
wire s0n15748,s1n15748,notn15748;
or (n15748,s0n15748,s1n15748);
not(notn15748,n42);
and (s0n15748,notn15748,1'b0);
and (s1n15748,n42,n15749);
wire s0n15749,s1n15749,notn15749;
or (n15749,s0n15749,s1n15749);
not(notn15749,n14375);
and (s0n15749,notn15749,n15750);
and (s1n15749,n14375,n15752);
wire s0n15750,s1n15750,notn15750;
or (n15750,s0n15750,s1n15750);
not(notn15750,n14409);
and (s0n15750,notn15750,n15751);
and (s1n15750,n14409,n15733);
wire s0n15751,s1n15751,notn15751;
or (n15751,s0n15751,s1n15751);
not(notn15751,n14401);
and (s0n15751,notn15751,1'b0);
and (s1n15751,n14401,n15729);
or (n15753,n15754,n15755,n15763,n15764);
and (n15754,n15643,n13907);
and (n15755,n15756,n14385);
wire s0n15756,s1n15756,notn15756;
or (n15756,s0n15756,s1n15756);
not(notn15756,n2799);
and (s0n15756,notn15756,1'b0);
and (s1n15756,n2799,n15757);
or (n15757,1'b0,n15758,n15759);
and (n15758,n15645,n13900);
and (n15759,n15760,n14131);
wire s0n15760,s1n15760,notn15760;
or (n15760,s0n15760,s1n15760);
not(notn15760,n14573);
and (s0n15760,notn15760,n15761);
and (s1n15760,n14573,1'b0);
wire s0n15761,s1n15761,notn15761;
or (n15761,s0n15761,s1n15761);
not(notn15761,n14374);
and (s0n15761,notn15761,1'b0);
and (s1n15761,n14374,n15762);
and (n15763,n15722,n14381);
and (n15764,n15656,n14192);
or (n15765,1'b0,n15766,n15771,n15786,n15854,n15885,n15891,n15899,n15900);
and (n15766,n15767,n14237);
or (n15767,1'b0,n15768,n15770);
and (n15768,n15769,n14235);
wire s0n15770,s1n15770,notn15770;
or (n15770,s0n15770,s1n15770);
not(notn15770,n14455);
and (s0n15770,notn15770,1'b0);
and (s1n15770,n14455,n15722);
and (n15771,n15772,n14137);
or (n15772,1'b0,n15773,n15784,n15785);
and (n15773,n15774,n13889);
wire s0n15774,s1n15774,notn15774;
or (n15774,s0n15774,s1n15774);
not(notn15774,n14227);
and (s0n15774,notn15774,1'b0);
and (s1n15774,n14227,n15775);
or (n15775,1'b0,n15776,n15777,n15778,n15779,n15780,n15783);
and (n15776,n15658,n14193);
and (n15777,n15700,n14199);
and (n15778,n15702,n2781);
and (n15779,n15695,n14205);
and (n15780,n15781,n2789);
wire s0n15781,s1n15781,notn15781;
or (n15781,s0n15781,s1n15781);
not(notn15781,n14210);
and (s0n15781,notn15781,n15668);
and (s1n15781,n14210,n15782);
and (n15783,n15782,n14225);
and (n15784,n15658,n14243);
and (n15785,n15690,n14131);
and (n15786,n15787,n14111);
or (n15787,1'b0,n15788,n15790,n15792,n15822);
and (n15788,n15789,n13889);
and (n15790,n15791,n13897);
and (n15792,n15793,n13900);
wire s0n15793,s1n15793,notn15793;
or (n15793,s0n15793,s1n15793);
not(notn15793,n42);
and (s0n15793,notn15793,1'b0);
and (s1n15793,n42,n15794);
wire s0n15794,s1n15794,notn15794;
or (n15794,s0n15794,s1n15794);
not(notn15794,n14422);
and (s0n15794,notn15794,n15795);
and (s1n15794,n14422,n15805);
wire s0n15795,s1n15795,notn15795;
or (n15795,s0n15795,s1n15795);
not(notn15795,n14362);
and (s0n15795,notn15795,1'b0);
and (s1n15795,n14362,n15796);
or (n15796,1'b0,n15797,n15799,n15801,n15803);
and (n15797,n15798,n14352);
and (n15799,n15800,n14355);
and (n15801,n15802,n14358);
and (n15803,n15804,n14361);
or (n15805,1'b0,n15806,n15809,n15810,n15816);
and (n15806,n15807,n14387);
wire s0n15807,s1n15807,notn15807;
or (n15807,s0n15807,s1n15807);
not(notn15807,n14374);
and (s0n15807,notn15807,1'b0);
and (s1n15807,n14374,n15808);
and (n15809,n15761,n14393);
and (n15810,n15811,n14412);
wire s0n15811,s1n15811,notn15811;
or (n15811,s0n15811,s1n15811);
not(notn15811,n42);
and (s0n15811,notn15811,1'b0);
and (s1n15811,n42,n15812);
wire s0n15812,s1n15812,notn15812;
or (n15812,s0n15812,s1n15812);
not(notn15812,n14375);
and (s0n15812,notn15812,n15813);
and (s1n15812,n14375,n15815);
wire s0n15813,s1n15813,notn15813;
or (n15813,s0n15813,s1n15813);
not(notn15813,n14409);
and (s0n15813,notn15813,n15814);
and (s1n15813,n14409,n15802);
wire s0n15814,s1n15814,notn15814;
or (n15814,s0n15814,s1n15814);
not(notn15814,n14401);
and (s0n15814,notn15814,1'b0);
and (s1n15814,n14401,n15798);
and (n15816,n15817,n14421);
wire s0n15817,s1n15817,notn15817;
or (n15817,s0n15817,s1n15817);
not(notn15817,n42);
and (s0n15817,notn15817,1'b0);
and (s1n15817,n42,n15818);
wire s0n15818,s1n15818,notn15818;
or (n15818,s0n15818,s1n15818);
not(notn15818,n14375);
and (s0n15818,notn15818,n15819);
and (s1n15818,n14375,n15821);
wire s0n15819,s1n15819,notn15819;
or (n15819,s0n15819,s1n15819);
not(notn15819,n14409);
and (s0n15819,notn15819,n15820);
and (s1n15819,n14409,n15804);
wire s0n15820,s1n15820,notn15820;
or (n15820,s0n15820,s1n15820);
not(notn15820,n14401);
and (s0n15820,notn15820,1'b0);
and (s1n15820,n14401,n15800);
wire s0n15822,s1n15822,notn15822;
or (n15822,s0n15822,s1n15822);
not(notn15822,n14131);
and (s0n15822,notn15822,1'b0);
and (s1n15822,n14131,n15823);
wire s0n15823,s1n15823,notn15823;
or (n15823,s0n15823,s1n15823);
not(notn15823,n42);
and (s0n15823,notn15823,1'b0);
and (s1n15823,n42,n15824);
wire s0n15824,s1n15824,notn15824;
or (n15824,s0n15824,s1n15824);
not(notn15824,n14422);
and (s0n15824,notn15824,n15825);
and (s1n15824,n14422,n15835);
wire s0n15825,s1n15825,notn15825;
or (n15825,s0n15825,s1n15825);
not(notn15825,n14362);
and (s0n15825,notn15825,1'b0);
and (s1n15825,n14362,n15826);
or (n15826,1'b0,n15827,n15829,n15831,n15833);
and (n15827,n15828,n14352);
and (n15829,n15830,n14355);
and (n15831,n15832,n14358);
and (n15833,n15834,n14361);
or (n15835,1'b0,n15836,n15839,n15842,n15848);
and (n15836,n15837,n14387);
wire s0n15837,s1n15837,notn15837;
or (n15837,s0n15837,s1n15837);
not(notn15837,n14374);
and (s0n15837,notn15837,1'b0);
and (s1n15837,n14374,n15838);
and (n15839,n15840,n14393);
wire s0n15840,s1n15840,notn15840;
or (n15840,s0n15840,s1n15840);
not(notn15840,n14374);
and (s0n15840,notn15840,1'b0);
and (s1n15840,n14374,n15841);
and (n15842,n15843,n14412);
wire s0n15843,s1n15843,notn15843;
or (n15843,s0n15843,s1n15843);
not(notn15843,n42);
and (s0n15843,notn15843,1'b0);
and (s1n15843,n42,n15844);
wire s0n15844,s1n15844,notn15844;
or (n15844,s0n15844,s1n15844);
not(notn15844,n14375);
and (s0n15844,notn15844,n15845);
and (s1n15844,n14375,n15847);
wire s0n15845,s1n15845,notn15845;
or (n15845,s0n15845,s1n15845);
not(notn15845,n14409);
and (s0n15845,notn15845,n15846);
and (s1n15845,n14409,n15832);
wire s0n15846,s1n15846,notn15846;
or (n15846,s0n15846,s1n15846);
not(notn15846,n14401);
and (s0n15846,notn15846,1'b0);
and (s1n15846,n14401,n15828);
and (n15848,n15849,n14421);
wire s0n15849,s1n15849,notn15849;
or (n15849,s0n15849,s1n15849);
not(notn15849,n42);
and (s0n15849,notn15849,1'b0);
and (s1n15849,n42,n15850);
wire s0n15850,s1n15850,notn15850;
or (n15850,s0n15850,s1n15850);
not(notn15850,n14375);
and (s0n15850,notn15850,n15851);
and (s1n15850,n14375,n15853);
wire s0n15851,s1n15851,notn15851;
or (n15851,s0n15851,s1n15851);
not(notn15851,n14409);
and (s0n15851,notn15851,n15852);
and (s1n15851,n14409,n15834);
wire s0n15852,s1n15852,notn15852;
or (n15852,s0n15852,s1n15852);
not(notn15852,n14401);
and (s0n15852,notn15852,1'b0);
and (s1n15852,n14401,n15830);
not (n15854,n15855);
nand (n15855,n15856,n14108);
or (n15856,1'b0,n15857,n15859,n15861,n15863);
and (n15857,n15858,n13889);
and (n15859,n15860,n13897);
and (n15861,n15862,n13900);
and (n15863,n15864,n14131);
wire s0n15864,s1n15864,notn15864;
or (n15864,s0n15864,s1n15864);
not(notn15864,n14123);
and (s0n15864,notn15864,1'b0);
and (s1n15864,n14123,n15865);
wire s0n15865,s1n15865,notn15865;
or (n15865,s0n15865,s1n15865);
not(notn15865,n555);
and (s0n15865,notn15865,n15866);
and (s1n15865,n555,n15881);
wire s0n15866,s1n15866,notn15866;
or (n15866,s0n15866,s1n15866);
not(notn15866,n13948);
and (s0n15866,notn15866,n15867);
and (s1n15866,n13948,n15869);
wire s0n15867,s1n15867,notn15867;
or (n15867,s0n15867,s1n15867);
not(notn15867,n13907);
and (s0n15867,notn15867,1'b0);
and (s1n15867,n13907,n15868);
or (n15869,n15870,n15872,n15874,n15876,n15878,n15880);
and (n15870,n15871,n13913);
and (n15872,n15873,n13920);
and (n15874,n15875,n13923);
and (n15876,n15877,n13928);
and (n15878,n15879,n13935);
and (n15880,n15868,n13941);
wire s0n15881,s1n15881,notn15881;
or (n15881,s0n15881,s1n15881);
not(notn15881,n14119);
and (s0n15881,notn15881,1'b0);
and (s1n15881,n14119,n15882);
wire s0n15882,s1n15882,notn15882;
or (n15882,s0n15882,s1n15882);
not(notn15882,n14116);
and (s0n15882,notn15882,n15883);
and (s1n15882,n14116,n15884);
and (n15885,n15886,n13950);
or (n15886,1'b0,n15887,n15888,n15889,n15890);
and (n15887,n15860,n13889);
and (n15888,n15862,n13897);
and (n15889,n15791,n13900);
wire s0n15890,s1n15890,notn15890;
or (n15890,s0n15890,s1n15890);
not(notn15890,n14131);
and (s0n15890,notn15890,1'b0);
and (s1n15890,n14131,n15793);
and (n15891,n15892,n14239);
or (n15892,1'b0,n15893,n15895,n15897,n15898);
and (n15893,n15894,n13889);
and (n15895,n15896,n13897);
and (n15897,n15769,n13900);
and (n15898,n15674,n14131);
and (n15899,n15722,n14448);
and (n15900,n15656,n14266);
wire s0n15901,s1n15901,notn15901;
or (n15901,s0n15901,s1n15901);
not(notn15901,n14631);
and (s0n15901,notn15901,n15902);
and (s1n15901,n14631,n15920);
wire s0n15902,s1n15902,notn15902;
or (n15902,s0n15902,s1n15902);
not(notn15902,n14271);
and (s0n15902,notn15902,n15903);
and (s1n15902,n14271,n15908);
wire s0n15903,s1n15903,notn15903;
or (n15903,s0n15903,s1n15903);
not(notn15903,n14279);
and (s0n15903,notn15903,1'b0);
and (s1n15903,n14279,n15904);
and (n15904,n15905,n14120);
wire s0n15905,s1n15905,notn15905;
or (n15905,s0n15905,s1n15905);
not(notn15905,n14125);
and (s0n15905,notn15905,1'b0);
and (s1n15905,n14125,n15906);
wire s0n15906,s1n15906,notn15906;
or (n15906,s0n15906,s1n15906);
not(notn15906,n14317);
and (s0n15906,notn15906,n15907);
and (s1n15906,n14317,n15573);
or (n15908,n15909,n15913,1'b0);
and (n15909,n15910,n13907);
wire s0n15910,s1n15910,notn15910;
or (n15910,s0n15910,s1n15910);
not(notn15910,n14125);
and (s0n15910,notn15910,1'b0);
and (s1n15910,n14125,n15911);
wire s0n15911,s1n15911,notn15911;
or (n15911,s0n15911,s1n15911);
not(notn15911,n14563);
and (s0n15911,notn15911,n15907);
and (s1n15911,n14563,n15912);
and (n15913,n15914,n14385);
wire s0n15914,s1n15914,notn15914;
or (n15914,s0n15914,s1n15914);
not(notn15914,n2799);
and (s0n15914,notn15914,1'b0);
and (s1n15914,n2799,n15915);
or (n15915,1'b0,n15916,n15918);
and (n15916,n15917,n13900);
wire s0n15917,s1n15917,notn15917;
or (n15917,s0n15917,s1n15917);
not(notn15917,n14570);
and (s0n15917,notn15917,n15702);
and (s1n15917,n14570,1'b0);
and (n15918,n15919,n14131);
wire s0n15919,s1n15919,notn15919;
or (n15919,s0n15919,s1n15919);
not(notn15919,n14573);
and (s0n15919,notn15919,n15840);
and (s1n15919,n14573,1'b0);
or (n15920,n15921,n15954,n15967,n15968,n15971,n15973,1'b0);
and (n15921,n15922,n14237);
wire s0n15922,s1n15922,notn15922;
or (n15922,s0n15922,s1n15922);
not(notn15922,n14455);
and (s0n15922,notn15922,1'b0);
and (s1n15922,n14455,n15923);
wire s0n15923,s1n15923,notn15923;
or (n15923,s0n15923,s1n15923);
not(notn15923,n42);
and (s0n15923,notn15923,1'b0);
and (s1n15923,n42,n15924);
wire s0n15924,s1n15924,notn15924;
or (n15924,s0n15924,s1n15924);
not(notn15924,n14422);
and (s0n15924,notn15924,n15925);
and (s1n15924,n14422,n15935);
wire s0n15925,s1n15925,notn15925;
or (n15925,s0n15925,s1n15925);
not(notn15925,n14362);
and (s0n15925,notn15925,1'b0);
and (s1n15925,n14362,n15926);
or (n15926,1'b0,n15927,n15929,n15931,n15933);
and (n15927,n15928,n14352);
and (n15929,n15930,n14355);
and (n15931,n15932,n14358);
and (n15933,n15934,n14361);
or (n15935,1'b0,n15936,n15939,n15942,n15948);
and (n15936,n15937,n14387);
wire s0n15937,s1n15937,notn15937;
or (n15937,s0n15937,s1n15937);
not(notn15937,n14374);
and (s0n15937,notn15937,1'b0);
and (s1n15937,n14374,n15938);
and (n15939,n15940,n14393);
wire s0n15940,s1n15940,notn15940;
or (n15940,s0n15940,s1n15940);
not(notn15940,n14374);
and (s0n15940,notn15940,1'b0);
and (s1n15940,n14374,n15941);
and (n15942,n15943,n14412);
wire s0n15943,s1n15943,notn15943;
or (n15943,s0n15943,s1n15943);
not(notn15943,n42);
and (s0n15943,notn15943,1'b0);
and (s1n15943,n42,n15944);
wire s0n15944,s1n15944,notn15944;
or (n15944,s0n15944,s1n15944);
not(notn15944,n14375);
and (s0n15944,notn15944,n15945);
and (s1n15944,n14375,n15947);
wire s0n15945,s1n15945,notn15945;
or (n15945,s0n15945,s1n15945);
not(notn15945,n14409);
and (s0n15945,notn15945,n15946);
and (s1n15945,n14409,n15932);
wire s0n15946,s1n15946,notn15946;
or (n15946,s0n15946,s1n15946);
not(notn15946,n14401);
and (s0n15946,notn15946,1'b0);
and (s1n15946,n14401,n15928);
and (n15948,n15949,n14421);
wire s0n15949,s1n15949,notn15949;
or (n15949,s0n15949,s1n15949);
not(notn15949,n42);
and (s0n15949,notn15949,1'b0);
and (s1n15949,n42,n15950);
wire s0n15950,s1n15950,notn15950;
or (n15950,s0n15950,s1n15950);
not(notn15950,n14375);
and (s0n15950,notn15950,n15951);
and (s1n15950,n14375,n15953);
wire s0n15951,s1n15951,notn15951;
or (n15951,s0n15951,s1n15951);
not(notn15951,n14409);
and (s0n15951,notn15951,n15952);
and (s1n15951,n14409,n15934);
wire s0n15952,s1n15952,notn15952;
or (n15952,s0n15952,s1n15952);
not(notn15952,n14401);
and (s0n15952,notn15952,1'b0);
and (s1n15952,n14401,n15930);
and (n15954,n15955,n14137);
or (n15955,1'b0,n15956,n15966);
and (n15956,n15957,n14235);
wire s0n15957,s1n15957,notn15957;
or (n15957,s0n15957,s1n15957);
not(notn15957,n14227);
and (s0n15957,notn15957,1'b0);
and (s1n15957,n14227,n15958);
or (n15958,1'b0,n15776,n15959,n15960,n15961,n15962,n15965);
and (n15959,n15716,n14199);
and (n15960,n15718,n2781);
and (n15961,n15711,n14205);
and (n15962,n15963,n2789);
wire s0n15963,s1n15963,notn15963;
or (n15963,s0n15963,s1n15963);
not(notn15963,n14210);
and (s0n15963,notn15963,n15668);
and (s1n15963,n14210,n15964);
and (n15965,n15964,n14225);
and (n15966,n15674,n14455);
and (n15967,n15770,n14111);
not (n15968,n15969);
or (n15969,n14626,n15970);
not (n15970,n15823);
and (n15971,n15972,n13950);
wire s0n15972,s1n15972,notn15972;
or (n15972,s0n15972,s1n15972);
not(notn15972,n14131);
and (s0n15972,notn15972,1'b0);
and (s1n15972,n14131,n15722);
and (n15973,n15974,n14239);
wire s0n15974,s1n15974,notn15974;
or (n15974,s0n15974,s1n15974);
not(notn15974,n14131);
and (s0n15974,notn15974,1'b0);
and (s1n15974,n14131,n15957);
and (n15975,n15901,n15976);
or (n15976,n15977,n16315,n17023);
and (n15977,n15978,n16241);
wire s0n15978,s1n15978,notn15978;
or (n15978,s0n15978,s1n15978);
not(notn15978,n14631);
and (s0n15978,notn15978,n15979);
and (s1n15978,n14631,n16105);
wire s0n15979,s1n15979,notn15979;
or (n15979,s0n15979,s1n15979);
not(notn15979,n14271);
and (s0n15979,notn15979,n15980);
and (s1n15979,n14271,n16093);
wire s0n15980,s1n15980,notn15980;
or (n15980,s0n15980,s1n15980);
not(notn15980,n14279);
and (s0n15980,notn15980,1'b0);
and (s1n15980,n14279,n15981);
or (n15981,1'b0,n15982,n15995,n16061);
and (n15982,n15983,n14120);
wire s0n15983,s1n15983,notn15983;
or (n15983,s0n15983,s1n15983);
not(notn15983,n14125);
and (s0n15983,notn15983,1'b0);
and (s1n15983,n14125,n15984);
wire s0n15984,s1n15984,notn15984;
or (n15984,s0n15984,s1n15984);
not(notn15984,n14317);
and (s0n15984,notn15984,n15985);
and (s1n15984,n14317,n15986);
wire s0n15986,s1n15986,notn15986;
or (n15986,s0n15986,s1n15986);
not(notn15986,n14326);
and (s0n15986,notn15986,n15987);
and (s1n15986,n14326,n15989);
wire s0n15987,s1n15987,notn15987;
or (n15987,s0n15987,s1n15987);
not(notn15987,n14315);
and (s0n15987,notn15987,1'b0);
and (s1n15987,n14315,n15988);
or (n15989,1'b0,n15990,n15992,n15994);
and (n15990,n15991,n14321);
and (n15992,n15993,n14324);
and (n15994,n15988,n14184);
and (n15995,n15996,n14718);
or (n15996,1'b0,n15997,n16013,n16029,n16045);
and (n15997,n15998,n13889);
wire s0n15998,s1n15998,notn15998;
or (n15998,s0n15998,s1n15998);
not(notn15998,n42);
and (s0n15998,notn15998,1'b0);
and (s1n15998,n42,n15999);
wire s0n15999,s1n15999,notn15999;
or (n15999,s0n15999,s1n15999);
not(notn15999,n14187);
and (s0n15999,notn15999,n16000);
and (s1n15999,n14187,n16006);
wire s0n16000,s1n16000,notn16000;
or (n16000,s0n16000,s1n16000);
not(notn16000,n14163);
and (s0n16000,notn16000,1'b0);
and (s1n16000,n14163,n16001);
or (n16001,1'b0,n16002,n16004);
and (n16002,n16003,n14147);
and (n16004,n16005,n14156);
or (n16006,1'b0,n16007,n16009,n16011,n16012);
and (n16007,n16008,n14171);
and (n16009,n16010,n14176);
and (n16011,n16003,n14180);
and (n16012,n16005,n14184);
and (n16013,n16014,n13897);
wire s0n16014,s1n16014,notn16014;
or (n16014,s0n16014,s1n16014);
not(notn16014,n42);
and (s0n16014,notn16014,1'b0);
and (s1n16014,n42,n16015);
wire s0n16015,s1n16015,notn16015;
or (n16015,s0n16015,s1n16015);
not(notn16015,n14187);
and (s0n16015,notn16015,n16016);
and (s1n16015,n14187,n16022);
wire s0n16016,s1n16016,notn16016;
or (n16016,s0n16016,s1n16016);
not(notn16016,n14163);
and (s0n16016,notn16016,1'b0);
and (s1n16016,n14163,n16017);
or (n16017,1'b0,n16018,n16020);
and (n16018,n16019,n14147);
and (n16020,n16021,n14156);
or (n16022,1'b0,n16023,n16025,n16027,n16028);
and (n16023,n16024,n14171);
and (n16025,n16026,n14176);
and (n16027,n16019,n14180);
and (n16028,n16021,n14184);
and (n16029,n16030,n13900);
wire s0n16030,s1n16030,notn16030;
or (n16030,s0n16030,s1n16030);
not(notn16030,n42);
and (s0n16030,notn16030,1'b0);
and (s1n16030,n42,n16031);
wire s0n16031,s1n16031,notn16031;
or (n16031,s0n16031,s1n16031);
not(notn16031,n14187);
and (s0n16031,notn16031,n16032);
and (s1n16031,n14187,n16038);
wire s0n16032,s1n16032,notn16032;
or (n16032,s0n16032,s1n16032);
not(notn16032,n14163);
and (s0n16032,notn16032,1'b0);
and (s1n16032,n14163,n16033);
or (n16033,1'b0,n16034,n16036);
and (n16034,n16035,n14147);
and (n16036,n16037,n14156);
or (n16038,1'b0,n16039,n16041,n16043,n16044);
and (n16039,n16040,n14171);
and (n16041,n16042,n14176);
and (n16043,n16035,n14180);
and (n16044,n16037,n14184);
and (n16045,n16046,n14131);
wire s0n16046,s1n16046,notn16046;
or (n16046,s0n16046,s1n16046);
not(notn16046,n42);
and (s0n16046,notn16046,1'b0);
and (s1n16046,n42,n16047);
wire s0n16047,s1n16047,notn16047;
or (n16047,s0n16047,s1n16047);
not(notn16047,n14187);
and (s0n16047,notn16047,n16048);
and (s1n16047,n14187,n16054);
wire s0n16048,s1n16048,notn16048;
or (n16048,s0n16048,s1n16048);
not(notn16048,n14163);
and (s0n16048,notn16048,1'b0);
and (s1n16048,n14163,n16049);
or (n16049,1'b0,n16050,n16052);
and (n16050,n16051,n14147);
and (n16052,n16053,n14156);
or (n16054,1'b0,n16055,n16057,n16059,n16060);
and (n16055,n16056,n14171);
and (n16057,n16058,n14176);
and (n16059,n16051,n14180);
and (n16060,n16053,n14184);
and (n16061,n16062,n14365);
wire s0n16062,s1n16062,notn16062;
or (n16062,s0n16062,s1n16062);
not(notn16062,n42);
and (s0n16062,notn16062,1'b0);
and (s1n16062,n42,n16063);
wire s0n16063,s1n16063,notn16063;
or (n16063,s0n16063,s1n16063);
not(notn16063,n14422);
and (s0n16063,notn16063,n16064);
and (s1n16063,n14422,n16074);
wire s0n16064,s1n16064,notn16064;
or (n16064,s0n16064,s1n16064);
not(notn16064,n14362);
and (s0n16064,notn16064,1'b0);
and (s1n16064,n14362,n16065);
or (n16065,1'b0,n16066,n16068,n16070,n16072);
and (n16066,n16067,n14352);
and (n16068,n16069,n14355);
and (n16070,n16071,n14358);
and (n16072,n16073,n14361);
or (n16074,1'b0,n16075,n16078,n16081,n16087);
and (n16075,n16076,n14387);
wire s0n16076,s1n16076,notn16076;
or (n16076,s0n16076,s1n16076);
not(notn16076,n14374);
and (s0n16076,notn16076,1'b0);
and (s1n16076,n14374,n16077);
and (n16078,n16079,n14393);
wire s0n16079,s1n16079,notn16079;
or (n16079,s0n16079,s1n16079);
not(notn16079,n14374);
and (s0n16079,notn16079,1'b0);
and (s1n16079,n14374,n16080);
and (n16081,n16082,n14412);
wire s0n16082,s1n16082,notn16082;
or (n16082,s0n16082,s1n16082);
not(notn16082,n42);
and (s0n16082,notn16082,1'b0);
and (s1n16082,n42,n16083);
wire s0n16083,s1n16083,notn16083;
or (n16083,s0n16083,s1n16083);
not(notn16083,n14375);
and (s0n16083,notn16083,n16084);
and (s1n16083,n14375,n16086);
wire s0n16084,s1n16084,notn16084;
or (n16084,s0n16084,s1n16084);
not(notn16084,n14409);
and (s0n16084,notn16084,n16085);
and (s1n16084,n14409,n16071);
wire s0n16085,s1n16085,notn16085;
or (n16085,s0n16085,s1n16085);
not(notn16085,n14401);
and (s0n16085,notn16085,1'b0);
and (s1n16085,n14401,n16067);
and (n16087,n16088,n14421);
wire s0n16088,s1n16088,notn16088;
or (n16088,s0n16088,s1n16088);
not(notn16088,n42);
and (s0n16088,notn16088,1'b0);
and (s1n16088,n42,n16089);
wire s0n16089,s1n16089,notn16089;
or (n16089,s0n16089,s1n16089);
not(notn16089,n14375);
and (s0n16089,notn16089,n16090);
and (s1n16089,n14375,n16092);
wire s0n16090,s1n16090,notn16090;
or (n16090,s0n16090,s1n16090);
not(notn16090,n14409);
and (s0n16090,notn16090,n16091);
and (s1n16090,n14409,n16073);
wire s0n16091,s1n16091,notn16091;
or (n16091,s0n16091,s1n16091);
not(notn16091,n14401);
and (s0n16091,notn16091,1'b0);
and (s1n16091,n14401,n16069);
or (n16093,n16094,n16095,n16103,n16104);
and (n16094,n15983,n13907);
and (n16095,n16096,n14385);
wire s0n16096,s1n16096,notn16096;
or (n16096,s0n16096,s1n16096);
not(notn16096,n2799);
and (s0n16096,notn16096,1'b0);
and (s1n16096,n2799,n16097);
or (n16097,1'b0,n16098,n16099);
and (n16098,n15985,n13900);
and (n16099,n16100,n14131);
wire s0n16100,s1n16100,notn16100;
or (n16100,s0n16100,s1n16100);
not(notn16100,n14573);
and (s0n16100,notn16100,n16101);
and (s1n16100,n14573,1'b0);
wire s0n16101,s1n16101,notn16101;
or (n16101,s0n16101,s1n16101);
not(notn16101,n14374);
and (s0n16101,notn16101,1'b0);
and (s1n16101,n14374,n16102);
and (n16103,n16062,n14381);
and (n16104,n15996,n14192);
or (n16105,1'b0,n16106,n16111,n16126,n16194,n16225,n16231,n16239,n16240);
and (n16106,n16107,n14237);
or (n16107,1'b0,n16108,n16110);
and (n16108,n16109,n14235);
wire s0n16110,s1n16110,notn16110;
or (n16110,s0n16110,s1n16110);
not(notn16110,n14455);
and (s0n16110,notn16110,1'b0);
and (s1n16110,n14455,n16062);
and (n16111,n16112,n14137);
or (n16112,1'b0,n16113,n16124,n16125);
and (n16113,n16114,n13889);
wire s0n16114,s1n16114,notn16114;
or (n16114,s0n16114,s1n16114);
not(notn16114,n14227);
and (s0n16114,notn16114,1'b0);
and (s1n16114,n14227,n16115);
or (n16115,1'b0,n16116,n16117,n16118,n16119,n16120,n16123);
and (n16116,n15998,n14193);
and (n16117,n16040,n14199);
and (n16118,n16042,n2781);
and (n16119,n16035,n14205);
and (n16120,n16121,n2789);
wire s0n16121,s1n16121,notn16121;
or (n16121,s0n16121,s1n16121);
not(notn16121,n14210);
and (s0n16121,notn16121,n16008);
and (s1n16121,n14210,n16122);
and (n16123,n16122,n14225);
and (n16124,n15998,n14243);
and (n16125,n16030,n14131);
and (n16126,n16127,n14111);
or (n16127,1'b0,n16128,n16130,n16132,n16162);
and (n16128,n16129,n13889);
and (n16130,n16131,n13897);
and (n16132,n16133,n13900);
wire s0n16133,s1n16133,notn16133;
or (n16133,s0n16133,s1n16133);
not(notn16133,n42);
and (s0n16133,notn16133,1'b0);
and (s1n16133,n42,n16134);
wire s0n16134,s1n16134,notn16134;
or (n16134,s0n16134,s1n16134);
not(notn16134,n14422);
and (s0n16134,notn16134,n16135);
and (s1n16134,n14422,n16145);
wire s0n16135,s1n16135,notn16135;
or (n16135,s0n16135,s1n16135);
not(notn16135,n14362);
and (s0n16135,notn16135,1'b0);
and (s1n16135,n14362,n16136);
or (n16136,1'b0,n16137,n16139,n16141,n16143);
and (n16137,n16138,n14352);
and (n16139,n16140,n14355);
and (n16141,n16142,n14358);
and (n16143,n16144,n14361);
or (n16145,1'b0,n16146,n16149,n16150,n16156);
and (n16146,n16147,n14387);
wire s0n16147,s1n16147,notn16147;
or (n16147,s0n16147,s1n16147);
not(notn16147,n14374);
and (s0n16147,notn16147,1'b0);
and (s1n16147,n14374,n16148);
and (n16149,n16101,n14393);
and (n16150,n16151,n14412);
wire s0n16151,s1n16151,notn16151;
or (n16151,s0n16151,s1n16151);
not(notn16151,n42);
and (s0n16151,notn16151,1'b0);
and (s1n16151,n42,n16152);
wire s0n16152,s1n16152,notn16152;
or (n16152,s0n16152,s1n16152);
not(notn16152,n14375);
and (s0n16152,notn16152,n16153);
and (s1n16152,n14375,n16155);
wire s0n16153,s1n16153,notn16153;
or (n16153,s0n16153,s1n16153);
not(notn16153,n14409);
and (s0n16153,notn16153,n16154);
and (s1n16153,n14409,n16142);
wire s0n16154,s1n16154,notn16154;
or (n16154,s0n16154,s1n16154);
not(notn16154,n14401);
and (s0n16154,notn16154,1'b0);
and (s1n16154,n14401,n16138);
and (n16156,n16157,n14421);
wire s0n16157,s1n16157,notn16157;
or (n16157,s0n16157,s1n16157);
not(notn16157,n42);
and (s0n16157,notn16157,1'b0);
and (s1n16157,n42,n16158);
wire s0n16158,s1n16158,notn16158;
or (n16158,s0n16158,s1n16158);
not(notn16158,n14375);
and (s0n16158,notn16158,n16159);
and (s1n16158,n14375,n16161);
wire s0n16159,s1n16159,notn16159;
or (n16159,s0n16159,s1n16159);
not(notn16159,n14409);
and (s0n16159,notn16159,n16160);
and (s1n16159,n14409,n16144);
wire s0n16160,s1n16160,notn16160;
or (n16160,s0n16160,s1n16160);
not(notn16160,n14401);
and (s0n16160,notn16160,1'b0);
and (s1n16160,n14401,n16140);
wire s0n16162,s1n16162,notn16162;
or (n16162,s0n16162,s1n16162);
not(notn16162,n14131);
and (s0n16162,notn16162,1'b0);
and (s1n16162,n14131,n16163);
wire s0n16163,s1n16163,notn16163;
or (n16163,s0n16163,s1n16163);
not(notn16163,n42);
and (s0n16163,notn16163,1'b0);
and (s1n16163,n42,n16164);
wire s0n16164,s1n16164,notn16164;
or (n16164,s0n16164,s1n16164);
not(notn16164,n14422);
and (s0n16164,notn16164,n16165);
and (s1n16164,n14422,n16175);
wire s0n16165,s1n16165,notn16165;
or (n16165,s0n16165,s1n16165);
not(notn16165,n14362);
and (s0n16165,notn16165,1'b0);
and (s1n16165,n14362,n16166);
or (n16166,1'b0,n16167,n16169,n16171,n16173);
and (n16167,n16168,n14352);
and (n16169,n16170,n14355);
and (n16171,n16172,n14358);
and (n16173,n16174,n14361);
or (n16175,1'b0,n16176,n16179,n16182,n16188);
and (n16176,n16177,n14387);
wire s0n16177,s1n16177,notn16177;
or (n16177,s0n16177,s1n16177);
not(notn16177,n14374);
and (s0n16177,notn16177,1'b0);
and (s1n16177,n14374,n16178);
and (n16179,n16180,n14393);
wire s0n16180,s1n16180,notn16180;
or (n16180,s0n16180,s1n16180);
not(notn16180,n14374);
and (s0n16180,notn16180,1'b0);
and (s1n16180,n14374,n16181);
and (n16182,n16183,n14412);
wire s0n16183,s1n16183,notn16183;
or (n16183,s0n16183,s1n16183);
not(notn16183,n42);
and (s0n16183,notn16183,1'b0);
and (s1n16183,n42,n16184);
wire s0n16184,s1n16184,notn16184;
or (n16184,s0n16184,s1n16184);
not(notn16184,n14375);
and (s0n16184,notn16184,n16185);
and (s1n16184,n14375,n16187);
wire s0n16185,s1n16185,notn16185;
or (n16185,s0n16185,s1n16185);
not(notn16185,n14409);
and (s0n16185,notn16185,n16186);
and (s1n16185,n14409,n16172);
wire s0n16186,s1n16186,notn16186;
or (n16186,s0n16186,s1n16186);
not(notn16186,n14401);
and (s0n16186,notn16186,1'b0);
and (s1n16186,n14401,n16168);
and (n16188,n16189,n14421);
wire s0n16189,s1n16189,notn16189;
or (n16189,s0n16189,s1n16189);
not(notn16189,n42);
and (s0n16189,notn16189,1'b0);
and (s1n16189,n42,n16190);
wire s0n16190,s1n16190,notn16190;
or (n16190,s0n16190,s1n16190);
not(notn16190,n14375);
and (s0n16190,notn16190,n16191);
and (s1n16190,n14375,n16193);
wire s0n16191,s1n16191,notn16191;
or (n16191,s0n16191,s1n16191);
not(notn16191,n14409);
and (s0n16191,notn16191,n16192);
and (s1n16191,n14409,n16174);
wire s0n16192,s1n16192,notn16192;
or (n16192,s0n16192,s1n16192);
not(notn16192,n14401);
and (s0n16192,notn16192,1'b0);
and (s1n16192,n14401,n16170);
not (n16194,n16195);
nand (n16195,n16196,n14108);
or (n16196,1'b0,n16197,n16199,n16201,n16203);
and (n16197,n16198,n13889);
and (n16199,n16200,n13897);
and (n16201,n16202,n13900);
and (n16203,n16204,n14131);
wire s0n16204,s1n16204,notn16204;
or (n16204,s0n16204,s1n16204);
not(notn16204,n14123);
and (s0n16204,notn16204,1'b0);
and (s1n16204,n14123,n16205);
wire s0n16205,s1n16205,notn16205;
or (n16205,s0n16205,s1n16205);
not(notn16205,n555);
and (s0n16205,notn16205,n16206);
and (s1n16205,n555,n16221);
wire s0n16206,s1n16206,notn16206;
or (n16206,s0n16206,s1n16206);
not(notn16206,n13948);
and (s0n16206,notn16206,n16207);
and (s1n16206,n13948,n16209);
wire s0n16207,s1n16207,notn16207;
or (n16207,s0n16207,s1n16207);
not(notn16207,n13907);
and (s0n16207,notn16207,1'b0);
and (s1n16207,n13907,n16208);
or (n16209,n16210,n16212,n16214,n16216,n16218,n16220);
and (n16210,n16211,n13913);
and (n16212,n16213,n13920);
and (n16214,n16215,n13923);
and (n16216,n16217,n13928);
and (n16218,n16219,n13935);
and (n16220,n16208,n13941);
wire s0n16221,s1n16221,notn16221;
or (n16221,s0n16221,s1n16221);
not(notn16221,n14119);
and (s0n16221,notn16221,1'b0);
and (s1n16221,n14119,n16222);
wire s0n16222,s1n16222,notn16222;
or (n16222,s0n16222,s1n16222);
not(notn16222,n14116);
and (s0n16222,notn16222,n16223);
and (s1n16222,n14116,n16224);
and (n16225,n16226,n13950);
or (n16226,1'b0,n16227,n16228,n16229,n16230);
and (n16227,n16200,n13889);
and (n16228,n16202,n13897);
and (n16229,n16131,n13900);
wire s0n16230,s1n16230,notn16230;
or (n16230,s0n16230,s1n16230);
not(notn16230,n14131);
and (s0n16230,notn16230,1'b0);
and (s1n16230,n14131,n16133);
and (n16231,n16232,n14239);
or (n16232,1'b0,n16233,n16235,n16237,n16238);
and (n16233,n16234,n13889);
and (n16235,n16236,n13897);
and (n16237,n16109,n13900);
and (n16238,n16014,n14131);
and (n16239,n16062,n14448);
and (n16240,n15996,n14266);
wire s0n16241,s1n16241,notn16241;
or (n16241,s0n16241,s1n16241);
not(notn16241,n14631);
and (s0n16241,notn16241,n16242);
and (s1n16241,n14631,n16260);
wire s0n16242,s1n16242,notn16242;
or (n16242,s0n16242,s1n16242);
not(notn16242,n14271);
and (s0n16242,notn16242,n16243);
and (s1n16242,n14271,n16248);
wire s0n16243,s1n16243,notn16243;
or (n16243,s0n16243,s1n16243);
not(notn16243,n14279);
and (s0n16243,notn16243,1'b0);
and (s1n16243,n14279,n16244);
and (n16244,n16245,n14120);
wire s0n16245,s1n16245,notn16245;
or (n16245,s0n16245,s1n16245);
not(notn16245,n14125);
and (s0n16245,notn16245,1'b0);
and (s1n16245,n14125,n16246);
wire s0n16246,s1n16246,notn16246;
or (n16246,s0n16246,s1n16246);
not(notn16246,n14317);
and (s0n16246,notn16246,n16247);
and (s1n16246,n14317,n15912);
or (n16248,n16249,n16253,1'b0);
and (n16249,n16250,n13907);
wire s0n16250,s1n16250,notn16250;
or (n16250,s0n16250,s1n16250);
not(notn16250,n14125);
and (s0n16250,notn16250,1'b0);
and (s1n16250,n14125,n16251);
wire s0n16251,s1n16251,notn16251;
or (n16251,s0n16251,s1n16251);
not(notn16251,n14563);
and (s0n16251,notn16251,n16247);
and (s1n16251,n14563,n16252);
and (n16253,n16254,n14385);
wire s0n16254,s1n16254,notn16254;
or (n16254,s0n16254,s1n16254);
not(notn16254,n2799);
and (s0n16254,notn16254,1'b0);
and (s1n16254,n2799,n16255);
or (n16255,1'b0,n16256,n16258);
and (n16256,n16257,n13900);
wire s0n16257,s1n16257,notn16257;
or (n16257,s0n16257,s1n16257);
not(notn16257,n14570);
and (s0n16257,notn16257,n16042);
and (s1n16257,n14570,1'b0);
and (n16258,n16259,n14131);
wire s0n16259,s1n16259,notn16259;
or (n16259,s0n16259,s1n16259);
not(notn16259,n14573);
and (s0n16259,notn16259,n16180);
and (s1n16259,n14573,1'b0);
or (n16260,n16261,n16294,n16307,n16308,n16311,n16313,1'b0);
and (n16261,n16262,n14237);
wire s0n16262,s1n16262,notn16262;
or (n16262,s0n16262,s1n16262);
not(notn16262,n14455);
and (s0n16262,notn16262,1'b0);
and (s1n16262,n14455,n16263);
wire s0n16263,s1n16263,notn16263;
or (n16263,s0n16263,s1n16263);
not(notn16263,n42);
and (s0n16263,notn16263,1'b0);
and (s1n16263,n42,n16264);
wire s0n16264,s1n16264,notn16264;
or (n16264,s0n16264,s1n16264);
not(notn16264,n14422);
and (s0n16264,notn16264,n16265);
and (s1n16264,n14422,n16275);
wire s0n16265,s1n16265,notn16265;
or (n16265,s0n16265,s1n16265);
not(notn16265,n14362);
and (s0n16265,notn16265,1'b0);
and (s1n16265,n14362,n16266);
or (n16266,1'b0,n16267,n16269,n16271,n16273);
and (n16267,n16268,n14352);
and (n16269,n16270,n14355);
and (n16271,n16272,n14358);
and (n16273,n16274,n14361);
or (n16275,1'b0,n16276,n16279,n16282,n16288);
and (n16276,n16277,n14387);
wire s0n16277,s1n16277,notn16277;
or (n16277,s0n16277,s1n16277);
not(notn16277,n14374);
and (s0n16277,notn16277,1'b0);
and (s1n16277,n14374,n16278);
and (n16279,n16280,n14393);
wire s0n16280,s1n16280,notn16280;
or (n16280,s0n16280,s1n16280);
not(notn16280,n14374);
and (s0n16280,notn16280,1'b0);
and (s1n16280,n14374,n16281);
and (n16282,n16283,n14412);
wire s0n16283,s1n16283,notn16283;
or (n16283,s0n16283,s1n16283);
not(notn16283,n42);
and (s0n16283,notn16283,1'b0);
and (s1n16283,n42,n16284);
wire s0n16284,s1n16284,notn16284;
or (n16284,s0n16284,s1n16284);
not(notn16284,n14375);
and (s0n16284,notn16284,n16285);
and (s1n16284,n14375,n16287);
wire s0n16285,s1n16285,notn16285;
or (n16285,s0n16285,s1n16285);
not(notn16285,n14409);
and (s0n16285,notn16285,n16286);
and (s1n16285,n14409,n16272);
wire s0n16286,s1n16286,notn16286;
or (n16286,s0n16286,s1n16286);
not(notn16286,n14401);
and (s0n16286,notn16286,1'b0);
and (s1n16286,n14401,n16268);
and (n16288,n16289,n14421);
wire s0n16289,s1n16289,notn16289;
or (n16289,s0n16289,s1n16289);
not(notn16289,n42);
and (s0n16289,notn16289,1'b0);
and (s1n16289,n42,n16290);
wire s0n16290,s1n16290,notn16290;
or (n16290,s0n16290,s1n16290);
not(notn16290,n14375);
and (s0n16290,notn16290,n16291);
and (s1n16290,n14375,n16293);
wire s0n16291,s1n16291,notn16291;
or (n16291,s0n16291,s1n16291);
not(notn16291,n14409);
and (s0n16291,notn16291,n16292);
and (s1n16291,n14409,n16274);
wire s0n16292,s1n16292,notn16292;
or (n16292,s0n16292,s1n16292);
not(notn16292,n14401);
and (s0n16292,notn16292,1'b0);
and (s1n16292,n14401,n16270);
and (n16294,n16295,n14137);
or (n16295,1'b0,n16296,n16306);
and (n16296,n16297,n14235);
wire s0n16297,s1n16297,notn16297;
or (n16297,s0n16297,s1n16297);
not(notn16297,n14227);
and (s0n16297,notn16297,1'b0);
and (s1n16297,n14227,n16298);
or (n16298,1'b0,n16116,n16299,n16300,n16301,n16302,n16305);
and (n16299,n16056,n14199);
and (n16300,n16058,n2781);
and (n16301,n16051,n14205);
and (n16302,n16303,n2789);
wire s0n16303,s1n16303,notn16303;
or (n16303,s0n16303,s1n16303);
not(notn16303,n14210);
and (s0n16303,notn16303,n16008);
and (s1n16303,n14210,n16304);
and (n16305,n16304,n14225);
and (n16306,n16014,n14455);
and (n16307,n16110,n14111);
not (n16308,n16309);
or (n16309,n14626,n16310);
not (n16310,n16163);
and (n16311,n16312,n13950);
wire s0n16312,s1n16312,notn16312;
or (n16312,s0n16312,s1n16312);
not(notn16312,n14131);
and (s0n16312,notn16312,1'b0);
and (s1n16312,n14131,n16062);
and (n16313,n16314,n14239);
wire s0n16314,s1n16314,notn16314;
or (n16314,s0n16314,s1n16314);
not(notn16314,n14131);
and (s0n16314,notn16314,1'b0);
and (s1n16314,n14131,n16297);
and (n16315,n16241,n16316);
or (n16316,n16317,n16684,n17022);
and (n16317,n16318,n16581);
wire s0n16318,s1n16318,notn16318;
or (n16318,s0n16318,s1n16318);
not(notn16318,n14631);
and (s0n16318,notn16318,n16319);
and (s1n16318,n14631,n16445);
wire s0n16319,s1n16319,notn16319;
or (n16319,s0n16319,s1n16319);
not(notn16319,n14271);
and (s0n16319,notn16319,n16320);
and (s1n16319,n14271,n16433);
wire s0n16320,s1n16320,notn16320;
or (n16320,s0n16320,s1n16320);
not(notn16320,n14279);
and (s0n16320,notn16320,1'b0);
and (s1n16320,n14279,n16321);
or (n16321,1'b0,n16322,n16335,n16401);
and (n16322,n16323,n14120);
wire s0n16323,s1n16323,notn16323;
or (n16323,s0n16323,s1n16323);
not(notn16323,n14125);
and (s0n16323,notn16323,1'b0);
and (s1n16323,n14125,n16324);
wire s0n16324,s1n16324,notn16324;
or (n16324,s0n16324,s1n16324);
not(notn16324,n14317);
and (s0n16324,notn16324,n16325);
and (s1n16324,n14317,n16326);
wire s0n16326,s1n16326,notn16326;
or (n16326,s0n16326,s1n16326);
not(notn16326,n14326);
and (s0n16326,notn16326,n16327);
and (s1n16326,n14326,n16329);
wire s0n16327,s1n16327,notn16327;
or (n16327,s0n16327,s1n16327);
not(notn16327,n14315);
and (s0n16327,notn16327,1'b0);
and (s1n16327,n14315,n16328);
or (n16329,1'b0,n16330,n16332,n16334);
and (n16330,n16331,n14321);
and (n16332,n16333,n14324);
and (n16334,n16328,n14184);
and (n16335,n16336,n14718);
or (n16336,1'b0,n16337,n16353,n16369,n16385);
and (n16337,n16338,n13889);
wire s0n16338,s1n16338,notn16338;
or (n16338,s0n16338,s1n16338);
not(notn16338,n42);
and (s0n16338,notn16338,1'b0);
and (s1n16338,n42,n16339);
wire s0n16339,s1n16339,notn16339;
or (n16339,s0n16339,s1n16339);
not(notn16339,n14187);
and (s0n16339,notn16339,n16340);
and (s1n16339,n14187,n16346);
wire s0n16340,s1n16340,notn16340;
or (n16340,s0n16340,s1n16340);
not(notn16340,n14163);
and (s0n16340,notn16340,1'b0);
and (s1n16340,n14163,n16341);
or (n16341,1'b0,n16342,n16344);
and (n16342,n16343,n14147);
and (n16344,n16345,n14156);
or (n16346,1'b0,n16347,n16349,n16351,n16352);
and (n16347,n16348,n14171);
and (n16349,n16350,n14176);
and (n16351,n16343,n14180);
and (n16352,n16345,n14184);
and (n16353,n16354,n13897);
wire s0n16354,s1n16354,notn16354;
or (n16354,s0n16354,s1n16354);
not(notn16354,n42);
and (s0n16354,notn16354,1'b0);
and (s1n16354,n42,n16355);
wire s0n16355,s1n16355,notn16355;
or (n16355,s0n16355,s1n16355);
not(notn16355,n14187);
and (s0n16355,notn16355,n16356);
and (s1n16355,n14187,n16362);
wire s0n16356,s1n16356,notn16356;
or (n16356,s0n16356,s1n16356);
not(notn16356,n14163);
and (s0n16356,notn16356,1'b0);
and (s1n16356,n14163,n16357);
or (n16357,1'b0,n16358,n16360);
and (n16358,n16359,n14147);
and (n16360,n16361,n14156);
or (n16362,1'b0,n16363,n16365,n16367,n16368);
and (n16363,n16364,n14171);
and (n16365,n16366,n14176);
and (n16367,n16359,n14180);
and (n16368,n16361,n14184);
and (n16369,n16370,n13900);
wire s0n16370,s1n16370,notn16370;
or (n16370,s0n16370,s1n16370);
not(notn16370,n42);
and (s0n16370,notn16370,1'b0);
and (s1n16370,n42,n16371);
wire s0n16371,s1n16371,notn16371;
or (n16371,s0n16371,s1n16371);
not(notn16371,n14187);
and (s0n16371,notn16371,n16372);
and (s1n16371,n14187,n16378);
wire s0n16372,s1n16372,notn16372;
or (n16372,s0n16372,s1n16372);
not(notn16372,n14163);
and (s0n16372,notn16372,1'b0);
and (s1n16372,n14163,n16373);
or (n16373,1'b0,n16374,n16376);
and (n16374,n16375,n14147);
and (n16376,n16377,n14156);
or (n16378,1'b0,n16379,n16381,n16383,n16384);
and (n16379,n16380,n14171);
and (n16381,n16382,n14176);
and (n16383,n16375,n14180);
and (n16384,n16377,n14184);
and (n16385,n16386,n14131);
wire s0n16386,s1n16386,notn16386;
or (n16386,s0n16386,s1n16386);
not(notn16386,n42);
and (s0n16386,notn16386,1'b0);
and (s1n16386,n42,n16387);
wire s0n16387,s1n16387,notn16387;
or (n16387,s0n16387,s1n16387);
not(notn16387,n14187);
and (s0n16387,notn16387,n16388);
and (s1n16387,n14187,n16394);
wire s0n16388,s1n16388,notn16388;
or (n16388,s0n16388,s1n16388);
not(notn16388,n14163);
and (s0n16388,notn16388,1'b0);
and (s1n16388,n14163,n16389);
or (n16389,1'b0,n16390,n16392);
and (n16390,n16391,n14147);
and (n16392,n16393,n14156);
or (n16394,1'b0,n16395,n16397,n16399,n16400);
and (n16395,n16396,n14171);
and (n16397,n16398,n14176);
and (n16399,n16391,n14180);
and (n16400,n16393,n14184);
and (n16401,n16402,n14365);
wire s0n16402,s1n16402,notn16402;
or (n16402,s0n16402,s1n16402);
not(notn16402,n42);
and (s0n16402,notn16402,1'b0);
and (s1n16402,n42,n16403);
wire s0n16403,s1n16403,notn16403;
or (n16403,s0n16403,s1n16403);
not(notn16403,n14422);
and (s0n16403,notn16403,n16404);
and (s1n16403,n14422,n16414);
wire s0n16404,s1n16404,notn16404;
or (n16404,s0n16404,s1n16404);
not(notn16404,n14362);
and (s0n16404,notn16404,1'b0);
and (s1n16404,n14362,n16405);
or (n16405,1'b0,n16406,n16408,n16410,n16412);
and (n16406,n16407,n14352);
and (n16408,n16409,n14355);
and (n16410,n16411,n14358);
and (n16412,n16413,n14361);
or (n16414,1'b0,n16415,n16418,n16421,n16427);
and (n16415,n16416,n14387);
wire s0n16416,s1n16416,notn16416;
or (n16416,s0n16416,s1n16416);
not(notn16416,n14374);
and (s0n16416,notn16416,1'b0);
and (s1n16416,n14374,n16417);
and (n16418,n16419,n14393);
wire s0n16419,s1n16419,notn16419;
or (n16419,s0n16419,s1n16419);
not(notn16419,n14374);
and (s0n16419,notn16419,1'b0);
and (s1n16419,n14374,n16420);
and (n16421,n16422,n14412);
wire s0n16422,s1n16422,notn16422;
or (n16422,s0n16422,s1n16422);
not(notn16422,n42);
and (s0n16422,notn16422,1'b0);
and (s1n16422,n42,n16423);
wire s0n16423,s1n16423,notn16423;
or (n16423,s0n16423,s1n16423);
not(notn16423,n14375);
and (s0n16423,notn16423,n16424);
and (s1n16423,n14375,n16426);
wire s0n16424,s1n16424,notn16424;
or (n16424,s0n16424,s1n16424);
not(notn16424,n14409);
and (s0n16424,notn16424,n16425);
and (s1n16424,n14409,n16411);
wire s0n16425,s1n16425,notn16425;
or (n16425,s0n16425,s1n16425);
not(notn16425,n14401);
and (s0n16425,notn16425,1'b0);
and (s1n16425,n14401,n16407);
and (n16427,n16428,n14421);
wire s0n16428,s1n16428,notn16428;
or (n16428,s0n16428,s1n16428);
not(notn16428,n42);
and (s0n16428,notn16428,1'b0);
and (s1n16428,n42,n16429);
wire s0n16429,s1n16429,notn16429;
or (n16429,s0n16429,s1n16429);
not(notn16429,n14375);
and (s0n16429,notn16429,n16430);
and (s1n16429,n14375,n16432);
wire s0n16430,s1n16430,notn16430;
or (n16430,s0n16430,s1n16430);
not(notn16430,n14409);
and (s0n16430,notn16430,n16431);
and (s1n16430,n14409,n16413);
wire s0n16431,s1n16431,notn16431;
or (n16431,s0n16431,s1n16431);
not(notn16431,n14401);
and (s0n16431,notn16431,1'b0);
and (s1n16431,n14401,n16409);
or (n16433,n16434,n16435,n16443,n16444);
and (n16434,n16323,n13907);
and (n16435,n16436,n14385);
wire s0n16436,s1n16436,notn16436;
or (n16436,s0n16436,s1n16436);
not(notn16436,n2799);
and (s0n16436,notn16436,1'b0);
and (s1n16436,n2799,n16437);
or (n16437,1'b0,n16438,n16439);
and (n16438,n16325,n13900);
and (n16439,n16440,n14131);
wire s0n16440,s1n16440,notn16440;
or (n16440,s0n16440,s1n16440);
not(notn16440,n14573);
and (s0n16440,notn16440,n16441);
and (s1n16440,n14573,1'b0);
wire s0n16441,s1n16441,notn16441;
or (n16441,s0n16441,s1n16441);
not(notn16441,n14374);
and (s0n16441,notn16441,1'b0);
and (s1n16441,n14374,n16442);
and (n16443,n16402,n14381);
and (n16444,n16336,n14192);
or (n16445,1'b0,n16446,n16451,n16466,n16534,n16565,n16571,n16579,n16580);
and (n16446,n16447,n14237);
or (n16447,1'b0,n16448,n16450);
and (n16448,n16449,n14235);
wire s0n16450,s1n16450,notn16450;
or (n16450,s0n16450,s1n16450);
not(notn16450,n14455);
and (s0n16450,notn16450,1'b0);
and (s1n16450,n14455,n16402);
and (n16451,n16452,n14137);
or (n16452,1'b0,n16453,n16464,n16465);
and (n16453,n16454,n13889);
wire s0n16454,s1n16454,notn16454;
or (n16454,s0n16454,s1n16454);
not(notn16454,n14227);
and (s0n16454,notn16454,1'b0);
and (s1n16454,n14227,n16455);
or (n16455,1'b0,n16456,n16457,n16458,n16459,n16460,n16463);
and (n16456,n16338,n14193);
and (n16457,n16380,n14199);
and (n16458,n16382,n2781);
and (n16459,n16375,n14205);
and (n16460,n16461,n2789);
wire s0n16461,s1n16461,notn16461;
or (n16461,s0n16461,s1n16461);
not(notn16461,n14210);
and (s0n16461,notn16461,n16348);
and (s1n16461,n14210,n16462);
and (n16463,n16462,n14225);
and (n16464,n16338,n14243);
and (n16465,n16370,n14131);
and (n16466,n16467,n14111);
or (n16467,1'b0,n16468,n16470,n16472,n16502);
and (n16468,n16469,n13889);
and (n16470,n16471,n13897);
and (n16472,n16473,n13900);
wire s0n16473,s1n16473,notn16473;
or (n16473,s0n16473,s1n16473);
not(notn16473,n42);
and (s0n16473,notn16473,1'b0);
and (s1n16473,n42,n16474);
wire s0n16474,s1n16474,notn16474;
or (n16474,s0n16474,s1n16474);
not(notn16474,n14422);
and (s0n16474,notn16474,n16475);
and (s1n16474,n14422,n16485);
wire s0n16475,s1n16475,notn16475;
or (n16475,s0n16475,s1n16475);
not(notn16475,n14362);
and (s0n16475,notn16475,1'b0);
and (s1n16475,n14362,n16476);
or (n16476,1'b0,n16477,n16479,n16481,n16483);
and (n16477,n16478,n14352);
and (n16479,n16480,n14355);
and (n16481,n16482,n14358);
and (n16483,n16484,n14361);
or (n16485,1'b0,n16486,n16489,n16490,n16496);
and (n16486,n16487,n14387);
wire s0n16487,s1n16487,notn16487;
or (n16487,s0n16487,s1n16487);
not(notn16487,n14374);
and (s0n16487,notn16487,1'b0);
and (s1n16487,n14374,n16488);
and (n16489,n16441,n14393);
and (n16490,n16491,n14412);
wire s0n16491,s1n16491,notn16491;
or (n16491,s0n16491,s1n16491);
not(notn16491,n42);
and (s0n16491,notn16491,1'b0);
and (s1n16491,n42,n16492);
wire s0n16492,s1n16492,notn16492;
or (n16492,s0n16492,s1n16492);
not(notn16492,n14375);
and (s0n16492,notn16492,n16493);
and (s1n16492,n14375,n16495);
wire s0n16493,s1n16493,notn16493;
or (n16493,s0n16493,s1n16493);
not(notn16493,n14409);
and (s0n16493,notn16493,n16494);
and (s1n16493,n14409,n16482);
wire s0n16494,s1n16494,notn16494;
or (n16494,s0n16494,s1n16494);
not(notn16494,n14401);
and (s0n16494,notn16494,1'b0);
and (s1n16494,n14401,n16478);
and (n16496,n16497,n14421);
wire s0n16497,s1n16497,notn16497;
or (n16497,s0n16497,s1n16497);
not(notn16497,n42);
and (s0n16497,notn16497,1'b0);
and (s1n16497,n42,n16498);
wire s0n16498,s1n16498,notn16498;
or (n16498,s0n16498,s1n16498);
not(notn16498,n14375);
and (s0n16498,notn16498,n16499);
and (s1n16498,n14375,n16501);
wire s0n16499,s1n16499,notn16499;
or (n16499,s0n16499,s1n16499);
not(notn16499,n14409);
and (s0n16499,notn16499,n16500);
and (s1n16499,n14409,n16484);
wire s0n16500,s1n16500,notn16500;
or (n16500,s0n16500,s1n16500);
not(notn16500,n14401);
and (s0n16500,notn16500,1'b0);
and (s1n16500,n14401,n16480);
wire s0n16502,s1n16502,notn16502;
or (n16502,s0n16502,s1n16502);
not(notn16502,n14131);
and (s0n16502,notn16502,1'b0);
and (s1n16502,n14131,n16503);
wire s0n16503,s1n16503,notn16503;
or (n16503,s0n16503,s1n16503);
not(notn16503,n42);
and (s0n16503,notn16503,1'b0);
and (s1n16503,n42,n16504);
wire s0n16504,s1n16504,notn16504;
or (n16504,s0n16504,s1n16504);
not(notn16504,n14422);
and (s0n16504,notn16504,n16505);
and (s1n16504,n14422,n16515);
wire s0n16505,s1n16505,notn16505;
or (n16505,s0n16505,s1n16505);
not(notn16505,n14362);
and (s0n16505,notn16505,1'b0);
and (s1n16505,n14362,n16506);
or (n16506,1'b0,n16507,n16509,n16511,n16513);
and (n16507,n16508,n14352);
and (n16509,n16510,n14355);
and (n16511,n16512,n14358);
and (n16513,n16514,n14361);
or (n16515,1'b0,n16516,n16519,n16522,n16528);
and (n16516,n16517,n14387);
wire s0n16517,s1n16517,notn16517;
or (n16517,s0n16517,s1n16517);
not(notn16517,n14374);
and (s0n16517,notn16517,1'b0);
and (s1n16517,n14374,n16518);
and (n16519,n16520,n14393);
wire s0n16520,s1n16520,notn16520;
or (n16520,s0n16520,s1n16520);
not(notn16520,n14374);
and (s0n16520,notn16520,1'b0);
and (s1n16520,n14374,n16521);
and (n16522,n16523,n14412);
wire s0n16523,s1n16523,notn16523;
or (n16523,s0n16523,s1n16523);
not(notn16523,n42);
and (s0n16523,notn16523,1'b0);
and (s1n16523,n42,n16524);
wire s0n16524,s1n16524,notn16524;
or (n16524,s0n16524,s1n16524);
not(notn16524,n14375);
and (s0n16524,notn16524,n16525);
and (s1n16524,n14375,n16527);
wire s0n16525,s1n16525,notn16525;
or (n16525,s0n16525,s1n16525);
not(notn16525,n14409);
and (s0n16525,notn16525,n16526);
and (s1n16525,n14409,n16512);
wire s0n16526,s1n16526,notn16526;
or (n16526,s0n16526,s1n16526);
not(notn16526,n14401);
and (s0n16526,notn16526,1'b0);
and (s1n16526,n14401,n16508);
and (n16528,n16529,n14421);
wire s0n16529,s1n16529,notn16529;
or (n16529,s0n16529,s1n16529);
not(notn16529,n42);
and (s0n16529,notn16529,1'b0);
and (s1n16529,n42,n16530);
wire s0n16530,s1n16530,notn16530;
or (n16530,s0n16530,s1n16530);
not(notn16530,n14375);
and (s0n16530,notn16530,n16531);
and (s1n16530,n14375,n16533);
wire s0n16531,s1n16531,notn16531;
or (n16531,s0n16531,s1n16531);
not(notn16531,n14409);
and (s0n16531,notn16531,n16532);
and (s1n16531,n14409,n16514);
wire s0n16532,s1n16532,notn16532;
or (n16532,s0n16532,s1n16532);
not(notn16532,n14401);
and (s0n16532,notn16532,1'b0);
and (s1n16532,n14401,n16510);
not (n16534,n16535);
nand (n16535,n16536,n14108);
or (n16536,1'b0,n16537,n16539,n16541,n16543);
and (n16537,n16538,n13889);
and (n16539,n16540,n13897);
and (n16541,n16542,n13900);
and (n16543,n16544,n14131);
wire s0n16544,s1n16544,notn16544;
or (n16544,s0n16544,s1n16544);
not(notn16544,n14123);
and (s0n16544,notn16544,1'b0);
and (s1n16544,n14123,n16545);
wire s0n16545,s1n16545,notn16545;
or (n16545,s0n16545,s1n16545);
not(notn16545,n555);
and (s0n16545,notn16545,n16546);
and (s1n16545,n555,n16561);
wire s0n16546,s1n16546,notn16546;
or (n16546,s0n16546,s1n16546);
not(notn16546,n13948);
and (s0n16546,notn16546,n16547);
and (s1n16546,n13948,n16549);
wire s0n16547,s1n16547,notn16547;
or (n16547,s0n16547,s1n16547);
not(notn16547,n13907);
and (s0n16547,notn16547,1'b0);
and (s1n16547,n13907,n16548);
or (n16549,n16550,n16552,n16554,n16556,n16558,n16560);
and (n16550,n16551,n13913);
and (n16552,n16553,n13920);
and (n16554,n16555,n13923);
and (n16556,n16557,n13928);
and (n16558,n16559,n13935);
and (n16560,n16548,n13941);
wire s0n16561,s1n16561,notn16561;
or (n16561,s0n16561,s1n16561);
not(notn16561,n14119);
and (s0n16561,notn16561,1'b0);
and (s1n16561,n14119,n16562);
wire s0n16562,s1n16562,notn16562;
or (n16562,s0n16562,s1n16562);
not(notn16562,n14116);
and (s0n16562,notn16562,n16563);
and (s1n16562,n14116,n16564);
and (n16565,n16566,n13950);
or (n16566,1'b0,n16567,n16568,n16569,n16570);
and (n16567,n16540,n13889);
and (n16568,n16542,n13897);
and (n16569,n16471,n13900);
wire s0n16570,s1n16570,notn16570;
or (n16570,s0n16570,s1n16570);
not(notn16570,n14131);
and (s0n16570,notn16570,1'b0);
and (s1n16570,n14131,n16473);
and (n16571,n16572,n14239);
or (n16572,1'b0,n16573,n16575,n16577,n16578);
and (n16573,n16574,n13889);
and (n16575,n16576,n13897);
and (n16577,n16449,n13900);
and (n16578,n16354,n14131);
and (n16579,n16402,n14448);
and (n16580,n16336,n14266);
wire s0n16581,s1n16581,notn16581;
or (n16581,s0n16581,s1n16581);
not(notn16581,n14631);
and (s0n16581,notn16581,n16582);
and (s1n16581,n14631,n16600);
wire s0n16582,s1n16582,notn16582;
or (n16582,s0n16582,s1n16582);
not(notn16582,n14271);
and (s0n16582,notn16582,n16583);
and (s1n16582,n14271,n16588);
wire s0n16583,s1n16583,notn16583;
or (n16583,s0n16583,s1n16583);
not(notn16583,n14279);
and (s0n16583,notn16583,1'b0);
and (s1n16583,n14279,n16584);
and (n16584,n16585,n14120);
wire s0n16585,s1n16585,notn16585;
or (n16585,s0n16585,s1n16585);
not(notn16585,n14125);
and (s0n16585,notn16585,1'b0);
and (s1n16585,n14125,n16586);
wire s0n16586,s1n16586,notn16586;
or (n16586,s0n16586,s1n16586);
not(notn16586,n14317);
and (s0n16586,notn16586,n16587);
and (s1n16586,n14317,n16252);
or (n16588,n16589,n16593,1'b0);
and (n16589,n16590,n13907);
wire s0n16590,s1n16590,notn16590;
or (n16590,s0n16590,s1n16590);
not(notn16590,n14125);
and (s0n16590,notn16590,1'b0);
and (s1n16590,n14125,n16591);
wire s0n16591,s1n16591,notn16591;
or (n16591,s0n16591,s1n16591);
not(notn16591,n14563);
and (s0n16591,notn16591,n16587);
and (s1n16591,n14563,n16592);
and (n16593,n16594,n14385);
wire s0n16594,s1n16594,notn16594;
or (n16594,s0n16594,s1n16594);
not(notn16594,n2799);
and (s0n16594,notn16594,1'b0);
and (s1n16594,n2799,n16595);
or (n16595,1'b0,n16596,n16598);
and (n16596,n16597,n13900);
wire s0n16597,s1n16597,notn16597;
or (n16597,s0n16597,s1n16597);
not(notn16597,n14570);
and (s0n16597,notn16597,n16382);
and (s1n16597,n14570,1'b0);
and (n16598,n16599,n14131);
wire s0n16599,s1n16599,notn16599;
or (n16599,s0n16599,s1n16599);
not(notn16599,n14573);
and (s0n16599,notn16599,n16520);
and (s1n16599,n14573,1'b0);
or (n16600,n16601,n16665,n16678,n16679,n16680,n16682,1'b0);
not (n16601,n16602);
or (n16602,n16603,n16664);
not (n16603,n16604);
nand (n16604,n16605,n16617,n16628,n16639);
nand (n16605,n16606,n16613);
wire s0n16606,s1n16606,notn16606;
or (n16606,s0n16606,s1n16606);
not(notn16606,n42);
and (s0n16606,notn16606,1'b0);
and (s1n16606,n42,n16607);
wire s0n16607,s1n16607,notn16607;
or (n16607,s0n16607,s1n16607);
not(notn16607,n14375);
and (s0n16607,notn16607,n16608);
and (s1n16607,n14375,n16612);
wire s0n16608,s1n16608,notn16608;
or (n16608,s0n16608,s1n16608);
not(notn16608,n14409);
and (s0n16608,notn16608,n16609);
and (s1n16608,n14409,n16611);
wire s0n16609,s1n16609,notn16609;
or (n16609,s0n16609,s1n16609);
not(notn16609,n14401);
and (s0n16609,notn16609,1'b0);
and (s1n16609,n14401,n16610);
nor (n16613,n16614,n16616);
nand (n16614,n14423,n16615);
not (n16615,n14230);
not (n16616,n14499);
nand (n16617,n16618,n16625);
wire s0n16618,s1n16618,notn16618;
or (n16618,s0n16618,s1n16618);
not(notn16618,n42);
and (s0n16618,notn16618,1'b0);
and (s1n16618,n42,n16619);
wire s0n16619,s1n16619,notn16619;
or (n16619,s0n16619,s1n16619);
not(notn16619,n14375);
and (s0n16619,notn16619,n16620);
and (s1n16619,n14375,n16624);
wire s0n16620,s1n16620,notn16620;
or (n16620,s0n16620,s1n16620);
not(notn16620,n14409);
and (s0n16620,notn16620,n16621);
and (s1n16620,n14409,n16623);
wire s0n16621,s1n16621,notn16621;
or (n16621,s0n16621,s1n16621);
not(notn16621,n14401);
and (s0n16621,notn16621,1'b0);
and (s1n16621,n14401,n16622);
nor (n16625,n16614,n16626);
nand (n16626,n29,n16627);
not (n16627,n582);
nor (n16628,n16629,n16634);
and (n16629,n16630,n16632);
wire s0n16630,s1n16630,notn16630;
or (n16630,s0n16630,s1n16630);
not(notn16630,n14374);
and (s0n16630,notn16630,1'b0);
and (s1n16630,n14374,n16631);
nor (n16632,n16614,n16633);
nand (n16633,n582,n2773);
and (n16634,n16635,n16637);
wire s0n16635,s1n16635,notn16635;
or (n16635,s0n16635,s1n16635);
not(notn16635,n14374);
and (s0n16635,notn16635,1'b0);
and (s1n16635,n14374,n16636);
nor (n16637,n16614,n16638);
nand (n16638,n29,n582);
and (n16639,n16640,n16655);
nor (n16640,n16641,n16650);
and (n16641,n16642,n16623);
not (n16642,n16643);
nand (n16643,n16644,n16649);
nor (n16644,n16645,n16646);
not (n16645,n14364);
nand (n16646,n16647,n585);
not (n16647,n16648);
nand (n16648,n42,n14363);
not (n16649,n16626);
and (n16650,n16651,n16610);
not (n16651,n16652);
nand (n16652,n16653,n16654);
nor (n16653,n16645,n16648);
nor (n16654,n16616,n585);
nor (n16655,n16656,n16659);
and (n16656,n16657,n16611);
not (n16657,n16658);
nand (n16658,n16644,n14499);
and (n16659,n16660,n16622);
not (n16660,n16661);
nand (n16661,n16653,n16662);
and (n16662,n16663,n16627);
nor (n16663,n2773,n585);
not (n16664,n14453);
and (n16665,n16666,n14137);
or (n16666,1'b0,n16667,n16677);
and (n16667,n16668,n14235);
wire s0n16668,s1n16668,notn16668;
or (n16668,s0n16668,s1n16668);
not(notn16668,n14227);
and (s0n16668,notn16668,1'b0);
and (s1n16668,n14227,n16669);
or (n16669,1'b0,n16456,n16670,n16671,n16672,n16673,n16676);
and (n16670,n16396,n14199);
and (n16671,n16398,n2781);
and (n16672,n16391,n14205);
and (n16673,n16674,n2789);
wire s0n16674,s1n16674,notn16674;
or (n16674,s0n16674,s1n16674);
not(notn16674,n14210);
and (s0n16674,notn16674,n16348);
and (s1n16674,n14210,n16675);
and (n16676,n16675,n14225);
and (n16677,n16354,n14455);
and (n16678,n16450,n14111);
and (n16679,n16502,n14108);
and (n16680,n16681,n13950);
wire s0n16681,s1n16681,notn16681;
or (n16681,s0n16681,s1n16681);
not(notn16681,n14131);
and (s0n16681,notn16681,1'b0);
and (s1n16681,n14131,n16402);
and (n16682,n16683,n14239);
wire s0n16683,s1n16683,notn16683;
or (n16683,s0n16683,s1n16683);
not(notn16683,n14131);
and (s0n16683,notn16683,1'b0);
and (s1n16683,n14131,n16668);
and (n16684,n16581,n16685);
and (n16685,n16686,n16949);
wire s0n16686,s1n16686,notn16686;
or (n16686,s0n16686,s1n16686);
not(notn16686,n14631);
and (s0n16686,notn16686,n16687);
and (s1n16686,n14631,n16813);
wire s0n16687,s1n16687,notn16687;
or (n16687,s0n16687,s1n16687);
not(notn16687,n14271);
and (s0n16687,notn16687,n16688);
and (s1n16687,n14271,n16801);
wire s0n16688,s1n16688,notn16688;
or (n16688,s0n16688,s1n16688);
not(notn16688,n14279);
and (s0n16688,notn16688,1'b0);
and (s1n16688,n14279,n16689);
or (n16689,1'b0,n16690,n16703,n16769);
and (n16690,n16691,n14120);
wire s0n16691,s1n16691,notn16691;
or (n16691,s0n16691,s1n16691);
not(notn16691,n14125);
and (s0n16691,notn16691,1'b0);
and (s1n16691,n14125,n16692);
wire s0n16692,s1n16692,notn16692;
or (n16692,s0n16692,s1n16692);
not(notn16692,n14317);
and (s0n16692,notn16692,n16693);
and (s1n16692,n14317,n16694);
wire s0n16694,s1n16694,notn16694;
or (n16694,s0n16694,s1n16694);
not(notn16694,n14326);
and (s0n16694,notn16694,n16695);
and (s1n16694,n14326,n16697);
wire s0n16695,s1n16695,notn16695;
or (n16695,s0n16695,s1n16695);
not(notn16695,n14315);
and (s0n16695,notn16695,1'b0);
and (s1n16695,n14315,n16696);
or (n16697,1'b0,n16698,n16700,n16702);
and (n16698,n16699,n14321);
and (n16700,n16701,n14324);
and (n16702,n16696,n14184);
and (n16703,n16704,n14718);
or (n16704,1'b0,n16705,n16721,n16737,n16753);
and (n16705,n16706,n13889);
wire s0n16706,s1n16706,notn16706;
or (n16706,s0n16706,s1n16706);
not(notn16706,n42);
and (s0n16706,notn16706,1'b0);
and (s1n16706,n42,n16707);
wire s0n16707,s1n16707,notn16707;
or (n16707,s0n16707,s1n16707);
not(notn16707,n14187);
and (s0n16707,notn16707,n16708);
and (s1n16707,n14187,n16714);
wire s0n16708,s1n16708,notn16708;
or (n16708,s0n16708,s1n16708);
not(notn16708,n14163);
and (s0n16708,notn16708,1'b0);
and (s1n16708,n14163,n16709);
or (n16709,1'b0,n16710,n16712);
and (n16710,n16711,n14147);
and (n16712,n16713,n14156);
or (n16714,1'b0,n16715,n16717,n16719,n16720);
and (n16715,n16716,n14171);
and (n16717,n16718,n14176);
and (n16719,n16711,n14180);
and (n16720,n16713,n14184);
and (n16721,n16722,n13897);
wire s0n16722,s1n16722,notn16722;
or (n16722,s0n16722,s1n16722);
not(notn16722,n42);
and (s0n16722,notn16722,1'b0);
and (s1n16722,n42,n16723);
wire s0n16723,s1n16723,notn16723;
or (n16723,s0n16723,s1n16723);
not(notn16723,n14187);
and (s0n16723,notn16723,n16724);
and (s1n16723,n14187,n16730);
wire s0n16724,s1n16724,notn16724;
or (n16724,s0n16724,s1n16724);
not(notn16724,n14163);
and (s0n16724,notn16724,1'b0);
and (s1n16724,n14163,n16725);
or (n16725,1'b0,n16726,n16728);
and (n16726,n16727,n14147);
and (n16728,n16729,n14156);
or (n16730,1'b0,n16731,n16733,n16735,n16736);
and (n16731,n16732,n14171);
and (n16733,n16734,n14176);
and (n16735,n16727,n14180);
and (n16736,n16729,n14184);
and (n16737,n16738,n13900);
wire s0n16738,s1n16738,notn16738;
or (n16738,s0n16738,s1n16738);
not(notn16738,n42);
and (s0n16738,notn16738,1'b0);
and (s1n16738,n42,n16739);
wire s0n16739,s1n16739,notn16739;
or (n16739,s0n16739,s1n16739);
not(notn16739,n14187);
and (s0n16739,notn16739,n16740);
and (s1n16739,n14187,n16746);
wire s0n16740,s1n16740,notn16740;
or (n16740,s0n16740,s1n16740);
not(notn16740,n14163);
and (s0n16740,notn16740,1'b0);
and (s1n16740,n14163,n16741);
or (n16741,1'b0,n16742,n16744);
and (n16742,n16743,n14147);
and (n16744,n16745,n14156);
or (n16746,1'b0,n16747,n16749,n16751,n16752);
and (n16747,n16748,n14171);
and (n16749,n16750,n14176);
and (n16751,n16743,n14180);
and (n16752,n16745,n14184);
and (n16753,n16754,n14131);
wire s0n16754,s1n16754,notn16754;
or (n16754,s0n16754,s1n16754);
not(notn16754,n42);
and (s0n16754,notn16754,1'b0);
and (s1n16754,n42,n16755);
wire s0n16755,s1n16755,notn16755;
or (n16755,s0n16755,s1n16755);
not(notn16755,n14187);
and (s0n16755,notn16755,n16756);
and (s1n16755,n14187,n16762);
wire s0n16756,s1n16756,notn16756;
or (n16756,s0n16756,s1n16756);
not(notn16756,n14163);
and (s0n16756,notn16756,1'b0);
and (s1n16756,n14163,n16757);
or (n16757,1'b0,n16758,n16760);
and (n16758,n16759,n14147);
and (n16760,n16761,n14156);
or (n16762,1'b0,n16763,n16765,n16767,n16768);
and (n16763,n16764,n14171);
and (n16765,n16766,n14176);
and (n16767,n16759,n14180);
and (n16768,n16761,n14184);
and (n16769,n16770,n14365);
wire s0n16770,s1n16770,notn16770;
or (n16770,s0n16770,s1n16770);
not(notn16770,n42);
and (s0n16770,notn16770,1'b0);
and (s1n16770,n42,n16771);
wire s0n16771,s1n16771,notn16771;
or (n16771,s0n16771,s1n16771);
not(notn16771,n14422);
and (s0n16771,notn16771,n16772);
and (s1n16771,n14422,n16782);
wire s0n16772,s1n16772,notn16772;
or (n16772,s0n16772,s1n16772);
not(notn16772,n14362);
and (s0n16772,notn16772,1'b0);
and (s1n16772,n14362,n16773);
or (n16773,1'b0,n16774,n16776,n16778,n16780);
and (n16774,n16775,n14352);
and (n16776,n16777,n14355);
and (n16778,n16779,n14358);
and (n16780,n16781,n14361);
or (n16782,1'b0,n16783,n16786,n16789,n16795);
and (n16783,n16784,n14387);
wire s0n16784,s1n16784,notn16784;
or (n16784,s0n16784,s1n16784);
not(notn16784,n14374);
and (s0n16784,notn16784,1'b0);
and (s1n16784,n14374,n16785);
and (n16786,n16787,n14393);
wire s0n16787,s1n16787,notn16787;
or (n16787,s0n16787,s1n16787);
not(notn16787,n14374);
and (s0n16787,notn16787,1'b0);
and (s1n16787,n14374,n16788);
and (n16789,n16790,n14412);
wire s0n16790,s1n16790,notn16790;
or (n16790,s0n16790,s1n16790);
not(notn16790,n42);
and (s0n16790,notn16790,1'b0);
and (s1n16790,n42,n16791);
wire s0n16791,s1n16791,notn16791;
or (n16791,s0n16791,s1n16791);
not(notn16791,n14375);
and (s0n16791,notn16791,n16792);
and (s1n16791,n14375,n16794);
wire s0n16792,s1n16792,notn16792;
or (n16792,s0n16792,s1n16792);
not(notn16792,n14409);
and (s0n16792,notn16792,n16793);
and (s1n16792,n14409,n16779);
wire s0n16793,s1n16793,notn16793;
or (n16793,s0n16793,s1n16793);
not(notn16793,n14401);
and (s0n16793,notn16793,1'b0);
and (s1n16793,n14401,n16775);
and (n16795,n16796,n14421);
wire s0n16796,s1n16796,notn16796;
or (n16796,s0n16796,s1n16796);
not(notn16796,n42);
and (s0n16796,notn16796,1'b0);
and (s1n16796,n42,n16797);
wire s0n16797,s1n16797,notn16797;
or (n16797,s0n16797,s1n16797);
not(notn16797,n14375);
and (s0n16797,notn16797,n16798);
and (s1n16797,n14375,n16800);
wire s0n16798,s1n16798,notn16798;
or (n16798,s0n16798,s1n16798);
not(notn16798,n14409);
and (s0n16798,notn16798,n16799);
and (s1n16798,n14409,n16781);
wire s0n16799,s1n16799,notn16799;
or (n16799,s0n16799,s1n16799);
not(notn16799,n14401);
and (s0n16799,notn16799,1'b0);
and (s1n16799,n14401,n16777);
or (n16801,n16802,n16803,n16811,n16812);
and (n16802,n16691,n13907);
and (n16803,n16804,n14385);
wire s0n16804,s1n16804,notn16804;
or (n16804,s0n16804,s1n16804);
not(notn16804,n2799);
and (s0n16804,notn16804,1'b0);
and (s1n16804,n2799,n16805);
or (n16805,1'b0,n16806,n16807);
and (n16806,n16693,n13900);
and (n16807,n16808,n14131);
wire s0n16808,s1n16808,notn16808;
or (n16808,s0n16808,s1n16808);
not(notn16808,n14573);
and (s0n16808,notn16808,n16809);
and (s1n16808,n14573,1'b0);
wire s0n16809,s1n16809,notn16809;
or (n16809,s0n16809,s1n16809);
not(notn16809,n14374);
and (s0n16809,notn16809,1'b0);
and (s1n16809,n14374,n16810);
and (n16811,n16770,n14381);
and (n16812,n16704,n14192);
or (n16813,1'b0,n16814,n16819,n16834,n16902,n16933,n16939,n16947,n16948);
and (n16814,n16815,n14237);
or (n16815,1'b0,n16816,n16818);
and (n16816,n16817,n14235);
wire s0n16818,s1n16818,notn16818;
or (n16818,s0n16818,s1n16818);
not(notn16818,n14455);
and (s0n16818,notn16818,1'b0);
and (s1n16818,n14455,n16770);
and (n16819,n16820,n14137);
or (n16820,1'b0,n16821,n16832,n16833);
and (n16821,n16822,n13889);
wire s0n16822,s1n16822,notn16822;
or (n16822,s0n16822,s1n16822);
not(notn16822,n14227);
and (s0n16822,notn16822,1'b0);
and (s1n16822,n14227,n16823);
or (n16823,1'b0,n16824,n16825,n16826,n16827,n16828,n16831);
and (n16824,n16706,n14193);
and (n16825,n16748,n14199);
and (n16826,n16750,n2781);
and (n16827,n16743,n14205);
and (n16828,n16829,n2789);
wire s0n16829,s1n16829,notn16829;
or (n16829,s0n16829,s1n16829);
not(notn16829,n14210);
and (s0n16829,notn16829,n16716);
and (s1n16829,n14210,n16830);
and (n16831,n16830,n14225);
and (n16832,n16706,n14243);
and (n16833,n16738,n14131);
and (n16834,n16835,n14111);
or (n16835,1'b0,n16836,n16838,n16840,n16870);
and (n16836,n16837,n13889);
and (n16838,n16839,n13897);
and (n16840,n16841,n13900);
wire s0n16841,s1n16841,notn16841;
or (n16841,s0n16841,s1n16841);
not(notn16841,n42);
and (s0n16841,notn16841,1'b0);
and (s1n16841,n42,n16842);
wire s0n16842,s1n16842,notn16842;
or (n16842,s0n16842,s1n16842);
not(notn16842,n14422);
and (s0n16842,notn16842,n16843);
and (s1n16842,n14422,n16853);
wire s0n16843,s1n16843,notn16843;
or (n16843,s0n16843,s1n16843);
not(notn16843,n14362);
and (s0n16843,notn16843,1'b0);
and (s1n16843,n14362,n16844);
or (n16844,1'b0,n16845,n16847,n16849,n16851);
and (n16845,n16846,n14352);
and (n16847,n16848,n14355);
and (n16849,n16850,n14358);
and (n16851,n16852,n14361);
or (n16853,1'b0,n16854,n16857,n16858,n16864);
and (n16854,n16855,n14387);
wire s0n16855,s1n16855,notn16855;
or (n16855,s0n16855,s1n16855);
not(notn16855,n14374);
and (s0n16855,notn16855,1'b0);
and (s1n16855,n14374,n16856);
and (n16857,n16809,n14393);
and (n16858,n16859,n14412);
wire s0n16859,s1n16859,notn16859;
or (n16859,s0n16859,s1n16859);
not(notn16859,n42);
and (s0n16859,notn16859,1'b0);
and (s1n16859,n42,n16860);
wire s0n16860,s1n16860,notn16860;
or (n16860,s0n16860,s1n16860);
not(notn16860,n14375);
and (s0n16860,notn16860,n16861);
and (s1n16860,n14375,n16863);
wire s0n16861,s1n16861,notn16861;
or (n16861,s0n16861,s1n16861);
not(notn16861,n14409);
and (s0n16861,notn16861,n16862);
and (s1n16861,n14409,n16850);
wire s0n16862,s1n16862,notn16862;
or (n16862,s0n16862,s1n16862);
not(notn16862,n14401);
and (s0n16862,notn16862,1'b0);
and (s1n16862,n14401,n16846);
and (n16864,n16865,n14421);
wire s0n16865,s1n16865,notn16865;
or (n16865,s0n16865,s1n16865);
not(notn16865,n42);
and (s0n16865,notn16865,1'b0);
and (s1n16865,n42,n16866);
wire s0n16866,s1n16866,notn16866;
or (n16866,s0n16866,s1n16866);
not(notn16866,n14375);
and (s0n16866,notn16866,n16867);
and (s1n16866,n14375,n16869);
wire s0n16867,s1n16867,notn16867;
or (n16867,s0n16867,s1n16867);
not(notn16867,n14409);
and (s0n16867,notn16867,n16868);
and (s1n16867,n14409,n16852);
wire s0n16868,s1n16868,notn16868;
or (n16868,s0n16868,s1n16868);
not(notn16868,n14401);
and (s0n16868,notn16868,1'b0);
and (s1n16868,n14401,n16848);
wire s0n16870,s1n16870,notn16870;
or (n16870,s0n16870,s1n16870);
not(notn16870,n14131);
and (s0n16870,notn16870,1'b0);
and (s1n16870,n14131,n16871);
wire s0n16871,s1n16871,notn16871;
or (n16871,s0n16871,s1n16871);
not(notn16871,n42);
and (s0n16871,notn16871,1'b0);
and (s1n16871,n42,n16872);
wire s0n16872,s1n16872,notn16872;
or (n16872,s0n16872,s1n16872);
not(notn16872,n14422);
and (s0n16872,notn16872,n16873);
and (s1n16872,n14422,n16883);
wire s0n16873,s1n16873,notn16873;
or (n16873,s0n16873,s1n16873);
not(notn16873,n14362);
and (s0n16873,notn16873,1'b0);
and (s1n16873,n14362,n16874);
or (n16874,1'b0,n16875,n16877,n16879,n16881);
and (n16875,n16876,n14352);
and (n16877,n16878,n14355);
and (n16879,n16880,n14358);
and (n16881,n16882,n14361);
or (n16883,1'b0,n16884,n16887,n16890,n16896);
and (n16884,n16885,n14387);
wire s0n16885,s1n16885,notn16885;
or (n16885,s0n16885,s1n16885);
not(notn16885,n14374);
and (s0n16885,notn16885,1'b0);
and (s1n16885,n14374,n16886);
and (n16887,n16888,n14393);
wire s0n16888,s1n16888,notn16888;
or (n16888,s0n16888,s1n16888);
not(notn16888,n14374);
and (s0n16888,notn16888,1'b0);
and (s1n16888,n14374,n16889);
and (n16890,n16891,n14412);
wire s0n16891,s1n16891,notn16891;
or (n16891,s0n16891,s1n16891);
not(notn16891,n42);
and (s0n16891,notn16891,1'b0);
and (s1n16891,n42,n16892);
wire s0n16892,s1n16892,notn16892;
or (n16892,s0n16892,s1n16892);
not(notn16892,n14375);
and (s0n16892,notn16892,n16893);
and (s1n16892,n14375,n16895);
wire s0n16893,s1n16893,notn16893;
or (n16893,s0n16893,s1n16893);
not(notn16893,n14409);
and (s0n16893,notn16893,n16894);
and (s1n16893,n14409,n16880);
wire s0n16894,s1n16894,notn16894;
or (n16894,s0n16894,s1n16894);
not(notn16894,n14401);
and (s0n16894,notn16894,1'b0);
and (s1n16894,n14401,n16876);
and (n16896,n16897,n14421);
wire s0n16897,s1n16897,notn16897;
or (n16897,s0n16897,s1n16897);
not(notn16897,n42);
and (s0n16897,notn16897,1'b0);
and (s1n16897,n42,n16898);
wire s0n16898,s1n16898,notn16898;
or (n16898,s0n16898,s1n16898);
not(notn16898,n14375);
and (s0n16898,notn16898,n16899);
and (s1n16898,n14375,n16901);
wire s0n16899,s1n16899,notn16899;
or (n16899,s0n16899,s1n16899);
not(notn16899,n14409);
and (s0n16899,notn16899,n16900);
and (s1n16899,n14409,n16882);
wire s0n16900,s1n16900,notn16900;
or (n16900,s0n16900,s1n16900);
not(notn16900,n14401);
and (s0n16900,notn16900,1'b0);
and (s1n16900,n14401,n16878);
not (n16902,n16903);
nand (n16903,n16904,n14108);
or (n16904,1'b0,n16905,n16907,n16909,n16911);
and (n16905,n16906,n13889);
and (n16907,n16908,n13897);
and (n16909,n16910,n13900);
and (n16911,n16912,n14131);
wire s0n16912,s1n16912,notn16912;
or (n16912,s0n16912,s1n16912);
not(notn16912,n14123);
and (s0n16912,notn16912,1'b0);
and (s1n16912,n14123,n16913);
wire s0n16913,s1n16913,notn16913;
or (n16913,s0n16913,s1n16913);
not(notn16913,n555);
and (s0n16913,notn16913,n16914);
and (s1n16913,n555,n16929);
wire s0n16914,s1n16914,notn16914;
or (n16914,s0n16914,s1n16914);
not(notn16914,n13948);
and (s0n16914,notn16914,n16915);
and (s1n16914,n13948,n16917);
wire s0n16915,s1n16915,notn16915;
or (n16915,s0n16915,s1n16915);
not(notn16915,n13907);
and (s0n16915,notn16915,1'b0);
and (s1n16915,n13907,n16916);
or (n16917,n16918,n16920,n16922,n16924,n16926,n16928);
and (n16918,n16919,n13913);
and (n16920,n16921,n13920);
and (n16922,n16923,n13923);
and (n16924,n16925,n13928);
and (n16926,n16927,n13935);
and (n16928,n16916,n13941);
wire s0n16929,s1n16929,notn16929;
or (n16929,s0n16929,s1n16929);
not(notn16929,n14119);
and (s0n16929,notn16929,1'b0);
and (s1n16929,n14119,n16930);
wire s0n16930,s1n16930,notn16930;
or (n16930,s0n16930,s1n16930);
not(notn16930,n14116);
and (s0n16930,notn16930,n16931);
and (s1n16930,n14116,n16932);
and (n16933,n16934,n13950);
or (n16934,1'b0,n16935,n16936,n16937,n16938);
and (n16935,n16908,n13889);
and (n16936,n16910,n13897);
and (n16937,n16839,n13900);
wire s0n16938,s1n16938,notn16938;
or (n16938,s0n16938,s1n16938);
not(notn16938,n14131);
and (s0n16938,notn16938,1'b0);
and (s1n16938,n14131,n16841);
and (n16939,n16940,n14239);
or (n16940,1'b0,n16941,n16943,n16945,n16946);
and (n16941,n16942,n13889);
and (n16943,n16944,n13897);
and (n16945,n16817,n13900);
and (n16946,n16722,n14131);
and (n16947,n16770,n14448);
and (n16948,n16704,n14266);
wire s0n16949,s1n16949,notn16949;
or (n16949,s0n16949,s1n16949);
not(notn16949,n14631);
and (s0n16949,notn16949,n16950);
and (s1n16949,n14631,n16967);
wire s0n16950,s1n16950,notn16950;
or (n16950,s0n16950,s1n16950);
not(notn16950,n14271);
and (s0n16950,notn16950,n16951);
and (s1n16950,n14271,n16956);
wire s0n16951,s1n16951,notn16951;
or (n16951,s0n16951,s1n16951);
not(notn16951,n14279);
and (s0n16951,notn16951,1'b0);
and (s1n16951,n14279,n16952);
and (n16952,n16953,n14120);
wire s0n16953,s1n16953,notn16953;
or (n16953,s0n16953,s1n16953);
not(notn16953,n14125);
and (s0n16953,notn16953,1'b0);
and (s1n16953,n14125,n16954);
wire s0n16954,s1n16954,notn16954;
or (n16954,s0n16954,s1n16954);
not(notn16954,n14317);
and (s0n16954,notn16954,n16955);
and (s1n16954,n14317,n16592);
or (n16956,n16957,n16960,1'b0);
and (n16957,n16958,n13907);
wire s0n16958,s1n16958,notn16958;
or (n16958,s0n16958,s1n16958);
not(notn16958,n14125);
and (s0n16958,notn16958,1'b0);
and (s1n16958,n14125,n16959);
wire s0n16959,s1n16959,notn16959;
or (n16959,s0n16959,s1n16959);
not(notn16959,n14563);
and (s0n16959,notn16959,n16955);
and (s1n16959,n14563,1'b0);
and (n16960,n16961,n14385);
wire s0n16961,s1n16961,notn16961;
or (n16961,s0n16961,s1n16961);
not(notn16961,n2799);
and (s0n16961,notn16961,1'b0);
and (s1n16961,n2799,n16962);
or (n16962,1'b0,n16963,n16965);
and (n16963,n16964,n13900);
wire s0n16964,s1n16964,notn16964;
or (n16964,s0n16964,s1n16964);
not(notn16964,n14570);
and (s0n16964,notn16964,n16750);
and (s1n16964,n14570,1'b0);
and (n16965,n16966,n14131);
wire s0n16966,s1n16966,notn16966;
or (n16966,s0n16966,s1n16966);
not(notn16966,n14573);
and (s0n16966,notn16966,n16888);
and (s1n16966,n14573,1'b0);
or (n16967,n16968,n17001,n17014,n17015,n17018,n17020,1'b0);
and (n16968,n16969,n14237);
wire s0n16969,s1n16969,notn16969;
or (n16969,s0n16969,s1n16969);
not(notn16969,n14455);
and (s0n16969,notn16969,1'b0);
and (s1n16969,n14455,n16970);
wire s0n16970,s1n16970,notn16970;
or (n16970,s0n16970,s1n16970);
not(notn16970,n42);
and (s0n16970,notn16970,1'b0);
and (s1n16970,n42,n16971);
wire s0n16971,s1n16971,notn16971;
or (n16971,s0n16971,s1n16971);
not(notn16971,n14422);
and (s0n16971,notn16971,n16972);
and (s1n16971,n14422,n16982);
wire s0n16972,s1n16972,notn16972;
or (n16972,s0n16972,s1n16972);
not(notn16972,n14362);
and (s0n16972,notn16972,1'b0);
and (s1n16972,n14362,n16973);
or (n16973,1'b0,n16974,n16976,n16978,n16980);
and (n16974,n16975,n14352);
and (n16976,n16977,n14355);
and (n16978,n16979,n14358);
and (n16980,n16981,n14361);
or (n16982,1'b0,n16983,n16986,n16989,n16995);
and (n16983,n16984,n14387);
wire s0n16984,s1n16984,notn16984;
or (n16984,s0n16984,s1n16984);
not(notn16984,n14374);
and (s0n16984,notn16984,1'b0);
and (s1n16984,n14374,n16985);
and (n16986,n16987,n14393);
wire s0n16987,s1n16987,notn16987;
or (n16987,s0n16987,s1n16987);
not(notn16987,n14374);
and (s0n16987,notn16987,1'b0);
and (s1n16987,n14374,n16988);
and (n16989,n16990,n14412);
wire s0n16990,s1n16990,notn16990;
or (n16990,s0n16990,s1n16990);
not(notn16990,n42);
and (s0n16990,notn16990,1'b0);
and (s1n16990,n42,n16991);
wire s0n16991,s1n16991,notn16991;
or (n16991,s0n16991,s1n16991);
not(notn16991,n14375);
and (s0n16991,notn16991,n16992);
and (s1n16991,n14375,n16994);
wire s0n16992,s1n16992,notn16992;
or (n16992,s0n16992,s1n16992);
not(notn16992,n14409);
and (s0n16992,notn16992,n16993);
and (s1n16992,n14409,n16979);
wire s0n16993,s1n16993,notn16993;
or (n16993,s0n16993,s1n16993);
not(notn16993,n14401);
and (s0n16993,notn16993,1'b0);
and (s1n16993,n14401,n16975);
and (n16995,n16996,n14421);
wire s0n16996,s1n16996,notn16996;
or (n16996,s0n16996,s1n16996);
not(notn16996,n42);
and (s0n16996,notn16996,1'b0);
and (s1n16996,n42,n16997);
wire s0n16997,s1n16997,notn16997;
or (n16997,s0n16997,s1n16997);
not(notn16997,n14375);
and (s0n16997,notn16997,n16998);
and (s1n16997,n14375,n17000);
wire s0n16998,s1n16998,notn16998;
or (n16998,s0n16998,s1n16998);
not(notn16998,n14409);
and (s0n16998,notn16998,n16999);
and (s1n16998,n14409,n16981);
wire s0n16999,s1n16999,notn16999;
or (n16999,s0n16999,s1n16999);
not(notn16999,n14401);
and (s0n16999,notn16999,1'b0);
and (s1n16999,n14401,n16977);
and (n17001,n17002,n14137);
or (n17002,1'b0,n17003,n17013);
and (n17003,n17004,n14235);
wire s0n17004,s1n17004,notn17004;
or (n17004,s0n17004,s1n17004);
not(notn17004,n14227);
and (s0n17004,notn17004,1'b0);
and (s1n17004,n14227,n17005);
or (n17005,1'b0,n16824,n17006,n17007,n17008,n17009,n17012);
and (n17006,n16764,n14199);
and (n17007,n16766,n2781);
and (n17008,n16759,n14205);
and (n17009,n17010,n2789);
wire s0n17010,s1n17010,notn17010;
or (n17010,s0n17010,s1n17010);
not(notn17010,n14210);
and (s0n17010,notn17010,n16716);
and (s1n17010,n14210,n17011);
and (n17012,n17011,n14225);
and (n17013,n16722,n14455);
and (n17014,n16818,n14111);
not (n17015,n17016);
or (n17016,n17017,n14626);
not (n17017,n16871);
and (n17018,n17019,n13950);
wire s0n17019,s1n17019,notn17019;
or (n17019,s0n17019,s1n17019);
not(notn17019,n14131);
and (s0n17019,notn17019,1'b0);
and (s1n17019,n14131,n16770);
and (n17020,n17021,n14239);
wire s0n17021,s1n17021,notn17021;
or (n17021,s0n17021,s1n17021);
not(notn17021,n14131);
and (s0n17021,notn17021,1'b0);
and (s1n17021,n14131,n17004);
and (n17022,n16318,n16685);
and (n17023,n15978,n16316);
and (n17024,n15638,n15976);
and (n17025,n15299,n15636);
and (n17026,n14973,n15297);
and (n17027,n14635,n14971);
wire s0n17028,s1n17028,notn17028;
or (n17028,s0n17028,s1n17028);
not(notn17028,n14631);
and (s0n17028,notn17028,n17029);
and (s1n17028,n14631,n17032);
wire s0n17029,s1n17029,notn17029;
or (n17029,s0n17029,s1n17029);
not(notn17029,n14271);
and (s0n17029,notn17029,n17030);
and (s1n17029,n14271,n14382);
and (n17030,n17031,n14279);
or (n17031,n14365,n14718);
or (n17032,1'b0,n17033,n17035,n17039);
and (n17033,n14235,n17034);
or (n17034,n14111,n14237);
and (n17035,n17036,n17037);
not (n17036,n14131);
or (n17037,n17038,n14108);
or (n17038,n14239,n13950);
or (n17039,n14266,n14448);
wire s0n17040,s1n17040,notn17040;
or (n17040,s0n17040,s1n17040);
not(notn17040,n17293);
and (s0n17040,notn17040,n17041);
and (s1n17040,n17293,n17082);
xor (n17041,n17042,n17080);
xor (n17042,n17043,n17076);
wire s0n17043,s1n17043,notn17043;
or (n17043,s0n17043,s1n17043);
not(notn17043,n14631);
and (s0n17043,notn17043,n17044);
and (s1n17043,n14631,n17065);
not (n17044,n17045);
nor (n17045,n17046,n17047,n17057);
and (n17046,n14473,n14511);
nand (n17047,n17048,n17052);
or (n17048,n17049,n17050);
not (n17049,n14292);
not (n17050,n17051);
nor (n17051,n14496,n14570);
nand (n17052,n17053,n14557);
and (n17053,n17054,n585);
nor (n17054,n17055,n17056);
not (n17055,n14317);
nand (n17056,n14271,n13907);
nand (n17057,n17058,n17061);
not (n17058,n17059);
and (n17059,n17060,n14562);
and (n17060,n17054,n581);
not (n17061,n17062);
wire s0n17062,s1n17062,notn17062;
or (n17062,s0n17062,s1n17062);
not(notn17062,n14279);
and (s0n17062,notn17062,1'b0);
and (s1n17062,n14279,n17063);
and (n17063,n17064,n14120);
wire s0n17064,s1n17064,notn17064;
or (n17064,s0n17064,s1n17064);
not(notn17064,n14317);
and (s0n17064,notn17064,1'b0);
and (s1n17064,n14317,n14557);
or (n17065,n17066,n17068,n17070,n17072,n17074,1'b0);
and (n17066,n14577,n17067);
and (n17067,n13900,n14237);
and (n17068,n17069,n14111);
wire s0n17069,s1n17069,notn17069;
or (n17069,s0n17069,s1n17069);
not(notn17069,n13900);
and (s0n17069,notn17069,1'b0);
and (s1n17069,n13900,n14346);
and (n17070,n17071,n14108);
wire s0n17071,s1n17071,notn17071;
or (n17071,s0n17071,s1n17071);
not(notn17071,n14131);
and (s0n17071,notn17071,1'b0);
and (s1n17071,n14131,n14519);
and (n17072,n17073,n13950);
wire s0n17073,s1n17073,notn17073;
or (n17073,s0n17073,s1n17073);
not(notn17073,n14131);
and (s0n17073,notn17073,1'b0);
and (s1n17073,n14131,n14346);
and (n17074,n17075,n14239);
wire s0n17075,s1n17075,notn17075;
or (n17075,s0n17075,s1n17075);
not(notn17075,n14131);
and (s0n17075,notn17075,1'b0);
and (s1n17075,n14131,n14141);
nand (n17076,n17077,n17079);
or (n17077,n17078,n17050);
not (n17078,n14175);
nand (n17079,n14594,n14511);
or (n17080,n17081,n17109,n17292);
and (n17081,n17082,n17105);
wire s0n17082,s1n17082,notn17082;
or (n17082,s0n17082,s1n17082);
not(notn17082,n14631);
and (s0n17082,notn17082,n17083);
and (s1n17082,n14631,n17097);
not (n17083,n17084);
nor (n17084,n17085,n17086,n17090);
and (n17085,n14737,n14511);
nand (n17086,n17087,n17089);
or (n17087,n17088,n17050);
not (n17088,n14683);
nand (n17089,n17053,n14562);
nand (n17090,n17091,n17093);
not (n17091,n17092);
and (n17092,n17060,n14909);
not (n17093,n17094);
wire s0n17094,s1n17094,notn17094;
or (n17094,s0n17094,s1n17094);
not(notn17094,n14279);
and (s0n17094,notn17094,1'b0);
and (s1n17094,n14279,n17095);
and (n17095,n17096,n14120);
wire s0n17096,s1n17096,notn17096;
or (n17096,s0n17096,s1n17096);
not(notn17096,n14317);
and (s0n17096,notn17096,1'b0);
and (s1n17096,n14317,n14562);
or (n17097,n17098,n17099,n17101,n17102,n17103,1'b0);
and (n17098,n14920,n17067);
and (n17099,n17100,n14111);
wire s0n17100,s1n17100,notn17100;
or (n17100,s0n17100,s1n17100);
not(notn17100,n13900);
and (s0n17100,notn17100,1'b0);
and (s1n17100,n13900,n14821);
and (n17101,n14887,n14108);
and (n17102,n14820,n13950);
and (n17103,n17104,n14239);
wire s0n17104,s1n17104,notn17104;
or (n17104,s0n17104,s1n17104);
not(notn17104,n14131);
and (s0n17104,notn17104,1'b0);
and (s1n17104,n14131,n14655);
nand (n17105,n17106,n17108);
or (n17106,n17107,n17050);
not (n17107,n14667);
nand (n17108,n14937,n14511);
and (n17109,n17105,n17110);
or (n17110,n17111,n17139,n17291);
and (n17111,n17112,n17135);
wire s0n17112,s1n17112,notn17112;
or (n17112,s0n17112,s1n17112);
not(notn17112,n14631);
and (s0n17112,notn17112,n17113);
and (s1n17112,n14631,n17126);
not (n17113,n17114);
nor (n17114,n17115,n17116,n17120);
and (n17115,n15168,n14511);
nand (n17116,n17117,n17119);
or (n17117,n17118,n17050);
not (n17118,n15051);
nand (n17119,n17053,n14909);
nand (n17120,n17121,n17122);
nand (n17121,n17060,n15233);
not (n17122,n17123);
wire s0n17123,s1n17123,notn17123;
or (n17123,s0n17123,s1n17123);
not(notn17123,n14279);
and (s0n17123,notn17123,1'b0);
and (s1n17123,n14279,n17124);
and (n17124,n17125,n14120);
wire s0n17125,s1n17125,notn17125;
or (n17125,s0n17125,s1n17125);
not(notn17125,n14317);
and (s0n17125,notn17125,1'b0);
and (s1n17125,n14317,n14909);
or (n17126,n17127,n17128,n17130,n17132,n17133,1'b0);
and (n17127,n15244,n17067);
and (n17128,n17129,n14111);
wire s0n17129,s1n17129,notn17129;
or (n17129,s0n17129,s1n17129);
not(notn17129,n13900);
and (s0n17129,notn17129,1'b0);
and (s1n17129,n13900,n15119);
and (n17130,n17131,n14108);
wire s0n17131,s1n17131,notn17131;
or (n17131,s0n17131,s1n17131);
not(notn17131,n14131);
and (s0n17131,notn17131,1'b0);
and (s1n17131,n14131,n15191);
and (n17132,n15291,n13950);
and (n17133,n17134,n14239);
wire s0n17134,s1n17134,notn17134;
or (n17134,s0n17134,s1n17134);
not(notn17134,n14131);
and (s0n17134,notn17134,1'b0);
and (s1n17134,n14131,n15056);
nand (n17135,n17136,n17138);
or (n17136,n17137,n17050);
not (n17137,n15068);
nand (n17138,n15261,n14511);
and (n17139,n17135,n17140);
or (n17140,n17141,n17171,n17290);
and (n17141,n17142,n17167);
wire s0n17142,s1n17142,notn17142;
or (n17142,s0n17142,s1n17142);
not(notn17142,n14631);
and (s0n17142,notn17142,n17143);
and (s1n17142,n14631,n17159);
not (n17143,n17144);
nor (n17144,n17145,n17146,n17150);
and (n17145,n15400,n14511);
nand (n17146,n17147,n17149);
or (n17147,n17148,n17050);
not (n17148,n15347);
nand (n17149,n17053,n15233);
nand (n17150,n17151,n17155);
not (n17151,n17152);
nor (n17152,n17153,n17154);
not (n17153,n17060);
not (n17154,n15573);
not (n17155,n17156);
wire s0n17156,s1n17156,notn17156;
or (n17156,s0n17156,s1n17156);
not(notn17156,n14279);
and (s0n17156,notn17156,1'b0);
and (s1n17156,n14279,n17157);
and (n17157,n17158,n14120);
wire s0n17158,s1n17158,notn17158;
or (n17158,s0n17158,s1n17158);
not(notn17158,n14317);
and (s0n17158,notn17158,1'b0);
and (s1n17158,n14317,n15233);
or (n17159,n17160,n17161,n17163,n17164,n17165,1'b0);
and (n17160,n15584,n17067);
and (n17161,n17162,n14111);
wire s0n17162,s1n17162,notn17162;
or (n17162,s0n17162,s1n17162);
not(notn17162,n13900);
and (s0n17162,notn17162,1'b0);
and (s1n17162,n13900,n15484);
and (n17163,n15551,n14108);
and (n17164,n15483,n13950);
and (n17165,n17166,n14239);
wire s0n17166,s1n17166,notn17166;
or (n17166,s0n17166,s1n17166);
not(notn17166,n14131);
and (s0n17166,notn17166,1'b0);
and (s1n17166,n14131,n15319);
nand (n17167,n17168,n17170);
or (n17168,n17169,n17050);
not (n17169,n15331);
nand (n17170,n15601,n14511);
and (n17171,n17167,n17172);
or (n17172,n17173,n17201,n17289);
and (n17173,n17174,n17197);
wire s0n17174,s1n17174,notn17174;
or (n17174,s0n17174,s1n17174);
not(notn17174,n14631);
and (s0n17174,notn17174,n17175);
and (s1n17174,n14631,n17189);
not (n17175,n17176);
nor (n17176,n17177,n17178,n17182);
and (n17177,n15739,n14511);
not (n17178,n17179);
nor (n17179,n17180,n17181);
and (n17180,n17051,n15686);
and (n17181,n17060,n15912);
nand (n17182,n17183,n17185);
or (n17183,n17184,n17154);
not (n17184,n17053);
not (n17185,n17186);
wire s0n17186,s1n17186,notn17186;
or (n17186,s0n17186,s1n17186);
not(notn17186,n14279);
and (s0n17186,notn17186,1'b0);
and (s1n17186,n14279,n17187);
and (n17187,n17188,n14120);
wire s0n17188,s1n17188,notn17188;
or (n17188,s0n17188,s1n17188);
not(notn17188,n14317);
and (s0n17188,notn17188,1'b0);
and (s1n17188,n14317,n15573);
or (n17189,n17190,n17191,n17193,n17194,n17195,1'b0);
and (n17190,n15923,n17067);
and (n17191,n17192,n14111);
wire s0n17192,s1n17192,notn17192;
or (n17192,s0n17192,s1n17192);
not(notn17192,n13900);
and (s0n17192,notn17192,1'b0);
and (s1n17192,n13900,n15823);
and (n17193,n15890,n14108);
and (n17194,n15822,n13950);
and (n17195,n17196,n14239);
wire s0n17196,s1n17196,notn17196;
or (n17196,s0n17196,s1n17196);
not(notn17196,n14131);
and (s0n17196,notn17196,1'b0);
and (s1n17196,n14131,n15658);
nand (n17197,n17198,n17200);
or (n17198,n17199,n17050);
not (n17199,n15670);
nand (n17200,n15940,n14511);
and (n17201,n17197,n17202);
or (n17202,n17203,n17230,n17288);
and (n17203,n17204,n17226);
wire s0n17204,s1n17204,notn17204;
or (n17204,s0n17204,s1n17204);
not(notn17204,n14631);
and (s0n17204,notn17204,n17205);
and (s1n17204,n14631,n17218);
not (n17205,n17206);
nor (n17206,n17207,n17208,n17212);
and (n17207,n16079,n14511);
not (n17208,n17209);
nor (n17209,n17210,n17211);
and (n17210,n17051,n16026);
and (n17211,n17060,n16252);
nand (n17212,n17213,n17214);
nand (n17213,n17053,n15912);
not (n17214,n17215);
wire s0n17215,s1n17215,notn17215;
or (n17215,s0n17215,s1n17215);
not(notn17215,n14279);
and (s0n17215,notn17215,1'b0);
and (s1n17215,n14279,n17216);
and (n17216,n17217,n14120);
wire s0n17217,s1n17217,notn17217;
or (n17217,s0n17217,s1n17217);
not(notn17217,n14317);
and (s0n17217,notn17217,1'b0);
and (s1n17217,n14317,n15912);
or (n17218,n17219,n17220,n17222,n17223,n17224,1'b0);
and (n17219,n16263,n17067);
and (n17220,n17221,n14111);
wire s0n17221,s1n17221,notn17221;
or (n17221,s0n17221,s1n17221);
not(notn17221,n13900);
and (s0n17221,notn17221,1'b0);
and (s1n17221,n13900,n16163);
and (n17222,n16230,n14108);
and (n17223,n16162,n13950);
and (n17224,n17225,n14239);
wire s0n17225,s1n17225,notn17225;
or (n17225,s0n17225,s1n17225);
not(notn17225,n14131);
and (s0n17225,notn17225,1'b0);
and (s1n17225,n14131,n15998);
nand (n17226,n17227,n17229);
or (n17227,n17228,n17050);
not (n17228,n16010);
nand (n17229,n16280,n14511);
and (n17230,n17226,n17231);
or (n17231,n17232,n17261,n17287);
and (n17232,n17233,n17257);
wire s0n17233,s1n17233,notn17233;
or (n17233,s0n17233,s1n17233);
not(notn17233,n14631);
and (s0n17233,notn17233,n17234);
and (s1n17233,n14631,n17249);
wire s0n17234,s1n17234,notn17234;
or (n17234,s0n17234,s1n17234);
not(notn17234,n14271);
and (s0n17234,notn17234,n17235);
and (s1n17234,n14271,n17238);
wire s0n17235,s1n17235,notn17235;
or (n17235,s0n17235,s1n17235);
not(notn17235,n14279);
and (s0n17235,notn17235,1'b0);
and (s1n17235,n14279,n17236);
and (n17236,n17237,n14120);
wire s0n17237,s1n17237,notn17237;
or (n17237,s0n17237,s1n17237);
not(notn17237,n14317);
and (s0n17237,notn17237,1'b0);
and (s1n17237,n14317,n16252);
or (n17238,n17239,n17242,1'b0);
and (n17239,n17240,n13907);
wire s0n17240,s1n17240,notn17240;
or (n17240,s0n17240,s1n17240);
not(notn17240,n14317);
and (s0n17240,notn17240,1'b0);
and (s1n17240,n14317,n17241);
wire s0n17241,s1n17241,notn17241;
or (n17241,s0n17241,s1n17241);
not(notn17241,n581);
and (s0n17241,notn17241,n16252);
and (s1n17241,n581,n16592);
and (n17242,n17243,n14385);
wire s0n17243,s1n17243,notn17243;
or (n17243,s0n17243,s1n17243);
not(notn17243,n2799);
and (s0n17243,notn17243,1'b0);
and (s1n17243,n2799,n17244);
or (n17244,1'b0,n17245,n17247);
and (n17245,n17246,n13900);
wire s0n17246,s1n17246,notn17246;
or (n17246,s0n17246,s1n17246);
not(notn17246,n14570);
and (s0n17246,notn17246,n16366);
and (s1n17246,n14570,1'b0);
and (n17247,n17248,n14131);
wire s0n17248,s1n17248,notn17248;
or (n17248,s0n17248,s1n17248);
not(notn17248,n14573);
and (s0n17248,notn17248,n16419);
and (s1n17248,n14573,1'b0);
or (n17249,n17250,n17251,n17253,n17254,n17255,1'b0);
and (n17250,n16604,n17067);
and (n17251,n17252,n14111);
wire s0n17252,s1n17252,notn17252;
or (n17252,s0n17252,s1n17252);
not(notn17252,n13900);
and (s0n17252,notn17252,1'b0);
and (s1n17252,n13900,n16503);
and (n17253,n16570,n14108);
and (n17254,n16502,n13950);
and (n17255,n17256,n14239);
wire s0n17256,s1n17256,notn17256;
or (n17256,s0n17256,s1n17256);
not(notn17256,n14131);
and (s0n17256,notn17256,1'b0);
and (s1n17256,n14131,n16338);
nand (n17257,n17258,n17260);
or (n17258,n17259,n17050);
not (n17259,n16350);
nand (n17260,n16630,n14511);
and (n17261,n17257,n17262);
and (n17262,n17263,n17283);
wire s0n17263,s1n17263,notn17263;
or (n17263,s0n17263,s1n17263);
not(notn17263,n14631);
and (s0n17263,notn17263,n17264);
and (s1n17263,n14631,n17275);
not (n17264,n17265);
nor (n17265,n17266,n17267,n17268);
and (n17266,n17051,n16734);
and (n17267,n16787,n14511);
not (n17268,n17269);
and (n17269,n17270,n17271);
nand (n17270,n17053,n16592);
not (n17271,n17272);
wire s0n17272,s1n17272,notn17272;
or (n17272,s0n17272,s1n17272);
not(notn17272,n14279);
and (s0n17272,notn17272,1'b0);
and (s1n17272,n14279,n17273);
and (n17273,n17274,n14120);
wire s0n17274,s1n17274,notn17274;
or (n17274,s0n17274,s1n17274);
not(notn17274,n14317);
and (s0n17274,notn17274,1'b0);
and (s1n17274,n14317,n16592);
or (n17275,n17276,n17277,n17279,n17280,n17281,1'b0);
and (n17276,n16970,n17067);
and (n17277,n17278,n14111);
wire s0n17278,s1n17278,notn17278;
or (n17278,s0n17278,s1n17278);
not(notn17278,n13900);
and (s0n17278,notn17278,1'b0);
and (s1n17278,n13900,n16871);
and (n17279,n16938,n14108);
and (n17280,n16870,n13950);
and (n17281,n17282,n14239);
wire s0n17282,s1n17282,notn17282;
or (n17282,s0n17282,s1n17282);
not(notn17282,n14131);
and (s0n17282,notn17282,1'b0);
and (s1n17282,n14131,n16706);
nand (n17283,n17284,n17286);
or (n17284,n17285,n17050);
not (n17285,n16718);
nand (n17286,n16987,n14511);
and (n17287,n17233,n17262);
and (n17288,n17204,n17231);
and (n17289,n17174,n17202);
and (n17290,n17142,n17172);
and (n17291,n17112,n17140);
and (n17292,n17082,n17110);
wire s0n17293,s1n17293,notn17293;
or (n17293,s0n17293,s1n17293);
not(notn17293,n14631);
and (s0n17293,notn17293,n14315);
and (s1n17293,n14631,n17294);
or (n17294,1'b0,n17295,n17296,n17297,1'b0);
and (n17295,n13900,n17034);
and (n17296,n14125,n13949);
and (n17297,n14131,n14239);
or (n17298,n17299,n17306,n17362);
and (n17299,n17300,n17303);
wire s0n17300,s1n17300,notn17300;
or (n17300,s0n17300,s1n17300);
not(notn17300,n17028);
and (s0n17300,notn17300,n17301);
and (s1n17300,n17028,1'b0);
xor (n17301,n17302,n14971);
xor (n17302,n14635,n14898);
wire s0n17303,s1n17303,notn17303;
or (n17303,s0n17303,s1n17303);
not(notn17303,n17293);
and (s0n17303,notn17303,n17304);
and (s1n17303,n17293,n17112);
xor (n17304,n17305,n17110);
xor (n17305,n17082,n17105);
and (n17306,n17303,n17307);
or (n17307,n17308,n17315,n17361);
and (n17308,n17309,n17312);
wire s0n17309,s1n17309,notn17309;
or (n17309,s0n17309,s1n17309);
not(notn17309,n17028);
and (s0n17309,notn17309,n17310);
and (s1n17309,n17028,1'b0);
xor (n17310,n17311,n15297);
xor (n17311,n14973,n15222);
wire s0n17312,s1n17312,notn17312;
or (n17312,s0n17312,s1n17312);
not(notn17312,n17293);
and (s0n17312,notn17312,n17313);
and (s1n17312,n17293,n17142);
xor (n17313,n17314,n17140);
xor (n17314,n17112,n17135);
and (n17315,n17312,n17316);
or (n17316,n17317,n17324,n17360);
and (n17317,n17318,n17321);
wire s0n17318,s1n17318,notn17318;
or (n17318,s0n17318,s1n17318);
not(notn17318,n17028);
and (s0n17318,notn17318,n17319);
and (s1n17318,n17028,1'b0);
xor (n17319,n17320,n15636);
xor (n17320,n15299,n15562);
wire s0n17321,s1n17321,notn17321;
or (n17321,s0n17321,s1n17321);
not(notn17321,n17293);
and (s0n17321,notn17321,n17322);
and (s1n17321,n17293,n17174);
xor (n17322,n17323,n17172);
xor (n17323,n17142,n17167);
and (n17324,n17321,n17325);
or (n17325,n17326,n17333,n17359);
and (n17326,n17327,n17330);
wire s0n17327,s1n17327,notn17327;
or (n17327,s0n17327,s1n17327);
not(notn17327,n17028);
and (s0n17327,notn17327,n17328);
and (s1n17327,n17028,1'b0);
xor (n17328,n17329,n15976);
xor (n17329,n15638,n15901);
wire s0n17330,s1n17330,notn17330;
or (n17330,s0n17330,s1n17330);
not(notn17330,n17293);
and (s0n17330,notn17330,n17331);
and (s1n17330,n17293,n17204);
xor (n17331,n17332,n17202);
xor (n17332,n17174,n17197);
and (n17333,n17330,n17334);
or (n17334,n17335,n17342,n17358);
and (n17335,n17336,n17339);
wire s0n17336,s1n17336,notn17336;
or (n17336,s0n17336,s1n17336);
not(notn17336,n17028);
and (s0n17336,notn17336,n17337);
and (s1n17336,n17028,1'b0);
xor (n17337,n17338,n16316);
xor (n17338,n15978,n16241);
wire s0n17339,s1n17339,notn17339;
or (n17339,s0n17339,s1n17339);
not(notn17339,n17293);
and (s0n17339,notn17339,n17340);
and (s1n17339,n17293,n17233);
xor (n17340,n17341,n17231);
xor (n17341,n17204,n17226);
and (n17342,n17339,n17343);
or (n17343,n17344,n17351,n17357);
and (n17344,n17345,n17348);
wire s0n17345,s1n17345,notn17345;
or (n17345,s0n17345,s1n17345);
not(notn17345,n17028);
and (s0n17345,notn17345,n17346);
and (s1n17345,n17028,1'b0);
xor (n17346,n17347,n16685);
xor (n17347,n16318,n16581);
wire s0n17348,s1n17348,notn17348;
or (n17348,s0n17348,s1n17348);
not(notn17348,n17293);
and (s0n17348,notn17348,n17349);
and (s1n17348,n17293,n17263);
xor (n17349,n17350,n17262);
xor (n17350,n17233,n17257);
and (n17351,n17348,n17352);
and (n17352,n17353,n17355);
wire s0n17353,s1n17353,notn17353;
or (n17353,s0n17353,s1n17353);
not(notn17353,n17028);
and (s0n17353,notn17353,n17354);
and (s1n17353,n17028,1'b0);
xor (n17354,n16686,n16949);
wire s0n17355,s1n17355,notn17355;
or (n17355,s0n17355,s1n17355);
not(notn17355,n17293);
and (s0n17355,notn17355,n17356);
and (s1n17355,n17293,1'b0);
xor (n17356,n17263,n17283);
and (n17357,n17345,n17352);
and (n17358,n17336,n17343);
and (n17359,n17327,n17334);
and (n17360,n17318,n17325);
and (n17361,n17309,n17316);
and (n17362,n17300,n17307);
and (n17363,n17364,n17366);
xor (n17364,n17365,n17307);
xor (n17365,n17300,n17303);
and (n17366,n17367,n17369);
xor (n17367,n17368,n17316);
xor (n17368,n17309,n17312);
or (n17369,n17370,n17373,n17391);
and (n17370,n17371,n14503);
xor (n17371,n17372,n17325);
xor (n17372,n17318,n17321);
and (n17373,n14503,n17374);
and (n17374,n17375,n17377);
xor (n17375,n17376,n17334);
xor (n17376,n17327,n17330);
and (n17377,n17378,n17380);
xor (n17378,n17379,n17343);
xor (n17379,n17336,n17339);
or (n17380,n17381,n17384,n17390);
and (n17381,n17382,n17294);
xor (n17382,n17383,n17352);
xor (n17383,n17345,n17348);
and (n17384,n17294,n17385);
and (n17385,n17386,n17387);
xor (n17386,n17353,n17355);
or (n17387,n17388,n17389,1'b0,1'b0,1'b0);
and (n17388,n14125,n14137);
and (n17389,n14131,n17034);
and (n17390,n17382,n17385);
and (n17391,n17371,n17374);
xor (n17392,n17393,n17442);
xor (n17393,n17394,n17438);
xor (n17394,n17395,n17425);
xor (n17395,n17396,n17421);
xor (n17396,n17397,n17411);
nand (n17397,n17398,n17401);
or (n17398,n17399,n14494);
not (n17399,n17400);
not (n17401,n17402);
wire s0n17402,s1n17402,notn17402;
or (n17402,s0n17402,s1n17402);
not(notn17402,n14326);
and (s0n17402,notn17402,n17403);
and (s1n17402,n14326,n17405);
wire s0n17403,s1n17403,notn17403;
or (n17403,s0n17403,s1n17403);
not(notn17403,n14315);
and (s0n17403,notn17403,1'b0);
and (s1n17403,n14315,n17404);
or (n17405,1'b0,n17406,n17408,n17410);
and (n17406,n17407,n14321);
and (n17408,n17409,n14324);
and (n17410,n17404,n14184);
wire s0n17411,s1n17411,notn17411;
or (n17411,s0n17411,s1n17411);
not(notn17411,n14271);
and (s0n17411,notn17411,n17412);
and (s1n17411,n14271,n17418);
wire s0n17412,s1n17412,notn17412;
or (n17412,s0n17412,s1n17412);
not(notn17412,n14279);
and (s0n17412,notn17412,1'b0);
and (s1n17412,n14279,n17413);
and (n17413,n17414,n14120);
wire s0n17414,s1n17414,notn17414;
or (n17414,s0n17414,s1n17414);
not(notn17414,n14125);
and (s0n17414,notn17414,1'b0);
and (s1n17414,n14125,n17415);
wire s0n17415,s1n17415,notn17415;
or (n17415,s0n17415,s1n17415);
not(notn17415,n14317);
and (s0n17415,notn17415,n17416);
and (s1n17415,n14317,n17417);
and (n17418,n17419,n13907);
wire s0n17419,s1n17419,notn17419;
or (n17419,s0n17419,s1n17419);
not(notn17419,n14125);
and (s0n17419,notn17419,1'b0);
and (s1n17419,n14125,n17420);
wire s0n17420,s1n17420,notn17420;
or (n17420,s0n17420,s1n17420);
not(notn17420,n14563);
and (s0n17420,notn17420,n17416);
and (s1n17420,n14563,n14557);
or (n17421,n17422,n17423,n17424);
and (n17422,n13883,n14550);
and (n17423,n14550,n14633);
and (n17424,n13883,n14633);
wire s0n17425,s1n17425,notn17425;
or (n17425,s0n17425,s1n17425);
not(notn17425,n17293);
and (s0n17425,notn17425,n17426);
and (s1n17425,n17293,n17043);
xor (n17426,n17427,n17434);
wire s0n17427,s1n17427,notn17427;
or (n17427,s0n17427,s1n17427);
not(notn17427,n14271);
and (s0n17427,notn17427,n17428);
and (s1n17427,n14271,n17431);
wire s0n17428,s1n17428,notn17428;
or (n17428,s0n17428,s1n17428);
not(notn17428,n14279);
and (s0n17428,notn17428,1'b0);
and (s1n17428,n14279,n17429);
and (n17429,n17430,n14120);
wire s0n17430,s1n17430,notn17430;
or (n17430,s0n17430,s1n17430);
not(notn17430,n14317);
and (s0n17430,notn17430,1'b0);
and (s1n17430,n14317,n17417);
and (n17431,n17432,n13907);
wire s0n17432,s1n17432,notn17432;
or (n17432,s0n17432,s1n17432);
not(notn17432,n14317);
and (s0n17432,notn17432,1'b0);
and (s1n17432,n14317,n17433);
wire s0n17433,s1n17433,notn17433;
or (n17433,s0n17433,s1n17433);
not(notn17433,n581);
and (s0n17433,notn17433,n17417);
and (s1n17433,n581,n14557);
or (n17434,n17435,n17436,n17437);
and (n17435,n17043,n17076);
and (n17436,n17076,n17080);
and (n17437,n17043,n17080);
or (n17438,n17439,n17440,n17441);
and (n17439,n13880,n17040);
and (n17440,n17040,n17298);
and (n17441,n13880,n17298);
and (n17442,n13878,n17363);
or (n17443,n17387,n14503);
wire s0n17444,s1n17444,notn17444;
or (n17444,s0n17444,s1n17444);
not(notn17444,n17443);
and (s0n17444,notn17444,n17445);
and (s1n17444,n17443,n17491);
xor (n17445,n17446,n17490);
xor (n17446,n17447,n17486);
xor (n17447,n17448,n17478);
xor (n17448,n17449,n17474);
xor (n17449,n17450,n17464);
nand (n17450,n17451,n17454);
or (n17451,n17452,n14494);
not (n17452,n17453);
not (n17454,n17455);
wire s0n17455,s1n17455,notn17455;
or (n17455,s0n17455,s1n17455);
not(notn17455,n14326);
and (s0n17455,notn17455,n17456);
and (s1n17455,n14326,n17458);
wire s0n17456,s1n17456,notn17456;
or (n17456,s0n17456,s1n17456);
not(notn17456,n14315);
and (s0n17456,notn17456,1'b0);
and (s1n17456,n14315,n17457);
or (n17458,1'b0,n17459,n17461,n17463);
and (n17459,n17460,n14321);
and (n17461,n17462,n14324);
and (n17463,n17457,n14184);
wire s0n17464,s1n17464,notn17464;
or (n17464,s0n17464,s1n17464);
not(notn17464,n14271);
and (s0n17464,notn17464,n17465);
and (s1n17464,n14271,n17471);
wire s0n17465,s1n17465,notn17465;
or (n17465,s0n17465,s1n17465);
not(notn17465,n14279);
and (s0n17465,notn17465,1'b0);
and (s1n17465,n14279,n17466);
and (n17466,n17467,n14120);
wire s0n17467,s1n17467,notn17467;
or (n17467,s0n17467,s1n17467);
not(notn17467,n14125);
and (s0n17467,notn17467,1'b0);
and (s1n17467,n14125,n17468);
wire s0n17468,s1n17468,notn17468;
or (n17468,s0n17468,s1n17468);
not(notn17468,n14317);
and (s0n17468,notn17468,n17469);
and (s1n17468,n14317,n17470);
and (n17471,n17472,n13907);
wire s0n17472,s1n17472,notn17472;
or (n17472,s0n17472,s1n17472);
not(notn17472,n14125);
and (s0n17472,notn17472,1'b0);
and (s1n17472,n14125,n17473);
wire s0n17473,s1n17473,notn17473;
or (n17473,s0n17473,s1n17473);
not(notn17473,n14563);
and (s0n17473,notn17473,n17469);
and (s1n17473,n14563,n17417);
or (n17474,n17475,n17476,n17477);
and (n17475,n17397,n17411);
and (n17476,n17411,n17421);
and (n17477,n17397,n17421);
wire s0n17478,s1n17478,notn17478;
or (n17478,s0n17478,s1n17478);
not(notn17478,n17293);
and (s0n17478,notn17478,n17479);
and (s1n17478,n17293,n17427);
wire s0n17479,s1n17479,notn17479;
or (n17479,s0n17479,s1n17479);
not(notn17479,n14271);
and (s0n17479,notn17479,n17480);
and (s1n17479,n14271,n17483);
wire s0n17480,s1n17480,notn17480;
or (n17480,s0n17480,s1n17480);
not(notn17480,n14279);
and (s0n17480,notn17480,1'b0);
and (s1n17480,n14279,n17481);
and (n17481,n17482,n14120);
wire s0n17482,s1n17482,notn17482;
or (n17482,s0n17482,s1n17482);
not(notn17482,n14317);
and (s0n17482,notn17482,1'b0);
and (s1n17482,n14317,n17470);
and (n17483,n17484,n13907);
wire s0n17484,s1n17484,notn17484;
or (n17484,s0n17484,s1n17484);
not(notn17484,n14317);
and (s0n17484,notn17484,1'b0);
and (s1n17484,n14317,n17485);
wire s0n17485,s1n17485,notn17485;
or (n17485,s0n17485,s1n17485);
not(notn17485,n581);
and (s0n17485,notn17485,n17470);
and (s1n17485,n581,n17417);
or (n17486,n17487,n17488,n17489);
and (n17487,n17395,n17425);
and (n17488,n17425,n17438);
and (n17489,n17395,n17438);
and (n17490,n17393,n17442);
xor (n17491,n17492,n17536);
xor (n17492,n17493,n17532);
xor (n17493,n17494,n17524);
xor (n17494,n17495,n17520);
xor (n17495,n17496,n17510);
nand (n17496,n17497,n17500);
or (n17497,n17498,n14494);
not (n17498,n17499);
not (n17500,n17501);
wire s0n17501,s1n17501,notn17501;
or (n17501,s0n17501,s1n17501);
not(notn17501,n14326);
and (s0n17501,notn17501,n17502);
and (s1n17501,n14326,n17504);
wire s0n17502,s1n17502,notn17502;
or (n17502,s0n17502,s1n17502);
not(notn17502,n14315);
and (s0n17502,notn17502,1'b0);
and (s1n17502,n14315,n17503);
or (n17504,1'b0,n17505,n17507,n17509);
and (n17505,n17506,n14321);
and (n17507,n17508,n14324);
and (n17509,n17503,n14184);
wire s0n17510,s1n17510,notn17510;
or (n17510,s0n17510,s1n17510);
not(notn17510,n14271);
and (s0n17510,notn17510,n17511);
and (s1n17510,n14271,n17517);
wire s0n17511,s1n17511,notn17511;
or (n17511,s0n17511,s1n17511);
not(notn17511,n14279);
and (s0n17511,notn17511,1'b0);
and (s1n17511,n14279,n17512);
and (n17512,n17513,n14120);
wire s0n17513,s1n17513,notn17513;
or (n17513,s0n17513,s1n17513);
not(notn17513,n14125);
and (s0n17513,notn17513,1'b0);
and (s1n17513,n14125,n17514);
wire s0n17514,s1n17514,notn17514;
or (n17514,s0n17514,s1n17514);
not(notn17514,n14317);
and (s0n17514,notn17514,n17515);
and (s1n17514,n14317,n17516);
and (n17517,n17518,n13907);
wire s0n17518,s1n17518,notn17518;
or (n17518,s0n17518,s1n17518);
not(notn17518,n14125);
and (s0n17518,notn17518,1'b0);
and (s1n17518,n14125,n17519);
wire s0n17519,s1n17519,notn17519;
or (n17519,s0n17519,s1n17519);
not(notn17519,n14563);
and (s0n17519,notn17519,n17515);
and (s1n17519,n14563,n17470);
or (n17520,n17521,n17522,n17523);
and (n17521,n17450,n17464);
and (n17522,n17464,n17474);
and (n17523,n17450,n17474);
wire s0n17524,s1n17524,notn17524;
or (n17524,s0n17524,s1n17524);
not(notn17524,n17293);
and (s0n17524,notn17524,n17525);
and (s1n17524,n17293,n17479);
wire s0n17525,s1n17525,notn17525;
or (n17525,s0n17525,s1n17525);
not(notn17525,n14271);
and (s0n17525,notn17525,n17526);
and (s1n17525,n14271,n17529);
wire s0n17526,s1n17526,notn17526;
or (n17526,s0n17526,s1n17526);
not(notn17526,n14279);
and (s0n17526,notn17526,1'b0);
and (s1n17526,n14279,n17527);
and (n17527,n17528,n14120);
wire s0n17528,s1n17528,notn17528;
or (n17528,s0n17528,s1n17528);
not(notn17528,n14317);
and (s0n17528,notn17528,1'b0);
and (s1n17528,n14317,n17516);
and (n17529,n17530,n13907);
wire s0n17530,s1n17530,notn17530;
or (n17530,s0n17530,s1n17530);
not(notn17530,n14317);
and (s0n17530,notn17530,1'b0);
and (s1n17530,n14317,n17531);
wire s0n17531,s1n17531,notn17531;
or (n17531,s0n17531,s1n17531);
not(notn17531,n581);
and (s0n17531,notn17531,n17516);
and (s1n17531,n581,n17470);
or (n17532,n17533,n17534,n17535);
and (n17533,n17448,n17478);
and (n17534,n17478,n17486);
and (n17535,n17448,n17486);
and (n17536,n17446,n17490);
wire s0n17537,s1n17537,notn17537;
or (n17537,s0n17537,s1n17537);
not(notn17537,n17443);
and (s0n17537,notn17537,n17538);
and (s1n17537,n17443,n17584);
xor (n17538,n17539,n17583);
xor (n17539,n17540,n17579);
xor (n17540,n17541,n17571);
xor (n17541,n17542,n17567);
xor (n17542,n17543,n17557);
nand (n17543,n17544,n17547);
or (n17544,n17545,n14494);
not (n17545,n17546);
not (n17547,n17548);
wire s0n17548,s1n17548,notn17548;
or (n17548,s0n17548,s1n17548);
not(notn17548,n14326);
and (s0n17548,notn17548,n17549);
and (s1n17548,n14326,n17551);
wire s0n17549,s1n17549,notn17549;
or (n17549,s0n17549,s1n17549);
not(notn17549,n14315);
and (s0n17549,notn17549,1'b0);
and (s1n17549,n14315,n17550);
or (n17551,1'b0,n17552,n17554,n17556);
and (n17552,n17553,n14321);
and (n17554,n17555,n14324);
and (n17556,n17550,n14184);
wire s0n17557,s1n17557,notn17557;
or (n17557,s0n17557,s1n17557);
not(notn17557,n14271);
and (s0n17557,notn17557,n17558);
and (s1n17557,n14271,n17564);
wire s0n17558,s1n17558,notn17558;
or (n17558,s0n17558,s1n17558);
not(notn17558,n14279);
and (s0n17558,notn17558,1'b0);
and (s1n17558,n14279,n17559);
and (n17559,n17560,n14120);
wire s0n17560,s1n17560,notn17560;
or (n17560,s0n17560,s1n17560);
not(notn17560,n14125);
and (s0n17560,notn17560,1'b0);
and (s1n17560,n14125,n17561);
wire s0n17561,s1n17561,notn17561;
or (n17561,s0n17561,s1n17561);
not(notn17561,n14317);
and (s0n17561,notn17561,n17562);
and (s1n17561,n14317,n17563);
and (n17564,n17565,n13907);
wire s0n17565,s1n17565,notn17565;
or (n17565,s0n17565,s1n17565);
not(notn17565,n14125);
and (s0n17565,notn17565,1'b0);
and (s1n17565,n14125,n17566);
wire s0n17566,s1n17566,notn17566;
or (n17566,s0n17566,s1n17566);
not(notn17566,n14563);
and (s0n17566,notn17566,n17562);
and (s1n17566,n14563,n17516);
or (n17567,n17568,n17569,n17570);
and (n17568,n17496,n17510);
and (n17569,n17510,n17520);
and (n17570,n17496,n17520);
wire s0n17571,s1n17571,notn17571;
or (n17571,s0n17571,s1n17571);
not(notn17571,n17293);
and (s0n17571,notn17571,n17572);
and (s1n17571,n17293,n17525);
wire s0n17572,s1n17572,notn17572;
or (n17572,s0n17572,s1n17572);
not(notn17572,n14271);
and (s0n17572,notn17572,n17573);
and (s1n17572,n14271,n17576);
wire s0n17573,s1n17573,notn17573;
or (n17573,s0n17573,s1n17573);
not(notn17573,n14279);
and (s0n17573,notn17573,1'b0);
and (s1n17573,n14279,n17574);
and (n17574,n17575,n14120);
wire s0n17575,s1n17575,notn17575;
or (n17575,s0n17575,s1n17575);
not(notn17575,n14317);
and (s0n17575,notn17575,1'b0);
and (s1n17575,n14317,n17563);
and (n17576,n17577,n13907);
wire s0n17577,s1n17577,notn17577;
or (n17577,s0n17577,s1n17577);
not(notn17577,n14317);
and (s0n17577,notn17577,1'b0);
and (s1n17577,n14317,n17578);
wire s0n17578,s1n17578,notn17578;
or (n17578,s0n17578,s1n17578);
not(notn17578,n581);
and (s0n17578,notn17578,n17563);
and (s1n17578,n581,n17516);
or (n17579,n17580,n17581,n17582);
and (n17580,n17494,n17524);
and (n17581,n17524,n17532);
and (n17582,n17494,n17532);
and (n17583,n17492,n17536);
xor (n17584,n17585,n17617);
xor (n17585,n17586,n17613);
xor (n17586,n17587,n17611);
xor (n17587,n17588,n17607);
xor (n17588,n17589,n17603);
nand (n17589,n17590,n17593);
or (n17590,n17591,n14494);
not (n17591,n17592);
not (n17593,n17594);
wire s0n17594,s1n17594,notn17594;
or (n17594,s0n17594,s1n17594);
not(notn17594,n14326);
and (s0n17594,notn17594,n17595);
and (s1n17594,n14326,n17597);
wire s0n17595,s1n17595,notn17595;
or (n17595,s0n17595,s1n17595);
not(notn17595,n14315);
and (s0n17595,notn17595,1'b0);
and (s1n17595,n14315,n17596);
or (n17597,1'b0,n17598,n17600,n17602);
and (n17598,n17599,n14321);
and (n17600,n17601,n14324);
and (n17602,n17596,n14184);
wire s0n17603,s1n17603,notn17603;
or (n17603,s0n17603,s1n17603);
not(notn17603,n14271);
and (s0n17603,notn17603,n17558);
and (s1n17603,n14271,n17604);
and (n17604,n17605,n13907);
wire s0n17605,s1n17605,notn17605;
or (n17605,s0n17605,s1n17605);
not(notn17605,n14125);
and (s0n17605,notn17605,1'b0);
and (s1n17605,n14125,n17606);
wire s0n17606,s1n17606,notn17606;
or (n17606,s0n17606,s1n17606);
not(notn17606,n14563);
and (s0n17606,notn17606,n17562);
and (s1n17606,n14563,n17563);
or (n17607,n17608,n17609,n17610);
and (n17608,n17543,n17557);
and (n17609,n17557,n17567);
and (n17610,n17543,n17567);
wire s0n17611,s1n17611,notn17611;
or (n17611,s0n17611,s1n17611);
not(notn17611,n14271);
and (s0n17611,notn17611,n17573);
and (s1n17611,n14271,n17612);
and (n17612,n17575,n13907);
or (n17613,n17614,n17615,n17616);
and (n17614,n17541,n17571);
and (n17615,n17571,n17579);
and (n17616,n17541,n17579);
and (n17617,n17539,n17583);
wire s0n17618,s1n17618,notn17618;
or (n17618,s0n17618,s1n17618);
not(notn17618,n17722);
and (s0n17618,notn17618,n17619);
and (s1n17618,n17722,1'b0);
wire s0n17619,s1n17619,notn17619;
or (n17619,s0n17619,s1n17619);
not(notn17619,n17620);
and (s0n17619,notn17619,1'b1);
and (s1n17619,n17620,n13874);
nor (n17620,n17621,n17654,n17685,n17715,n17718,n17720,n17721,n17722);
wire s0n17621,s1n17621,notn17621;
or (n17621,s0n17621,s1n17621);
not(notn17621,n14503);
and (s0n17621,notn17621,n17622);
and (s1n17621,n14503,n17625);
wire s0n17622,s1n17622,notn17622;
or (n17622,s0n17622,s1n17622);
not(notn17622,n17294);
and (s0n17622,notn17622,n17623);
and (s1n17622,n17294,n17624);
wire s0n17623,s1n17623,notn17623;
or (n17623,s0n17623,s1n17623);
not(notn17623,n17443);
and (s0n17623,notn17623,n17392);
and (s1n17623,n17443,n17445);
wire s0n17624,s1n17624,notn17624;
or (n17624,s0n17624,s1n17624);
not(notn17624,n17443);
and (s0n17624,notn17624,n17491);
and (s1n17624,n17443,n17538);
wire s0n17625,s1n17625,notn17625;
or (n17625,s0n17625,s1n17625);
not(notn17625,n17443);
and (s0n17625,notn17625,n17584);
and (s1n17625,n17443,n17626);
xor (n17626,n17627,n17653);
xor (n17627,n17628,n17649);
xor (n17628,n17629,n17611);
xor (n17629,n17630,n17645);
xor (n17630,n17631,n17603);
nand (n17631,n17632,n17635);
or (n17632,n17633,n14494);
not (n17633,n17634);
not (n17635,n17636);
wire s0n17636,s1n17636,notn17636;
or (n17636,s0n17636,s1n17636);
not(notn17636,n14326);
and (s0n17636,notn17636,n17637);
and (s1n17636,n14326,n17639);
wire s0n17637,s1n17637,notn17637;
or (n17637,s0n17637,s1n17637);
not(notn17637,n14315);
and (s0n17637,notn17637,1'b0);
and (s1n17637,n14315,n17638);
or (n17639,1'b0,n17640,n17642,n17644);
and (n17640,n17641,n14321);
and (n17642,n17643,n14324);
and (n17644,n17638,n14184);
or (n17645,n17646,n17647,n17648);
and (n17646,n17589,n17603);
and (n17647,n17603,n17607);
and (n17648,n17589,n17607);
or (n17649,n17650,n17651,n17652);
and (n17650,n17587,n17611);
and (n17651,n17611,n17613);
and (n17652,n17587,n17613);
and (n17653,n17585,n17617);
wire s0n17654,s1n17654,notn17654;
or (n17654,s0n17654,s1n17654);
not(notn17654,n14503);
and (s0n17654,notn17654,n17655);
and (s1n17654,n14503,n17656);
wire s0n17655,s1n17655,notn17655;
or (n17655,s0n17655,s1n17655);
not(notn17655,n17294);
and (s0n17655,notn17655,n17444);
and (s1n17655,n17294,n17537);
wire s0n17656,s1n17656,notn17656;
or (n17656,s0n17656,s1n17656);
not(notn17656,n17443);
and (s0n17656,notn17656,n17626);
and (s1n17656,n17443,n17657);
xor (n17657,n17658,n17684);
xor (n17658,n17659,n17680);
xor (n17659,n17660,n17611);
xor (n17660,n17661,n17676);
xor (n17661,n17662,n17603);
nand (n17662,n17663,n17666);
or (n17663,n17664,n14494);
not (n17664,n17665);
not (n17666,n17667);
wire s0n17667,s1n17667,notn17667;
or (n17667,s0n17667,s1n17667);
not(notn17667,n14326);
and (s0n17667,notn17667,n17668);
and (s1n17667,n14326,n17670);
wire s0n17668,s1n17668,notn17668;
or (n17668,s0n17668,s1n17668);
not(notn17668,n14315);
and (s0n17668,notn17668,1'b0);
and (s1n17668,n14315,n17669);
or (n17670,1'b0,n17671,n17673,n17675);
and (n17671,n17672,n14321);
and (n17673,n17674,n14324);
and (n17675,n17669,n14184);
or (n17676,n17677,n17678,n17679);
and (n17677,n17631,n17603);
and (n17678,n17603,n17645);
and (n17679,n17631,n17645);
or (n17680,n17681,n17682,n17683);
and (n17681,n17629,n17611);
and (n17682,n17611,n17649);
and (n17683,n17629,n17649);
and (n17684,n17627,n17653);
wire s0n17685,s1n17685,notn17685;
or (n17685,s0n17685,s1n17685);
not(notn17685,n14503);
and (s0n17685,notn17685,n17624);
and (s1n17685,n14503,n17686);
wire s0n17686,s1n17686,notn17686;
or (n17686,s0n17686,s1n17686);
not(notn17686,n17443);
and (s0n17686,notn17686,n17657);
and (s1n17686,n17443,n17687);
xor (n17687,n17688,n17714);
xor (n17688,n17689,n17710);
xor (n17689,n17690,n17611);
xor (n17690,n17691,n17706);
xor (n17691,n17692,n17603);
nand (n17692,n17693,n17696);
or (n17693,n17694,n14494);
not (n17694,n17695);
not (n17696,n17697);
wire s0n17697,s1n17697,notn17697;
or (n17697,s0n17697,s1n17697);
not(notn17697,n14326);
and (s0n17697,notn17697,n17698);
and (s1n17697,n14326,n17700);
wire s0n17698,s1n17698,notn17698;
or (n17698,s0n17698,s1n17698);
not(notn17698,n14315);
and (s0n17698,notn17698,1'b0);
and (s1n17698,n14315,n17699);
or (n17700,1'b0,n17701,n17703,n17705);
and (n17701,n17702,n14321);
and (n17703,n17704,n14324);
and (n17705,n17699,n14184);
or (n17706,n17707,n17708,n17709);
and (n17707,n17662,n17603);
and (n17708,n17603,n17676);
and (n17709,n17662,n17676);
or (n17710,n17711,n17712,n17713);
and (n17711,n17660,n17611);
and (n17712,n17611,n17680);
and (n17713,n17660,n17680);
and (n17714,n17658,n17684);
wire s0n17715,s1n17715,notn17715;
or (n17715,s0n17715,s1n17715);
not(notn17715,n14503);
and (s0n17715,notn17715,n17537);
and (s1n17715,n14503,n17716);
wire s0n17716,s1n17716,notn17716;
or (n17716,s0n17716,s1n17716);
not(notn17716,n17443);
and (s0n17716,notn17716,n17687);
and (s1n17716,n17443,n17717);
and (n17717,n17688,n17714);
and (n17718,n17584,n17719);
not (n17719,n17443);
and (n17720,n17626,n17719);
wire s0n17721,s1n17721,notn17721;
or (n17721,s0n17721,s1n17721);
not(notn17721,n14503);
and (s0n17721,notn17721,n17686);
and (s1n17721,n14503,1'b0);
wire s0n17722,s1n17722,notn17722;
or (n17722,s0n17722,s1n17722);
not(notn17722,n14503);
and (s0n17722,notn17722,n17716);
and (s1n17722,n14503,1'b0);
and (n17723,n3,n17036);
wire s0n17724,s1n17724,notn17724;
or (n17724,s0n17724,s1n17724);
not(notn17724,n19716);
and (s0n17724,notn17724,n3);
and (s1n17724,n19716,n17725);
wire s0n17725,s1n17725,notn17725;
or (n17725,s0n17725,s1n17725);
not(notn17725,n18690);
and (s0n17725,notn17725,n17726);
and (s1n17725,n18690,n17736);
wire s0n17726,s1n17726,notn17726;
or (n17726,s0n17726,s1n17726);
not(notn17726,n14503);
and (s0n17726,notn17726,n17727);
and (s1n17726,n14503,n19717);
wire s0n17727,s1n17727,notn17727;
or (n17727,s0n17727,s1n17727);
not(notn17727,n19713);
and (s0n17727,notn17727,n17728);
and (s1n17727,n19713,n19430);
wire s0n17728,s1n17728,notn17728;
or (n17728,s0n17728,s1n17728);
not(notn17728,n19421);
and (s0n17728,notn17728,n17729);
and (s1n17728,n19421,n19274);
wire s0n17729,s1n17729,notn17729;
or (n17729,s0n17729,s1n17729);
not(notn17729,n19269);
and (s0n17729,notn17729,n17730);
and (s1n17729,n19269,n19195);
xor (n17730,n17731,n19128);
xor (n17731,n17732,n19063);
xor (n17732,n17733,n18707);
wire s0n17733,s1n17733,notn17733;
or (n17733,s0n17733,s1n17733);
not(notn17733,n18690);
and (s0n17733,notn17733,n17734);
and (s1n17733,n18690,1'b0);
xor (n17734,n17735,n17879);
xor (n17735,n17736,n17837);
wire s0n17736,s1n17736,notn17736;
or (n17736,s0n17736,s1n17736);
not(notn17736,n14631);
and (s0n17736,notn17736,n17737);
and (s1n17736,n14631,n17780);
wire s0n17737,s1n17737,notn17737;
or (n17737,s0n17737,s1n17737);
not(notn17737,n14271);
and (s0n17737,notn17737,n17738);
and (s1n17737,n14271,n17768);
wire s0n17738,s1n17738,notn17738;
or (n17738,s0n17738,s1n17738);
not(notn17738,n14279);
and (s0n17738,notn17738,1'b0);
and (s1n17738,n14279,n17739);
or (n17739,n17740,n17744,n17750,n17751);
and (n17740,n17741,n14120);
wire s0n17741,s1n17741,notn17741;
or (n17741,s0n17741,s1n17741);
not(notn17741,n14125);
and (s0n17741,notn17741,1'b0);
and (s1n17741,n14125,n17742);
wire s0n17742,s1n17742,notn17742;
or (n17742,s0n17742,s1n17742);
not(notn17742,n14317);
and (s0n17742,notn17742,n17743);
and (s1n17742,n14317,n14312);
and (n17744,n17745,n14718);
or (n17745,1'b0,n17746,n17747,n17748,n17749);
and (n17746,n14141,n13889);
and (n17747,n14280,n13897);
and (n17748,n14247,n13900);
and (n17749,n14297,n14131);
and (n17750,n14519,n14365);
and (n17751,n17752,n14367);
or (n17752,n17753,n17759,n17763,n17766);
and (n17753,n17754,n17758);
wire s0n17754,s1n17754,notn17754;
or (n17754,s0n17754,s1n17754);
not(notn17754,n14131);
and (s0n17754,notn17754,n17755);
and (s1n17754,n14131,n17756);
wire s0n17755,s1n17755,notn17755;
or (n17755,s0n17755,s1n17755);
not(notn17755,n13900);
and (s0n17755,notn17755,1'b0);
and (s1n17755,n13900,n17743);
wire s0n17756,s1n17756,notn17756;
or (n17756,s0n17756,s1n17756);
not(notn17756,n17757);
and (s0n17756,notn17756,n14297);
and (s1n17756,n17757,1'b0);
or (n17757,n14160,n14162);
and (n17758,n14211,n14368);
and (n17759,n17760,n17762);
wire s0n17760,s1n17760,notn17760;
or (n17760,s0n17760,s1n17760);
not(notn17760,n13900);
and (s0n17760,notn17760,1'b0);
and (s1n17760,n13900,n17761);
and (n17762,n14570,n14368);
and (n17763,n17764,n17765);
wire s0n17764,s1n17764,notn17764;
or (n17764,s0n17764,s1n17764);
not(notn17764,n14131);
and (s0n17764,notn17764,n17755);
and (s1n17764,n14131,n14297);
nor (n17765,n14570,n14368);
and (n17766,n13900,n17767);
nor (n17767,n14211,n14368);
or (n17768,n17769,n17770,n17778,n17779);
and (n17769,n17741,n13907);
and (n17770,n17771,n14385);
wire s0n17771,s1n17771,notn17771;
or (n17771,s0n17771,s1n17771);
not(notn17771,n2799);
and (s0n17771,notn17771,1'b0);
and (s1n17771,n2799,n17772);
or (n17772,1'b0,n17773,n17775,n17776);
and (n17773,n17774,n13889);
wire s0n17774,s1n17774,notn17774;
or (n17774,s0n17774,s1n17774);
not(notn17774,n17767);
and (s0n17774,notn17774,n17743);
and (s1n17774,n17767,1'b1);
and (n17775,n17743,n14243);
and (n17776,n17777,n14131);
wire s0n17777,s1n17777,notn17777;
or (n17777,s0n17777,s1n17777);
not(notn17777,n14573);
and (s0n17777,notn17777,n14543);
and (s1n17777,n14573,1'b0);
and (n17778,n14519,n14381);
and (n17779,n17745,n14192);
or (n17780,1'b0,n17781,n17786,n17793,n17797,n17801,n17807,n17812,n17835,n17836);
and (n17781,n17782,n14237);
or (n17782,1'b0,n17783,n17784,n17785);
and (n17783,n14436,n13889);
and (n17784,n14341,n13897);
and (n17785,n14519,n14455);
and (n17786,n17787,n14137);
or (n17787,1'b0,n17788,n17790,n17792,n17749);
and (n17788,n17789,n13889);
and (n17790,n17791,n13897);
and (n17792,n3,n13900);
and (n17793,n17794,n14111);
or (n17794,1'b0,n17795,n17796,n17785);
and (n17795,n14297,n13889);
and (n17796,n13902,n13897);
and (n17797,n17798,n14108);
or (n17798,1'b0,n17799,n17800);
and (n17799,n14280,n14235);
and (n17800,n14297,n14455);
and (n17801,n17802,n13950);
or (n17802,1'b0,n17803,n17804,n17805);
and (n17803,n14247,n13889);
and (n17804,n13902,n13900);
and (n17805,n14297,n17806);
or (n17806,n14131,n13897);
and (n17807,n17808,n14239);
or (n17808,1'b0,n17809,n17810,n17811,n17749);
and (n17809,n14240,n13889);
and (n17810,n3,n13897);
and (n17811,n14341,n13900);
and (n17812,n17813,n17820);
or (n17813,1'b0,n17814,n17833);
and (n17814,n17815,n13900);
or (n17815,n17816,n17827,n17832);
and (n17816,n17743,n17817);
and (n17817,n17818,n17823);
not (n17818,n17819);
and (n17819,n17820,n17821);
nor (n17820,n13951,n14109,n14040,n14074);
and (n17821,n14184,n17822);
not (n17822,n14369);
not (n17823,n17824);
and (n17824,n17820,n17825);
and (n17825,n14421,n17826);
not (n17826,n14212);
and (n17827,n17828,n17829);
wire s0n17828,s1n17828,notn17828;
or (n17828,s0n17828,s1n17828);
not(notn17828,n17823);
and (s0n17828,notn17828,1'b0);
and (s1n17828,n17823,n17743);
or (n17829,n17830,n17831);
and (n17830,n17818,n17824);
nor (n17831,n17818,n17824);
nor (n17832,n17818,n17823);
and (n17833,n17834,n14131);
wire s0n17834,s1n17834,notn17834;
or (n17834,s0n17834,s1n17834);
not(notn17834,n17823);
and (s0n17834,notn17834,1'b0);
and (s1n17834,n17823,n14297);
and (n17835,n14519,n14448);
and (n17836,n17745,n14266);
wire s0n17837,s1n17837,notn17837;
or (n17837,s0n17837,s1n17837);
not(notn17837,n14631);
and (s0n17837,notn17837,n17838);
and (s1n17837,n14631,n17859);
wire s0n17838,s1n17838,notn17838;
or (n17838,s0n17838,s1n17838);
not(notn17838,n14271);
and (s0n17838,notn17838,n17839);
and (s1n17838,n14271,n17847);
wire s0n17839,s1n17839,notn17839;
or (n17839,s0n17839,s1n17839);
not(notn17839,n14279);
and (s0n17839,notn17839,1'b0);
and (s1n17839,n14279,n17840);
or (n17840,n14553,1'b0,n17841);
and (n17841,n17842,n14367);
or (n17842,n17843,n17846,1'b0);
and (n17843,n17844,n17758);
wire s0n17844,s1n17844,notn17844;
or (n17844,s0n17844,s1n17844);
not(notn17844,n14131);
and (s0n17844,notn17844,n17760);
and (s1n17844,n14131,n17845);
wire s0n17845,s1n17845,notn17845;
or (n17845,s0n17845,s1n17845);
not(notn17845,n17757);
and (s0n17845,notn17845,n14247);
and (s1n17845,n17757,1'b0);
and (n17846,n14246,n17765);
or (n17847,n17848,n17851,1'b0);
and (n17848,n17849,n13907);
wire s0n17849,s1n17849,notn17849;
or (n17849,s0n17849,s1n17849);
not(notn17849,n14125);
and (s0n17849,notn17849,1'b0);
and (s1n17849,n14125,n17850);
wire s0n17850,s1n17850,notn17850;
or (n17850,s0n17850,s1n17850);
not(notn17850,n14563);
and (s0n17850,notn17850,n14556);
and (s1n17850,n14563,n14557);
and (n17851,n17852,n14385);
wire s0n17852,s1n17852,notn17852;
or (n17852,s0n17852,s1n17852);
not(notn17852,n2799);
and (s0n17852,notn17852,1'b0);
and (s1n17852,n2799,n17853);
or (n17853,1'b0,n17854,n17855,n17857);
and (n17854,n17761,n14235);
and (n17855,n17856,n13900);
wire s0n17856,s1n17856,notn17856;
or (n17856,s0n17856,s1n17856);
not(notn17856,n14570);
and (s0n17856,notn17856,n14253);
and (s1n17856,n14570,1'b0);
and (n17857,n17858,n14131);
wire s0n17858,s1n17858,notn17858;
or (n17858,s0n17858,s1n17858);
not(notn17858,n14573);
and (s0n17858,notn17858,n14416);
and (s1n17858,n14573,1'b0);
or (n17859,n17860,n14245,n17863,n17868,n17871,n14548,n17873,1'b0);
and (n17860,n17861,n14237);
or (n17861,1'b0,n17862,n17073);
and (n17862,n14456,n13900);
and (n17863,n17864,n14111);
or (n17864,1'b0,n17865,n17866,n17867,n13901);
and (n17865,n14280,n13889);
and (n17866,n14247,n13897);
and (n17867,n14297,n13900);
and (n17868,n17869,n14108);
or (n17869,1'b0,n17746,n17870,n13901);
and (n17870,n14247,n14243);
and (n17871,n17872,n13950);
or (n17872,1'b0,n17746,n17747,n17748,n17071);
and (n17873,n17874,n17820);
or (n17874,1'b0,n17875,n17877);
and (n17875,n17876,n13900);
wire s0n17876,s1n17876,notn17876;
or (n17876,s0n17876,s1n17876);
not(notn17876,n17818);
and (s0n17876,notn17876,1'b0);
and (s1n17876,n17818,n17761);
and (n17877,n17878,n14131);
wire s0n17878,s1n17878,notn17878;
or (n17878,s0n17878,s1n17878);
not(notn17878,n17823);
and (s0n17878,notn17878,1'b0);
and (s1n17878,n17823,n14247);
or (n17879,n17880,n17992,n18689);
and (n17880,n17881,n17948);
wire s0n17881,s1n17881,notn17881;
or (n17881,s0n17881,s1n17881);
not(notn17881,n14631);
and (s0n17881,notn17881,n17882);
and (s1n17881,n14631,n17912);
wire s0n17882,s1n17882,notn17882;
or (n17882,s0n17882,s1n17882);
not(notn17882,n14271);
and (s0n17882,notn17882,n17883);
and (s1n17882,n14271,n17901);
wire s0n17883,s1n17883,notn17883;
or (n17883,s0n17883,s1n17883);
not(notn17883,n14279);
and (s0n17883,notn17883,1'b0);
and (s1n17883,n14279,n17884);
or (n17884,n17885,n14652,n17889,n17890);
and (n17885,n17886,n14120);
wire s0n17886,s1n17886,notn17886;
or (n17886,s0n17886,s1n17886);
not(notn17886,n14125);
and (s0n17886,notn17886,1'b0);
and (s1n17886,n14125,n17887);
wire s0n17887,s1n17887,notn17887;
or (n17887,s0n17887,s1n17887);
not(notn17887,n14317);
and (s0n17887,notn17887,n17888);
and (s1n17887,n14317,n14643);
and (n17889,n14791,n14365);
and (n17890,n17891,n14367);
or (n17891,n17892,n17896,n17899,1'b0);
and (n17892,n17893,n17758);
wire s0n17893,s1n17893,notn17893;
or (n17893,s0n17893,s1n17893);
not(notn17893,n14131);
and (s0n17893,notn17893,n17894);
and (s1n17893,n14131,n17895);
wire s0n17894,s1n17894,notn17894;
or (n17894,s0n17894,s1n17894);
not(notn17894,n13900);
and (s0n17894,notn17894,1'b0);
and (s1n17894,n13900,n17888);
wire s0n17895,s1n17895,notn17895;
or (n17895,s0n17895,s1n17895);
not(notn17895,n17757);
and (s0n17895,notn17895,n14703);
and (s1n17895,n17757,1'b0);
and (n17896,n17897,n17762);
wire s0n17897,s1n17897,notn17897;
or (n17897,s0n17897,s1n17897);
not(notn17897,n13900);
and (s0n17897,notn17897,1'b0);
and (s1n17897,n13900,n17898);
and (n17899,n17900,n17765);
wire s0n17900,s1n17900,notn17900;
or (n17900,s0n17900,s1n17900);
not(notn17900,n14131);
and (s0n17900,notn17900,n17894);
and (s1n17900,n14131,n14703);
or (n17901,n17902,n17903,n17911,n14762);
and (n17902,n17886,n13907);
and (n17903,n17904,n14385);
wire s0n17904,s1n17904,notn17904;
or (n17904,s0n17904,s1n17904);
not(notn17904,n2799);
and (s0n17904,notn17904,1'b0);
and (s1n17904,n2799,n17905);
or (n17905,1'b0,n17906,n17908,n17909);
and (n17906,n17907,n13889);
wire s0n17907,s1n17907,notn17907;
or (n17907,s0n17907,s1n17907);
not(notn17907,n17767);
and (s0n17907,notn17907,n17888);
and (s1n17907,n17767,1'b0);
and (n17908,n17888,n14243);
and (n17909,n17910,n14131);
wire s0n17910,s1n17910,notn17910;
or (n17910,s0n17910,s1n17910);
not(notn17910,n14573);
and (s0n17910,notn17910,n14815);
and (s1n17910,n14573,1'b0);
and (n17911,n14791,n14381);
or (n17912,1'b0,n17913,n17916,n17924,n17928,n17932,n17937,n17941,n17947,n14897);
and (n17913,n17914,n14237);
or (n17914,1'b0,n14786,n14788,n17915);
and (n17915,n14791,n14455);
and (n17916,n17917,n14137);
or (n17917,1'b0,n17918,n17920,n17922,n14702);
and (n17918,n17919,n13889);
and (n17920,n17921,n13897);
and (n17922,n17923,n13900);
and (n17924,n17925,n14111);
or (n17925,1'b0,n17926,n17927,n17915);
and (n17926,n14703,n13889);
and (n17927,n14861,n13897);
and (n17928,n17929,n14108);
or (n17929,1'b0,n17930,n17931);
and (n17930,n14671,n14235);
and (n17931,n14703,n14455);
and (n17932,n17933,n13950);
or (n17933,1'b0,n17934,n17935,n17936);
and (n17934,n14687,n13889);
and (n17935,n14861,n13900);
and (n17936,n14703,n17806);
and (n17937,n17938,n14239);
or (n17938,1'b0,n17939,n17940,n14886,n14702);
and (n17939,n14767,n13889);
and (n17940,n17923,n13897);
and (n17941,n17942,n17820);
or (n17942,1'b0,n17943,n17945);
and (n17943,n17944,n13900);
wire s0n17944,s1n17944,notn17944;
or (n17944,s0n17944,s1n17944);
not(notn17944,n17823);
and (s0n17944,notn17944,1'b0);
and (s1n17944,n17823,n17888);
and (n17945,n17946,n14131);
wire s0n17946,s1n17946,notn17946;
or (n17946,s0n17946,s1n17946);
not(notn17946,n17823);
and (s0n17946,notn17946,1'b0);
and (s1n17946,n17823,n14703);
and (n17947,n14791,n14448);
wire s0n17948,s1n17948,notn17948;
or (n17948,s0n17948,s1n17948);
not(notn17948,n14631);
and (s0n17948,notn17948,n17949);
and (s1n17948,n14631,n17970);
wire s0n17949,s1n17949,notn17949;
or (n17949,s0n17949,s1n17949);
not(notn17949,n14271);
and (s0n17949,notn17949,n17950);
and (s1n17949,n14271,n17958);
wire s0n17950,s1n17950,notn17950;
or (n17950,s0n17950,s1n17950);
not(notn17950,n14279);
and (s0n17950,notn17950,1'b0);
and (s1n17950,n14279,n17951);
or (n17951,n14901,1'b0,n17952);
and (n17952,n17953,n14367);
or (n17953,n17954,n17957,1'b0);
and (n17954,n17955,n17758);
wire s0n17955,s1n17955,notn17955;
or (n17955,s0n17955,s1n17955);
not(notn17955,n14131);
and (s0n17955,notn17955,n17897);
and (s1n17955,n14131,n17956);
wire s0n17956,s1n17956,notn17956;
or (n17956,s0n17956,s1n17956);
not(notn17956,n17757);
and (s0n17956,notn17956,n14687);
and (s1n17956,n17757,1'b0);
and (n17957,n14783,n17765);
or (n17958,n17959,n17962,1'b0);
and (n17959,n17960,n13907);
wire s0n17960,s1n17960,notn17960;
or (n17960,s0n17960,s1n17960);
not(notn17960,n14125);
and (s0n17960,notn17960,1'b0);
and (s1n17960,n14125,n17961);
wire s0n17961,s1n17961,notn17961;
or (n17961,s0n17961,s1n17961);
not(notn17961,n14563);
and (s0n17961,notn17961,n14904);
and (s1n17961,n14563,n14562);
and (n17962,n17963,n14385);
wire s0n17963,s1n17963,notn17963;
or (n17963,s0n17963,s1n17963);
not(notn17963,n2799);
and (s0n17963,notn17963,1'b0);
and (s1n17963,n2799,n17964);
or (n17964,1'b0,n17965,n17966,n17968);
and (n17965,n17898,n14235);
and (n17966,n17967,n13900);
wire s0n17967,s1n17967,notn17967;
or (n17967,s0n17967,s1n17967);
not(notn17967,n14570);
and (s0n17967,notn17967,n14694);
and (s1n17967,n14570,1'b0);
and (n17968,n17969,n14131);
wire s0n17969,s1n17969,notn17969;
or (n17969,s0n17969,s1n17969);
not(notn17969,n14573);
and (s0n17969,notn17969,n14847);
and (s1n17969,n14573,1'b0);
or (n17970,n17971,n17974,n17975,n17980,n17983,n17985,n17986,1'b0);
and (n17971,n17972,n14237);
or (n17972,1'b0,n17973,n14820);
and (n17973,n14720,n13900);
and (n17974,n14783,n14137);
and (n17975,n17976,n14111);
or (n17976,1'b0,n17977,n17978,n17979,n14860);
and (n17977,n14671,n13889);
and (n17978,n14687,n13897);
and (n17979,n14703,n13900);
and (n17980,n17981,n14108);
or (n17981,1'b0,n14654,n17982,n14860);
and (n17982,n14687,n14243);
and (n17983,n17984,n13950);
or (n17984,1'b0,n14654,n14670,n14686,n14887);
and (n17985,n14895,n14239);
and (n17986,n17987,n17820);
or (n17987,1'b0,n17988,n17990);
and (n17988,n17989,n13900);
wire s0n17989,s1n17989,notn17989;
or (n17989,s0n17989,s1n17989);
not(notn17989,n17818);
and (s0n17989,notn17989,1'b0);
and (s1n17989,n17818,n17898);
and (n17990,n17991,n14131);
wire s0n17991,s1n17991,notn17991;
or (n17991,s0n17991,s1n17991);
not(notn17991,n17823);
and (s0n17991,notn17991,1'b0);
and (s1n17991,n17823,n14687);
and (n17992,n17948,n17993);
or (n17993,n17994,n18115,n18688);
and (n17994,n17995,n18073);
wire s0n17995,s1n17995,notn17995;
or (n17995,s0n17995,s1n17995);
not(notn17995,n14631);
and (s0n17995,notn17995,n17996);
and (s1n17995,n14631,n18033);
wire s0n17996,s1n17996,notn17996;
or (n17996,s0n17996,s1n17996);
not(notn17996,n14271);
and (s0n17996,notn17996,n17997);
and (s1n17996,n14271,n18021);
wire s0n17997,s1n17997,notn17997;
or (n17997,s0n17997,s1n17997);
not(notn17997,n14279);
and (s0n17997,notn17997,1'b0);
and (s1n17997,n14279,n17998);
or (n17998,n17999,n18003,n18009,n18010);
and (n17999,n18000,n14120);
wire s0n18000,s1n18000,notn18000;
or (n18000,s0n18000,s1n18000);
not(notn18000,n14125);
and (s0n18000,notn18000,1'b0);
and (s1n18000,n14125,n18001);
wire s0n18001,s1n18001,notn18001;
or (n18001,s0n18001,s1n18001);
not(notn18001,n14317);
and (s0n18001,notn18001,n18002);
and (s1n18001,n14317,n15029);
and (n18003,n18004,n14718);
or (n18004,1'b0,n18005,n18006,n18007,n18008);
and (n18005,n15056,n13889);
and (n18006,n15039,n13897);
and (n18007,n15072,n13900);
and (n18008,n15012,n14131);
and (n18009,n15191,n14365);
and (n18010,n18011,n14367);
or (n18011,n18012,n18016,n18019,1'b0);
and (n18012,n18013,n17758);
wire s0n18013,s1n18013,notn18013;
or (n18013,s0n18013,s1n18013);
not(notn18013,n14131);
and (s0n18013,notn18013,n18014);
and (s1n18013,n14131,n18015);
wire s0n18014,s1n18014,notn18014;
or (n18014,s0n18014,s1n18014);
not(notn18014,n13900);
and (s0n18014,notn18014,1'b0);
and (s1n18014,n13900,n18002);
wire s0n18015,s1n18015,notn18015;
or (n18015,s0n18015,s1n18015);
not(notn18015,n17757);
and (s0n18015,notn18015,n15012);
and (s1n18015,n17757,1'b0);
and (n18016,n18017,n17762);
wire s0n18017,s1n18017,notn18017;
or (n18017,s0n18017,s1n18017);
not(notn18017,n13900);
and (s0n18017,notn18017,1'b0);
and (s1n18017,n13900,n18018);
and (n18019,n18020,n17765);
wire s0n18020,s1n18020,notn18020;
or (n18020,s0n18020,s1n18020);
not(notn18020,n14131);
and (s0n18020,notn18020,n18014);
and (s1n18020,n14131,n15012);
or (n18021,n18022,n18023,n18031,n18032);
and (n18022,n18000,n13907);
and (n18023,n18024,n14385);
wire s0n18024,s1n18024,notn18024;
or (n18024,s0n18024,s1n18024);
not(notn18024,n2799);
and (s0n18024,notn18024,1'b0);
and (s1n18024,n2799,n18025);
or (n18025,1'b0,n18026,n18028,n18029);
and (n18026,n18027,n13889);
wire s0n18027,s1n18027,notn18027;
or (n18027,s0n18027,s1n18027);
not(notn18027,n17767);
and (s0n18027,notn18027,n18002);
and (s1n18027,n17767,1'b0);
and (n18028,n18002,n14243);
and (n18029,n18030,n14131);
wire s0n18030,s1n18030,notn18030;
or (n18030,s0n18030,s1n18030);
not(notn18030,n14573);
and (s0n18030,notn18030,n15215);
and (s1n18030,n14573,1'b0);
and (n18031,n15191,n14381);
and (n18032,n18004,n14192);
or (n18033,1'b0,n18034,n18039,n18047,n18051,n18055,n18060,n18065,n18071,n18072);
and (n18034,n18035,n14237);
or (n18035,1'b0,n18036,n18037,n18038);
and (n18036,n15117,n13889);
and (n18037,n15107,n13897);
and (n18038,n15191,n14455);
and (n18039,n18040,n14137);
or (n18040,1'b0,n18041,n18043,n18045,n18008);
and (n18041,n18042,n13889);
and (n18043,n18044,n13897);
and (n18045,n18046,n13900);
and (n18047,n18048,n14111);
or (n18048,1'b0,n18049,n18050,n18038);
and (n18049,n15012,n13889);
and (n18050,n14984,n13897);
and (n18051,n18052,n14108);
or (n18052,1'b0,n18053,n18054);
and (n18053,n15039,n14235);
and (n18054,n15012,n14455);
and (n18055,n18056,n13950);
or (n18056,1'b0,n18057,n18058,n18059);
and (n18057,n15072,n13889);
and (n18058,n14984,n13900);
and (n18059,n15012,n17806);
and (n18060,n18061,n14239);
or (n18061,1'b0,n18062,n18063,n18064,n18008);
and (n18062,n15100,n13889);
and (n18063,n18046,n13897);
and (n18064,n15107,n13900);
and (n18065,n18066,n17820);
or (n18066,1'b0,n18067,n18069);
and (n18067,n18068,n13900);
wire s0n18068,s1n18068,notn18068;
or (n18068,s0n18068,s1n18068);
not(notn18068,n17823);
and (s0n18068,notn18068,1'b0);
and (s1n18068,n17823,n18002);
and (n18069,n18070,n14131);
wire s0n18070,s1n18070,notn18070;
or (n18070,s0n18070,s1n18070);
not(notn18070,n17823);
and (s0n18070,notn18070,1'b0);
and (s1n18070,n17823,n15012);
and (n18071,n15191,n14448);
and (n18072,n18004,n14266);
wire s0n18073,s1n18073,notn18073;
or (n18073,s0n18073,s1n18073);
not(notn18073,n14631);
and (s0n18073,notn18073,n18074);
and (s1n18073,n14631,n18095);
wire s0n18074,s1n18074,notn18074;
or (n18074,s0n18074,s1n18074);
not(notn18074,n14271);
and (s0n18074,notn18074,n18075);
and (s1n18074,n14271,n18083);
wire s0n18075,s1n18075,notn18075;
or (n18075,s0n18075,s1n18075);
not(notn18075,n14279);
and (s0n18075,notn18075,1'b0);
and (s1n18075,n14279,n18076);
or (n18076,n15225,1'b0,n18077);
and (n18077,n18078,n14367);
or (n18078,n18079,n18082,1'b0);
and (n18079,n18080,n17758);
wire s0n18080,s1n18080,notn18080;
or (n18080,s0n18080,s1n18080);
not(notn18080,n14131);
and (s0n18080,notn18080,n18017);
and (s1n18080,n14131,n18081);
wire s0n18081,s1n18081,notn18081;
or (n18081,s0n18081,s1n18081);
not(notn18081,n17757);
and (s0n18081,notn18081,n15072);
and (s1n18081,n17757,1'b0);
and (n18082,n15104,n17765);
or (n18083,n18084,n18087,1'b0);
and (n18084,n18085,n13907);
wire s0n18085,s1n18085,notn18085;
or (n18085,s0n18085,s1n18085);
not(notn18085,n14125);
and (s0n18085,notn18085,1'b0);
and (s1n18085,n14125,n18086);
wire s0n18086,s1n18086,notn18086;
or (n18086,s0n18086,s1n18086);
not(notn18086,n14563);
and (s0n18086,notn18086,n15228);
and (s1n18086,n14563,n14909);
and (n18087,n18088,n14385);
wire s0n18088,s1n18088,notn18088;
or (n18088,s0n18088,s1n18088);
not(notn18088,n2799);
and (s0n18088,notn18088,1'b0);
and (s1n18088,n2799,n18089);
or (n18089,1'b0,n18090,n18091,n18093);
and (n18090,n18018,n14235);
and (n18091,n18092,n13900);
wire s0n18092,s1n18092,notn18092;
or (n18092,s0n18092,s1n18092);
not(notn18092,n14570);
and (s0n18092,notn18092,n15079);
and (s1n18092,n14570,1'b0);
and (n18093,n18094,n14131);
wire s0n18094,s1n18094,notn18094;
or (n18094,s0n18094,s1n18094);
not(notn18094,n14573);
and (s0n18094,notn18094,n15145);
and (s1n18094,n14573,1'b0);
or (n18095,n18096,n15103,n18099,n18104,n18107,n15220,n18109,1'b0);
and (n18096,n18097,n14237);
or (n18097,1'b0,n18098,n15291);
and (n18098,n15151,n13900);
and (n18099,n18100,n14111);
or (n18100,1'b0,n18101,n18102,n18103,n14983);
and (n18101,n15039,n13889);
and (n18102,n15072,n13897);
and (n18103,n15012,n13900);
and (n18104,n18105,n14108);
or (n18105,1'b0,n18005,n18106,n14983);
and (n18106,n15072,n14243);
and (n18107,n18108,n13950);
or (n18108,1'b0,n18005,n18006,n18007,n17131);
and (n18109,n18110,n17820);
or (n18110,1'b0,n18111,n18113);
and (n18111,n18112,n13900);
wire s0n18112,s1n18112,notn18112;
or (n18112,s0n18112,s1n18112);
not(notn18112,n17818);
and (s0n18112,notn18112,1'b0);
and (s1n18112,n17818,n18018);
and (n18113,n18114,n14131);
wire s0n18114,s1n18114,notn18114;
or (n18114,s0n18114,s1n18114);
not(notn18114,n17823);
and (s0n18114,notn18114,1'b0);
and (s1n18114,n17823,n15072);
and (n18115,n18073,n18116);
or (n18116,n18117,n18229,n18687);
and (n18117,n18118,n18185);
wire s0n18118,s1n18118,notn18118;
or (n18118,s0n18118,s1n18118);
not(notn18118,n14631);
and (s0n18118,notn18118,n18119);
and (s1n18118,n14631,n18149);
wire s0n18119,s1n18119,notn18119;
or (n18119,s0n18119,s1n18119);
not(notn18119,n14271);
and (s0n18119,notn18119,n18120);
and (s1n18119,n14271,n18138);
wire s0n18120,s1n18120,notn18120;
or (n18120,s0n18120,s1n18120);
not(notn18120,n14279);
and (s0n18120,notn18120,1'b0);
and (s1n18120,n14279,n18121);
or (n18121,n18122,n15316,n18126,n18127);
and (n18122,n18123,n14120);
wire s0n18123,s1n18123,notn18123;
or (n18123,s0n18123,s1n18123);
not(notn18123,n14125);
and (s0n18123,notn18123,1'b0);
and (s1n18123,n14125,n18124);
wire s0n18124,s1n18124,notn18124;
or (n18124,s0n18124,s1n18124);
not(notn18124,n14317);
and (s0n18124,notn18124,n18125);
and (s1n18124,n14317,n15307);
and (n18126,n15454,n14365);
and (n18127,n18128,n14367);
or (n18128,n18129,n18133,n18136,1'b0);
and (n18129,n18130,n17758);
wire s0n18130,s1n18130,notn18130;
or (n18130,s0n18130,s1n18130);
not(notn18130,n14131);
and (s0n18130,notn18130,n18131);
and (s1n18130,n14131,n18132);
wire s0n18131,s1n18131,notn18131;
or (n18131,s0n18131,s1n18131);
not(notn18131,n13900);
and (s0n18131,notn18131,1'b0);
and (s1n18131,n13900,n18125);
wire s0n18132,s1n18132,notn18132;
or (n18132,s0n18132,s1n18132);
not(notn18132,n17757);
and (s0n18132,notn18132,n15367);
and (s1n18132,n17757,1'b0);
and (n18133,n18134,n17762);
wire s0n18134,s1n18134,notn18134;
or (n18134,s0n18134,s1n18134);
not(notn18134,n13900);
and (s0n18134,notn18134,1'b0);
and (s1n18134,n13900,n18135);
and (n18136,n18137,n17765);
wire s0n18137,s1n18137,notn18137;
or (n18137,s0n18137,s1n18137);
not(notn18137,n14131);
and (s0n18137,notn18137,n18131);
and (s1n18137,n14131,n15367);
or (n18138,n18139,n18140,n18148,n15425);
and (n18139,n18123,n13907);
and (n18140,n18141,n14385);
wire s0n18141,s1n18141,notn18141;
or (n18141,s0n18141,s1n18141);
not(notn18141,n2799);
and (s0n18141,notn18141,1'b0);
and (s1n18141,n2799,n18142);
or (n18142,1'b0,n18143,n18145,n18146);
and (n18143,n18144,n13889);
wire s0n18144,s1n18144,notn18144;
or (n18144,s0n18144,s1n18144);
not(notn18144,n17767);
and (s0n18144,notn18144,n18125);
and (s1n18144,n17767,1'b0);
and (n18145,n18125,n14243);
and (n18146,n18147,n14131);
wire s0n18147,s1n18147,notn18147;
or (n18147,s0n18147,s1n18147);
not(notn18147,n14573);
and (s0n18147,notn18147,n15478);
and (s1n18147,n14573,1'b0);
and (n18148,n15454,n14381);
or (n18149,1'b0,n18150,n18153,n18161,n18165,n18169,n18174,n18178,n18184,n15561);
and (n18150,n18151,n14237);
or (n18151,1'b0,n15449,n15451,n18152);
and (n18152,n15454,n14455);
and (n18153,n18154,n14137);
or (n18154,1'b0,n18155,n18157,n18159,n15366);
and (n18155,n18156,n13889);
and (n18157,n18158,n13897);
and (n18159,n18160,n13900);
and (n18161,n18162,n14111);
or (n18162,1'b0,n18163,n18164,n18152);
and (n18163,n15367,n13889);
and (n18164,n15525,n13897);
and (n18165,n18166,n14108);
or (n18166,1'b0,n18167,n18168);
and (n18167,n15335,n14235);
and (n18168,n15367,n14455);
and (n18169,n18170,n13950);
or (n18170,1'b0,n18171,n18172,n18173);
and (n18171,n15351,n13889);
and (n18172,n15525,n13900);
and (n18173,n15367,n17806);
and (n18174,n18175,n14239);
or (n18175,1'b0,n18176,n18177,n15550,n15366);
and (n18176,n15430,n13889);
and (n18177,n18160,n13897);
and (n18178,n18179,n17820);
or (n18179,1'b0,n18180,n18182);
and (n18180,n18181,n13900);
wire s0n18181,s1n18181,notn18181;
or (n18181,s0n18181,s1n18181);
not(notn18181,n17823);
and (s0n18181,notn18181,1'b0);
and (s1n18181,n17823,n18125);
and (n18182,n18183,n14131);
wire s0n18183,s1n18183,notn18183;
or (n18183,s0n18183,s1n18183);
not(notn18183,n17823);
and (s0n18183,notn18183,1'b0);
and (s1n18183,n17823,n15367);
and (n18184,n15454,n14448);
wire s0n18185,s1n18185,notn18185;
or (n18185,s0n18185,s1n18185);
not(notn18185,n14631);
and (s0n18185,notn18185,n18186);
and (s1n18185,n14631,n18207);
wire s0n18186,s1n18186,notn18186;
or (n18186,s0n18186,s1n18186);
not(notn18186,n14271);
and (s0n18186,notn18186,n18187);
and (s1n18186,n14271,n18195);
wire s0n18187,s1n18187,notn18187;
or (n18187,s0n18187,s1n18187);
not(notn18187,n14279);
and (s0n18187,notn18187,1'b0);
and (s1n18187,n14279,n18188);
or (n18188,n15565,1'b0,n18189);
and (n18189,n18190,n14367);
or (n18190,n18191,n18194,1'b0);
and (n18191,n18192,n17758);
wire s0n18192,s1n18192,notn18192;
or (n18192,s0n18192,s1n18192);
not(notn18192,n14131);
and (s0n18192,notn18192,n18134);
and (s1n18192,n14131,n18193);
wire s0n18193,s1n18193,notn18193;
or (n18193,s0n18193,s1n18193);
not(notn18193,n17757);
and (s0n18193,notn18193,n15351);
and (s1n18193,n17757,1'b0);
and (n18194,n15446,n17765);
or (n18195,n18196,n18199,1'b0);
and (n18196,n18197,n13907);
wire s0n18197,s1n18197,notn18197;
or (n18197,s0n18197,s1n18197);
not(notn18197,n14125);
and (s0n18197,notn18197,1'b0);
and (s1n18197,n14125,n18198);
wire s0n18198,s1n18198,notn18198;
or (n18198,s0n18198,s1n18198);
not(notn18198,n14563);
and (s0n18198,notn18198,n15568);
and (s1n18198,n14563,n15233);
and (n18199,n18200,n14385);
wire s0n18200,s1n18200,notn18200;
or (n18200,s0n18200,s1n18200);
not(notn18200,n2799);
and (s0n18200,notn18200,1'b0);
and (s1n18200,n2799,n18201);
or (n18201,1'b0,n18202,n18203,n18205);
and (n18202,n18135,n14235);
and (n18203,n18204,n13900);
wire s0n18204,s1n18204,notn18204;
or (n18204,s0n18204,s1n18204);
not(notn18204,n14570);
and (s0n18204,notn18204,n15358);
and (s1n18204,n14570,1'b0);
and (n18205,n18206,n14131);
wire s0n18206,s1n18206,notn18206;
or (n18206,s0n18206,s1n18206);
not(notn18206,n14573);
and (s0n18206,notn18206,n15510);
and (s1n18206,n14573,1'b0);
or (n18207,n18208,n18211,n18212,n18217,n18220,n18222,n18223,1'b0);
and (n18208,n18209,n14237);
or (n18209,1'b0,n18210,n15483);
and (n18210,n15383,n13900);
and (n18211,n15446,n14137);
and (n18212,n18213,n14111);
or (n18213,1'b0,n18214,n18215,n18216,n15524);
and (n18214,n15335,n13889);
and (n18215,n15351,n13897);
and (n18216,n15367,n13900);
and (n18217,n18218,n14108);
or (n18218,1'b0,n15318,n18219,n15524);
and (n18219,n15351,n14243);
and (n18220,n18221,n13950);
or (n18221,1'b0,n15318,n15334,n15350,n15551);
and (n18222,n15559,n14239);
and (n18223,n18224,n17820);
or (n18224,1'b0,n18225,n18227);
and (n18225,n18226,n13900);
wire s0n18226,s1n18226,notn18226;
or (n18226,s0n18226,s1n18226);
not(notn18226,n17818);
and (s0n18226,notn18226,1'b0);
and (s1n18226,n17818,n18135);
and (n18227,n18228,n14131);
wire s0n18228,s1n18228,notn18228;
or (n18228,s0n18228,s1n18228);
not(notn18228,n17823);
and (s0n18228,notn18228,1'b0);
and (s1n18228,n17823,n15351);
and (n18229,n18185,n18230);
or (n18230,n18231,n18343,n18686);
and (n18231,n18232,n18299);
wire s0n18232,s1n18232,notn18232;
or (n18232,s0n18232,s1n18232);
not(notn18232,n14631);
and (s0n18232,notn18232,n18233);
and (s1n18232,n14631,n18263);
wire s0n18233,s1n18233,notn18233;
or (n18233,s0n18233,s1n18233);
not(notn18233,n14271);
and (s0n18233,notn18233,n18234);
and (s1n18233,n14271,n18252);
wire s0n18234,s1n18234,notn18234;
or (n18234,s0n18234,s1n18234);
not(notn18234,n14279);
and (s0n18234,notn18234,1'b0);
and (s1n18234,n14279,n18235);
or (n18235,n18236,n15655,n18240,n18241);
and (n18236,n18237,n14120);
wire s0n18237,s1n18237,notn18237;
or (n18237,s0n18237,s1n18237);
not(notn18237,n14125);
and (s0n18237,notn18237,1'b0);
and (s1n18237,n14125,n18238);
wire s0n18238,s1n18238,notn18238;
or (n18238,s0n18238,s1n18238);
not(notn18238,n14317);
and (s0n18238,notn18238,n18239);
and (s1n18238,n14317,n15646);
and (n18240,n15793,n14365);
and (n18241,n18242,n14367);
or (n18242,n18243,n18247,n18250,1'b0);
and (n18243,n18244,n17758);
wire s0n18244,s1n18244,notn18244;
or (n18244,s0n18244,s1n18244);
not(notn18244,n14131);
and (s0n18244,notn18244,n18245);
and (s1n18244,n14131,n18246);
wire s0n18245,s1n18245,notn18245;
or (n18245,s0n18245,s1n18245);
not(notn18245,n13900);
and (s0n18245,notn18245,1'b0);
and (s1n18245,n13900,n18239);
wire s0n18246,s1n18246,notn18246;
or (n18246,s0n18246,s1n18246);
not(notn18246,n17757);
and (s0n18246,notn18246,n15706);
and (s1n18246,n17757,1'b0);
and (n18247,n18248,n17762);
wire s0n18248,s1n18248,notn18248;
or (n18248,s0n18248,s1n18248);
not(notn18248,n13900);
and (s0n18248,notn18248,1'b0);
and (s1n18248,n13900,n18249);
and (n18250,n18251,n17765);
wire s0n18251,s1n18251,notn18251;
or (n18251,s0n18251,s1n18251);
not(notn18251,n14131);
and (s0n18251,notn18251,n18245);
and (s1n18251,n14131,n15706);
or (n18252,n18253,n18254,n18262,n15764);
and (n18253,n18237,n13907);
and (n18254,n18255,n14385);
wire s0n18255,s1n18255,notn18255;
or (n18255,s0n18255,s1n18255);
not(notn18255,n2799);
and (s0n18255,notn18255,1'b0);
and (s1n18255,n2799,n18256);
or (n18256,1'b0,n18257,n18259,n18260);
and (n18257,n18258,n13889);
wire s0n18258,s1n18258,notn18258;
or (n18258,s0n18258,s1n18258);
not(notn18258,n17767);
and (s0n18258,notn18258,n18239);
and (s1n18258,n17767,1'b0);
and (n18259,n18239,n14243);
and (n18260,n18261,n14131);
wire s0n18261,s1n18261,notn18261;
or (n18261,s0n18261,s1n18261);
not(notn18261,n14573);
and (s0n18261,notn18261,n15817);
and (s1n18261,n14573,1'b0);
and (n18262,n15793,n14381);
or (n18263,1'b0,n18264,n18267,n18275,n18279,n18283,n18288,n18292,n18298,n15900);
and (n18264,n18265,n14237);
or (n18265,1'b0,n15788,n15790,n18266);
and (n18266,n15793,n14455);
and (n18267,n18268,n14137);
or (n18268,1'b0,n18269,n18271,n18273,n15705);
and (n18269,n18270,n13889);
and (n18271,n18272,n13897);
and (n18273,n18274,n13900);
and (n18275,n18276,n14111);
or (n18276,1'b0,n18277,n18278,n18266);
and (n18277,n15706,n13889);
and (n18278,n15864,n13897);
and (n18279,n18280,n14108);
or (n18280,1'b0,n18281,n18282);
and (n18281,n15674,n14235);
and (n18282,n15706,n14455);
and (n18283,n18284,n13950);
or (n18284,1'b0,n18285,n18286,n18287);
and (n18285,n15690,n13889);
and (n18286,n15864,n13900);
and (n18287,n15706,n17806);
and (n18288,n18289,n14239);
or (n18289,1'b0,n18290,n18291,n15889,n15705);
and (n18290,n15769,n13889);
and (n18291,n18274,n13897);
and (n18292,n18293,n17820);
or (n18293,1'b0,n18294,n18296);
and (n18294,n18295,n13900);
wire s0n18295,s1n18295,notn18295;
or (n18295,s0n18295,s1n18295);
not(notn18295,n17823);
and (s0n18295,notn18295,1'b0);
and (s1n18295,n17823,n18239);
and (n18296,n18297,n14131);
wire s0n18297,s1n18297,notn18297;
or (n18297,s0n18297,s1n18297);
not(notn18297,n17823);
and (s0n18297,notn18297,1'b0);
and (s1n18297,n17823,n15706);
and (n18298,n15793,n14448);
wire s0n18299,s1n18299,notn18299;
or (n18299,s0n18299,s1n18299);
not(notn18299,n14631);
and (s0n18299,notn18299,n18300);
and (s1n18299,n14631,n18321);
wire s0n18300,s1n18300,notn18300;
or (n18300,s0n18300,s1n18300);
not(notn18300,n14271);
and (s0n18300,notn18300,n18301);
and (s1n18300,n14271,n18309);
wire s0n18301,s1n18301,notn18301;
or (n18301,s0n18301,s1n18301);
not(notn18301,n14279);
and (s0n18301,notn18301,1'b0);
and (s1n18301,n14279,n18302);
or (n18302,n15904,1'b0,n18303);
and (n18303,n18304,n14367);
or (n18304,n18305,n18308,1'b0);
and (n18305,n18306,n17758);
wire s0n18306,s1n18306,notn18306;
or (n18306,s0n18306,s1n18306);
not(notn18306,n14131);
and (s0n18306,notn18306,n18248);
and (s1n18306,n14131,n18307);
wire s0n18307,s1n18307,notn18307;
or (n18307,s0n18307,s1n18307);
not(notn18307,n17757);
and (s0n18307,notn18307,n15690);
and (s1n18307,n17757,1'b0);
and (n18308,n15785,n17765);
or (n18309,n18310,n18313,1'b0);
and (n18310,n18311,n13907);
wire s0n18311,s1n18311,notn18311;
or (n18311,s0n18311,s1n18311);
not(notn18311,n14125);
and (s0n18311,notn18311,1'b0);
and (s1n18311,n14125,n18312);
wire s0n18312,s1n18312,notn18312;
or (n18312,s0n18312,s1n18312);
not(notn18312,n14563);
and (s0n18312,notn18312,n15907);
and (s1n18312,n14563,n15573);
and (n18313,n18314,n14385);
wire s0n18314,s1n18314,notn18314;
or (n18314,s0n18314,s1n18314);
not(notn18314,n2799);
and (s0n18314,notn18314,1'b0);
and (s1n18314,n2799,n18315);
or (n18315,1'b0,n18316,n18317,n18319);
and (n18316,n18249,n14235);
and (n18317,n18318,n13900);
wire s0n18318,s1n18318,notn18318;
or (n18318,s0n18318,s1n18318);
not(notn18318,n14570);
and (s0n18318,notn18318,n15697);
and (s1n18318,n14570,1'b0);
and (n18319,n18320,n14131);
wire s0n18320,s1n18320,notn18320;
or (n18320,s0n18320,s1n18320);
not(notn18320,n14573);
and (s0n18320,notn18320,n15849);
and (s1n18320,n14573,1'b0);
or (n18321,n18322,n18325,n18326,n18331,n18334,n18336,n18337,1'b0);
and (n18322,n18323,n14237);
or (n18323,1'b0,n18324,n15822);
and (n18324,n15722,n13900);
and (n18325,n15785,n14137);
and (n18326,n18327,n14111);
or (n18327,1'b0,n18328,n18329,n18330,n15863);
and (n18328,n15674,n13889);
and (n18329,n15690,n13897);
and (n18330,n15706,n13900);
and (n18331,n18332,n14108);
or (n18332,1'b0,n15657,n18333,n15863);
and (n18333,n15690,n14243);
and (n18334,n18335,n13950);
or (n18335,1'b0,n15657,n15673,n15689,n15890);
and (n18336,n15898,n14239);
and (n18337,n18338,n17820);
or (n18338,1'b0,n18339,n18341);
and (n18339,n18340,n13900);
wire s0n18340,s1n18340,notn18340;
or (n18340,s0n18340,s1n18340);
not(notn18340,n17818);
and (s0n18340,notn18340,1'b0);
and (s1n18340,n17818,n18249);
and (n18341,n18342,n14131);
wire s0n18342,s1n18342,notn18342;
or (n18342,s0n18342,s1n18342);
not(notn18342,n17823);
and (s0n18342,notn18342,1'b0);
and (s1n18342,n17823,n15690);
and (n18343,n18299,n18344);
or (n18344,n18345,n18457,n18685);
and (n18345,n18346,n18413);
wire s0n18346,s1n18346,notn18346;
or (n18346,s0n18346,s1n18346);
not(notn18346,n14631);
and (s0n18346,notn18346,n18347);
and (s1n18346,n14631,n18377);
wire s0n18347,s1n18347,notn18347;
or (n18347,s0n18347,s1n18347);
not(notn18347,n14271);
and (s0n18347,notn18347,n18348);
and (s1n18347,n14271,n18366);
wire s0n18348,s1n18348,notn18348;
or (n18348,s0n18348,s1n18348);
not(notn18348,n14279);
and (s0n18348,notn18348,1'b0);
and (s1n18348,n14279,n18349);
or (n18349,n18350,n15995,n18354,n18355);
and (n18350,n18351,n14120);
wire s0n18351,s1n18351,notn18351;
or (n18351,s0n18351,s1n18351);
not(notn18351,n14125);
and (s0n18351,notn18351,1'b0);
and (s1n18351,n14125,n18352);
wire s0n18352,s1n18352,notn18352;
or (n18352,s0n18352,s1n18352);
not(notn18352,n14317);
and (s0n18352,notn18352,n18353);
and (s1n18352,n14317,n15986);
and (n18354,n16133,n14365);
and (n18355,n18356,n14367);
or (n18356,n18357,n18361,n18364,1'b0);
and (n18357,n18358,n17758);
wire s0n18358,s1n18358,notn18358;
or (n18358,s0n18358,s1n18358);
not(notn18358,n14131);
and (s0n18358,notn18358,n18359);
and (s1n18358,n14131,n18360);
wire s0n18359,s1n18359,notn18359;
or (n18359,s0n18359,s1n18359);
not(notn18359,n13900);
and (s0n18359,notn18359,1'b0);
and (s1n18359,n13900,n18353);
wire s0n18360,s1n18360,notn18360;
or (n18360,s0n18360,s1n18360);
not(notn18360,n17757);
and (s0n18360,notn18360,n16046);
and (s1n18360,n17757,1'b0);
and (n18361,n18362,n17762);
wire s0n18362,s1n18362,notn18362;
or (n18362,s0n18362,s1n18362);
not(notn18362,n13900);
and (s0n18362,notn18362,1'b0);
and (s1n18362,n13900,n18363);
and (n18364,n18365,n17765);
wire s0n18365,s1n18365,notn18365;
or (n18365,s0n18365,s1n18365);
not(notn18365,n14131);
and (s0n18365,notn18365,n18359);
and (s1n18365,n14131,n16046);
or (n18366,n18367,n18368,n18376,n16104);
and (n18367,n18351,n13907);
and (n18368,n18369,n14385);
wire s0n18369,s1n18369,notn18369;
or (n18369,s0n18369,s1n18369);
not(notn18369,n2799);
and (s0n18369,notn18369,1'b0);
and (s1n18369,n2799,n18370);
or (n18370,1'b0,n18371,n18373,n18374);
and (n18371,n18372,n13889);
wire s0n18372,s1n18372,notn18372;
or (n18372,s0n18372,s1n18372);
not(notn18372,n17767);
and (s0n18372,notn18372,n18353);
and (s1n18372,n17767,1'b0);
and (n18373,n18353,n14243);
and (n18374,n18375,n14131);
wire s0n18375,s1n18375,notn18375;
or (n18375,s0n18375,s1n18375);
not(notn18375,n14573);
and (s0n18375,notn18375,n16157);
and (s1n18375,n14573,1'b0);
and (n18376,n16133,n14381);
or (n18377,1'b0,n18378,n18381,n18389,n18393,n18397,n18402,n18406,n18412,n16240);
and (n18378,n18379,n14237);
or (n18379,1'b0,n16128,n16130,n18380);
and (n18380,n16133,n14455);
and (n18381,n18382,n14137);
or (n18382,1'b0,n18383,n18385,n18387,n16045);
and (n18383,n18384,n13889);
and (n18385,n18386,n13897);
and (n18387,n18388,n13900);
and (n18389,n18390,n14111);
or (n18390,1'b0,n18391,n18392,n18380);
and (n18391,n16046,n13889);
and (n18392,n16204,n13897);
and (n18393,n18394,n14108);
or (n18394,1'b0,n18395,n18396);
and (n18395,n16014,n14235);
and (n18396,n16046,n14455);
and (n18397,n18398,n13950);
or (n18398,1'b0,n18399,n18400,n18401);
and (n18399,n16030,n13889);
and (n18400,n16204,n13900);
and (n18401,n16046,n17806);
and (n18402,n18403,n14239);
or (n18403,1'b0,n18404,n18405,n16229,n16045);
and (n18404,n16109,n13889);
and (n18405,n18388,n13897);
and (n18406,n18407,n17820);
or (n18407,1'b0,n18408,n18410);
and (n18408,n18409,n13900);
wire s0n18409,s1n18409,notn18409;
or (n18409,s0n18409,s1n18409);
not(notn18409,n17823);
and (s0n18409,notn18409,1'b0);
and (s1n18409,n17823,n18353);
and (n18410,n18411,n14131);
wire s0n18411,s1n18411,notn18411;
or (n18411,s0n18411,s1n18411);
not(notn18411,n17823);
and (s0n18411,notn18411,1'b0);
and (s1n18411,n17823,n16046);
and (n18412,n16133,n14448);
wire s0n18413,s1n18413,notn18413;
or (n18413,s0n18413,s1n18413);
not(notn18413,n14631);
and (s0n18413,notn18413,n18414);
and (s1n18413,n14631,n18435);
wire s0n18414,s1n18414,notn18414;
or (n18414,s0n18414,s1n18414);
not(notn18414,n14271);
and (s0n18414,notn18414,n18415);
and (s1n18414,n14271,n18423);
wire s0n18415,s1n18415,notn18415;
or (n18415,s0n18415,s1n18415);
not(notn18415,n14279);
and (s0n18415,notn18415,1'b0);
and (s1n18415,n14279,n18416);
or (n18416,n16244,1'b0,n18417);
and (n18417,n18418,n14367);
or (n18418,n18419,n18422,1'b0);
and (n18419,n18420,n17758);
wire s0n18420,s1n18420,notn18420;
or (n18420,s0n18420,s1n18420);
not(notn18420,n14131);
and (s0n18420,notn18420,n18362);
and (s1n18420,n14131,n18421);
wire s0n18421,s1n18421,notn18421;
or (n18421,s0n18421,s1n18421);
not(notn18421,n17757);
and (s0n18421,notn18421,n16030);
and (s1n18421,n17757,1'b0);
and (n18422,n16125,n17765);
or (n18423,n18424,n18427,1'b0);
and (n18424,n18425,n13907);
wire s0n18425,s1n18425,notn18425;
or (n18425,s0n18425,s1n18425);
not(notn18425,n14125);
and (s0n18425,notn18425,1'b0);
and (s1n18425,n14125,n18426);
wire s0n18426,s1n18426,notn18426;
or (n18426,s0n18426,s1n18426);
not(notn18426,n14563);
and (s0n18426,notn18426,n16247);
and (s1n18426,n14563,n15912);
and (n18427,n18428,n14385);
wire s0n18428,s1n18428,notn18428;
or (n18428,s0n18428,s1n18428);
not(notn18428,n2799);
and (s0n18428,notn18428,1'b0);
and (s1n18428,n2799,n18429);
or (n18429,1'b0,n18430,n18431,n18433);
and (n18430,n18363,n14235);
and (n18431,n18432,n13900);
wire s0n18432,s1n18432,notn18432;
or (n18432,s0n18432,s1n18432);
not(notn18432,n14570);
and (s0n18432,notn18432,n16037);
and (s1n18432,n14570,1'b0);
and (n18433,n18434,n14131);
wire s0n18434,s1n18434,notn18434;
or (n18434,s0n18434,s1n18434);
not(notn18434,n14573);
and (s0n18434,notn18434,n16189);
and (s1n18434,n14573,1'b0);
or (n18435,n18436,n18439,n18440,n18445,n18448,n18450,n18451,1'b0);
and (n18436,n18437,n14237);
or (n18437,1'b0,n18438,n16162);
and (n18438,n16062,n13900);
and (n18439,n16125,n14137);
and (n18440,n18441,n14111);
or (n18441,1'b0,n18442,n18443,n18444,n16203);
and (n18442,n16014,n13889);
and (n18443,n16030,n13897);
and (n18444,n16046,n13900);
and (n18445,n18446,n14108);
or (n18446,1'b0,n15997,n18447,n16203);
and (n18447,n16030,n14243);
and (n18448,n18449,n13950);
or (n18449,1'b0,n15997,n16013,n16029,n16230);
and (n18450,n16238,n14239);
and (n18451,n18452,n17820);
or (n18452,1'b0,n18453,n18455);
and (n18453,n18454,n13900);
wire s0n18454,s1n18454,notn18454;
or (n18454,s0n18454,s1n18454);
not(notn18454,n17818);
and (s0n18454,notn18454,1'b0);
and (s1n18454,n17818,n18363);
and (n18455,n18456,n14131);
wire s0n18456,s1n18456,notn18456;
or (n18456,s0n18456,s1n18456);
not(notn18456,n17823);
and (s0n18456,notn18456,1'b0);
and (s1n18456,n17823,n16030);
and (n18457,n18413,n18458);
or (n18458,n18459,n18571,n18684);
and (n18459,n18460,n18527);
wire s0n18460,s1n18460,notn18460;
or (n18460,s0n18460,s1n18460);
not(notn18460,n14631);
and (s0n18460,notn18460,n18461);
and (s1n18460,n14631,n18491);
wire s0n18461,s1n18461,notn18461;
or (n18461,s0n18461,s1n18461);
not(notn18461,n14271);
and (s0n18461,notn18461,n18462);
and (s1n18461,n14271,n18480);
wire s0n18462,s1n18462,notn18462;
or (n18462,s0n18462,s1n18462);
not(notn18462,n14279);
and (s0n18462,notn18462,1'b0);
and (s1n18462,n14279,n18463);
or (n18463,n18464,n16335,n18468,n18469);
and (n18464,n18465,n14120);
wire s0n18465,s1n18465,notn18465;
or (n18465,s0n18465,s1n18465);
not(notn18465,n14125);
and (s0n18465,notn18465,1'b0);
and (s1n18465,n14125,n18466);
wire s0n18466,s1n18466,notn18466;
or (n18466,s0n18466,s1n18466);
not(notn18466,n14317);
and (s0n18466,notn18466,n18467);
and (s1n18466,n14317,n16326);
and (n18468,n16473,n14365);
and (n18469,n18470,n14367);
or (n18470,n18471,n18475,n18478,1'b0);
and (n18471,n18472,n17758);
wire s0n18472,s1n18472,notn18472;
or (n18472,s0n18472,s1n18472);
not(notn18472,n14131);
and (s0n18472,notn18472,n18473);
and (s1n18472,n14131,n18474);
wire s0n18473,s1n18473,notn18473;
or (n18473,s0n18473,s1n18473);
not(notn18473,n13900);
and (s0n18473,notn18473,1'b0);
and (s1n18473,n13900,n18467);
wire s0n18474,s1n18474,notn18474;
or (n18474,s0n18474,s1n18474);
not(notn18474,n17757);
and (s0n18474,notn18474,n16386);
and (s1n18474,n17757,1'b0);
and (n18475,n18476,n17762);
wire s0n18476,s1n18476,notn18476;
or (n18476,s0n18476,s1n18476);
not(notn18476,n13900);
and (s0n18476,notn18476,1'b0);
and (s1n18476,n13900,n18477);
and (n18478,n18479,n17765);
wire s0n18479,s1n18479,notn18479;
or (n18479,s0n18479,s1n18479);
not(notn18479,n14131);
and (s0n18479,notn18479,n18473);
and (s1n18479,n14131,n16386);
or (n18480,n18481,n18482,n18490,n16444);
and (n18481,n18465,n13907);
and (n18482,n18483,n14385);
wire s0n18483,s1n18483,notn18483;
or (n18483,s0n18483,s1n18483);
not(notn18483,n2799);
and (s0n18483,notn18483,1'b0);
and (s1n18483,n2799,n18484);
or (n18484,1'b0,n18485,n18487,n18488);
and (n18485,n18486,n13889);
wire s0n18486,s1n18486,notn18486;
or (n18486,s0n18486,s1n18486);
not(notn18486,n17767);
and (s0n18486,notn18486,n18467);
and (s1n18486,n17767,1'b0);
and (n18487,n18467,n14243);
and (n18488,n18489,n14131);
wire s0n18489,s1n18489,notn18489;
or (n18489,s0n18489,s1n18489);
not(notn18489,n14573);
and (s0n18489,notn18489,n16497);
and (s1n18489,n14573,1'b0);
and (n18490,n16473,n14381);
or (n18491,1'b0,n18492,n18495,n18503,n18507,n18511,n18516,n18520,n18526,n16580);
and (n18492,n18493,n14237);
or (n18493,1'b0,n16468,n16470,n18494);
and (n18494,n16473,n14455);
and (n18495,n18496,n14137);
or (n18496,1'b0,n18497,n18499,n18501,n16385);
and (n18497,n18498,n13889);
and (n18499,n18500,n13897);
and (n18501,n18502,n13900);
and (n18503,n18504,n14111);
or (n18504,1'b0,n18505,n18506,n18494);
and (n18505,n16386,n13889);
and (n18506,n16544,n13897);
and (n18507,n18508,n14108);
or (n18508,1'b0,n18509,n18510);
and (n18509,n16354,n14235);
and (n18510,n16386,n14455);
and (n18511,n18512,n13950);
or (n18512,1'b0,n18513,n18514,n18515);
and (n18513,n16370,n13889);
and (n18514,n16544,n13900);
and (n18515,n16386,n17806);
and (n18516,n18517,n14239);
or (n18517,1'b0,n18518,n18519,n16569,n16385);
and (n18518,n16449,n13889);
and (n18519,n18502,n13897);
and (n18520,n18521,n17820);
or (n18521,1'b0,n18522,n18524);
and (n18522,n18523,n13900);
wire s0n18523,s1n18523,notn18523;
or (n18523,s0n18523,s1n18523);
not(notn18523,n17823);
and (s0n18523,notn18523,1'b0);
and (s1n18523,n17823,n18467);
and (n18524,n18525,n14131);
wire s0n18525,s1n18525,notn18525;
or (n18525,s0n18525,s1n18525);
not(notn18525,n17823);
and (s0n18525,notn18525,1'b0);
and (s1n18525,n17823,n16386);
and (n18526,n16473,n14448);
wire s0n18527,s1n18527,notn18527;
or (n18527,s0n18527,s1n18527);
not(notn18527,n14631);
and (s0n18527,notn18527,n18528);
and (s1n18527,n14631,n18549);
wire s0n18528,s1n18528,notn18528;
or (n18528,s0n18528,s1n18528);
not(notn18528,n14271);
and (s0n18528,notn18528,n18529);
and (s1n18528,n14271,n18537);
wire s0n18529,s1n18529,notn18529;
or (n18529,s0n18529,s1n18529);
not(notn18529,n14279);
and (s0n18529,notn18529,1'b0);
and (s1n18529,n14279,n18530);
or (n18530,n16584,1'b0,n18531);
and (n18531,n18532,n14367);
or (n18532,n18533,n18536,1'b0);
and (n18533,n18534,n17758);
wire s0n18534,s1n18534,notn18534;
or (n18534,s0n18534,s1n18534);
not(notn18534,n14131);
and (s0n18534,notn18534,n18476);
and (s1n18534,n14131,n18535);
wire s0n18535,s1n18535,notn18535;
or (n18535,s0n18535,s1n18535);
not(notn18535,n17757);
and (s0n18535,notn18535,n16370);
and (s1n18535,n17757,1'b0);
and (n18536,n16465,n17765);
or (n18537,n18538,n18541,1'b0);
and (n18538,n18539,n13907);
wire s0n18539,s1n18539,notn18539;
or (n18539,s0n18539,s1n18539);
not(notn18539,n14125);
and (s0n18539,notn18539,1'b0);
and (s1n18539,n14125,n18540);
wire s0n18540,s1n18540,notn18540;
or (n18540,s0n18540,s1n18540);
not(notn18540,n14563);
and (s0n18540,notn18540,n16587);
and (s1n18540,n14563,n16252);
and (n18541,n18542,n14385);
wire s0n18542,s1n18542,notn18542;
or (n18542,s0n18542,s1n18542);
not(notn18542,n2799);
and (s0n18542,notn18542,1'b0);
and (s1n18542,n2799,n18543);
or (n18543,1'b0,n18544,n18545,n18547);
and (n18544,n18477,n14235);
and (n18545,n18546,n13900);
wire s0n18546,s1n18546,notn18546;
or (n18546,s0n18546,s1n18546);
not(notn18546,n14570);
and (s0n18546,notn18546,n16377);
and (s1n18546,n14570,1'b0);
and (n18547,n18548,n14131);
wire s0n18548,s1n18548,notn18548;
or (n18548,s0n18548,s1n18548);
not(notn18548,n14573);
and (s0n18548,notn18548,n16529);
and (s1n18548,n14573,1'b0);
or (n18549,n18550,n18553,n18554,n18559,n18562,n18564,n18565,1'b0);
and (n18550,n18551,n14237);
or (n18551,1'b0,n18552,n16502);
and (n18552,n16402,n13900);
and (n18553,n16465,n14137);
and (n18554,n18555,n14111);
or (n18555,1'b0,n18556,n18557,n18558,n16543);
and (n18556,n16354,n13889);
and (n18557,n16370,n13897);
and (n18558,n16386,n13900);
and (n18559,n18560,n14108);
or (n18560,1'b0,n16337,n18561,n16543);
and (n18561,n16370,n14243);
and (n18562,n18563,n13950);
or (n18563,1'b0,n16337,n16353,n16369,n16570);
and (n18564,n16578,n14239);
and (n18565,n18566,n17820);
or (n18566,1'b0,n18567,n18569);
and (n18567,n18568,n13900);
wire s0n18568,s1n18568,notn18568;
or (n18568,s0n18568,s1n18568);
not(notn18568,n17818);
and (s0n18568,notn18568,1'b0);
and (s1n18568,n17818,n18477);
and (n18569,n18570,n14131);
wire s0n18570,s1n18570,notn18570;
or (n18570,s0n18570,s1n18570);
not(notn18570,n17823);
and (s0n18570,notn18570,1'b0);
and (s1n18570,n17823,n16370);
and (n18571,n18527,n18572);
and (n18572,n18573,n18640);
wire s0n18573,s1n18573,notn18573;
or (n18573,s0n18573,s1n18573);
not(notn18573,n14631);
and (s0n18573,notn18573,n18574);
and (s1n18573,n14631,n18604);
wire s0n18574,s1n18574,notn18574;
or (n18574,s0n18574,s1n18574);
not(notn18574,n14271);
and (s0n18574,notn18574,n18575);
and (s1n18574,n14271,n18593);
wire s0n18575,s1n18575,notn18575;
or (n18575,s0n18575,s1n18575);
not(notn18575,n14279);
and (s0n18575,notn18575,1'b0);
and (s1n18575,n14279,n18576);
or (n18576,n18577,n16703,n18581,n18582);
and (n18577,n18578,n14120);
wire s0n18578,s1n18578,notn18578;
or (n18578,s0n18578,s1n18578);
not(notn18578,n14125);
and (s0n18578,notn18578,1'b0);
and (s1n18578,n14125,n18579);
wire s0n18579,s1n18579,notn18579;
or (n18579,s0n18579,s1n18579);
not(notn18579,n14317);
and (s0n18579,notn18579,n18580);
and (s1n18579,n14317,n16694);
and (n18581,n16841,n14365);
and (n18582,n18583,n14367);
or (n18583,n18584,n18588,n18591,1'b0);
and (n18584,n18585,n17758);
wire s0n18585,s1n18585,notn18585;
or (n18585,s0n18585,s1n18585);
not(notn18585,n14131);
and (s0n18585,notn18585,n18586);
and (s1n18585,n14131,n18587);
wire s0n18586,s1n18586,notn18586;
or (n18586,s0n18586,s1n18586);
not(notn18586,n13900);
and (s0n18586,notn18586,1'b0);
and (s1n18586,n13900,n18580);
wire s0n18587,s1n18587,notn18587;
or (n18587,s0n18587,s1n18587);
not(notn18587,n17757);
and (s0n18587,notn18587,n16754);
and (s1n18587,n17757,1'b0);
and (n18588,n18589,n17762);
wire s0n18589,s1n18589,notn18589;
or (n18589,s0n18589,s1n18589);
not(notn18589,n13900);
and (s0n18589,notn18589,1'b0);
and (s1n18589,n13900,n18590);
and (n18591,n18592,n17765);
wire s0n18592,s1n18592,notn18592;
or (n18592,s0n18592,s1n18592);
not(notn18592,n14131);
and (s0n18592,notn18592,n18586);
and (s1n18592,n14131,n16754);
or (n18593,n18594,n18595,n18603,n16812);
and (n18594,n18578,n13907);
and (n18595,n18596,n14385);
wire s0n18596,s1n18596,notn18596;
or (n18596,s0n18596,s1n18596);
not(notn18596,n2799);
and (s0n18596,notn18596,1'b0);
and (s1n18596,n2799,n18597);
or (n18597,1'b0,n18598,n18600,n18601);
and (n18598,n18599,n13889);
wire s0n18599,s1n18599,notn18599;
or (n18599,s0n18599,s1n18599);
not(notn18599,n17767);
and (s0n18599,notn18599,n18580);
and (s1n18599,n17767,1'b0);
and (n18600,n18580,n14243);
and (n18601,n18602,n14131);
wire s0n18602,s1n18602,notn18602;
or (n18602,s0n18602,s1n18602);
not(notn18602,n14573);
and (s0n18602,notn18602,n16865);
and (s1n18602,n14573,1'b0);
and (n18603,n16841,n14381);
or (n18604,1'b0,n18605,n18608,n18616,n18620,n18624,n18629,n18633,n18639,n16948);
and (n18605,n18606,n14237);
or (n18606,1'b0,n16836,n16838,n18607);
and (n18607,n16841,n14455);
and (n18608,n18609,n14137);
or (n18609,1'b0,n18610,n18612,n18614,n16753);
and (n18610,n18611,n13889);
and (n18612,n18613,n13897);
and (n18614,n18615,n13900);
and (n18616,n18617,n14111);
or (n18617,1'b0,n18618,n18619,n18607);
and (n18618,n16754,n13889);
and (n18619,n16912,n13897);
and (n18620,n18621,n14108);
or (n18621,1'b0,n18622,n18623);
and (n18622,n16722,n14235);
and (n18623,n16754,n14455);
and (n18624,n18625,n13950);
or (n18625,1'b0,n18626,n18627,n18628);
and (n18626,n16738,n13889);
and (n18627,n16912,n13900);
and (n18628,n16754,n17806);
and (n18629,n18630,n14239);
or (n18630,1'b0,n18631,n18632,n16937,n16753);
and (n18631,n16817,n13889);
and (n18632,n18615,n13897);
and (n18633,n18634,n17820);
or (n18634,1'b0,n18635,n18637);
and (n18635,n18636,n13900);
wire s0n18636,s1n18636,notn18636;
or (n18636,s0n18636,s1n18636);
not(notn18636,n17823);
and (s0n18636,notn18636,1'b0);
and (s1n18636,n17823,n18580);
and (n18637,n18638,n14131);
wire s0n18638,s1n18638,notn18638;
or (n18638,s0n18638,s1n18638);
not(notn18638,n17823);
and (s0n18638,notn18638,1'b0);
and (s1n18638,n17823,n16754);
and (n18639,n16841,n14448);
wire s0n18640,s1n18640,notn18640;
or (n18640,s0n18640,s1n18640);
not(notn18640,n14631);
and (s0n18640,notn18640,n18641);
and (s1n18640,n14631,n18662);
wire s0n18641,s1n18641,notn18641;
or (n18641,s0n18641,s1n18641);
not(notn18641,n14271);
and (s0n18641,notn18641,n18642);
and (s1n18641,n14271,n18650);
wire s0n18642,s1n18642,notn18642;
or (n18642,s0n18642,s1n18642);
not(notn18642,n14279);
and (s0n18642,notn18642,1'b0);
and (s1n18642,n14279,n18643);
or (n18643,n16952,1'b0,n18644);
and (n18644,n18645,n14367);
or (n18645,n18646,n18649,1'b0);
and (n18646,n18647,n17758);
wire s0n18647,s1n18647,notn18647;
or (n18647,s0n18647,s1n18647);
not(notn18647,n14131);
and (s0n18647,notn18647,n18589);
and (s1n18647,n14131,n18648);
wire s0n18648,s1n18648,notn18648;
or (n18648,s0n18648,s1n18648);
not(notn18648,n17757);
and (s0n18648,notn18648,n16738);
and (s1n18648,n17757,1'b0);
and (n18649,n16833,n17765);
or (n18650,n18651,n18654,1'b0);
and (n18651,n18652,n13907);
wire s0n18652,s1n18652,notn18652;
or (n18652,s0n18652,s1n18652);
not(notn18652,n14125);
and (s0n18652,notn18652,1'b0);
and (s1n18652,n14125,n18653);
wire s0n18653,s1n18653,notn18653;
or (n18653,s0n18653,s1n18653);
not(notn18653,n14563);
and (s0n18653,notn18653,n16955);
and (s1n18653,n14563,n16592);
and (n18654,n18655,n14385);
wire s0n18655,s1n18655,notn18655;
or (n18655,s0n18655,s1n18655);
not(notn18655,n2799);
and (s0n18655,notn18655,1'b0);
and (s1n18655,n2799,n18656);
or (n18656,1'b0,n18657,n18658,n18660);
and (n18657,n18590,n14235);
and (n18658,n18659,n13900);
wire s0n18659,s1n18659,notn18659;
or (n18659,s0n18659,s1n18659);
not(notn18659,n14570);
and (s0n18659,notn18659,n16745);
and (s1n18659,n14570,1'b0);
and (n18660,n18661,n14131);
wire s0n18661,s1n18661,notn18661;
or (n18661,s0n18661,s1n18661);
not(notn18661,n14573);
and (s0n18661,notn18661,n16897);
and (s1n18661,n14573,1'b0);
or (n18662,n18663,n18666,n18667,n18672,n18675,n18677,n18678,1'b0);
and (n18663,n18664,n14237);
or (n18664,1'b0,n18665,n16870);
and (n18665,n16770,n13900);
and (n18666,n16833,n14137);
and (n18667,n18668,n14111);
or (n18668,1'b0,n18669,n18670,n18671,n16911);
and (n18669,n16722,n13889);
and (n18670,n16738,n13897);
and (n18671,n16754,n13900);
and (n18672,n18673,n14108);
or (n18673,1'b0,n16705,n18674,n16911);
and (n18674,n16738,n14243);
and (n18675,n18676,n13950);
or (n18676,1'b0,n16705,n16721,n16737,n16938);
and (n18677,n16946,n14239);
and (n18678,n18679,n17820);
or (n18679,1'b0,n18680,n18682);
and (n18680,n18681,n13900);
wire s0n18681,s1n18681,notn18681;
or (n18681,s0n18681,s1n18681);
not(notn18681,n17818);
and (s0n18681,notn18681,1'b0);
and (s1n18681,n17818,n18590);
and (n18682,n18683,n14131);
wire s0n18683,s1n18683,notn18683;
or (n18683,s0n18683,s1n18683);
not(notn18683,n17823);
and (s0n18683,notn18683,1'b0);
and (s1n18683,n17823,n16738);
and (n18684,n18460,n18572);
and (n18685,n18346,n18458);
and (n18686,n18232,n18344);
and (n18687,n18118,n18230);
and (n18688,n17995,n18116);
and (n18689,n17881,n17993);
wire s0n18690,s1n18690,notn18690;
or (n18690,s0n18690,s1n18690);
not(notn18690,n14631);
and (s0n18690,notn18690,n18691);
and (s1n18690,n14631,n18699);
wire s0n18691,s1n18691,notn18691;
or (n18691,s0n18691,s1n18691);
not(notn18691,n14271);
and (s0n18691,notn18691,n18692);
and (s1n18691,n14271,n18695);
and (n18692,n18693,n14279);
or (n18693,1'b0,n17031,n18694);
and (n18694,n17766,n14367);
or (n18695,1'b0,n18696,n14382);
and (n18696,n18697,n14385);
and (n18697,n18698,n2799);
and (n18698,n17767,n13889);
or (n18699,n18700,1'b0,n18701,n18703,n17039);
and (n18700,n14454,n14237);
and (n18701,n17036,n18702);
or (n18702,n14239,n14137);
and (n18703,n18704,n17820);
or (n18704,n14454,n18705,n18706);
and (n18705,n17832,n13900);
and (n18706,n17824,n14131);
wire s0n18707,s1n18707,notn18707;
or (n18707,s0n18707,s1n18707);
not(notn18707,n19059);
and (s0n18707,notn18707,n18708);
and (s1n18707,n19059,n18756);
xor (n18708,n18709,n18754);
xor (n18709,n18710,n18737);
wire s0n18710,s1n18710,notn18710;
or (n18710,s0n18710,s1n18710);
not(notn18710,n14631);
and (s0n18710,notn18710,n18711);
and (s1n18710,n14631,n18727);
wire s0n18711,s1n18711,notn18711;
or (n18711,s0n18711,s1n18711);
not(notn18711,n14271);
and (s0n18711,notn18711,n18712);
and (s1n18711,n14271,n18719);
wire s0n18712,s1n18712,notn18712;
or (n18712,s0n18712,s1n18712);
not(notn18712,n14279);
and (s0n18712,notn18712,1'b0);
and (s1n18712,n14279,n18713);
and (n18713,n18714,n14367);
wire s0n18714,s1n18714,notn18714;
or (n18714,s0n18714,s1n18714);
not(notn18714,n18715);
and (s0n18714,notn18714,1'b0);
and (s1n18714,n18715,n14280);
and (n18715,n14211,n18716);
and (n18716,n14131,n18717);
not (n18717,n18718);
and (n18718,n17757,n14368);
and (n18719,n18720,n14385);
wire s0n18720,s1n18720,notn18720;
or (n18720,s0n18720,s1n18720);
not(notn18720,n2799);
and (s0n18720,notn18720,1'b0);
and (s1n18720,n2799,n18721);
or (n18721,1'b0,n18722,n18723,n18725);
and (n18722,n14507,n13897);
and (n18723,n18724,n13900);
wire s0n18724,s1n18724,notn18724;
or (n18724,s0n18724,s1n18724);
not(notn18724,n14570);
and (s0n18724,notn18724,n14287);
and (s1n18724,n14570,1'b0);
and (n18725,n18726,n14131);
wire s0n18726,s1n18726,notn18726;
or (n18726,s0n18726,s1n18726);
not(notn18726,n14573);
and (s0n18726,notn18726,n14482);
and (s1n18726,n14573,1'b0);
or (n18727,n18728,n18729,n18732,n18733,n18734,1'b0);
and (n18728,n17069,n14237);
and (n18729,n18730,n14111);
or (n18730,n17803,n18731,n17804,1'b0);
and (n18731,n14297,n13897);
and (n18732,n17864,n13950);
and (n18733,n14246,n14239);
and (n18734,n18735,n17820);
and (n18735,n18736,n14131);
wire s0n18736,s1n18736,notn18736;
or (n18736,s0n18736,s1n18736);
not(notn18736,n17823);
and (s0n18736,notn18736,1'b0);
and (s1n18736,n17823,n14280);
wire s0n18737,s1n18737,notn18737;
or (n18737,s0n18737,s1n18737);
not(notn18737,n14631);
and (s0n18737,notn18737,n18738);
and (s1n18737,n14631,n18751);
wire s0n18738,s1n18738,notn18738;
or (n18738,s0n18738,s1n18738);
not(notn18738,n14271);
and (s0n18738,notn18738,n18739);
and (s1n18738,n14271,n18742);
wire s0n18739,s1n18739,notn18739;
or (n18739,s0n18739,s1n18739);
not(notn18739,n14279);
and (s0n18739,notn18739,1'b0);
and (s1n18739,n14279,n18740);
and (n18740,n18741,n14367);
wire s0n18741,s1n18741,notn18741;
or (n18741,s0n18741,s1n18741);
not(notn18741,n18715);
and (s0n18741,notn18741,1'b0);
and (s1n18741,n18715,n14141);
and (n18742,n18743,n14385);
wire s0n18743,s1n18743,notn18743;
or (n18743,s0n18743,s1n18743);
not(notn18743,n2799);
and (s0n18743,notn18743,1'b0);
and (s1n18743,n2799,n18744);
or (n18744,1'b0,n18745,n18747,n18749);
and (n18745,n18746,n13897);
and (n18747,n18748,n13900);
wire s0n18748,s1n18748,notn18748;
or (n18748,s0n18748,s1n18748);
not(notn18748,n14570);
and (s0n18748,notn18748,n14155);
and (s1n18748,n14570,1'b0);
and (n18749,n18750,n14131);
wire s0n18750,s1n18750,notn18750;
or (n18750,s0n18750,s1n18750);
not(notn18750,n14573);
and (s0n18750,notn18750,n14603);
and (s1n18750,n14573,1'b0);
and (n18751,n18752,n17820);
and (n18752,n18753,n14131);
wire s0n18753,s1n18753,notn18753;
or (n18753,s0n18753,s1n18753);
not(notn18753,n17823);
and (s0n18753,notn18753,1'b0);
and (s1n18753,n17823,n14141);
or (n18754,n18755,n18796,n19058);
and (n18755,n18756,n18779);
wire s0n18756,s1n18756,notn18756;
or (n18756,s0n18756,s1n18756);
not(notn18756,n14631);
and (s0n18756,notn18756,n18757);
and (s1n18756,n14631,n18769);
wire s0n18757,s1n18757,notn18757;
or (n18757,s0n18757,s1n18757);
not(notn18757,n14271);
and (s0n18757,notn18757,n18758);
and (s1n18757,n14271,n18761);
wire s0n18758,s1n18758,notn18758;
or (n18758,s0n18758,s1n18758);
not(notn18758,n14279);
and (s0n18758,notn18758,1'b0);
and (s1n18758,n14279,n18759);
and (n18759,n18760,n14367);
wire s0n18760,s1n18760,notn18760;
or (n18760,s0n18760,s1n18760);
not(notn18760,n18715);
and (s0n18760,notn18760,1'b0);
and (s1n18760,n18715,n14671);
and (n18761,n18762,n14385);
wire s0n18762,s1n18762,notn18762;
or (n18762,s0n18762,s1n18762);
not(notn18762,n2799);
and (s0n18762,notn18762,1'b0);
and (s1n18762,n2799,n18763);
or (n18763,1'b0,n18764,n18765,n18767);
and (n18764,n14642,n13897);
and (n18765,n18766,n13900);
wire s0n18766,s1n18766,notn18766;
or (n18766,s0n18766,s1n18766);
not(notn18766,n14570);
and (s0n18766,notn18766,n14678);
and (s1n18766,n14570,1'b0);
and (n18767,n18768,n14131);
wire s0n18768,s1n18768,notn18768;
or (n18768,s0n18768,s1n18768);
not(notn18768,n14573);
and (s0n18768,notn18768,n14746);
and (s1n18768,n14573,1'b0);
or (n18769,n18770,n18771,n18774,n18775,n18776,1'b0);
and (n18770,n17100,n14237);
and (n18771,n18772,n14111);
or (n18772,n17934,n18773,n17935,1'b0);
and (n18773,n14703,n13897);
and (n18774,n17976,n13950);
and (n18775,n14783,n14239);
and (n18776,n18777,n17820);
and (n18777,n18778,n14131);
wire s0n18778,s1n18778,notn18778;
or (n18778,s0n18778,s1n18778);
not(notn18778,n17823);
and (s0n18778,notn18778,1'b0);
and (s1n18778,n17823,n14671);
wire s0n18779,s1n18779,notn18779;
or (n18779,s0n18779,s1n18779);
not(notn18779,n14631);
and (s0n18779,notn18779,n18780);
and (s1n18779,n14631,n18793);
wire s0n18780,s1n18780,notn18780;
or (n18780,s0n18780,s1n18780);
not(notn18780,n14271);
and (s0n18780,notn18780,n18781);
and (s1n18780,n14271,n18784);
wire s0n18781,s1n18781,notn18781;
or (n18781,s0n18781,s1n18781);
not(notn18781,n14279);
and (s0n18781,notn18781,1'b0);
and (s1n18781,n14279,n18782);
and (n18782,n18783,n14367);
wire s0n18783,s1n18783,notn18783;
or (n18783,s0n18783,s1n18783);
not(notn18783,n18715);
and (s0n18783,notn18783,1'b0);
and (s1n18783,n18715,n14655);
and (n18784,n18785,n14385);
wire s0n18785,s1n18785,notn18785;
or (n18785,s0n18785,s1n18785);
not(notn18785,n2799);
and (s0n18785,notn18785,1'b0);
and (s1n18785,n2799,n18786);
or (n18786,1'b0,n18787,n18789,n18791);
and (n18787,n18788,n13897);
and (n18789,n18790,n13900);
wire s0n18790,s1n18790,notn18790;
or (n18790,s0n18790,s1n18790);
not(notn18790,n14570);
and (s0n18790,notn18790,n14662);
and (s1n18790,n14570,1'b0);
and (n18791,n18792,n14131);
wire s0n18792,s1n18792,notn18792;
or (n18792,s0n18792,s1n18792);
not(notn18792,n14573);
and (s0n18792,notn18792,n14946);
and (s1n18792,n14573,1'b0);
and (n18793,n18794,n17820);
and (n18794,n18795,n14131);
wire s0n18795,s1n18795,notn18795;
or (n18795,s0n18795,s1n18795);
not(notn18795,n17823);
and (s0n18795,notn18795,1'b0);
and (s1n18795,n17823,n14655);
and (n18796,n18779,n18797);
or (n18797,n18798,n18839,n19057);
and (n18798,n18799,n18822);
wire s0n18799,s1n18799,notn18799;
or (n18799,s0n18799,s1n18799);
not(notn18799,n14631);
and (s0n18799,notn18799,n18800);
and (s1n18799,n14631,n18812);
wire s0n18800,s1n18800,notn18800;
or (n18800,s0n18800,s1n18800);
not(notn18800,n14271);
and (s0n18800,notn18800,n18801);
and (s1n18800,n14271,n18804);
wire s0n18801,s1n18801,notn18801;
or (n18801,s0n18801,s1n18801);
not(notn18801,n14279);
and (s0n18801,notn18801,1'b0);
and (s1n18801,n14279,n18802);
and (n18802,n18803,n14367);
wire s0n18803,s1n18803,notn18803;
or (n18803,s0n18803,s1n18803);
not(notn18803,n18715);
and (s0n18803,notn18803,1'b0);
and (s1n18803,n18715,n15039);
and (n18804,n18805,n14385);
wire s0n18805,s1n18805,notn18805;
or (n18805,s0n18805,s1n18805);
not(notn18805,n2799);
and (s0n18805,notn18805,1'b0);
and (s1n18805,n2799,n18806);
or (n18806,1'b0,n18807,n18808,n18810);
and (n18807,n15185,n13897);
and (n18808,n18809,n13900);
wire s0n18809,s1n18809,notn18809;
or (n18809,s0n18809,s1n18809);
not(notn18809,n14570);
and (s0n18809,notn18809,n15046);
and (s1n18809,n14570,1'b0);
and (n18810,n18811,n14131);
wire s0n18811,s1n18811,notn18811;
or (n18811,s0n18811,s1n18811);
not(notn18811,n14573);
and (s0n18811,notn18811,n15177);
and (s1n18811,n14573,1'b0);
or (n18812,n18813,n18814,n18817,n18818,n18819,1'b0);
and (n18813,n17129,n14237);
and (n18814,n18815,n14111);
or (n18815,n18057,n18816,n18058,1'b0);
and (n18816,n15012,n13897);
and (n18817,n18100,n13950);
and (n18818,n15104,n14239);
and (n18819,n18820,n17820);
and (n18820,n18821,n14131);
wire s0n18821,s1n18821,notn18821;
or (n18821,s0n18821,s1n18821);
not(notn18821,n17823);
and (s0n18821,notn18821,1'b0);
and (s1n18821,n17823,n15039);
wire s0n18822,s1n18822,notn18822;
or (n18822,s0n18822,s1n18822);
not(notn18822,n14631);
and (s0n18822,notn18822,n18823);
and (s1n18822,n14631,n18836);
wire s0n18823,s1n18823,notn18823;
or (n18823,s0n18823,s1n18823);
not(notn18823,n14271);
and (s0n18823,notn18823,n18824);
and (s1n18823,n14271,n18827);
wire s0n18824,s1n18824,notn18824;
or (n18824,s0n18824,s1n18824);
not(notn18824,n14279);
and (s0n18824,notn18824,1'b0);
and (s1n18824,n14279,n18825);
and (n18825,n18826,n14367);
wire s0n18826,s1n18826,notn18826;
or (n18826,s0n18826,s1n18826);
not(notn18826,n18715);
and (s0n18826,notn18826,1'b0);
and (s1n18826,n18715,n15056);
and (n18827,n18828,n14385);
wire s0n18828,s1n18828,notn18828;
or (n18828,s0n18828,s1n18828);
not(notn18828,n2799);
and (s0n18828,notn18828,1'b0);
and (s1n18828,n2799,n18829);
or (n18829,1'b0,n18830,n18832,n18834);
and (n18830,n18831,n13897);
and (n18832,n18833,n13900);
wire s0n18833,s1n18833,notn18833;
or (n18833,s0n18833,s1n18833);
not(notn18833,n14570);
and (s0n18833,notn18833,n15063);
and (s1n18833,n14570,1'b0);
and (n18834,n18835,n14131);
wire s0n18835,s1n18835,notn18835;
or (n18835,s0n18835,s1n18835);
not(notn18835,n14573);
and (s0n18835,notn18835,n15270);
and (s1n18835,n14573,1'b0);
and (n18836,n18837,n17820);
and (n18837,n18838,n14131);
wire s0n18838,s1n18838,notn18838;
or (n18838,s0n18838,s1n18838);
not(notn18838,n17823);
and (s0n18838,notn18838,1'b0);
and (s1n18838,n17823,n15056);
and (n18839,n18822,n18840);
or (n18840,n18841,n18882,n19056);
and (n18841,n18842,n18865);
wire s0n18842,s1n18842,notn18842;
or (n18842,s0n18842,s1n18842);
not(notn18842,n14631);
and (s0n18842,notn18842,n18843);
and (s1n18842,n14631,n18855);
wire s0n18843,s1n18843,notn18843;
or (n18843,s0n18843,s1n18843);
not(notn18843,n14271);
and (s0n18843,notn18843,n18844);
and (s1n18843,n14271,n18847);
wire s0n18844,s1n18844,notn18844;
or (n18844,s0n18844,s1n18844);
not(notn18844,n14279);
and (s0n18844,notn18844,1'b0);
and (s1n18844,n14279,n18845);
and (n18845,n18846,n14367);
wire s0n18846,s1n18846,notn18846;
or (n18846,s0n18846,s1n18846);
not(notn18846,n18715);
and (s0n18846,notn18846,1'b0);
and (s1n18846,n18715,n15335);
and (n18847,n18848,n14385);
wire s0n18848,s1n18848,notn18848;
or (n18848,s0n18848,s1n18848);
not(notn18848,n2799);
and (s0n18848,notn18848,1'b0);
and (s1n18848,n2799,n18849);
or (n18849,1'b0,n18850,n18851,n18853);
and (n18850,n15306,n13897);
and (n18851,n18852,n13900);
wire s0n18852,s1n18852,notn18852;
or (n18852,s0n18852,s1n18852);
not(notn18852,n14570);
and (s0n18852,notn18852,n15342);
and (s1n18852,n14570,1'b0);
and (n18853,n18854,n14131);
wire s0n18854,s1n18854,notn18854;
or (n18854,s0n18854,s1n18854);
not(notn18854,n14573);
and (s0n18854,notn18854,n15409);
and (s1n18854,n14573,1'b0);
or (n18855,n18856,n18857,n18860,n18861,n18862,1'b0);
and (n18856,n17162,n14237);
and (n18857,n18858,n14111);
or (n18858,n18171,n18859,n18172,1'b0);
and (n18859,n15367,n13897);
and (n18860,n18213,n13950);
and (n18861,n15446,n14239);
and (n18862,n18863,n17820);
and (n18863,n18864,n14131);
wire s0n18864,s1n18864,notn18864;
or (n18864,s0n18864,s1n18864);
not(notn18864,n17823);
and (s0n18864,notn18864,1'b0);
and (s1n18864,n17823,n15335);
wire s0n18865,s1n18865,notn18865;
or (n18865,s0n18865,s1n18865);
not(notn18865,n14631);
and (s0n18865,notn18865,n18866);
and (s1n18865,n14631,n18879);
wire s0n18866,s1n18866,notn18866;
or (n18866,s0n18866,s1n18866);
not(notn18866,n14271);
and (s0n18866,notn18866,n18867);
and (s1n18866,n14271,n18870);
wire s0n18867,s1n18867,notn18867;
or (n18867,s0n18867,s1n18867);
not(notn18867,n14279);
and (s0n18867,notn18867,1'b0);
and (s1n18867,n14279,n18868);
and (n18868,n18869,n14367);
wire s0n18869,s1n18869,notn18869;
or (n18869,s0n18869,s1n18869);
not(notn18869,n18715);
and (s0n18869,notn18869,1'b0);
and (s1n18869,n18715,n15319);
and (n18870,n18871,n14385);
wire s0n18871,s1n18871,notn18871;
or (n18871,s0n18871,s1n18871);
not(notn18871,n2799);
and (s0n18871,notn18871,1'b0);
and (s1n18871,n2799,n18872);
or (n18872,1'b0,n18873,n18875,n18877);
and (n18873,n18874,n13897);
and (n18875,n18876,n13900);
wire s0n18876,s1n18876,notn18876;
or (n18876,s0n18876,s1n18876);
not(notn18876,n14570);
and (s0n18876,notn18876,n15326);
and (s1n18876,n14570,1'b0);
and (n18877,n18878,n14131);
wire s0n18878,s1n18878,notn18878;
or (n18878,s0n18878,s1n18878);
not(notn18878,n14573);
and (s0n18878,notn18878,n15610);
and (s1n18878,n14573,1'b0);
and (n18879,n18880,n17820);
and (n18880,n18881,n14131);
wire s0n18881,s1n18881,notn18881;
or (n18881,s0n18881,s1n18881);
not(notn18881,n17823);
and (s0n18881,notn18881,1'b0);
and (s1n18881,n17823,n15319);
and (n18882,n18865,n18883);
or (n18883,n18884,n18925,n19055);
and (n18884,n18885,n18908);
wire s0n18885,s1n18885,notn18885;
or (n18885,s0n18885,s1n18885);
not(notn18885,n14631);
and (s0n18885,notn18885,n18886);
and (s1n18885,n14631,n18898);
wire s0n18886,s1n18886,notn18886;
or (n18886,s0n18886,s1n18886);
not(notn18886,n14271);
and (s0n18886,notn18886,n18887);
and (s1n18886,n14271,n18890);
wire s0n18887,s1n18887,notn18887;
or (n18887,s0n18887,s1n18887);
not(notn18887,n14279);
and (s0n18887,notn18887,1'b0);
and (s1n18887,n14279,n18888);
and (n18888,n18889,n14367);
wire s0n18889,s1n18889,notn18889;
or (n18889,s0n18889,s1n18889);
not(notn18889,n18715);
and (s0n18889,notn18889,1'b0);
and (s1n18889,n18715,n15674);
and (n18890,n18891,n14385);
wire s0n18891,s1n18891,notn18891;
or (n18891,s0n18891,s1n18891);
not(notn18891,n2799);
and (s0n18891,notn18891,1'b0);
and (s1n18891,n2799,n18892);
or (n18892,1'b0,n18893,n18894,n18896);
and (n18893,n15645,n13897);
and (n18894,n18895,n13900);
wire s0n18895,s1n18895,notn18895;
or (n18895,s0n18895,s1n18895);
not(notn18895,n14570);
and (s0n18895,notn18895,n15681);
and (s1n18895,n14570,1'b0);
and (n18896,n18897,n14131);
wire s0n18897,s1n18897,notn18897;
or (n18897,s0n18897,s1n18897);
not(notn18897,n14573);
and (s0n18897,notn18897,n15748);
and (s1n18897,n14573,1'b0);
or (n18898,n18899,n18900,n18903,n18904,n18905,1'b0);
and (n18899,n17192,n14237);
and (n18900,n18901,n14111);
or (n18901,n18285,n18902,n18286,1'b0);
and (n18902,n15706,n13897);
and (n18903,n18327,n13950);
and (n18904,n15785,n14239);
and (n18905,n18906,n17820);
and (n18906,n18907,n14131);
wire s0n18907,s1n18907,notn18907;
or (n18907,s0n18907,s1n18907);
not(notn18907,n17823);
and (s0n18907,notn18907,1'b0);
and (s1n18907,n17823,n15674);
wire s0n18908,s1n18908,notn18908;
or (n18908,s0n18908,s1n18908);
not(notn18908,n14631);
and (s0n18908,notn18908,n18909);
and (s1n18908,n14631,n18922);
wire s0n18909,s1n18909,notn18909;
or (n18909,s0n18909,s1n18909);
not(notn18909,n14271);
and (s0n18909,notn18909,n18910);
and (s1n18909,n14271,n18913);
wire s0n18910,s1n18910,notn18910;
or (n18910,s0n18910,s1n18910);
not(notn18910,n14279);
and (s0n18910,notn18910,1'b0);
and (s1n18910,n14279,n18911);
and (n18911,n18912,n14367);
wire s0n18912,s1n18912,notn18912;
or (n18912,s0n18912,s1n18912);
not(notn18912,n18715);
and (s0n18912,notn18912,1'b0);
and (s1n18912,n18715,n15658);
and (n18913,n18914,n14385);
wire s0n18914,s1n18914,notn18914;
or (n18914,s0n18914,s1n18914);
not(notn18914,n2799);
and (s0n18914,notn18914,1'b0);
and (s1n18914,n2799,n18915);
or (n18915,1'b0,n18916,n18918,n18920);
and (n18916,n18917,n13897);
and (n18918,n18919,n13900);
wire s0n18919,s1n18919,notn18919;
or (n18919,s0n18919,s1n18919);
not(notn18919,n14570);
and (s0n18919,notn18919,n15665);
and (s1n18919,n14570,1'b0);
and (n18920,n18921,n14131);
wire s0n18921,s1n18921,notn18921;
or (n18921,s0n18921,s1n18921);
not(notn18921,n14573);
and (s0n18921,notn18921,n15949);
and (s1n18921,n14573,1'b0);
and (n18922,n18923,n17820);
and (n18923,n18924,n14131);
wire s0n18924,s1n18924,notn18924;
or (n18924,s0n18924,s1n18924);
not(notn18924,n17823);
and (s0n18924,notn18924,1'b0);
and (s1n18924,n17823,n15658);
and (n18925,n18908,n18926);
or (n18926,n18927,n18968,n19054);
and (n18927,n18928,n18951);
wire s0n18928,s1n18928,notn18928;
or (n18928,s0n18928,s1n18928);
not(notn18928,n14631);
and (s0n18928,notn18928,n18929);
and (s1n18928,n14631,n18941);
wire s0n18929,s1n18929,notn18929;
or (n18929,s0n18929,s1n18929);
not(notn18929,n14271);
and (s0n18929,notn18929,n18930);
and (s1n18929,n14271,n18933);
wire s0n18930,s1n18930,notn18930;
or (n18930,s0n18930,s1n18930);
not(notn18930,n14279);
and (s0n18930,notn18930,1'b0);
and (s1n18930,n14279,n18931);
and (n18931,n18932,n14367);
wire s0n18932,s1n18932,notn18932;
or (n18932,s0n18932,s1n18932);
not(notn18932,n18715);
and (s0n18932,notn18932,1'b0);
and (s1n18932,n18715,n16014);
and (n18933,n18934,n14385);
wire s0n18934,s1n18934,notn18934;
or (n18934,s0n18934,s1n18934);
not(notn18934,n2799);
and (s0n18934,notn18934,1'b0);
and (s1n18934,n2799,n18935);
or (n18935,1'b0,n18936,n18937,n18939);
and (n18936,n15985,n13897);
and (n18937,n18938,n13900);
wire s0n18938,s1n18938,notn18938;
or (n18938,s0n18938,s1n18938);
not(notn18938,n14570);
and (s0n18938,notn18938,n16021);
and (s1n18938,n14570,1'b0);
and (n18939,n18940,n14131);
wire s0n18940,s1n18940,notn18940;
or (n18940,s0n18940,s1n18940);
not(notn18940,n14573);
and (s0n18940,notn18940,n16088);
and (s1n18940,n14573,1'b0);
or (n18941,n18942,n18943,n18946,n18947,n18948,1'b0);
and (n18942,n17221,n14237);
and (n18943,n18944,n14111);
or (n18944,n18399,n18945,n18400,1'b0);
and (n18945,n16046,n13897);
and (n18946,n18441,n13950);
and (n18947,n16125,n14239);
and (n18948,n18949,n17820);
and (n18949,n18950,n14131);
wire s0n18950,s1n18950,notn18950;
or (n18950,s0n18950,s1n18950);
not(notn18950,n17823);
and (s0n18950,notn18950,1'b0);
and (s1n18950,n17823,n16014);
wire s0n18951,s1n18951,notn18951;
or (n18951,s0n18951,s1n18951);
not(notn18951,n14631);
and (s0n18951,notn18951,n18952);
and (s1n18951,n14631,n18965);
wire s0n18952,s1n18952,notn18952;
or (n18952,s0n18952,s1n18952);
not(notn18952,n14271);
and (s0n18952,notn18952,n18953);
and (s1n18952,n14271,n18956);
wire s0n18953,s1n18953,notn18953;
or (n18953,s0n18953,s1n18953);
not(notn18953,n14279);
and (s0n18953,notn18953,1'b0);
and (s1n18953,n14279,n18954);
and (n18954,n18955,n14367);
wire s0n18955,s1n18955,notn18955;
or (n18955,s0n18955,s1n18955);
not(notn18955,n18715);
and (s0n18955,notn18955,1'b0);
and (s1n18955,n18715,n15998);
and (n18956,n18957,n14385);
wire s0n18957,s1n18957,notn18957;
or (n18957,s0n18957,s1n18957);
not(notn18957,n2799);
and (s0n18957,notn18957,1'b0);
and (s1n18957,n2799,n18958);
or (n18958,1'b0,n18959,n18961,n18963);
and (n18959,n18960,n13897);
and (n18961,n18962,n13900);
wire s0n18962,s1n18962,notn18962;
or (n18962,s0n18962,s1n18962);
not(notn18962,n14570);
and (s0n18962,notn18962,n16005);
and (s1n18962,n14570,1'b0);
and (n18963,n18964,n14131);
wire s0n18964,s1n18964,notn18964;
or (n18964,s0n18964,s1n18964);
not(notn18964,n14573);
and (s0n18964,notn18964,n16289);
and (s1n18964,n14573,1'b0);
and (n18965,n18966,n17820);
and (n18966,n18967,n14131);
wire s0n18967,s1n18967,notn18967;
or (n18967,s0n18967,s1n18967);
not(notn18967,n17823);
and (s0n18967,notn18967,1'b0);
and (s1n18967,n17823,n15998);
and (n18968,n18951,n18969);
or (n18969,n18970,n19011,n19053);
and (n18970,n18971,n18994);
wire s0n18971,s1n18971,notn18971;
or (n18971,s0n18971,s1n18971);
not(notn18971,n14631);
and (s0n18971,notn18971,n18972);
and (s1n18971,n14631,n18984);
wire s0n18972,s1n18972,notn18972;
or (n18972,s0n18972,s1n18972);
not(notn18972,n14271);
and (s0n18972,notn18972,n18973);
and (s1n18972,n14271,n18976);
wire s0n18973,s1n18973,notn18973;
or (n18973,s0n18973,s1n18973);
not(notn18973,n14279);
and (s0n18973,notn18973,1'b0);
and (s1n18973,n14279,n18974);
and (n18974,n18975,n14367);
wire s0n18975,s1n18975,notn18975;
or (n18975,s0n18975,s1n18975);
not(notn18975,n18715);
and (s0n18975,notn18975,1'b0);
and (s1n18975,n18715,n16354);
and (n18976,n18977,n14385);
wire s0n18977,s1n18977,notn18977;
or (n18977,s0n18977,s1n18977);
not(notn18977,n2799);
and (s0n18977,notn18977,1'b0);
and (s1n18977,n2799,n18978);
or (n18978,1'b0,n18979,n18980,n18982);
and (n18979,n16325,n13897);
and (n18980,n18981,n13900);
wire s0n18981,s1n18981,notn18981;
or (n18981,s0n18981,s1n18981);
not(notn18981,n14570);
and (s0n18981,notn18981,n16361);
and (s1n18981,n14570,1'b0);
and (n18982,n18983,n14131);
wire s0n18983,s1n18983,notn18983;
or (n18983,s0n18983,s1n18983);
not(notn18983,n14573);
and (s0n18983,notn18983,n16428);
and (s1n18983,n14573,1'b0);
or (n18984,n18985,n18986,n18989,n18990,n18991,1'b0);
and (n18985,n17252,n14237);
and (n18986,n18987,n14111);
or (n18987,n18513,n18988,n18514,1'b0);
and (n18988,n16386,n13897);
and (n18989,n18555,n13950);
and (n18990,n16465,n14239);
and (n18991,n18992,n17820);
and (n18992,n18993,n14131);
wire s0n18993,s1n18993,notn18993;
or (n18993,s0n18993,s1n18993);
not(notn18993,n17823);
and (s0n18993,notn18993,1'b0);
and (s1n18993,n17823,n16354);
wire s0n18994,s1n18994,notn18994;
or (n18994,s0n18994,s1n18994);
not(notn18994,n14631);
and (s0n18994,notn18994,n18995);
and (s1n18994,n14631,n19008);
wire s0n18995,s1n18995,notn18995;
or (n18995,s0n18995,s1n18995);
not(notn18995,n14271);
and (s0n18995,notn18995,n18996);
and (s1n18995,n14271,n18999);
wire s0n18996,s1n18996,notn18996;
or (n18996,s0n18996,s1n18996);
not(notn18996,n14279);
and (s0n18996,notn18996,1'b0);
and (s1n18996,n14279,n18997);
and (n18997,n18998,n14367);
wire s0n18998,s1n18998,notn18998;
or (n18998,s0n18998,s1n18998);
not(notn18998,n18715);
and (s0n18998,notn18998,1'b0);
and (s1n18998,n18715,n16338);
and (n18999,n19000,n14385);
wire s0n19000,s1n19000,notn19000;
or (n19000,s0n19000,s1n19000);
not(notn19000,n2799);
and (s0n19000,notn19000,1'b0);
and (s1n19000,n2799,n19001);
or (n19001,1'b0,n19002,n19004,n19006);
and (n19002,n19003,n13897);
and (n19004,n19005,n13900);
wire s0n19005,s1n19005,notn19005;
or (n19005,s0n19005,s1n19005);
not(notn19005,n14570);
and (s0n19005,notn19005,n16345);
and (s1n19005,n14570,1'b0);
and (n19006,n19007,n14131);
wire s0n19007,s1n19007,notn19007;
or (n19007,s0n19007,s1n19007);
not(notn19007,n14573);
and (s0n19007,notn19007,n16606);
and (s1n19007,n14573,1'b0);
and (n19008,n19009,n17820);
and (n19009,n19010,n14131);
wire s0n19010,s1n19010,notn19010;
or (n19010,s0n19010,s1n19010);
not(notn19010,n17823);
and (s0n19010,notn19010,1'b0);
and (s1n19010,n17823,n16338);
and (n19011,n18994,n19012);
and (n19012,n19013,n19036);
wire s0n19013,s1n19013,notn19013;
or (n19013,s0n19013,s1n19013);
not(notn19013,n14631);
and (s0n19013,notn19013,n19014);
and (s1n19013,n14631,n19026);
wire s0n19014,s1n19014,notn19014;
or (n19014,s0n19014,s1n19014);
not(notn19014,n14271);
and (s0n19014,notn19014,n19015);
and (s1n19014,n14271,n19018);
wire s0n19015,s1n19015,notn19015;
or (n19015,s0n19015,s1n19015);
not(notn19015,n14279);
and (s0n19015,notn19015,1'b0);
and (s1n19015,n14279,n19016);
and (n19016,n19017,n14367);
wire s0n19017,s1n19017,notn19017;
or (n19017,s0n19017,s1n19017);
not(notn19017,n18715);
and (s0n19017,notn19017,1'b0);
and (s1n19017,n18715,n16722);
and (n19018,n19019,n14385);
wire s0n19019,s1n19019,notn19019;
or (n19019,s0n19019,s1n19019);
not(notn19019,n2799);
and (s0n19019,notn19019,1'b0);
and (s1n19019,n2799,n19020);
or (n19020,1'b0,n19021,n19022,n19024);
and (n19021,n16693,n13897);
and (n19022,n19023,n13900);
wire s0n19023,s1n19023,notn19023;
or (n19023,s0n19023,s1n19023);
not(notn19023,n14570);
and (s0n19023,notn19023,n16729);
and (s1n19023,n14570,1'b0);
and (n19024,n19025,n14131);
wire s0n19025,s1n19025,notn19025;
or (n19025,s0n19025,s1n19025);
not(notn19025,n14573);
and (s0n19025,notn19025,n16796);
and (s1n19025,n14573,1'b0);
or (n19026,n19027,n19028,n19031,n19032,n19033,1'b0);
and (n19027,n17278,n14237);
and (n19028,n19029,n14111);
or (n19029,n18626,n19030,n18627,1'b0);
and (n19030,n16754,n13897);
and (n19031,n18668,n13950);
and (n19032,n16833,n14239);
and (n19033,n19034,n17820);
and (n19034,n19035,n14131);
wire s0n19035,s1n19035,notn19035;
or (n19035,s0n19035,s1n19035);
not(notn19035,n17823);
and (s0n19035,notn19035,1'b0);
and (s1n19035,n17823,n16722);
wire s0n19036,s1n19036,notn19036;
or (n19036,s0n19036,s1n19036);
not(notn19036,n14631);
and (s0n19036,notn19036,n19037);
and (s1n19036,n14631,n19050);
wire s0n19037,s1n19037,notn19037;
or (n19037,s0n19037,s1n19037);
not(notn19037,n14271);
and (s0n19037,notn19037,n19038);
and (s1n19037,n14271,n19041);
wire s0n19038,s1n19038,notn19038;
or (n19038,s0n19038,s1n19038);
not(notn19038,n14279);
and (s0n19038,notn19038,1'b0);
and (s1n19038,n14279,n19039);
and (n19039,n19040,n14367);
wire s0n19040,s1n19040,notn19040;
or (n19040,s0n19040,s1n19040);
not(notn19040,n18715);
and (s0n19040,notn19040,1'b0);
and (s1n19040,n18715,n16706);
and (n19041,n19042,n14385);
wire s0n19042,s1n19042,notn19042;
or (n19042,s0n19042,s1n19042);
not(notn19042,n2799);
and (s0n19042,notn19042,1'b0);
and (s1n19042,n2799,n19043);
or (n19043,1'b0,n19044,n19046,n19048);
and (n19044,n19045,n13897);
and (n19046,n19047,n13900);
wire s0n19047,s1n19047,notn19047;
or (n19047,s0n19047,s1n19047);
not(notn19047,n14570);
and (s0n19047,notn19047,n16713);
and (s1n19047,n14570,1'b0);
and (n19048,n19049,n14131);
wire s0n19049,s1n19049,notn19049;
or (n19049,s0n19049,s1n19049);
not(notn19049,n14573);
and (s0n19049,notn19049,n16996);
and (s1n19049,n14573,1'b0);
and (n19050,n19051,n17820);
and (n19051,n19052,n14131);
wire s0n19052,s1n19052,notn19052;
or (n19052,s0n19052,s1n19052);
not(notn19052,n17823);
and (s0n19052,notn19052,1'b0);
and (s1n19052,n17823,n16706);
and (n19053,n18971,n19012);
and (n19054,n18928,n18969);
and (n19055,n18885,n18926);
and (n19056,n18842,n18883);
and (n19057,n18799,n18840);
and (n19058,n18756,n18797);
or (n19059,n17067,n19060,n19062,n17297,1'b0,1'b0);
and (n19060,n19061,n14111);
or (n19061,n14243,n13889);
and (n19062,n14125,n13950);
or (n19063,n19064,n19071,n19127);
and (n19064,n19065,n19068);
wire s0n19065,s1n19065,notn19065;
or (n19065,s0n19065,s1n19065);
not(notn19065,n18690);
and (s0n19065,notn19065,n19066);
and (s1n19065,n18690,1'b0);
xor (n19066,n19067,n17993);
xor (n19067,n17881,n17948);
wire s0n19068,s1n19068,notn19068;
or (n19068,s0n19068,s1n19068);
not(notn19068,n19059);
and (s0n19068,notn19068,n19069);
and (s1n19068,n19059,n18799);
xor (n19069,n19070,n18797);
xor (n19070,n18756,n18779);
and (n19071,n19068,n19072);
or (n19072,n19073,n19080,n19126);
and (n19073,n19074,n19077);
wire s0n19074,s1n19074,notn19074;
or (n19074,s0n19074,s1n19074);
not(notn19074,n18690);
and (s0n19074,notn19074,n19075);
and (s1n19074,n18690,1'b0);
xor (n19075,n19076,n18116);
xor (n19076,n17995,n18073);
wire s0n19077,s1n19077,notn19077;
or (n19077,s0n19077,s1n19077);
not(notn19077,n19059);
and (s0n19077,notn19077,n19078);
and (s1n19077,n19059,n18842);
xor (n19078,n19079,n18840);
xor (n19079,n18799,n18822);
and (n19080,n19077,n19081);
or (n19081,n19082,n19089,n19125);
and (n19082,n19083,n19086);
wire s0n19083,s1n19083,notn19083;
or (n19083,s0n19083,s1n19083);
not(notn19083,n18690);
and (s0n19083,notn19083,n19084);
and (s1n19083,n18690,1'b0);
xor (n19084,n19085,n18230);
xor (n19085,n18118,n18185);
wire s0n19086,s1n19086,notn19086;
or (n19086,s0n19086,s1n19086);
not(notn19086,n19059);
and (s0n19086,notn19086,n19087);
and (s1n19086,n19059,n18885);
xor (n19087,n19088,n18883);
xor (n19088,n18842,n18865);
and (n19089,n19086,n19090);
or (n19090,n19091,n19098,n19124);
and (n19091,n19092,n19095);
wire s0n19092,s1n19092,notn19092;
or (n19092,s0n19092,s1n19092);
not(notn19092,n18690);
and (s0n19092,notn19092,n19093);
and (s1n19092,n18690,1'b0);
xor (n19093,n19094,n18344);
xor (n19094,n18232,n18299);
wire s0n19095,s1n19095,notn19095;
or (n19095,s0n19095,s1n19095);
not(notn19095,n19059);
and (s0n19095,notn19095,n19096);
and (s1n19095,n19059,n18928);
xor (n19096,n19097,n18926);
xor (n19097,n18885,n18908);
and (n19098,n19095,n19099);
or (n19099,n19100,n19107,n19123);
and (n19100,n19101,n19104);
wire s0n19101,s1n19101,notn19101;
or (n19101,s0n19101,s1n19101);
not(notn19101,n18690);
and (s0n19101,notn19101,n19102);
and (s1n19101,n18690,1'b0);
xor (n19102,n19103,n18458);
xor (n19103,n18346,n18413);
wire s0n19104,s1n19104,notn19104;
or (n19104,s0n19104,s1n19104);
not(notn19104,n19059);
and (s0n19104,notn19104,n19105);
and (s1n19104,n19059,n18971);
xor (n19105,n19106,n18969);
xor (n19106,n18928,n18951);
and (n19107,n19104,n19108);
or (n19108,n19109,n19116,n19122);
and (n19109,n19110,n19113);
wire s0n19110,s1n19110,notn19110;
or (n19110,s0n19110,s1n19110);
not(notn19110,n18690);
and (s0n19110,notn19110,n19111);
and (s1n19110,n18690,1'b0);
xor (n19111,n19112,n18572);
xor (n19112,n18460,n18527);
wire s0n19113,s1n19113,notn19113;
or (n19113,s0n19113,s1n19113);
not(notn19113,n19059);
and (s0n19113,notn19113,n19114);
and (s1n19113,n19059,n19013);
xor (n19114,n19115,n19012);
xor (n19115,n18971,n18994);
and (n19116,n19113,n19117);
and (n19117,n19118,n19120);
wire s0n19118,s1n19118,notn19118;
or (n19118,s0n19118,s1n19118);
not(notn19118,n18690);
and (s0n19118,notn19118,n19119);
and (s1n19118,n18690,1'b0);
xor (n19119,n18573,n18640);
wire s0n19120,s1n19120,notn19120;
or (n19120,s0n19120,s1n19120);
not(notn19120,n19059);
and (s0n19120,notn19120,n19121);
and (s1n19120,n19059,1'b0);
xor (n19121,n19013,n19036);
and (n19122,n19110,n19117);
and (n19123,n19101,n19108);
and (n19124,n19092,n19099);
and (n19125,n19083,n19090);
and (n19126,n19074,n19081);
and (n19127,n19065,n19072);
and (n19128,n19129,n19131);
xor (n19129,n19130,n19072);
xor (n19130,n19065,n19068);
and (n19131,n19132,n19134);
xor (n19132,n19133,n19081);
xor (n19133,n19074,n19077);
or (n19134,n19135,n19143,n19194);
and (n19135,n19136,n19138);
xor (n19136,n19137,n19090);
xor (n19137,n19083,n19086);
wire s0n19138,s1n19138,notn19138;
or (n19138,s0n19138,s1n19138);
not(notn19138,n14271);
and (s0n19138,notn19138,n14504);
and (s1n19138,n14271,n19139);
or (n19139,n14506,n19140,1'b0);
and (n19140,n19141,n14385);
wire s0n19141,s1n19141,notn19141;
or (n19141,s0n19141,s1n19141);
not(notn19141,n2799);
and (s0n19141,notn19141,1'b0);
and (s1n19141,n2799,n19142);
and (n19142,n17758,n13889);
and (n19143,n19138,n19144);
or (n19144,n19145,n19153,n19193);
and (n19145,n19146,n19148);
xor (n19146,n19147,n19099);
xor (n19147,n19092,n19095);
wire s0n19148,s1n19148,notn19148;
or (n19148,s0n19148,s1n19148);
not(notn19148,n14271);
and (s0n19148,notn19148,1'b0);
and (s1n19148,n14271,n19149);
and (n19149,n19150,n14385);
wire s0n19150,s1n19150,notn19150;
or (n19150,s0n19150,s1n19150);
not(notn19150,n2799);
and (s0n19150,notn19150,1'b0);
and (s1n19150,n2799,n19151);
and (n19151,n19152,n13889);
not (n19152,n17758);
and (n19153,n19148,n19154);
or (n19154,n19155,n19167,n19192);
and (n19155,n19156,n19158);
xor (n19156,n19157,n19108);
xor (n19157,n19101,n19104);
wire s0n19158,s1n19158,notn19158;
or (n19158,s0n19158,s1n19158);
not(notn19158,n14631);
and (s0n19158,notn19158,n19159);
and (s1n19158,n14631,n19165);
and (n19159,n19160,n14367);
and (n19160,n19161,n17758);
wire s0n19161,s1n19161,notn19161;
or (n19161,s0n19161,s1n19161);
not(notn19161,n13900);
and (s0n19161,notn19161,1'b0);
and (s1n19161,n13900,n19162);
or (n19162,n19163,n14153);
or (n19163,n19164,n14161);
or (n19164,n14159,n14151);
and (n19165,n19166,n17820);
and (n19166,n17817,n13900);
and (n19167,n19158,n19168);
or (n19168,n19169,n19184,n19191);
and (n19169,n19170,n19172);
xor (n19170,n19171,n19117);
xor (n19171,n19110,n19113);
wire s0n19172,s1n19172,notn19172;
or (n19172,s0n19172,s1n19172);
not(notn19172,n14631);
and (s0n19172,notn19172,n19173);
and (s1n19172,n14631,n19181);
wire s0n19173,s1n19173,notn19173;
or (n19173,s0n19173,s1n19173);
not(notn19173,n14279);
and (s0n19173,notn19173,1'b0);
and (s1n19173,n14279,n19174);
and (n19174,n19175,n14367);
or (n19175,n19176,n19179,1'b0);
and (n19176,n19177,n17758);
wire s0n19177,s1n19177,notn19177;
or (n19177,s0n19177,s1n19177);
not(notn19177,n13900);
and (s0n19177,notn19177,1'b0);
and (s1n19177,n13900,n19178);
not (n19178,n19162);
and (n19179,n13900,n19180);
or (n19180,n17765,n17762);
or (n19181,n17067,1'b0,n19060,1'b0,n19062,n17297,n19182,1'b0);
and (n19182,n19183,n17820);
and (n19183,n17829,n13900);
and (n19184,n19172,n19185);
and (n19185,n19186,n19187);
xor (n19186,n19118,n19120);
or (n19187,n19188,n19189,n14345,n19190,1'b0,1'b0,1'b0,1'b0);
and (n19188,n14131,n14237);
and (n19189,n14131,n14137);
and (n19190,n14125,n14108);
and (n19191,n19170,n19185);
and (n19192,n19156,n19168);
and (n19193,n19146,n19154);
and (n19194,n19136,n19144);
xor (n19195,n19196,n19268);
xor (n19196,n19197,n19264);
xor (n19197,n19198,n19248);
wire s0n19198,s1n19198,notn19198;
or (n19198,s0n19198,s1n19198);
not(notn19198,n18690);
and (s0n19198,notn19198,n19199);
and (s1n19198,n18690,1'b0);
xor (n19199,n19200,n19244);
xor (n19200,n19201,n19228);
wire s0n19201,s1n19201,notn19201;
or (n19201,s0n19201,s1n19201);
not(notn19201,n14631);
and (s0n19201,notn19201,n19202);
and (s1n19201,n14631,n19225);
wire s0n19202,s1n19202,notn19202;
or (n19202,s0n19202,s1n19202);
not(notn19202,n14271);
and (s0n19202,notn19202,n19203);
and (s1n19202,n14271,n19217);
wire s0n19203,s1n19203,notn19203;
or (n19203,s0n19203,s1n19203);
not(notn19203,n14279);
and (s0n19203,notn19203,1'b0);
and (s1n19203,n14279,n19204);
or (n19204,n19205,1'b0,1'b0,n19209);
and (n19205,n19206,n14120);
wire s0n19206,s1n19206,notn19206;
or (n19206,s0n19206,s1n19206);
not(notn19206,n14125);
and (s0n19206,notn19206,1'b0);
and (s1n19206,n14125,n19207);
wire s0n19207,s1n19207,notn19207;
or (n19207,s0n19207,s1n19207);
not(notn19207,n14317);
and (s0n19207,notn19207,n19208);
and (s1n19207,n14317,n17402);
and (n19209,n19210,n14367);
or (n19210,n19211,n19213,n19216,1'b0);
and (n19211,n19212,n17758);
wire s0n19212,s1n19212,notn19212;
or (n19212,s0n19212,s1n19212);
not(notn19212,n13900);
and (s0n19212,notn19212,1'b0);
and (s1n19212,n13900,n19208);
and (n19213,n19214,n17762);
wire s0n19214,s1n19214,notn19214;
or (n19214,s0n19214,s1n19214);
not(notn19214,n13900);
and (s0n19214,notn19214,1'b0);
and (s1n19214,n13900,n19215);
and (n19216,n19212,n17765);
or (n19217,n19218,n19219,1'b0,1'b0);
and (n19218,n19206,n13907);
and (n19219,n19220,n14385);
wire s0n19220,s1n19220,notn19220;
or (n19220,s0n19220,s1n19220);
not(notn19220,n2799);
and (s0n19220,notn19220,1'b0);
and (s1n19220,n2799,n19221);
or (n19221,1'b0,n19222,n19224,1'b0);
and (n19222,n19223,n13889);
wire s0n19223,s1n19223,notn19223;
or (n19223,s0n19223,s1n19223);
not(notn19223,n17767);
and (s0n19223,notn19223,n19208);
and (s1n19223,n17767,1'b0);
and (n19224,n19208,n14243);
and (n19225,n19226,n17820);
and (n19226,n19227,n13900);
wire s0n19227,s1n19227,notn19227;
or (n19227,s0n19227,s1n19227);
not(notn19227,n17823);
and (s0n19227,notn19227,1'b0);
and (s1n19227,n17823,n19208);
wire s0n19228,s1n19228,notn19228;
or (n19228,s0n19228,s1n19228);
not(notn19228,n14631);
and (s0n19228,notn19228,n19229);
and (s1n19228,n14631,n19241);
wire s0n19229,s1n19229,notn19229;
or (n19229,s0n19229,s1n19229);
not(notn19229,n14271);
and (s0n19229,notn19229,n19230);
and (s1n19229,n14271,n19234);
wire s0n19230,s1n19230,notn19230;
or (n19230,s0n19230,s1n19230);
not(notn19230,n14279);
and (s0n19230,notn19230,1'b0);
and (s1n19230,n14279,n19231);
or (n19231,n17413,1'b0,n19232);
and (n19232,n19233,n14367);
and (n19233,n19214,n17758);
or (n19234,n19235,n19238,1'b0);
and (n19235,n19236,n13907);
wire s0n19236,s1n19236,notn19236;
or (n19236,s0n19236,s1n19236);
not(notn19236,n14125);
and (s0n19236,notn19236,1'b0);
and (s1n19236,n14125,n19237);
wire s0n19237,s1n19237,notn19237;
or (n19237,s0n19237,s1n19237);
not(notn19237,n14563);
and (s0n19237,notn19237,n17416);
and (s1n19237,n14563,n17417);
and (n19238,n19239,n14385);
wire s0n19239,s1n19239,notn19239;
or (n19239,s0n19239,s1n19239);
not(notn19239,n2799);
and (s0n19239,notn19239,1'b0);
and (s1n19239,n2799,n19240);
and (n19240,n19215,n14235);
and (n19241,n19242,n17820);
and (n19242,n19243,n13900);
wire s0n19243,s1n19243,notn19243;
or (n19243,s0n19243,s1n19243);
not(notn19243,n17818);
and (s0n19243,notn19243,1'b0);
and (s1n19243,n17818,n19215);
or (n19244,n19245,n19246,n19247);
and (n19245,n17736,n17837);
and (n19246,n17837,n17879);
and (n19247,n17736,n17879);
wire s0n19248,s1n19248,notn19248;
or (n19248,s0n19248,s1n19248);
not(notn19248,n19059);
and (s0n19248,notn19248,n19249);
and (s1n19248,n19059,n18710);
xor (n19249,n19250,n19260);
xor (n19250,n19251,n19255);
wire s0n19251,s1n19251,notn19251;
or (n19251,s0n19251,s1n19251);
not(notn19251,n14271);
and (s0n19251,notn19251,1'b0);
and (s1n19251,n14271,n19252);
and (n19252,n19253,n14385);
wire s0n19253,s1n19253,notn19253;
or (n19253,s0n19253,s1n19253);
not(notn19253,n2799);
and (s0n19253,notn19253,1'b0);
and (s1n19253,n2799,n19254);
and (n19254,n17400,n13897);
wire s0n19255,s1n19255,notn19255;
or (n19255,s0n19255,s1n19255);
not(notn19255,n14271);
and (s0n19255,notn19255,1'b0);
and (s1n19255,n14271,n19256);
and (n19256,n19257,n14385);
wire s0n19257,s1n19257,notn19257;
or (n19257,s0n19257,s1n19257);
not(notn19257,n2799);
and (s0n19257,notn19257,1'b0);
and (s1n19257,n2799,n19258);
and (n19258,n19259,n13897);
or (n19260,n19261,n19262,n19263);
and (n19261,n18710,n18737);
and (n19262,n18737,n18754);
and (n19263,n18710,n18754);
or (n19264,n19265,n19266,n19267);
and (n19265,n17733,n18707);
and (n19266,n18707,n19063);
and (n19267,n17733,n19063);
and (n19268,n17731,n19128);
wire s0n19269,s1n19269,notn19269;
or (n19269,s0n19269,s1n19269);
not(notn19269,n14631);
and (s0n19269,notn19269,n19270);
and (s1n19269,n14631,n19273);
wire s0n19270,s1n19270,notn19270;
or (n19270,s0n19270,s1n19270);
not(notn19270,n14271);
and (s0n19270,notn19270,n19271);
and (s1n19270,n14271,n19139);
wire s0n19271,s1n19271,notn19271;
or (n19271,s0n19271,s1n19271);
not(notn19271,n14279);
and (s0n19271,notn19271,1'b0);
and (s1n19271,n14279,n19272);
or (n19272,n14505,1'b0,n19159);
or (n19273,n19188,n19189,n14345,n19190,1'b0,1'b0,n19165,1'b0);
wire s0n19274,s1n19274,notn19274;
or (n19274,s0n19274,s1n19274);
not(notn19274,n19269);
and (s0n19274,notn19274,n19275);
and (s1n19274,n19269,n19348);
xor (n19275,n19276,n19347);
xor (n19276,n19277,n19343);
xor (n19277,n19278,n19328);
wire s0n19278,s1n19278,notn19278;
or (n19278,s0n19278,s1n19278);
not(notn19278,n18690);
and (s0n19278,notn19278,n19279);
and (s1n19278,n18690,1'b0);
xor (n19279,n19280,n19324);
xor (n19280,n19281,n19308);
wire s0n19281,s1n19281,notn19281;
or (n19281,s0n19281,s1n19281);
not(notn19281,n14631);
and (s0n19281,notn19281,n19282);
and (s1n19281,n14631,n19305);
wire s0n19282,s1n19282,notn19282;
or (n19282,s0n19282,s1n19282);
not(notn19282,n14271);
and (s0n19282,notn19282,n19283);
and (s1n19282,n14271,n19297);
wire s0n19283,s1n19283,notn19283;
or (n19283,s0n19283,s1n19283);
not(notn19283,n14279);
and (s0n19283,notn19283,1'b0);
and (s1n19283,n14279,n19284);
or (n19284,n19285,1'b0,1'b0,n19289);
and (n19285,n19286,n14120);
wire s0n19286,s1n19286,notn19286;
or (n19286,s0n19286,s1n19286);
not(notn19286,n14125);
and (s0n19286,notn19286,1'b0);
and (s1n19286,n14125,n19287);
wire s0n19287,s1n19287,notn19287;
or (n19287,s0n19287,s1n19287);
not(notn19287,n14317);
and (s0n19287,notn19287,n19288);
and (s1n19287,n14317,n17455);
and (n19289,n19290,n14367);
or (n19290,n19291,n19293,n19296,1'b0);
and (n19291,n19292,n17758);
wire s0n19292,s1n19292,notn19292;
or (n19292,s0n19292,s1n19292);
not(notn19292,n13900);
and (s0n19292,notn19292,1'b0);
and (s1n19292,n13900,n19288);
and (n19293,n19294,n17762);
wire s0n19294,s1n19294,notn19294;
or (n19294,s0n19294,s1n19294);
not(notn19294,n13900);
and (s0n19294,notn19294,1'b0);
and (s1n19294,n13900,n19295);
and (n19296,n19292,n17765);
or (n19297,n19298,n19299,1'b0,1'b0);
and (n19298,n19286,n13907);
and (n19299,n19300,n14385);
wire s0n19300,s1n19300,notn19300;
or (n19300,s0n19300,s1n19300);
not(notn19300,n2799);
and (s0n19300,notn19300,1'b0);
and (s1n19300,n2799,n19301);
or (n19301,1'b0,n19302,n19304,1'b0);
and (n19302,n19303,n13889);
wire s0n19303,s1n19303,notn19303;
or (n19303,s0n19303,s1n19303);
not(notn19303,n17767);
and (s0n19303,notn19303,n19288);
and (s1n19303,n17767,1'b0);
and (n19304,n19288,n14243);
and (n19305,n19306,n17820);
and (n19306,n19307,n13900);
wire s0n19307,s1n19307,notn19307;
or (n19307,s0n19307,s1n19307);
not(notn19307,n17823);
and (s0n19307,notn19307,1'b0);
and (s1n19307,n17823,n19288);
wire s0n19308,s1n19308,notn19308;
or (n19308,s0n19308,s1n19308);
not(notn19308,n14631);
and (s0n19308,notn19308,n19309);
and (s1n19308,n14631,n19321);
wire s0n19309,s1n19309,notn19309;
or (n19309,s0n19309,s1n19309);
not(notn19309,n14271);
and (s0n19309,notn19309,n19310);
and (s1n19309,n14271,n19314);
wire s0n19310,s1n19310,notn19310;
or (n19310,s0n19310,s1n19310);
not(notn19310,n14279);
and (s0n19310,notn19310,1'b0);
and (s1n19310,n14279,n19311);
or (n19311,n17466,1'b0,n19312);
and (n19312,n19313,n14367);
and (n19313,n19294,n17758);
or (n19314,n19315,n19318,1'b0);
and (n19315,n19316,n13907);
wire s0n19316,s1n19316,notn19316;
or (n19316,s0n19316,s1n19316);
not(notn19316,n14125);
and (s0n19316,notn19316,1'b0);
and (s1n19316,n14125,n19317);
wire s0n19317,s1n19317,notn19317;
or (n19317,s0n19317,s1n19317);
not(notn19317,n14563);
and (s0n19317,notn19317,n17469);
and (s1n19317,n14563,n17470);
and (n19318,n19319,n14385);
wire s0n19319,s1n19319,notn19319;
or (n19319,s0n19319,s1n19319);
not(notn19319,n2799);
and (s0n19319,notn19319,1'b0);
and (s1n19319,n2799,n19320);
and (n19320,n19295,n14235);
and (n19321,n19322,n17820);
and (n19322,n19323,n13900);
wire s0n19323,s1n19323,notn19323;
or (n19323,s0n19323,s1n19323);
not(notn19323,n17818);
and (s0n19323,notn19323,1'b0);
and (s1n19323,n17818,n19295);
or (n19324,n19325,n19326,n19327);
and (n19325,n19201,n19228);
and (n19326,n19228,n19244);
and (n19327,n19201,n19244);
xor (n19328,n19329,n19339);
xor (n19329,n19330,n19334);
wire s0n19330,s1n19330,notn19330;
or (n19330,s0n19330,s1n19330);
not(notn19330,n14271);
and (s0n19330,notn19330,1'b0);
and (s1n19330,n14271,n19331);
and (n19331,n19332,n14385);
wire s0n19332,s1n19332,notn19332;
or (n19332,s0n19332,s1n19332);
not(notn19332,n2799);
and (s0n19332,notn19332,1'b0);
and (s1n19332,n2799,n19333);
and (n19333,n17453,n13897);
wire s0n19334,s1n19334,notn19334;
or (n19334,s0n19334,s1n19334);
not(notn19334,n14271);
and (s0n19334,notn19334,1'b0);
and (s1n19334,n14271,n19335);
and (n19335,n19336,n14385);
wire s0n19336,s1n19336,notn19336;
or (n19336,s0n19336,s1n19336);
not(notn19336,n2799);
and (s0n19336,notn19336,1'b0);
and (s1n19336,n2799,n19337);
and (n19337,n19338,n13897);
or (n19339,n19340,n19341,n19342);
and (n19340,n19251,n19255);
and (n19341,n19255,n19260);
and (n19342,n19251,n19260);
or (n19343,n19344,n19345,n19346);
and (n19344,n19198,n19248);
and (n19345,n19248,n19264);
and (n19346,n19198,n19264);
and (n19347,n19196,n19268);
xor (n19348,n19349,n19420);
xor (n19349,n19350,n19416);
xor (n19350,n19351,n19401);
wire s0n19351,s1n19351,notn19351;
or (n19351,s0n19351,s1n19351);
not(notn19351,n18690);
and (s0n19351,notn19351,n19352);
and (s1n19351,n18690,1'b0);
xor (n19352,n19353,n19397);
xor (n19353,n19354,n19381);
wire s0n19354,s1n19354,notn19354;
or (n19354,s0n19354,s1n19354);
not(notn19354,n14631);
and (s0n19354,notn19354,n19355);
and (s1n19354,n14631,n19378);
wire s0n19355,s1n19355,notn19355;
or (n19355,s0n19355,s1n19355);
not(notn19355,n14271);
and (s0n19355,notn19355,n19356);
and (s1n19355,n14271,n19370);
wire s0n19356,s1n19356,notn19356;
or (n19356,s0n19356,s1n19356);
not(notn19356,n14279);
and (s0n19356,notn19356,1'b0);
and (s1n19356,n14279,n19357);
or (n19357,n19358,1'b0,1'b0,n19362);
and (n19358,n19359,n14120);
wire s0n19359,s1n19359,notn19359;
or (n19359,s0n19359,s1n19359);
not(notn19359,n14125);
and (s0n19359,notn19359,1'b0);
and (s1n19359,n14125,n19360);
wire s0n19360,s1n19360,notn19360;
or (n19360,s0n19360,s1n19360);
not(notn19360,n14317);
and (s0n19360,notn19360,n19361);
and (s1n19360,n14317,n17501);
and (n19362,n19363,n14367);
or (n19363,n19364,n19366,n19369,1'b0);
and (n19364,n19365,n17758);
wire s0n19365,s1n19365,notn19365;
or (n19365,s0n19365,s1n19365);
not(notn19365,n13900);
and (s0n19365,notn19365,1'b0);
and (s1n19365,n13900,n19361);
and (n19366,n19367,n17762);
wire s0n19367,s1n19367,notn19367;
or (n19367,s0n19367,s1n19367);
not(notn19367,n13900);
and (s0n19367,notn19367,1'b0);
and (s1n19367,n13900,n19368);
and (n19369,n19365,n17765);
or (n19370,n19371,n19372,1'b0,1'b0);
and (n19371,n19359,n13907);
and (n19372,n19373,n14385);
wire s0n19373,s1n19373,notn19373;
or (n19373,s0n19373,s1n19373);
not(notn19373,n2799);
and (s0n19373,notn19373,1'b0);
and (s1n19373,n2799,n19374);
or (n19374,1'b0,n19375,n19377,1'b0);
and (n19375,n19376,n13889);
wire s0n19376,s1n19376,notn19376;
or (n19376,s0n19376,s1n19376);
not(notn19376,n17767);
and (s0n19376,notn19376,n19361);
and (s1n19376,n17767,1'b0);
and (n19377,n19361,n14243);
and (n19378,n19379,n17820);
and (n19379,n19380,n13900);
wire s0n19380,s1n19380,notn19380;
or (n19380,s0n19380,s1n19380);
not(notn19380,n17823);
and (s0n19380,notn19380,1'b0);
and (s1n19380,n17823,n19361);
wire s0n19381,s1n19381,notn19381;
or (n19381,s0n19381,s1n19381);
not(notn19381,n14631);
and (s0n19381,notn19381,n19382);
and (s1n19381,n14631,n19394);
wire s0n19382,s1n19382,notn19382;
or (n19382,s0n19382,s1n19382);
not(notn19382,n14271);
and (s0n19382,notn19382,n19383);
and (s1n19382,n14271,n19387);
wire s0n19383,s1n19383,notn19383;
or (n19383,s0n19383,s1n19383);
not(notn19383,n14279);
and (s0n19383,notn19383,1'b0);
and (s1n19383,n14279,n19384);
or (n19384,n17512,1'b0,n19385);
and (n19385,n19386,n14367);
and (n19386,n19367,n17758);
or (n19387,n19388,n19391,1'b0);
and (n19388,n19389,n13907);
wire s0n19389,s1n19389,notn19389;
or (n19389,s0n19389,s1n19389);
not(notn19389,n14125);
and (s0n19389,notn19389,1'b0);
and (s1n19389,n14125,n19390);
wire s0n19390,s1n19390,notn19390;
or (n19390,s0n19390,s1n19390);
not(notn19390,n14563);
and (s0n19390,notn19390,n17515);
and (s1n19390,n14563,n17516);
and (n19391,n19392,n14385);
wire s0n19392,s1n19392,notn19392;
or (n19392,s0n19392,s1n19392);
not(notn19392,n2799);
and (s0n19392,notn19392,1'b0);
and (s1n19392,n2799,n19393);
and (n19393,n19368,n14235);
and (n19394,n19395,n17820);
and (n19395,n19396,n13900);
wire s0n19396,s1n19396,notn19396;
or (n19396,s0n19396,s1n19396);
not(notn19396,n17818);
and (s0n19396,notn19396,1'b0);
and (s1n19396,n17818,n19368);
or (n19397,n19398,n19399,n19400);
and (n19398,n19281,n19308);
and (n19399,n19308,n19324);
and (n19400,n19281,n19324);
xor (n19401,n19402,n19412);
xor (n19402,n19403,n19407);
wire s0n19403,s1n19403,notn19403;
or (n19403,s0n19403,s1n19403);
not(notn19403,n14271);
and (s0n19403,notn19403,1'b0);
and (s1n19403,n14271,n19404);
and (n19404,n19405,n14385);
wire s0n19405,s1n19405,notn19405;
or (n19405,s0n19405,s1n19405);
not(notn19405,n2799);
and (s0n19405,notn19405,1'b0);
and (s1n19405,n2799,n19406);
and (n19406,n17499,n13897);
wire s0n19407,s1n19407,notn19407;
or (n19407,s0n19407,s1n19407);
not(notn19407,n14271);
and (s0n19407,notn19407,1'b0);
and (s1n19407,n14271,n19408);
and (n19408,n19409,n14385);
wire s0n19409,s1n19409,notn19409;
or (n19409,s0n19409,s1n19409);
not(notn19409,n2799);
and (s0n19409,notn19409,1'b0);
and (s1n19409,n2799,n19410);
and (n19410,n19411,n13897);
or (n19412,n19413,n19414,n19415);
and (n19413,n19330,n19334);
and (n19414,n19334,n19339);
and (n19415,n19330,n19339);
or (n19416,n19417,n19418,n19419);
and (n19417,n19278,n19328);
and (n19418,n19328,n19343);
and (n19419,n19278,n19343);
and (n19420,n19276,n19347);
wire s0n19421,s1n19421,notn19421;
or (n19421,s0n19421,s1n19421);
not(notn19421,n14631);
and (s0n19421,notn19421,n19422);
and (s1n19421,n14631,n19426);
wire s0n19422,s1n19422,notn19422;
or (n19422,s0n19422,s1n19422);
not(notn19422,n14279);
and (s0n19422,notn19422,1'b0);
and (s1n19422,n14279,n19423);
and (n19423,n19424,n14367);
or (n19424,n19425,n19179,1'b0);
and (n19425,n13900,n17758);
or (n19426,n17067,1'b0,n19060,1'b0,n19062,n17297,n19427,1'b0);
and (n19427,n19428,n17820);
and (n19428,n19429,n13900);
not (n19429,n17832);
wire s0n19430,s1n19430,notn19430;
or (n19430,s0n19430,s1n19430);
not(notn19430,n19421);
and (s0n19430,notn19430,n19431);
and (s1n19430,n19421,n19572);
wire s0n19431,s1n19431,notn19431;
or (n19431,s0n19431,s1n19431);
not(notn19431,n19269);
and (s0n19431,notn19431,n19432);
and (s1n19431,n19269,n19502);
xor (n19432,n19433,n19501);
xor (n19433,n19434,n19497);
xor (n19434,n19435,n19482);
wire s0n19435,s1n19435,notn19435;
or (n19435,s0n19435,s1n19435);
not(notn19435,n18690);
and (s0n19435,notn19435,n19436);
and (s1n19435,n18690,1'b0);
xor (n19436,n19437,n19478);
xor (n19437,n19438,n19465);
wire s0n19438,s1n19438,notn19438;
or (n19438,s0n19438,s1n19438);
not(notn19438,n14631);
and (s0n19438,notn19438,n19439);
and (s1n19438,n14631,n19462);
wire s0n19439,s1n19439,notn19439;
or (n19439,s0n19439,s1n19439);
not(notn19439,n14271);
and (s0n19439,notn19439,n19440);
and (s1n19439,n14271,n19454);
wire s0n19440,s1n19440,notn19440;
or (n19440,s0n19440,s1n19440);
not(notn19440,n14279);
and (s0n19440,notn19440,1'b0);
and (s1n19440,n14279,n19441);
or (n19441,n19442,1'b0,1'b0,n19446);
and (n19442,n19443,n14120);
wire s0n19443,s1n19443,notn19443;
or (n19443,s0n19443,s1n19443);
not(notn19443,n14125);
and (s0n19443,notn19443,1'b0);
and (s1n19443,n14125,n19444);
wire s0n19444,s1n19444,notn19444;
or (n19444,s0n19444,s1n19444);
not(notn19444,n14317);
and (s0n19444,notn19444,n19445);
and (s1n19444,n14317,n17548);
and (n19446,n19447,n14367);
or (n19447,n19448,n19450,n19453,1'b0);
and (n19448,n19449,n17758);
wire s0n19449,s1n19449,notn19449;
or (n19449,s0n19449,s1n19449);
not(notn19449,n13900);
and (s0n19449,notn19449,1'b0);
and (s1n19449,n13900,n19445);
and (n19450,n19451,n17762);
wire s0n19451,s1n19451,notn19451;
or (n19451,s0n19451,s1n19451);
not(notn19451,n13900);
and (s0n19451,notn19451,1'b0);
and (s1n19451,n13900,n19452);
and (n19453,n19449,n17765);
or (n19454,n19455,n19456,1'b0,1'b0);
and (n19455,n19443,n13907);
and (n19456,n19457,n14385);
wire s0n19457,s1n19457,notn19457;
or (n19457,s0n19457,s1n19457);
not(notn19457,n2799);
and (s0n19457,notn19457,1'b0);
and (s1n19457,n2799,n19458);
or (n19458,1'b0,n19459,n19461,1'b0);
and (n19459,n19460,n13889);
wire s0n19460,s1n19460,notn19460;
or (n19460,s0n19460,s1n19460);
not(notn19460,n17767);
and (s0n19460,notn19460,n19445);
and (s1n19460,n17767,1'b0);
and (n19461,n19445,n14243);
and (n19462,n19463,n17820);
and (n19463,n19464,n13900);
wire s0n19464,s1n19464,notn19464;
or (n19464,s0n19464,s1n19464);
not(notn19464,n17823);
and (s0n19464,notn19464,1'b0);
and (s1n19464,n17823,n19445);
wire s0n19465,s1n19465,notn19465;
or (n19465,s0n19465,s1n19465);
not(notn19465,n14631);
and (s0n19465,notn19465,n19466);
and (s1n19465,n14631,n19475);
wire s0n19466,s1n19466,notn19466;
or (n19466,s0n19466,s1n19466);
not(notn19466,n14271);
and (s0n19466,notn19466,n19467);
and (s1n19466,n14271,n19471);
wire s0n19467,s1n19467,notn19467;
or (n19467,s0n19467,s1n19467);
not(notn19467,n14279);
and (s0n19467,notn19467,1'b0);
and (s1n19467,n14279,n19468);
or (n19468,n17559,1'b0,n19469);
and (n19469,n19470,n14367);
and (n19470,n19451,n17758);
or (n19471,n17604,n19472,1'b0);
and (n19472,n19473,n14385);
wire s0n19473,s1n19473,notn19473;
or (n19473,s0n19473,s1n19473);
not(notn19473,n2799);
and (s0n19473,notn19473,1'b0);
and (s1n19473,n2799,n19474);
and (n19474,n19452,n14235);
and (n19475,n19476,n17820);
and (n19476,n19477,n13900);
wire s0n19477,s1n19477,notn19477;
or (n19477,s0n19477,s1n19477);
not(notn19477,n17818);
and (s0n19477,notn19477,1'b0);
and (s1n19477,n17818,n19452);
or (n19478,n19479,n19480,n19481);
and (n19479,n19354,n19381);
and (n19480,n19381,n19397);
and (n19481,n19354,n19397);
xor (n19482,n19483,n19493);
xor (n19483,n19484,n19488);
wire s0n19484,s1n19484,notn19484;
or (n19484,s0n19484,s1n19484);
not(notn19484,n14271);
and (s0n19484,notn19484,1'b0);
and (s1n19484,n14271,n19485);
and (n19485,n19486,n14385);
wire s0n19486,s1n19486,notn19486;
or (n19486,s0n19486,s1n19486);
not(notn19486,n2799);
and (s0n19486,notn19486,1'b0);
and (s1n19486,n2799,n19487);
and (n19487,n17546,n13897);
wire s0n19488,s1n19488,notn19488;
or (n19488,s0n19488,s1n19488);
not(notn19488,n14271);
and (s0n19488,notn19488,1'b0);
and (s1n19488,n14271,n19489);
and (n19489,n19490,n14385);
wire s0n19490,s1n19490,notn19490;
or (n19490,s0n19490,s1n19490);
not(notn19490,n2799);
and (s0n19490,notn19490,1'b0);
and (s1n19490,n2799,n19491);
and (n19491,n19492,n13897);
or (n19493,n19494,n19495,n19496);
and (n19494,n19403,n19407);
and (n19495,n19407,n19412);
and (n19496,n19403,n19412);
or (n19497,n19498,n19499,n19500);
and (n19498,n19351,n19401);
and (n19499,n19401,n19416);
and (n19500,n19351,n19416);
and (n19501,n19349,n19420);
xor (n19502,n19503,n19571);
xor (n19503,n19504,n19567);
xor (n19504,n19505,n19552);
wire s0n19505,s1n19505,notn19505;
or (n19505,s0n19505,s1n19505);
not(notn19505,n18690);
and (s0n19505,notn19505,n19506);
and (s1n19505,n18690,1'b0);
xor (n19506,n19507,n19548);
xor (n19507,n19508,n19535);
wire s0n19508,s1n19508,notn19508;
or (n19508,s0n19508,s1n19508);
not(notn19508,n14631);
and (s0n19508,notn19508,n19509);
and (s1n19508,n14631,n19532);
wire s0n19509,s1n19509,notn19509;
or (n19509,s0n19509,s1n19509);
not(notn19509,n14271);
and (s0n19509,notn19509,n19510);
and (s1n19509,n14271,n19524);
wire s0n19510,s1n19510,notn19510;
or (n19510,s0n19510,s1n19510);
not(notn19510,n14279);
and (s0n19510,notn19510,1'b0);
and (s1n19510,n14279,n19511);
or (n19511,n19512,1'b0,1'b0,n19516);
and (n19512,n19513,n14120);
wire s0n19513,s1n19513,notn19513;
or (n19513,s0n19513,s1n19513);
not(notn19513,n14125);
and (s0n19513,notn19513,1'b0);
and (s1n19513,n14125,n19514);
wire s0n19514,s1n19514,notn19514;
or (n19514,s0n19514,s1n19514);
not(notn19514,n14317);
and (s0n19514,notn19514,n19515);
and (s1n19514,n14317,n17594);
and (n19516,n19517,n14367);
or (n19517,n19518,n19520,n19523,1'b0);
and (n19518,n19519,n17758);
wire s0n19519,s1n19519,notn19519;
or (n19519,s0n19519,s1n19519);
not(notn19519,n13900);
and (s0n19519,notn19519,1'b0);
and (s1n19519,n13900,n19515);
and (n19520,n19521,n17762);
wire s0n19521,s1n19521,notn19521;
or (n19521,s0n19521,s1n19521);
not(notn19521,n13900);
and (s0n19521,notn19521,1'b0);
and (s1n19521,n13900,n19522);
and (n19523,n19519,n17765);
or (n19524,n19525,n19526,1'b0,1'b0);
and (n19525,n19513,n13907);
and (n19526,n19527,n14385);
wire s0n19527,s1n19527,notn19527;
or (n19527,s0n19527,s1n19527);
not(notn19527,n2799);
and (s0n19527,notn19527,1'b0);
and (s1n19527,n2799,n19528);
or (n19528,1'b0,n19529,n19531,1'b0);
and (n19529,n19530,n13889);
wire s0n19530,s1n19530,notn19530;
or (n19530,s0n19530,s1n19530);
not(notn19530,n17767);
and (s0n19530,notn19530,n19515);
and (s1n19530,n17767,1'b0);
and (n19531,n19515,n14243);
and (n19532,n19533,n17820);
and (n19533,n19534,n13900);
wire s0n19534,s1n19534,notn19534;
or (n19534,s0n19534,s1n19534);
not(notn19534,n17823);
and (s0n19534,notn19534,1'b0);
and (s1n19534,n17823,n19515);
wire s0n19535,s1n19535,notn19535;
or (n19535,s0n19535,s1n19535);
not(notn19535,n14631);
and (s0n19535,notn19535,n19536);
and (s1n19535,n14631,n19545);
wire s0n19536,s1n19536,notn19536;
or (n19536,s0n19536,s1n19536);
not(notn19536,n14271);
and (s0n19536,notn19536,n19537);
and (s1n19536,n14271,n19541);
wire s0n19537,s1n19537,notn19537;
or (n19537,s0n19537,s1n19537);
not(notn19537,n14279);
and (s0n19537,notn19537,1'b0);
and (s1n19537,n14279,n19538);
or (n19538,n17559,1'b0,n19539);
and (n19539,n19540,n14367);
and (n19540,n19521,n17758);
or (n19541,n17604,n19542,1'b0);
and (n19542,n19543,n14385);
wire s0n19543,s1n19543,notn19543;
or (n19543,s0n19543,s1n19543);
not(notn19543,n2799);
and (s0n19543,notn19543,1'b0);
and (s1n19543,n2799,n19544);
and (n19544,n19522,n14235);
and (n19545,n19546,n17820);
and (n19546,n19547,n13900);
wire s0n19547,s1n19547,notn19547;
or (n19547,s0n19547,s1n19547);
not(notn19547,n17818);
and (s0n19547,notn19547,1'b0);
and (s1n19547,n17818,n19522);
or (n19548,n19549,n19550,n19551);
and (n19549,n19438,n19465);
and (n19550,n19465,n19478);
and (n19551,n19438,n19478);
xor (n19552,n19553,n19563);
xor (n19553,n19554,n19558);
wire s0n19554,s1n19554,notn19554;
or (n19554,s0n19554,s1n19554);
not(notn19554,n14271);
and (s0n19554,notn19554,1'b0);
and (s1n19554,n14271,n19555);
and (n19555,n19556,n14385);
wire s0n19556,s1n19556,notn19556;
or (n19556,s0n19556,s1n19556);
not(notn19556,n2799);
and (s0n19556,notn19556,1'b0);
and (s1n19556,n2799,n19557);
and (n19557,n17592,n13897);
wire s0n19558,s1n19558,notn19558;
or (n19558,s0n19558,s1n19558);
not(notn19558,n14271);
and (s0n19558,notn19558,1'b0);
and (s1n19558,n14271,n19559);
and (n19559,n19560,n14385);
wire s0n19560,s1n19560,notn19560;
or (n19560,s0n19560,s1n19560);
not(notn19560,n2799);
and (s0n19560,notn19560,1'b0);
and (s1n19560,n2799,n19561);
and (n19561,n19562,n13897);
or (n19563,n19564,n19565,n19566);
and (n19564,n19484,n19488);
and (n19565,n19488,n19493);
and (n19566,n19484,n19493);
or (n19567,n19568,n19569,n19570);
and (n19568,n19435,n19482);
and (n19569,n19482,n19497);
and (n19570,n19435,n19497);
and (n19571,n19433,n19501);
wire s0n19572,s1n19572,notn19572;
or (n19572,s0n19572,s1n19572);
not(notn19572,n19269);
and (s0n19572,notn19572,n19573);
and (s1n19572,n19269,n19643);
xor (n19573,n19574,n19642);
xor (n19574,n19575,n19638);
xor (n19575,n19576,n19623);
wire s0n19576,s1n19576,notn19576;
or (n19576,s0n19576,s1n19576);
not(notn19576,n18690);
and (s0n19576,notn19576,n19577);
and (s1n19576,n18690,1'b0);
xor (n19577,n19578,n19619);
xor (n19578,n19579,n19606);
wire s0n19579,s1n19579,notn19579;
or (n19579,s0n19579,s1n19579);
not(notn19579,n14631);
and (s0n19579,notn19579,n19580);
and (s1n19579,n14631,n19603);
wire s0n19580,s1n19580,notn19580;
or (n19580,s0n19580,s1n19580);
not(notn19580,n14271);
and (s0n19580,notn19580,n19581);
and (s1n19580,n14271,n19595);
wire s0n19581,s1n19581,notn19581;
or (n19581,s0n19581,s1n19581);
not(notn19581,n14279);
and (s0n19581,notn19581,1'b0);
and (s1n19581,n14279,n19582);
or (n19582,n19583,1'b0,1'b0,n19587);
and (n19583,n19584,n14120);
wire s0n19584,s1n19584,notn19584;
or (n19584,s0n19584,s1n19584);
not(notn19584,n14125);
and (s0n19584,notn19584,1'b0);
and (s1n19584,n14125,n19585);
wire s0n19585,s1n19585,notn19585;
or (n19585,s0n19585,s1n19585);
not(notn19585,n14317);
and (s0n19585,notn19585,n19586);
and (s1n19585,n14317,n17636);
and (n19587,n19588,n14367);
or (n19588,n19589,n19591,n19594,1'b0);
and (n19589,n19590,n17758);
wire s0n19590,s1n19590,notn19590;
or (n19590,s0n19590,s1n19590);
not(notn19590,n13900);
and (s0n19590,notn19590,1'b0);
and (s1n19590,n13900,n19586);
and (n19591,n19592,n17762);
wire s0n19592,s1n19592,notn19592;
or (n19592,s0n19592,s1n19592);
not(notn19592,n13900);
and (s0n19592,notn19592,1'b0);
and (s1n19592,n13900,n19593);
and (n19594,n19590,n17765);
or (n19595,n19596,n19597,1'b0,1'b0);
and (n19596,n19584,n13907);
and (n19597,n19598,n14385);
wire s0n19598,s1n19598,notn19598;
or (n19598,s0n19598,s1n19598);
not(notn19598,n2799);
and (s0n19598,notn19598,1'b0);
and (s1n19598,n2799,n19599);
or (n19599,1'b0,n19600,n19602,1'b0);
and (n19600,n19601,n13889);
wire s0n19601,s1n19601,notn19601;
or (n19601,s0n19601,s1n19601);
not(notn19601,n17767);
and (s0n19601,notn19601,n19586);
and (s1n19601,n17767,1'b0);
and (n19602,n19586,n14243);
and (n19603,n19604,n17820);
and (n19604,n19605,n13900);
wire s0n19605,s1n19605,notn19605;
or (n19605,s0n19605,s1n19605);
not(notn19605,n17823);
and (s0n19605,notn19605,1'b0);
and (s1n19605,n17823,n19586);
wire s0n19606,s1n19606,notn19606;
or (n19606,s0n19606,s1n19606);
not(notn19606,n14631);
and (s0n19606,notn19606,n19607);
and (s1n19606,n14631,n19616);
wire s0n19607,s1n19607,notn19607;
or (n19607,s0n19607,s1n19607);
not(notn19607,n14271);
and (s0n19607,notn19607,n19608);
and (s1n19607,n14271,n19612);
wire s0n19608,s1n19608,notn19608;
or (n19608,s0n19608,s1n19608);
not(notn19608,n14279);
and (s0n19608,notn19608,1'b0);
and (s1n19608,n14279,n19609);
or (n19609,n17559,1'b0,n19610);
and (n19610,n19611,n14367);
and (n19611,n19592,n17758);
or (n19612,n17604,n19613,1'b0);
and (n19613,n19614,n14385);
wire s0n19614,s1n19614,notn19614;
or (n19614,s0n19614,s1n19614);
not(notn19614,n2799);
and (s0n19614,notn19614,1'b0);
and (s1n19614,n2799,n19615);
and (n19615,n19593,n14235);
and (n19616,n19617,n17820);
and (n19617,n19618,n13900);
wire s0n19618,s1n19618,notn19618;
or (n19618,s0n19618,s1n19618);
not(notn19618,n17818);
and (s0n19618,notn19618,1'b0);
and (s1n19618,n17818,n19593);
or (n19619,n19620,n19621,n19622);
and (n19620,n19508,n19535);
and (n19621,n19535,n19548);
and (n19622,n19508,n19548);
xor (n19623,n19624,n19634);
xor (n19624,n19625,n19629);
wire s0n19625,s1n19625,notn19625;
or (n19625,s0n19625,s1n19625);
not(notn19625,n14271);
and (s0n19625,notn19625,1'b0);
and (s1n19625,n14271,n19626);
and (n19626,n19627,n14385);
wire s0n19627,s1n19627,notn19627;
or (n19627,s0n19627,s1n19627);
not(notn19627,n2799);
and (s0n19627,notn19627,1'b0);
and (s1n19627,n2799,n19628);
and (n19628,n17634,n13897);
wire s0n19629,s1n19629,notn19629;
or (n19629,s0n19629,s1n19629);
not(notn19629,n14271);
and (s0n19629,notn19629,1'b0);
and (s1n19629,n14271,n19630);
and (n19630,n19631,n14385);
wire s0n19631,s1n19631,notn19631;
or (n19631,s0n19631,s1n19631);
not(notn19631,n2799);
and (s0n19631,notn19631,1'b0);
and (s1n19631,n2799,n19632);
and (n19632,n19633,n13897);
or (n19634,n19635,n19636,n19637);
and (n19635,n19554,n19558);
and (n19636,n19558,n19563);
and (n19637,n19554,n19563);
or (n19638,n19639,n19640,n19641);
and (n19639,n19505,n19552);
and (n19640,n19552,n19567);
and (n19641,n19505,n19567);
and (n19642,n19503,n19571);
xor (n19643,n19644,n19712);
xor (n19644,n19645,n19708);
xor (n19645,n19646,n19693);
wire s0n19646,s1n19646,notn19646;
or (n19646,s0n19646,s1n19646);
not(notn19646,n18690);
and (s0n19646,notn19646,n19647);
and (s1n19646,n18690,1'b0);
xor (n19647,n19648,n19689);
xor (n19648,n19649,n19676);
wire s0n19649,s1n19649,notn19649;
or (n19649,s0n19649,s1n19649);
not(notn19649,n14631);
and (s0n19649,notn19649,n19650);
and (s1n19649,n14631,n19673);
wire s0n19650,s1n19650,notn19650;
or (n19650,s0n19650,s1n19650);
not(notn19650,n14271);
and (s0n19650,notn19650,n19651);
and (s1n19650,n14271,n19665);
wire s0n19651,s1n19651,notn19651;
or (n19651,s0n19651,s1n19651);
not(notn19651,n14279);
and (s0n19651,notn19651,1'b0);
and (s1n19651,n14279,n19652);
or (n19652,n19653,1'b0,1'b0,n19657);
and (n19653,n19654,n14120);
wire s0n19654,s1n19654,notn19654;
or (n19654,s0n19654,s1n19654);
not(notn19654,n14125);
and (s0n19654,notn19654,1'b0);
and (s1n19654,n14125,n19655);
wire s0n19655,s1n19655,notn19655;
or (n19655,s0n19655,s1n19655);
not(notn19655,n14317);
and (s0n19655,notn19655,n19656);
and (s1n19655,n14317,n17667);
and (n19657,n19658,n14367);
or (n19658,n19659,n19661,n19664,1'b0);
and (n19659,n19660,n17758);
wire s0n19660,s1n19660,notn19660;
or (n19660,s0n19660,s1n19660);
not(notn19660,n13900);
and (s0n19660,notn19660,1'b0);
and (s1n19660,n13900,n19656);
and (n19661,n19662,n17762);
wire s0n19662,s1n19662,notn19662;
or (n19662,s0n19662,s1n19662);
not(notn19662,n13900);
and (s0n19662,notn19662,1'b0);
and (s1n19662,n13900,n19663);
and (n19664,n19660,n17765);
or (n19665,n19666,n19667,1'b0,1'b0);
and (n19666,n19654,n13907);
and (n19667,n19668,n14385);
wire s0n19668,s1n19668,notn19668;
or (n19668,s0n19668,s1n19668);
not(notn19668,n2799);
and (s0n19668,notn19668,1'b0);
and (s1n19668,n2799,n19669);
or (n19669,1'b0,n19670,n19672,1'b0);
and (n19670,n19671,n13889);
wire s0n19671,s1n19671,notn19671;
or (n19671,s0n19671,s1n19671);
not(notn19671,n17767);
and (s0n19671,notn19671,n19656);
and (s1n19671,n17767,1'b0);
and (n19672,n19656,n14243);
and (n19673,n19674,n17820);
and (n19674,n19675,n13900);
wire s0n19675,s1n19675,notn19675;
or (n19675,s0n19675,s1n19675);
not(notn19675,n17823);
and (s0n19675,notn19675,1'b0);
and (s1n19675,n17823,n19656);
wire s0n19676,s1n19676,notn19676;
or (n19676,s0n19676,s1n19676);
not(notn19676,n14631);
and (s0n19676,notn19676,n19677);
and (s1n19676,n14631,n19686);
wire s0n19677,s1n19677,notn19677;
or (n19677,s0n19677,s1n19677);
not(notn19677,n14271);
and (s0n19677,notn19677,n19678);
and (s1n19677,n14271,n19682);
wire s0n19678,s1n19678,notn19678;
or (n19678,s0n19678,s1n19678);
not(notn19678,n14279);
and (s0n19678,notn19678,1'b0);
and (s1n19678,n14279,n19679);
or (n19679,n17559,1'b0,n19680);
and (n19680,n19681,n14367);
and (n19681,n19662,n17758);
or (n19682,n17604,n19683,1'b0);
and (n19683,n19684,n14385);
wire s0n19684,s1n19684,notn19684;
or (n19684,s0n19684,s1n19684);
not(notn19684,n2799);
and (s0n19684,notn19684,1'b0);
and (s1n19684,n2799,n19685);
and (n19685,n19663,n14235);
and (n19686,n19687,n17820);
and (n19687,n19688,n13900);
wire s0n19688,s1n19688,notn19688;
or (n19688,s0n19688,s1n19688);
not(notn19688,n17818);
and (s0n19688,notn19688,1'b0);
and (s1n19688,n17818,n19663);
or (n19689,n19690,n19691,n19692);
and (n19690,n19579,n19606);
and (n19691,n19606,n19619);
and (n19692,n19579,n19619);
xor (n19693,n19694,n19704);
xor (n19694,n19695,n19699);
wire s0n19695,s1n19695,notn19695;
or (n19695,s0n19695,s1n19695);
not(notn19695,n14271);
and (s0n19695,notn19695,1'b0);
and (s1n19695,n14271,n19696);
and (n19696,n19697,n14385);
wire s0n19697,s1n19697,notn19697;
or (n19697,s0n19697,s1n19697);
not(notn19697,n2799);
and (s0n19697,notn19697,1'b0);
and (s1n19697,n2799,n19698);
and (n19698,n17665,n13897);
wire s0n19699,s1n19699,notn19699;
or (n19699,s0n19699,s1n19699);
not(notn19699,n14271);
and (s0n19699,notn19699,1'b0);
and (s1n19699,n14271,n19700);
and (n19700,n19701,n14385);
wire s0n19701,s1n19701,notn19701;
or (n19701,s0n19701,s1n19701);
not(notn19701,n2799);
and (s0n19701,notn19701,1'b0);
and (s1n19701,n2799,n19702);
and (n19702,n19703,n13897);
or (n19704,n19705,n19706,n19707);
and (n19705,n19625,n19629);
and (n19706,n19629,n19634);
and (n19707,n19625,n19634);
or (n19708,n19709,n19710,n19711);
and (n19709,n19576,n19623);
and (n19710,n19623,n19638);
and (n19711,n19576,n19638);
and (n19712,n19574,n19642);
wire s0n19713,s1n19713,notn19713;
or (n19713,s0n19713,s1n19713);
not(notn19713,n14271);
and (s0n19713,notn19713,n14504);
and (s1n19713,n14271,n19714);
or (n19714,n14506,n19715,1'b0);
and (n19715,n19716,n14385);
wire s0n19716,s1n19716,notn19716;
or (n19716,s0n19716,s1n19716);
not(notn19716,n2799);
and (s0n19716,notn19716,1'b0);
and (s1n19716,n2799,n13889);
wire s0n19717,s1n19717,notn19717;
or (n19717,s0n19717,s1n19717);
not(notn19717,n19812);
and (s0n19717,notn19717,n19718);
and (s1n19717,n19812,1'b0);
wire s0n19718,s1n19718,notn19718;
or (n19718,s0n19718,s1n19718);
not(notn19718,n19719);
and (s0n19718,notn19718,1'b1);
and (s1n19718,n19719,n17727);
nor (n19719,n19720,n19797,n19802,n19806,n19808,n19810,n19811,n19812);
wire s0n19720,s1n19720,notn19720;
or (n19720,s0n19720,s1n19720);
not(notn19720,n19713);
and (s0n19720,notn19720,n19721);
and (s1n19720,n19713,n19724);
wire s0n19721,s1n19721,notn19721;
or (n19721,s0n19721,s1n19721);
not(notn19721,n19421);
and (s0n19721,notn19721,n19722);
and (s1n19721,n19421,n19723);
wire s0n19722,s1n19722,notn19722;
or (n19722,s0n19722,s1n19722);
not(notn19722,n19269);
and (s0n19722,notn19722,n19195);
and (s1n19722,n19269,n19275);
wire s0n19723,s1n19723,notn19723;
or (n19723,s0n19723,s1n19723);
not(notn19723,n19269);
and (s0n19723,notn19723,n19348);
and (s1n19723,n19269,n19432);
wire s0n19724,s1n19724,notn19724;
or (n19724,s0n19724,s1n19724);
not(notn19724,n19421);
and (s0n19724,notn19724,n19725);
and (s1n19724,n19421,n19726);
wire s0n19725,s1n19725,notn19725;
or (n19725,s0n19725,s1n19725);
not(notn19725,n19269);
and (s0n19725,notn19725,n19502);
and (s1n19725,n19269,n19573);
wire s0n19726,s1n19726,notn19726;
or (n19726,s0n19726,s1n19726);
not(notn19726,n19269);
and (s0n19726,notn19726,n19643);
and (s1n19726,n19269,n19727);
xor (n19727,n19728,n19796);
xor (n19728,n19729,n19792);
xor (n19729,n19730,n19777);
wire s0n19730,s1n19730,notn19730;
or (n19730,s0n19730,s1n19730);
not(notn19730,n18690);
and (s0n19730,notn19730,n19731);
and (s1n19730,n18690,1'b0);
xor (n19731,n19732,n19773);
xor (n19732,n19733,n19760);
wire s0n19733,s1n19733,notn19733;
or (n19733,s0n19733,s1n19733);
not(notn19733,n14631);
and (s0n19733,notn19733,n19734);
and (s1n19733,n14631,n19757);
wire s0n19734,s1n19734,notn19734;
or (n19734,s0n19734,s1n19734);
not(notn19734,n14271);
and (s0n19734,notn19734,n19735);
and (s1n19734,n14271,n19749);
wire s0n19735,s1n19735,notn19735;
or (n19735,s0n19735,s1n19735);
not(notn19735,n14279);
and (s0n19735,notn19735,1'b0);
and (s1n19735,n14279,n19736);
or (n19736,n19737,1'b0,1'b0,n19741);
and (n19737,n19738,n14120);
wire s0n19738,s1n19738,notn19738;
or (n19738,s0n19738,s1n19738);
not(notn19738,n14125);
and (s0n19738,notn19738,1'b0);
and (s1n19738,n14125,n19739);
wire s0n19739,s1n19739,notn19739;
or (n19739,s0n19739,s1n19739);
not(notn19739,n14317);
and (s0n19739,notn19739,n19740);
and (s1n19739,n14317,n17697);
and (n19741,n19742,n14367);
or (n19742,n19743,n19745,n19748,1'b0);
and (n19743,n19744,n17758);
wire s0n19744,s1n19744,notn19744;
or (n19744,s0n19744,s1n19744);
not(notn19744,n13900);
and (s0n19744,notn19744,1'b0);
and (s1n19744,n13900,n19740);
and (n19745,n19746,n17762);
wire s0n19746,s1n19746,notn19746;
or (n19746,s0n19746,s1n19746);
not(notn19746,n13900);
and (s0n19746,notn19746,1'b0);
and (s1n19746,n13900,n19747);
and (n19748,n19744,n17765);
or (n19749,n19750,n19751,1'b0,1'b0);
and (n19750,n19738,n13907);
and (n19751,n19752,n14385);
wire s0n19752,s1n19752,notn19752;
or (n19752,s0n19752,s1n19752);
not(notn19752,n2799);
and (s0n19752,notn19752,1'b0);
and (s1n19752,n2799,n19753);
or (n19753,1'b0,n19754,n19756,1'b0);
and (n19754,n19755,n13889);
wire s0n19755,s1n19755,notn19755;
or (n19755,s0n19755,s1n19755);
not(notn19755,n17767);
and (s0n19755,notn19755,n19740);
and (s1n19755,n17767,1'b0);
and (n19756,n19740,n14243);
and (n19757,n19758,n17820);
and (n19758,n19759,n13900);
wire s0n19759,s1n19759,notn19759;
or (n19759,s0n19759,s1n19759);
not(notn19759,n17823);
and (s0n19759,notn19759,1'b0);
and (s1n19759,n17823,n19740);
wire s0n19760,s1n19760,notn19760;
or (n19760,s0n19760,s1n19760);
not(notn19760,n14631);
and (s0n19760,notn19760,n19761);
and (s1n19760,n14631,n19770);
wire s0n19761,s1n19761,notn19761;
or (n19761,s0n19761,s1n19761);
not(notn19761,n14271);
and (s0n19761,notn19761,n19762);
and (s1n19761,n14271,n19766);
wire s0n19762,s1n19762,notn19762;
or (n19762,s0n19762,s1n19762);
not(notn19762,n14279);
and (s0n19762,notn19762,1'b0);
and (s1n19762,n14279,n19763);
or (n19763,n17559,1'b0,n19764);
and (n19764,n19765,n14367);
and (n19765,n19746,n17758);
or (n19766,n17604,n19767,1'b0);
and (n19767,n19768,n14385);
wire s0n19768,s1n19768,notn19768;
or (n19768,s0n19768,s1n19768);
not(notn19768,n2799);
and (s0n19768,notn19768,1'b0);
and (s1n19768,n2799,n19769);
and (n19769,n19747,n14235);
and (n19770,n19771,n17820);
and (n19771,n19772,n13900);
wire s0n19772,s1n19772,notn19772;
or (n19772,s0n19772,s1n19772);
not(notn19772,n17818);
and (s0n19772,notn19772,1'b0);
and (s1n19772,n17818,n19747);
or (n19773,n19774,n19775,n19776);
and (n19774,n19649,n19676);
and (n19775,n19676,n19689);
and (n19776,n19649,n19689);
xor (n19777,n19778,n19788);
xor (n19778,n19779,n19783);
wire s0n19779,s1n19779,notn19779;
or (n19779,s0n19779,s1n19779);
not(notn19779,n14271);
and (s0n19779,notn19779,1'b0);
and (s1n19779,n14271,n19780);
and (n19780,n19781,n14385);
wire s0n19781,s1n19781,notn19781;
or (n19781,s0n19781,s1n19781);
not(notn19781,n2799);
and (s0n19781,notn19781,1'b0);
and (s1n19781,n2799,n19782);
and (n19782,n17695,n13897);
wire s0n19783,s1n19783,notn19783;
or (n19783,s0n19783,s1n19783);
not(notn19783,n14271);
and (s0n19783,notn19783,1'b0);
and (s1n19783,n14271,n19784);
and (n19784,n19785,n14385);
wire s0n19785,s1n19785,notn19785;
or (n19785,s0n19785,s1n19785);
not(notn19785,n2799);
and (s0n19785,notn19785,1'b0);
and (s1n19785,n2799,n19786);
and (n19786,n19787,n13897);
or (n19788,n19789,n19790,n19791);
and (n19789,n19695,n19699);
and (n19790,n19699,n19704);
and (n19791,n19695,n19704);
or (n19792,n19793,n19794,n19795);
and (n19793,n19646,n19693);
and (n19794,n19693,n19708);
and (n19795,n19646,n19708);
and (n19796,n19644,n19712);
wire s0n19797,s1n19797,notn19797;
or (n19797,s0n19797,s1n19797);
not(notn19797,n19713);
and (s0n19797,notn19797,n19798);
and (s1n19797,n19713,n19799);
wire s0n19798,s1n19798,notn19798;
or (n19798,s0n19798,s1n19798);
not(notn19798,n19421);
and (s0n19798,notn19798,n19274);
and (s1n19798,n19421,n19431);
wire s0n19799,s1n19799,notn19799;
or (n19799,s0n19799,s1n19799);
not(notn19799,n19421);
and (s0n19799,notn19799,n19572);
and (s1n19799,n19421,n19800);
wire s0n19800,s1n19800,notn19800;
or (n19800,s0n19800,s1n19800);
not(notn19800,n19269);
and (s0n19800,notn19800,n19727);
and (s1n19800,n19269,n19801);
and (n19801,n19728,n19796);
wire s0n19802,s1n19802,notn19802;
or (n19802,s0n19802,s1n19802);
not(notn19802,n19713);
and (s0n19802,notn19802,n19803);
and (s1n19802,n19713,n19804);
wire s0n19803,s1n19803,notn19803;
or (n19803,s0n19803,s1n19803);
not(notn19803,n19421);
and (s0n19803,notn19803,n19723);
and (s1n19803,n19421,n19725);
wire s0n19804,s1n19804,notn19804;
or (n19804,s0n19804,s1n19804);
not(notn19804,n19421);
and (s0n19804,notn19804,n19726);
and (s1n19804,n19421,n19805);
wire s0n19805,s1n19805,notn19805;
or (n19805,s0n19805,s1n19805);
not(notn19805,n19269);
and (s0n19805,notn19805,n19801);
and (s1n19805,n19269,1'b0);
wire s0n19806,s1n19806,notn19806;
or (n19806,s0n19806,s1n19806);
not(notn19806,n19713);
and (s0n19806,notn19806,n19430);
and (s1n19806,n19713,n19807);
wire s0n19807,s1n19807,notn19807;
or (n19807,s0n19807,s1n19807);
not(notn19807,n19421);
and (s0n19807,notn19807,n19800);
and (s1n19807,n19421,1'b0);
wire s0n19808,s1n19808,notn19808;
or (n19808,s0n19808,s1n19808);
not(notn19808,n19713);
and (s0n19808,notn19808,n19724);
and (s1n19808,n19713,n19809);
wire s0n19809,s1n19809,notn19809;
or (n19809,s0n19809,s1n19809);
not(notn19809,n19421);
and (s0n19809,notn19809,n19805);
and (s1n19809,n19421,1'b0);
wire s0n19810,s1n19810,notn19810;
or (n19810,s0n19810,s1n19810);
not(notn19810,n19713);
and (s0n19810,notn19810,n19799);
and (s1n19810,n19713,1'b0);
wire s0n19811,s1n19811,notn19811;
or (n19811,s0n19811,s1n19811);
not(notn19811,n19713);
and (s0n19811,notn19811,n19804);
and (s1n19811,n19713,1'b0);
wire s0n19812,s1n19812,notn19812;
or (n19812,s0n19812,s1n19812);
not(notn19812,n19713);
and (s0n19812,notn19812,n19807);
and (s1n19812,n19713,1'b0);
and (n19813,n14271,n14385);
wire s0n19814,s1n19814,notn19814;
or (n19814,s0n19814,s1n19814);
not(notn19814,n13900);
and (s0n19814,notn19814,n3);
and (s1n19814,n13900,n17725);
or (n19815,n17820,n19816);
and (n19816,n14279,n14367);
or (n19817,n19818,n19853);
and (n19818,n19819,n3);
and (n19819,n19820,n19846);
nor (n19820,n19821,n19827);
and (n19821,n19822,n19825,n559);
and (n19822,n2907,n19823,n558);
nor (n19823,n19824,n561);
not (n19824,n560);
and (n19825,n8689,n19826);
not (n19826,n14125);
nand (n19827,n19828,n19831,n19837);
or (n19828,n19829,n13863);
nand (n19829,n19830,n19825);
not (n19830,n2907);
or (n19831,n19832,n19833);
or (n19832,n13890,n13892);
not (n19833,n19834);
nor (n19834,n19835,n19826);
not (n19835,n19836);
nor (n19836,n19815,n19813);
nand (n19837,n19838,n14125);
nand (n19838,n19839,n19841);
or (n19839,n19840,n14338);
not (n19840,n19815);
nand (n19841,n19842,n19813,n19844,n19845);
not (n19842,n19843);
or (n19843,n13894,n13892);
nor (n19844,n29,n581);
nor (n19845,n28,n582);
nand (n19846,n19847,n19849);
nor (n19847,n19848,n8689,n14125);
not (n19848,n8696);
nand (n19849,n19850,n19851);
or (n19850,n577,n8691);
nand (n19851,n19852,n577,n604);
not (n19852,n605);
and (n19853,n19854,n19855);
not (n19854,n19819);
nand (n19855,n19856,n20689);
or (n19856,n19857,n19858);
not (n19857,n19847);
not (n19858,n19859);
nand (n19859,n19860,n19861);
not (n19860,n2881);
nor (n19861,n2700,n19862);
and (n19862,n19863,n20688);
nand (n19863,n19864,n20661);
not (n19864,n19865);
or (n19865,n19866,n20660);
and (n19866,n19867,n20255);
xor (n19867,n19868,n20197);
xor (n19868,n19869,n20146);
xor (n19869,n19870,n20121);
or (n19870,n19871,n20120);
and (n19871,n19872,n19991);
xor (n19872,n19873,n19966);
xor (n19873,n19874,n19907);
xor (n19874,n19875,n19877);
xor (n19875,n19876,n1160);
xor (n19876,n1083,n2011);
xor (n19877,n19878,n2265);
xor (n19878,n19879,n19905);
or (n19879,n19880,n19904);
and (n19880,n19881,n2423);
xor (n19881,n19882,n1511);
and (n19882,n19883,n1519);
xor (n19883,n1518,n19884);
xor (n19884,n19885,n19892);
xor (n19885,n19886,n19891);
xor (n19886,n19887,n19890);
xor (n19887,n19888,n19889);
and (n19888,n2081,n1027);
and (n19889,n1245,n1027);
and (n19890,n19889,n1261);
and (n19891,n19888,n2097);
or (n19892,n19893,n19903);
and (n19893,n19894,n19902);
xor (n19894,n19895,n19896);
nor (n19895,n2287,n1026);
and (n19896,n19897,n1027);
nand (n19897,n19898,n19900);
or (n19898,n19899,n1376);
not (n19899,n1258);
or (n19900,n19901,n1258);
not (n19901,n1376);
and (n19902,n2278,n1027);
and (n19903,n19895,n19896);
and (n19904,n19882,n1511);
xor (n19905,n19906,n1504);
xor (n19906,n1428,n1503);
or (n19907,n19908,n19965);
and (n19908,n19909,n19915);
xor (n19909,n19910,n19914);
or (n19910,n19911,n19913);
and (n19911,n19912,n1175);
xor (n19912,n1895,n2022);
and (n19913,n1895,n2022);
xor (n19914,n19881,n2423);
and (n19915,n19916,n1092);
xor (n19916,n1174,n19917);
or (n19917,n19918,n19964);
and (n19918,n19919,n19943);
xor (n19919,n2435,n19920);
and (n19920,n19921,n19942);
or (n19921,n19922,n19941);
and (n19922,n19923,n19932);
xor (n19923,n19924,n19925);
and (n19924,n2311,n1027);
nor (n19925,n1026,n19926);
nor (n19926,n1292,n19927);
nor (n19927,n19928,n19931);
and (n19928,n19929,n19930);
not (n19929,n1305);
not (n19930,n1293);
not (n19931,n1393);
nor (n19932,n19933,n1026);
nor (n19933,n19934,n19939);
and (n19934,n19935,n1277);
not (n19935,n19936);
xor (n19936,n19937,n19938);
not (n19937,n1387);
not (n19938,n1289);
and (n19939,n19936,n19940);
not (n19940,n1277);
and (n19941,n19924,n19925);
and (n19942,n2293,n1027);
or (n19943,n19944,n19963);
and (n19944,n19945,n2441);
xor (n19945,n1535,n19946);
xor (n19946,n19947,n19955);
xor (n19947,n19948,n19954);
and (n19948,n19949,n1027);
nand (n19949,n19950,n19952,n19953);
or (n19950,n19951,n19930);
not (n19951,n1381);
not (n19952,n1276);
or (n19953,n19937,n19938);
and (n19954,n2298,n1027);
and (n19955,n19956,n1027);
nor (n19956,n19957,n19960);
and (n19957,n19958,n1261);
xor (n19958,n19959,n19951);
not (n19959,n1273);
and (n19960,n19961,n19962);
not (n19961,n19958);
not (n19962,n1261);
and (n19963,n1535,n19946);
and (n19964,n2435,n19920);
and (n19965,n19910,n19914);
xor (n19966,n19967,n19987);
xor (n19967,n19968,n19977);
xor (n19968,n19969,n2418);
xor (n19969,n1159,n19970);
and (n19970,n19971,n19974);
or (n19971,n19972,n19973);
and (n19972,n19885,n19892);
and (n19973,n19886,n19891);
or (n19974,n19975,n19976);
and (n19975,n19887,n19890);
and (n19976,n19888,n19889);
or (n19977,n19978,n19986);
and (n19978,n19979,n1167);
xor (n19979,n19980,n2016);
or (n19980,n19981,n19985);
and (n19981,n19982,n2275);
xor (n19982,n19983,n19984);
xor (n19983,n19883,n1519);
and (n19984,n1525,n1443);
and (n19985,n19983,n19984);
and (n19986,n19980,n2016);
or (n19987,n19988,n19990);
and (n19988,n19989,n1087);
xor (n19989,n1088,n1891);
and (n19990,n1088,n1891);
or (n19991,n19992,n20119);
and (n19992,n19993,n20018);
xor (n19993,n19994,n19995);
xor (n19994,n19909,n19915);
or (n19995,n19996,n20017);
and (n19996,n19997,n20004);
xor (n19997,n19998,n19999);
xor (n19998,n19916,n1092);
or (n19999,n20000,n20003);
and (n20000,n20001,n1956);
xor (n20001,n1183,n20002);
xor (n20002,n19919,n19943);
and (n20003,n1183,n20002);
or (n20004,n20005,n20016);
and (n20005,n20006,n1099);
xor (n20006,n1952,n20007);
or (n20007,n20008,n20015);
and (n20008,n20009,n1190);
xor (n20009,n20010,n20012);
xor (n20010,n20011,n1534);
xor (n20011,n19921,n19942);
and (n20012,n20013,n2447);
xor (n20013,n20014,n1542);
xor (n20014,n19923,n19932);
and (n20015,n20010,n20012);
and (n20016,n1952,n20007);
and (n20017,n19998,n19999);
or (n20018,n20019,n20118);
and (n20019,n20020,n20100);
xor (n20020,n20021,n20099);
or (n20021,n20022,n20098);
and (n20022,n20023,n1102);
xor (n20023,n20024,n20042);
or (n20024,n20025,n20041);
and (n20025,n20026,n2034);
xor (n20026,n20027,n20028);
xor (n20027,n19945,n2441);
or (n20028,n20029,n20040);
and (n20029,n20030,n2376);
xor (n20030,n1457,n20031);
or (n20031,n20032,n20039);
and (n20032,n20033,n1551);
xor (n20033,n20034,n20035);
and (n20034,n2328,n1027);
and (n20035,n20036,n1027);
nand (n20036,n20037,n20038);
or (n20037,n19931,n1395);
nand (n20038,n1395,n19931);
and (n20039,n20034,n20035);
and (n20040,n1457,n20031);
and (n20041,n20027,n20028);
or (n20042,n20043,n20097);
and (n20043,n20044,n1191);
xor (n20044,n20045,n20061);
xor (n20045,n20046,n2369);
xor (n20046,n1450,n20047);
or (n20047,n20048,n20060);
and (n20048,n20049,n1543);
xor (n20049,n20050,n20059);
or (n20050,n20051,n20058);
and (n20051,n20052,n1027);
nand (n20052,n20053,n20055,n20057);
or (n20053,n19937,n20054);
not (n20054,n1353);
or (n20055,n19931,n20056);
not (n20056,n1325);
not (n20057,n1308);
and (n20058,n2322,n1027);
nor (n20059,n2308,n1026);
and (n20060,n20050,n20059);
and (n20061,n20062,n20096);
xor (n20062,n20063,n20094);
or (n20063,n20064,n20093);
and (n20064,n20065,n2453);
xor (n20065,n20066,n20075);
and (n20066,n20067,n20074);
xor (n20067,n20068,n1558);
and (n20068,n20069,n20071);
nor (n20069,n20070,n2341);
not (n20070,n2565);
and (n20071,n20072,n1027);
nor (n20072,n20073,n20054);
not (n20073,n1410);
and (n20074,n2340,n1027);
or (n20075,n20076,n20092);
and (n20076,n20077,n20086);
xor (n20077,n20078,n20085);
and (n20078,n20079,n1027);
nand (n20079,n20080,n20082,n20084);
or (n20080,n20081,n20056);
not (n20081,n1405);
or (n20082,n19931,n20083);
not (n20083,n1368);
not (n20084,n1324);
and (n20085,n2334,n1027);
and (n20086,n20087,n1027);
xor (n20087,n20088,n20089);
not (n20088,n1309);
xnor (n20089,n20090,n20091);
not (n20090,n1399);
not (n20091,n1321);
and (n20092,n20078,n20085);
and (n20093,n20066,n20075);
and (n20094,n20095,n1464);
xor (n20095,n2382,n1550);
xor (n20096,n20013,n2447);
and (n20097,n20045,n20061);
and (n20098,n20024,n20042);
xor (n20099,n19912,n1175);
xor (n20100,n20101,n1095);
xor (n20101,n1948,n20102);
xor (n20102,n20103,n2429);
xor (n20103,n1436,n20104);
or (n20104,n20105,n20117);
and (n20105,n20106,n20114);
xor (n20106,n20107,n20108);
xor (n20107,n19894,n19902);
and (n20108,n20109,n1027);
nand (n20109,n20110,n20112);
or (n20110,n20111,n19962);
and (n20111,n19959,n19951);
or (n20112,n19929,n20113);
not (n20113,n1245);
or (n20114,n20115,n20116);
and (n20115,n19947,n19955);
and (n20116,n19948,n19954);
and (n20117,n20107,n20108);
and (n20118,n20021,n20099);
and (n20119,n19994,n19995);
and (n20120,n19873,n19966);
xor (n20121,n20122,n20139);
xor (n20122,n20123,n20126);
or (n20123,n20124,n20125);
and (n20124,n19967,n19987);
and (n20125,n19968,n19977);
and (n20126,n20127,n20134);
xor (n20127,n20128,n1886);
or (n20128,n20129,n20133);
and (n20129,n20130,n1889);
xor (n20130,n1431,n20131);
xor (n20131,n20132,n1510);
xor (n20132,n19971,n19974);
and (n20133,n1431,n20131);
and (n20134,n20135,n2268);
xor (n20135,n1166,n20136);
or (n20136,n20137,n20138);
and (n20137,n20103,n2429);
and (n20138,n1436,n20104);
xor (n20139,n20140,n20143);
xor (n20140,n20141,n20142);
and (n20141,n19969,n2418);
and (n20142,n19906,n1504);
or (n20143,n20144,n20145);
and (n20144,n19876,n1160);
and (n20145,n1083,n2011);
xor (n20146,n20147,n20159);
xor (n20147,n20148,n20151);
or (n20148,n20149,n20150);
and (n20149,n19874,n19907);
and (n20150,n19875,n19877);
xor (n20151,n20152,n20157);
xor (n20152,n20153,n20156);
or (n20153,n20154,n20155);
and (n20154,n19878,n2265);
and (n20155,n19879,n19905);
xor (n20156,n1422,n1077);
xor (n20157,n20158,n1080);
xor (n20158,n1684,n2078);
or (n20159,n20160,n20196);
and (n20160,n20161,n20172);
xor (n20161,n20162,n20171);
or (n20162,n20163,n20170);
and (n20163,n20164,n20167);
xor (n20164,n20165,n20166);
xor (n20165,n19979,n1167);
xor (n20166,n20130,n1889);
or (n20167,n20168,n20169);
and (n20168,n20101,n1095);
and (n20169,n1948,n20102);
and (n20170,n20165,n20166);
xor (n20171,n20127,n20134);
or (n20172,n20173,n20195);
and (n20173,n20174,n20194);
xor (n20174,n20175,n20176);
xor (n20175,n20135,n2268);
or (n20176,n20177,n20193);
and (n20177,n20178,n20188);
xor (n20178,n20179,n20180);
xor (n20179,n19982,n2275);
or (n20180,n20181,n20187);
and (n20181,n20182,n2363);
xor (n20182,n20183,n20186);
or (n20183,n20184,n20185);
and (n20184,n20046,n2369);
and (n20185,n1450,n20047);
xor (n20186,n20106,n20114);
and (n20187,n20183,n20186);
or (n20188,n20189,n20192);
and (n20189,n20190,n2028);
xor (n20190,n1182,n20191);
xor (n20191,n1525,n1443);
and (n20192,n1182,n20191);
and (n20193,n20179,n20180);
xor (n20194,n19989,n1087);
and (n20195,n20175,n20176);
and (n20196,n20162,n20171);
or (n20197,n20198,n20254);
and (n20198,n20199,n20253);
xor (n20199,n20200,n20201);
xor (n20200,n20161,n20172);
or (n20201,n20202,n20252);
and (n20202,n20203,n20206);
xor (n20203,n20204,n20205);
xor (n20204,n20174,n20194);
xor (n20205,n20164,n20167);
or (n20206,n20207,n20251);
and (n20207,n20208,n20241);
xor (n20208,n20209,n20240);
or (n20209,n20210,n20239);
and (n20210,n20211,n20214);
xor (n20211,n20212,n20213);
xor (n20212,n20190,n2028);
xor (n20213,n20182,n2363);
or (n20214,n20215,n20238);
and (n20215,n20216,n1963);
xor (n20216,n20217,n20235);
or (n20217,n20218,n20234);
and (n20218,n20219,n1199);
xor (n20219,n20220,n20221);
xor (n20220,n20030,n2376);
or (n20221,n20222,n20233);
and (n20222,n20223,n20229);
xor (n20223,n20224,n20225);
xor (n20224,n20033,n1551);
nand (n20225,n20226,n20050);
or (n20226,n20227,n20228);
not (n20227,n20058);
not (n20228,n20051);
or (n20229,n20230,n20232);
and (n20230,n20231,n1471);
xor (n20231,n1559,n2459);
and (n20232,n1559,n2459);
and (n20233,n20224,n20225);
and (n20234,n20220,n20221);
and (n20235,n20236,n2040);
xor (n20236,n1198,n20237);
xor (n20237,n20049,n1543);
and (n20238,n20217,n20235);
and (n20239,n20212,n20213);
xor (n20240,n20178,n20188);
or (n20241,n20242,n20250);
and (n20242,n20243,n20249);
xor (n20243,n20244,n20245);
xor (n20244,n20001,n1956);
or (n20245,n20246,n20248);
and (n20246,n20247,n1109);
xor (n20247,n1106,n1960);
and (n20248,n1106,n1960);
xor (n20249,n20006,n1099);
and (n20250,n20244,n20245);
and (n20251,n20209,n20240);
and (n20252,n20204,n20205);
xor (n20253,n19872,n19991);
and (n20254,n20200,n20201);
or (n20255,n20256,n20659);
and (n20256,n20257,n20315);
xor (n20257,n20258,n20259);
xor (n20258,n20199,n20253);
or (n20259,n20260,n20314);
and (n20260,n20261,n20313);
xor (n20261,n20262,n20263);
xor (n20262,n19993,n20018);
or (n20263,n20264,n20312);
and (n20264,n20265,n20268);
xor (n20265,n20266,n20267);
xor (n20266,n19997,n20004);
xor (n20267,n20020,n20100);
or (n20268,n20269,n20311);
and (n20269,n20270,n20295);
xor (n20270,n20271,n20272);
xor (n20271,n20023,n1102);
or (n20272,n20273,n20294);
and (n20273,n20274,n20277);
xor (n20274,n20275,n20276);
xor (n20275,n20026,n2034);
xor (n20276,n20009,n1190);
or (n20277,n20278,n20293);
and (n20278,n20279,n1967);
xor (n20279,n20280,n1113);
and (n20280,n20281,n20282);
xor (n20281,n20065,n2453);
or (n20282,n20283,n20292);
and (n20283,n20284,n2388);
xor (n20284,n20285,n20291);
or (n20285,n20286,n20290);
and (n20286,n20287,n20289);
xor (n20287,n2465,n20288);
and (n20288,n2470,n2063);
and (n20289,n2346,n1027);
and (n20290,n2465,n20288);
xor (n20291,n20077,n20086);
and (n20292,n20285,n20291);
and (n20293,n20280,n1113);
and (n20294,n20275,n20276);
or (n20295,n20296,n20310);
and (n20296,n20297,n20309);
xor (n20297,n20298,n20299);
xor (n20298,n20044,n1191);
or (n20299,n20300,n20308);
and (n20300,n20301,n1116);
xor (n20301,n20302,n20307);
or (n20302,n20303,n20306);
and (n20303,n20304,n1207);
xor (n20304,n20305,n2046);
xor (n20305,n20095,n1464);
and (n20306,n20305,n2046);
xor (n20307,n20062,n20096);
and (n20308,n20302,n20307);
xor (n20309,n20247,n1109);
and (n20310,n20298,n20299);
and (n20311,n20271,n20272);
and (n20312,n20266,n20267);
xor (n20313,n20203,n20206);
and (n20314,n20262,n20263);
or (n20315,n20316,n20658);
and (n20316,n20317,n20422);
xor (n20317,n20318,n20319);
xor (n20318,n20261,n20313);
or (n20319,n20320,n20421);
and (n20320,n20321,n20420);
xor (n20321,n20322,n20323);
xor (n20322,n20208,n20241);
or (n20323,n20324,n20419);
and (n20324,n20325,n20418);
xor (n20325,n20326,n20327);
xor (n20326,n20211,n20214);
or (n20327,n20328,n20417);
and (n20328,n20329,n20360);
xor (n20329,n20330,n20359);
or (n20330,n20331,n20358);
and (n20331,n20332,n20334);
xor (n20332,n20333,n1970);
xor (n20333,n20236,n2040);
or (n20334,n20335,n20357);
and (n20335,n20336,n1120);
xor (n20336,n20337,n20344);
or (n20337,n20338,n20343);
and (n20338,n20339,n1215);
xor (n20339,n2052,n20340);
and (n20340,n20341,n2394);
xor (n20341,n20342,n1566);
xor (n20342,n20069,n20071);
and (n20343,n2052,n20340);
or (n20344,n20345,n20356);
and (n20345,n20346,n1214);
xor (n20346,n20347,n20348);
xor (n20347,n20067,n20074);
and (n20348,n20349,n1567);
xor (n20349,n20350,n1222);
and (n20350,n20351,n1027);
xnor (n20351,n20352,n20056);
nand (n20352,n20353,n20355);
or (n20353,n1405,n20354);
not (n20354,n1337);
nand (n20355,n1405,n20354);
and (n20356,n20347,n20348);
and (n20357,n20337,n20344);
and (n20358,n20333,n1970);
xor (n20359,n20216,n1963);
or (n20360,n20361,n20416);
and (n20361,n20362,n20415);
xor (n20362,n20363,n20414);
or (n20363,n20364,n20413);
and (n20364,n20365,n1974);
xor (n20365,n20366,n20367);
xor (n20366,n20223,n20229);
or (n20367,n20368,n20412);
and (n20368,n20369,n20392);
xor (n20369,n20370,n20371);
xor (n20370,n20231,n1471);
or (n20371,n20372,n20391);
and (n20372,n20373,n1478);
xor (n20373,n20374,n20383);
or (n20374,n20375,n20382);
and (n20375,n20376,n20378);
xor (n20376,n2400,n20377);
xor (n20377,n2470,n2063);
and (n20378,n20379,n1027);
nand (n20379,n20380,n20381);
or (n20380,n1353,n20073);
or (n20381,n1410,n20054);
and (n20382,n2400,n20377);
or (n20383,n20384,n20390);
and (n20384,n20385,n20388);
xor (n20385,n20386,n20387);
and (n20386,n1341,n1027);
and (n20387,n2177,n1027);
and (n20388,n20389,n1027);
not (n20389,n2352);
and (n20390,n20386,n20387);
and (n20391,n20374,n20383);
or (n20392,n20393,n20411);
and (n20393,n20394,n2058);
xor (n20394,n20395,n20396);
xor (n20395,n20287,n20289);
or (n20396,n20397,n20410);
and (n20397,n20398,n1228);
xor (n20398,n20399,n20405);
or (n20399,n20400,n20404);
and (n20400,n20401,n20403);
xor (n20401,n20402,n2405);
nor (n20402,n20083,n1026);
nor (n20403,n2338,n1026);
and (n20404,n20402,n2405);
and (n20405,n20406,n20408);
nor (n20406,n20407,n1026);
not (n20407,n1356);
nor (n20408,n20409,n1026);
not (n20409,n2193);
and (n20410,n20399,n20405);
and (n20411,n20395,n20396);
and (n20412,n20370,n20371);
and (n20413,n20366,n20367);
xor (n20414,n20219,n1199);
xor (n20415,n20279,n1967);
and (n20416,n20363,n20414);
and (n20417,n20330,n20359);
xor (n20418,n20243,n20249);
and (n20419,n20326,n20327);
xor (n20420,n20265,n20268);
and (n20421,n20322,n20323);
or (n20422,n20423,n20657);
and (n20423,n20424,n20474);
xor (n20424,n20425,n20426);
xor (n20425,n20321,n20420);
or (n20426,n20427,n20473);
and (n20427,n20428,n20472);
xor (n20428,n20429,n20430);
xor (n20429,n20270,n20295);
or (n20430,n20431,n20471);
and (n20431,n20432,n20470);
xor (n20432,n20433,n20434);
xor (n20433,n20274,n20277);
or (n20434,n20435,n20469);
and (n20435,n20436,n20468);
xor (n20436,n20437,n20443);
or (n20437,n20438,n20442);
and (n20438,n20439,n1977);
xor (n20439,n20440,n1123);
xor (n20440,n20441,n1206);
xor (n20441,n20281,n20282);
and (n20442,n20440,n1123);
or (n20443,n20444,n20467);
and (n20444,n20445,n20462);
xor (n20445,n20446,n20461);
or (n20446,n20447,n20460);
and (n20447,n20448,n1127);
xor (n20448,n20449,n20450);
xor (n20449,n20346,n1214);
or (n20450,n20451,n20459);
and (n20451,n20452,n20458);
xor (n20452,n1223,n20453);
or (n20453,n20454,n20457);
and (n20454,n20455,n1572);
xor (n20455,n20456,n1484);
xor (n20456,n20385,n20388);
and (n20457,n20456,n1484);
xor (n20458,n20341,n2394);
and (n20459,n1223,n20453);
and (n20460,n20449,n20450);
xor (n20461,n20304,n1207);
or (n20462,n20463,n20466);
and (n20463,n20464,n1130);
xor (n20464,n1981,n20465);
xor (n20465,n20284,n2388);
and (n20466,n1981,n20465);
and (n20467,n20446,n20461);
xor (n20468,n20301,n1116);
and (n20469,n20437,n20443);
xor (n20470,n20297,n20309);
and (n20471,n20433,n20434);
xor (n20472,n20325,n20418);
and (n20473,n20429,n20430);
or (n20474,n20475,n20656);
and (n20475,n20476,n20506);
xor (n20476,n20477,n20505);
or (n20477,n20478,n20504);
and (n20478,n20479,n20503);
xor (n20479,n20480,n20502);
or (n20480,n20481,n20501);
and (n20481,n20482,n20500);
xor (n20482,n20483,n20499);
or (n20483,n20484,n20498);
and (n20484,n20485,n20488);
xor (n20485,n20486,n20487);
xor (n20486,n20336,n1120);
xor (n20487,n20365,n1974);
or (n20488,n20489,n20497);
and (n20489,n20490,n1983);
xor (n20490,n20491,n20492);
xor (n20491,n20339,n1215);
or (n20492,n20493,n20496);
and (n20493,n20494,n1134);
xor (n20494,n20495,n1987);
xor (n20495,n20349,n1567);
and (n20496,n20495,n1987);
and (n20497,n20491,n20492);
and (n20498,n20486,n20487);
xor (n20499,n20332,n20334);
xor (n20500,n20362,n20415);
and (n20501,n20483,n20499);
xor (n20502,n20329,n20360);
xor (n20503,n20432,n20470);
and (n20504,n20480,n20502);
xor (n20505,n20428,n20472);
or (n20506,n20507,n20655);
and (n20507,n20508,n20564);
xor (n20508,n20509,n20563);
or (n20509,n20510,n20562);
and (n20510,n20511,n20561);
xor (n20511,n20512,n20560);
or (n20512,n20513,n20559);
and (n20513,n20514,n20552);
xor (n20514,n20515,n20551);
or (n20515,n20516,n20550);
and (n20516,n20517,n20536);
xor (n20517,n20518,n20535);
or (n20518,n20519,n20534);
and (n20519,n20520,n20533);
xor (n20520,n20521,n20532);
or (n20521,n20522,n20531);
and (n20522,n20523,n1140);
xor (n20523,n20524,n20525);
xor (n20524,n20376,n20378);
or (n20525,n20526,n20530);
and (n20526,n20527,n20529);
xor (n20527,n20528,n1998);
and (n20528,n1667,n2564);
xor (n20529,n20406,n20408);
and (n20530,n20528,n1998);
and (n20531,n20524,n20525);
xor (n20532,n20373,n1478);
xor (n20533,n20394,n2058);
and (n20534,n20521,n20532);
xor (n20535,n20369,n20392);
or (n20536,n20537,n20549);
and (n20537,n20538,n1136);
xor (n20538,n20539,n1989);
or (n20539,n20540,n20548);
and (n20540,n20541,n20547);
xor (n20541,n1993,n20542);
or (n20542,n20543,n20546);
and (n20543,n20544,n1489);
xor (n20544,n1145,n20545);
xor (n20545,n20401,n20403);
and (n20546,n1145,n20545);
xor (n20547,n20455,n1572);
and (n20548,n1993,n20542);
and (n20549,n20539,n1989);
and (n20550,n20518,n20535);
xor (n20551,n20439,n1977);
or (n20552,n20553,n20558);
and (n20553,n20554,n20557);
xor (n20554,n20555,n20556);
xor (n20555,n20448,n1127);
xor (n20556,n20464,n1130);
xor (n20557,n20490,n1983);
and (n20558,n20555,n20556);
and (n20559,n20515,n20551);
xor (n20560,n20436,n20468);
xor (n20561,n20482,n20500);
and (n20562,n20512,n20560);
xor (n20563,n20479,n20503);
or (n20564,n20565,n20654);
and (n20565,n20566,n20653);
xor (n20566,n20567,n20606);
or (n20567,n20568,n20605);
and (n20568,n20569,n20604);
xor (n20569,n20570,n20603);
or (n20570,n20571,n20602);
and (n20571,n20572,n20585);
xor (n20572,n20573,n20584);
or (n20573,n20574,n20583);
and (n20574,n20575,n20582);
xor (n20575,n20576,n20581);
or (n20576,n20577,n20580);
and (n20577,n20578,n1142);
xor (n20578,n1995,n20579);
xor (n20579,n20398,n1228);
and (n20580,n1995,n20579);
xor (n20581,n20452,n20458);
xor (n20582,n20494,n1134);
and (n20583,n20576,n20581);
xor (n20584,n20517,n20536);
or (n20585,n20586,n20601);
and (n20586,n20587,n20600);
xor (n20587,n20588,n20589);
xor (n20588,n20520,n20533);
or (n20589,n20590,n20599);
and (n20590,n20591,n20598);
xor (n20591,n20592,n20597);
or (n20592,n20593,n20596);
and (n20593,n20594,n2000);
xor (n20594,n1147,n20595);
xor (n20595,n20527,n20529);
and (n20596,n1147,n20595);
xor (n20597,n20523,n1140);
xor (n20598,n20541,n20547);
and (n20599,n20592,n20597);
xor (n20600,n20538,n1136);
and (n20601,n20588,n20589);
and (n20602,n20573,n20584);
xor (n20603,n20445,n20462);
xor (n20604,n20485,n20488);
and (n20605,n20570,n20603);
nand (n20606,n20607,n20649);
or (n20607,n20608,n20647);
not (n20608,n20609);
nand (n20609,n20610,n20612,n20646);
not (n20610,n20611);
xor (n20611,n20514,n20552);
nand (n20612,n20613,n20645);
or (n20613,n20614,n20615);
xor (n20614,n20572,n20585);
nand (n20615,n20616,n20642);
or (n20616,n20617,n20640);
not (n20617,n20618);
nand (n20618,n20619,n20637);
or (n20619,n20620,n20635);
not (n20620,n20621);
nand (n20621,n20622,n20632);
or (n20622,n20623,n20630);
not (n20623,n20624);
nand (n20624,n20625,n20627);
or (n20625,n20070,n20626);
not (n20626,n1666);
nand (n20627,n20628,n20629);
or (n20628,n1666,n2565);
xor (n20629,n1667,n2564);
not (n20630,n20631);
xor (n20631,n20544,n1489);
nand (n20632,n20633,n20634);
or (n20633,n20631,n20624);
xor (n20634,n20594,n2000);
not (n20635,n20636);
xor (n20636,n20578,n1142);
nand (n20637,n20638,n20639);
or (n20638,n20636,n20621);
xor (n20639,n20591,n20598);
not (n20640,n20641);
xor (n20641,n20575,n20582);
nand (n20642,n20643,n20644);
or (n20643,n20641,n20618);
xor (n20644,n20587,n20600);
xor (n20645,n20554,n20557);
nand (n20646,n20614,n20615);
not (n20647,n20648);
xor (n20648,n20569,n20604);
nand (n20649,n20650,n20611);
or (n20650,n20651,n20652);
not (n20651,n20646);
not (n20652,n20612);
xor (n20653,n20511,n20561);
and (n20654,n20567,n20606);
and (n20655,n20509,n20563);
and (n20656,n20477,n20505);
and (n20657,n20425,n20426);
and (n20658,n20318,n20319);
and (n20659,n20258,n20259);
and (n20660,n19868,n20197);
nor (n20661,n20662,n20685);
not (n20662,n20663);
nor (n20663,n20664,n20682);
not (n20664,n20665);
nor (n20665,n20666,n20679);
not (n20666,n20667);
nor (n20667,n20668,n20676);
not (n20668,n20669);
nor (n20669,n20670,n20671);
and (n20670,n20158,n1080);
not (n20671,n20672);
nor (n20672,n20673,n20674);
and (n20673,n1422,n1077);
not (n20674,n20675);
xnor (n20675,n15,n1242);
or (n20676,n20677,n20678);
and (n20677,n20152,n20157);
and (n20678,n20153,n20156);
or (n20679,n20680,n20681);
and (n20680,n20122,n20139);
and (n20681,n20123,n20126);
or (n20682,n20683,n20684);
and (n20683,n20147,n20159);
and (n20684,n20148,n20151);
or (n20685,n20686,n20687);
and (n20686,n19869,n20146);
and (n20687,n19870,n20121);
nor (n20688,n19848,n2705);
nor (n20689,n20690,n21494);
and (n20690,n20691,n19825);
nand (n20691,n20692,n20693);
not (n20692,n9932);
nor (n20693,n9900,n20694);
and (n20694,n20695,n20688);
nand (n20695,n20696,n21469);
not (n20696,n20697);
or (n20697,n20698,n21468);
and (n20698,n20699,n21076);
xor (n20699,n20700,n21019);
xor (n20700,n20701,n20968);
xor (n20701,n20702,n20943);
or (n20702,n20703,n20942);
and (n20703,n20704,n20819);
xor (n20704,n20705,n20794);
xor (n20705,n20706,n20747);
xor (n20706,n20707,n20709);
xor (n20707,n20708,n8766);
xor (n20708,n8715,n9329);
xor (n20709,n20710,n9543);
xor (n20710,n20711,n20745);
or (n20711,n20712,n20744);
and (n20712,n20713,n9624);
xor (n20713,n20714,n8913);
and (n20714,n20715,n8921);
xor (n20715,n8920,n20716);
xor (n20716,n20717,n20725);
xor (n20717,n20718,n20722);
xor (n20718,n20719,n19891);
xor (n20719,n20720,n19888);
nor (n20720,n20721,n1026);
not (n20721,n9399);
and (n20722,n20720,n20723);
not (n20723,n20724);
not (n20724,n9411);
or (n20725,n20726,n20743);
and (n20726,n20727,n20735);
xor (n20727,n19895,n20728);
and (n20728,n20729,n1027);
nand (n20729,n20730,n20734);
or (n20730,n20731,n20732);
not (n20731,n9408);
not (n20732,n20733);
not (n20733,n9498);
or (n20734,n20733,n9408);
and (n20735,n20736,n1027);
or (n20736,n20737,n20741);
nor (n20737,n20738,n20724);
and (n20738,n20739,n20740);
not (n20739,n9503);
not (n20740,n9419);
nor (n20741,n20742,n20721);
not (n20742,n9443);
and (n20743,n19895,n20728);
and (n20744,n20714,n8913);
xor (n20745,n20746,n8906);
xor (n20746,n8855,n8905);
or (n20747,n20748,n20793);
and (n20748,n20749,n20755);
xor (n20749,n20750,n20754);
or (n20750,n20751,n20753);
and (n20751,n20752,n8781);
xor (n20752,n9340,n9269);
and (n20753,n9340,n9269);
xor (n20754,n20713,n9624);
and (n20755,n20756,n8722);
xor (n20756,n8780,n20757);
or (n20757,n20758,n20792);
and (n20758,n20759,n20779);
xor (n20759,n9636,n20760);
and (n20760,n20761,n20773);
or (n20761,n20762,n20772);
and (n20762,n20763,n20059);
xor (n20763,n20764,n19924);
and (n20764,n20765,n1027);
nand (n20765,n20766,n20768,n20771);
or (n20766,n20767,n20739);
not (n20767,n9467);
or (n20768,n20769,n20770);
not (n20769,n9509);
not (n20770,n9447);
not (n20771,n9434);
and (n20772,n20764,n19924);
and (n20773,n20774,n1027);
nor (n20774,n20775,n20777);
and (n20775,n20776,n20723);
xor (n20776,n20739,n20740);
and (n20777,n20778,n20724);
not (n20778,n20776);
or (n20779,n20780,n20791);
and (n20780,n20781,n9642);
xor (n20781,n8937,n20782);
xor (n20782,n20783,n19942);
xor (n20783,n19954,n20784);
and (n20784,n20785,n1027);
nand (n20785,n20786,n20790);
or (n20786,n20787,n20769);
and (n20787,n20788,n20789);
not (n20788,n9423);
not (n20789,n9431);
not (n20790,n9422);
and (n20791,n8937,n20782);
and (n20792,n9636,n20760);
and (n20793,n20750,n20754);
xor (n20794,n20795,n20815);
xor (n20795,n20796,n20805);
xor (n20796,n20797,n9619);
xor (n20797,n8765,n20798);
and (n20798,n20799,n20802);
or (n20799,n20800,n20801);
and (n20800,n20717,n20725);
and (n20801,n20718,n20722);
or (n20802,n20803,n20804);
and (n20803,n20719,n19891);
and (n20804,n20720,n19888);
or (n20805,n20806,n20814);
and (n20806,n20807,n8773);
xor (n20807,n20808,n9334);
or (n20808,n20809,n20813);
and (n20809,n20810,n9553);
xor (n20810,n20811,n20812);
xor (n20811,n20715,n8921);
and (n20812,n8927,n8866);
and (n20813,n20811,n20812);
and (n20814,n20808,n9334);
or (n20815,n20816,n20818);
and (n20816,n20817,n8718);
xor (n20817,n1891,n9265);
and (n20818,n1891,n9265);
or (n20819,n20820,n20941);
and (n20820,n20821,n20846);
xor (n20821,n20822,n20823);
xor (n20822,n20749,n20755);
or (n20823,n20824,n20845);
and (n20824,n20825,n20832);
xor (n20825,n20826,n20831);
or (n20826,n20827,n20830);
and (n20827,n20828,n9277);
xor (n20828,n8789,n20829);
xor (n20829,n20759,n20779);
and (n20830,n8789,n20829);
xor (n20831,n20756,n8722);
or (n20832,n20833,n20844);
and (n20833,n20834,n8726);
xor (n20834,n9275,n20835);
or (n20835,n20836,n20843);
and (n20836,n20837,n8796);
xor (n20837,n20838,n20840);
xor (n20838,n20839,n8936);
xor (n20839,n20761,n20773);
and (n20840,n20841,n9648);
xor (n20841,n20842,n8944);
xor (n20842,n20763,n20059);
and (n20843,n20838,n20840);
and (n20844,n9275,n20835);
and (n20845,n20826,n20831);
or (n20846,n20847,n20940);
and (n20847,n20848,n20928);
xor (n20848,n20849,n20927);
or (n20849,n20850,n20926);
and (n20850,n20851,n1956);
xor (n20851,n20852,n20903);
or (n20852,n20853,n20902);
and (n20853,n20854,n8797);
xor (n20854,n20855,n20874);
xor (n20855,n20856,n9567);
xor (n20856,n8870,n20857);
or (n20857,n20858,n20873);
and (n20858,n20859,n8945);
xor (n20859,n20860,n20871);
or (n20860,n20058,n20861);
and (n20861,n20862,n1027);
nand (n20862,n20863,n20864);
not (n20863,n9446);
nand (n20864,n20865,n20869);
or (n20865,n20866,n20867);
not (n20866,n20770);
not (n20867,n20868);
not (n20868,n9455);
not (n20869,n20870);
not (n20870,n9521);
nor (n20871,n1026,n20872);
xor (n20872,n9511,n20769);
and (n20873,n20860,n20871);
and (n20874,n20875,n20901);
xor (n20875,n20876,n20899);
or (n20876,n20877,n20898);
and (n20877,n20878,n9654);
xor (n20878,n20879,n20885);
and (n20879,n20880,n20883);
xor (n20880,n20881,n8960);
and (n20881,n20882,n1027);
xnor (n20882,n20870,n9523);
and (n20883,n20884,n20069);
and (n20884,n9766,n20869);
or (n20885,n20886,n20897);
and (n20886,n20887,n20074);
xor (n20887,n20888,n20085);
and (n20888,n20889,n1027);
not (n20889,n20890);
nor (n20890,n20891,n20892);
and (n20891,n20869,n9471);
and (n20892,n20893,n20896);
nand (n20893,n20894,n20895);
not (n20894,n9527);
not (n20895,n9459);
not (n20896,n20767);
and (n20897,n20888,n20085);
and (n20898,n20879,n20885);
and (n20899,n20900,n8878);
xor (n20900,n9581,n8952);
xor (n20901,n20841,n9648);
and (n20902,n20855,n20874);
or (n20903,n20904,n20925);
and (n20904,n20905,n9352);
xor (n20905,n20906,n20907);
xor (n20906,n20781,n9642);
or (n20907,n20908,n20924);
and (n20908,n20909,n9574);
xor (n20909,n8874,n20910);
or (n20910,n20911,n20923);
and (n20911,n20912,n8953);
xor (n20912,n20913,n20034);
and (n20913,n20914,n1027);
not (n20914,n20915);
nor (n20915,n20916,n20922);
and (n20916,n20917,n20920);
not (n20917,n20918);
xor (n20918,n20742,n20919);
not (n20919,n9515);
not (n20920,n20921);
not (n20921,n9435);
and (n20922,n20918,n20921);
and (n20923,n20913,n20034);
and (n20924,n8874,n20910);
and (n20925,n20906,n20907);
and (n20926,n20852,n20903);
xor (n20927,n20752,n8781);
xor (n20928,n20929,n1948);
xor (n20929,n9271,n20930);
xor (n20930,n20931,n9630);
xor (n20931,n8862,n20932);
or (n20932,n20933,n20939);
and (n20933,n20934,n20936);
xor (n20934,n20935,n19902);
xor (n20935,n20727,n20735);
or (n20936,n20937,n20938);
and (n20937,n20783,n19942);
and (n20938,n19954,n20784);
and (n20939,n20935,n19902);
and (n20940,n20849,n20927);
and (n20941,n20822,n20823);
and (n20942,n20705,n20794);
xor (n20943,n20944,n20965);
xor (n20944,n20945,n20952);
xor (n20945,n20946,n20949);
xor (n20946,n20947,n20948);
and (n20947,n20797,n9619);
and (n20948,n20746,n8906);
or (n20949,n20950,n20951);
and (n20950,n20708,n8766);
and (n20951,n8715,n9329);
and (n20952,n20953,n20960);
xor (n20953,n20954,n9260);
or (n20954,n20955,n20959);
and (n20955,n20956,n9263);
xor (n20956,n8858,n20957);
xor (n20957,n20958,n8912);
xor (n20958,n20799,n20802);
and (n20959,n8858,n20957);
and (n20960,n20961,n9546);
xor (n20961,n8772,n20962);
or (n20962,n20963,n20964);
and (n20963,n20931,n9630);
and (n20964,n8862,n20932);
or (n20965,n20966,n20967);
and (n20966,n20795,n20815);
and (n20967,n20796,n20805);
xor (n20968,n20969,n20981);
xor (n20969,n20970,n20973);
or (n20970,n20971,n20972);
and (n20971,n20706,n20747);
and (n20972,n20707,n20709);
xor (n20973,n20974,n20979);
xor (n20974,n20975,n20978);
or (n20975,n20976,n20977);
and (n20976,n20710,n9543);
and (n20977,n20711,n20745);
xor (n20978,n8851,n8712);
xor (n20979,n20980,n8713);
xor (n20980,n9083,n9396);
or (n20981,n20982,n21018);
and (n20982,n20983,n20994);
xor (n20983,n20984,n20993);
or (n20984,n20985,n20992);
and (n20985,n20986,n20991);
xor (n20986,n20987,n20990);
or (n20987,n20988,n20989);
and (n20988,n20929,n1948);
and (n20989,n9271,n20930);
xor (n20990,n20956,n9263);
xor (n20991,n20807,n8773);
and (n20992,n20987,n20990);
xor (n20993,n20953,n20960);
or (n20994,n20995,n21017);
and (n20995,n20996,n21016);
xor (n20996,n20997,n20998);
xor (n20997,n20961,n9546);
or (n20998,n20999,n21015);
and (n20999,n21000,n21010);
xor (n21000,n21001,n21002);
xor (n21001,n20810,n9553);
or (n21002,n21003,n21009);
and (n21003,n21004,n9560);
xor (n21004,n21005,n21008);
or (n21005,n21006,n21007);
and (n21006,n20856,n9567);
and (n21007,n8870,n20857);
xor (n21008,n20934,n20936);
and (n21009,n21005,n21008);
or (n21010,n21011,n21014);
and (n21011,n21012,n9346);
xor (n21012,n8788,n21013);
xor (n21013,n8927,n8866);
and (n21014,n8788,n21013);
and (n21015,n21001,n21002);
xor (n21016,n20817,n8718);
and (n21017,n20997,n20998);
and (n21018,n20984,n20993);
or (n21019,n21020,n21075);
and (n21020,n21021,n21074);
xor (n21021,n21022,n21073);
or (n21022,n21023,n21072);
and (n21023,n21024,n21027);
xor (n21024,n21025,n21026);
xor (n21025,n20996,n21016);
xor (n21026,n20986,n20991);
or (n21027,n21028,n21071);
and (n21028,n21029,n21061);
xor (n21029,n21030,n21060);
or (n21030,n21031,n21059);
and (n21031,n21032,n21035);
xor (n21032,n21033,n21034);
xor (n21033,n21012,n9346);
xor (n21034,n21004,n9560);
or (n21035,n21036,n21058);
and (n21036,n21037,n9283);
xor (n21037,n21038,n21041);
and (n21038,n21039,n9358);
xor (n21039,n8804,n21040);
xor (n21040,n20859,n8945);
or (n21041,n21042,n21057);
and (n21042,n21043,n8805);
xor (n21043,n21044,n21045);
xor (n21044,n20909,n9574);
or (n21045,n21046,n21056);
and (n21046,n21047,n21052);
xor (n21047,n21048,n21049);
xor (n21048,n20912,n8953);
nand (n21049,n21050,n20860);
or (n21050,n21051,n20227);
not (n21051,n20861);
or (n21052,n21053,n21055);
and (n21053,n21054,n8882);
xor (n21054,n8961,n9660);
and (n21055,n8961,n9660);
and (n21056,n21048,n21049);
and (n21057,n21044,n21045);
and (n21058,n21038,n21041);
and (n21059,n21033,n21034);
xor (n21060,n21000,n21010);
or (n21061,n21062,n21070);
and (n21062,n21063,n21069);
xor (n21063,n21064,n21065);
xor (n21064,n20828,n9277);
or (n21065,n21066,n21068);
and (n21066,n21067,n1963);
xor (n21067,n8730,n9281);
and (n21068,n8730,n9281);
xor (n21069,n20834,n8726);
and (n21070,n21064,n21065);
and (n21071,n21030,n21060);
and (n21072,n21025,n21026);
xor (n21073,n20983,n20994);
xor (n21074,n20704,n20819);
and (n21075,n21022,n21073);
or (n21076,n21077,n21467);
and (n21077,n21078,n21148);
xor (n21078,n21079,n21080);
xor (n21079,n21021,n21074);
or (n21080,n21081,n21147);
and (n21081,n21082,n21146);
xor (n21082,n21083,n21145);
or (n21083,n21084,n21144);
and (n21084,n21085,n21143);
xor (n21085,n21086,n21087);
xor (n21086,n20825,n20832);
or (n21087,n21088,n21142);
and (n21088,n21089,n21119);
xor (n21089,n21090,n21091);
xor (n21090,n20851,n1956);
or (n21091,n21092,n21118);
and (n21092,n21093,n21096);
xor (n21093,n21094,n21095);
xor (n21094,n20837,n8796);
xor (n21095,n20905,n9352);
or (n21096,n21097,n21117);
and (n21097,n21098,n9287);
xor (n21098,n21099,n8734);
and (n21099,n21100,n21116);
and (n21100,n21101,n21106);
or (n21101,n21102,n21105);
and (n21102,n21103,n9595);
xor (n21103,n8969,n21104);
xor (n21104,n20884,n20069);
and (n21105,n8969,n21104);
and (n21106,n21107,n20289);
xor (n21107,n21108,n8828);
and (n21108,n21109,n1027);
nand (n21109,n21110,n21115);
or (n21110,n20895,n21111);
nand (n21111,n21112,n21114);
or (n21112,n21113,n20767);
not (n21113,n20894);
nand (n21114,n21113,n20767);
nand (n21115,n21111,n20895);
xor (n21116,n20878,n9654);
and (n21117,n21099,n8734);
and (n21118,n21094,n21095);
or (n21119,n21120,n21141);
and (n21120,n21121,n21140);
xor (n21121,n21122,n21139);
or (n21122,n21123,n21138);
and (n21123,n21124,n1970);
xor (n21124,n21125,n21137);
or (n21125,n21126,n21136);
and (n21126,n21127,n8813);
xor (n21127,n21128,n21129);
xor (n21128,n20900,n8878);
or (n21129,n21130,n21135);
and (n21130,n21131,n9588);
xor (n21131,n21132,n21133);
xor (n21132,n20887,n20074);
and (n21133,n9666,n21134);
and (n21134,n9671,n9381);
and (n21135,n21132,n21133);
and (n21136,n21128,n21129);
xor (n21137,n20875,n20901);
and (n21138,n21125,n21137);
xor (n21139,n20854,n8797);
xor (n21140,n21067,n1963);
and (n21141,n21122,n21139);
and (n21142,n21090,n21091);
xor (n21143,n20848,n20928);
and (n21144,n21086,n21087);
xor (n21145,n20821,n20846);
xor (n21146,n21024,n21027);
and (n21147,n21083,n21145);
or (n21148,n21149,n21466);
and (n21149,n21150,n21235);
xor (n21150,n21151,n21152);
xor (n21151,n21082,n21146);
or (n21152,n21153,n21234);
and (n21153,n21154,n21233);
xor (n21154,n21155,n21156);
xor (n21155,n21029,n21061);
or (n21156,n21157,n21232);
and (n21157,n21158,n21231);
xor (n21158,n21159,n21160);
xor (n21159,n21032,n21035);
or (n21160,n21161,n21230);
and (n21161,n21162,n21178);
xor (n21162,n21163,n21177);
or (n21163,n21164,n21176);
and (n21164,n21165,n21167);
xor (n21165,n9289,n21166);
xor (n21166,n21039,n9358);
or (n21167,n21168,n21175);
and (n21168,n21169,n8738);
xor (n21169,n21170,n9364);
or (n21170,n21171,n21174);
and (n21171,n21172,n8821);
xor (n21172,n9370,n21173);
xor (n21173,n20880,n20883);
and (n21174,n9370,n21173);
and (n21175,n21170,n9364);
and (n21176,n9289,n21166);
xor (n21177,n21037,n9283);
or (n21178,n21179,n21229);
and (n21179,n21180,n21228);
xor (n21180,n21181,n21182);
xor (n21181,n21043,n8805);
or (n21182,n21183,n21227);
and (n21183,n21184,n9295);
xor (n21184,n9293,n21185);
or (n21185,n21186,n21226);
and (n21186,n21187,n21207);
xor (n21187,n21188,n21189);
xor (n21188,n21054,n8882);
or (n21189,n21190,n21206);
and (n21190,n21191,n8886);
xor (n21191,n21192,n21197);
or (n21192,n21193,n21196);
and (n21193,n21194,n20388);
xor (n21194,n21195,n9601);
xor (n21195,n9671,n9381);
and (n21196,n21195,n9601);
or (n21197,n21198,n21205);
and (n21198,n21199,n21201);
xor (n21199,n20387,n21200);
and (n21200,n9471,n1027);
and (n21201,n21202,n1027);
xor (n21202,n21203,n21204);
not (n21203,n9479);
not (n21204,n9532);
and (n21205,n20387,n21200);
and (n21206,n21192,n21197);
or (n21207,n21208,n21225);
and (n21208,n21209,n9376);
xor (n21209,n21210,n21223);
or (n21210,n21211,n21222);
and (n21211,n21212,n8834);
xor (n21212,n21213,n21219);
or (n21213,n21214,n21218);
and (n21214,n21215,n21216);
xor (n21215,n20403,n9606);
nor (n21216,n21217,n1026);
not (n21217,n9490);
and (n21218,n20403,n9606);
and (n21219,n20408,n21220);
nor (n21220,n21221,n1026);
not (n21221,n9482);
and (n21222,n21213,n21219);
xor (n21223,n21224,n8968);
xor (n21224,n9666,n21134);
and (n21225,n21210,n21223);
and (n21226,n21188,n21189);
and (n21227,n9293,n21185);
xor (n21228,n21098,n9287);
and (n21229,n21181,n21182);
and (n21230,n21163,n21177);
xor (n21231,n21063,n21069);
and (n21232,n21159,n21160);
xor (n21233,n21085,n21143);
and (n21234,n21155,n21156);
or (n21235,n21236,n21465);
and (n21236,n21237,n21289);
xor (n21237,n21238,n21288);
or (n21238,n21239,n21287);
and (n21239,n21240,n21286);
xor (n21240,n21241,n21285);
or (n21241,n21242,n21284);
and (n21242,n21243,n21283);
xor (n21243,n21244,n21282);
or (n21244,n21245,n21281);
and (n21245,n21246,n21280);
xor (n21246,n21247,n21274);
or (n21247,n21248,n21273);
and (n21248,n21249,n21268);
xor (n21249,n21250,n21252);
xor (n21250,n21251,n8812);
xor (n21251,n21100,n21116);
or (n21252,n21253,n21267);
and (n21253,n21254,n8742);
xor (n21254,n21255,n21265);
or (n21255,n21256,n21264);
and (n21256,n21257,n21263);
xor (n21257,n8829,n21258);
or (n21258,n21259,n21262);
and (n21259,n21260,n8974);
xor (n21260,n21261,n8890);
xor (n21261,n21199,n21201);
and (n21262,n21261,n8890);
xor (n21263,n21103,n9595);
and (n21264,n8829,n21258);
xor (n21265,n21266,n8820);
xor (n21266,n21101,n21106);
and (n21267,n21255,n21265);
or (n21268,n21269,n21272);
and (n21269,n21270,n1983);
xor (n21270,n9299,n21271);
xor (n21271,n21131,n9588);
and (n21272,n9299,n21271);
and (n21273,n21250,n21252);
or (n21274,n21275,n21279);
and (n21275,n21276,n1977);
xor (n21276,n21277,n21278);
xor (n21277,n21047,n21052);
xor (n21278,n21127,n8813);
and (n21279,n21277,n21278);
xor (n21280,n21124,n1970);
and (n21281,n21247,n21274);
xor (n21282,n21093,n21096);
xor (n21283,n21121,n21140);
and (n21284,n21244,n21282);
xor (n21285,n21089,n21119);
xor (n21286,n21158,n21231);
and (n21287,n21241,n21285);
xor (n21288,n21154,n21233);
or (n21289,n21290,n21464);
and (n21290,n21291,n21356);
xor (n21291,n21292,n21355);
or (n21292,n21293,n21354);
and (n21293,n21294,n21353);
xor (n21294,n21295,n21296);
xor (n21295,n21162,n21178);
or (n21296,n21297,n21352);
and (n21297,n21298,n21351);
xor (n21298,n21299,n21300);
xor (n21299,n21165,n21167);
or (n21300,n21301,n21350);
and (n21301,n21302,n21314);
xor (n21302,n21303,n21304);
xor (n21303,n21169,n8738);
or (n21304,n21305,n21313);
and (n21305,n21306,n9301);
xor (n21306,n21307,n21308);
xor (n21307,n21172,n8821);
or (n21308,n21309,n21312);
and (n21309,n21310,n8746);
xor (n21310,n9305,n21311);
xor (n21311,n21107,n20289);
and (n21312,n9305,n21311);
and (n21313,n21307,n21308);
or (n21314,n21315,n21349);
and (n21315,n21316,n21334);
xor (n21316,n21317,n21318);
xor (n21317,n21187,n21207);
or (n21318,n21319,n21333);
and (n21319,n21320,n9307);
xor (n21320,n21321,n21332);
or (n21321,n21322,n21331);
and (n21322,n21323,n8750);
xor (n21323,n21324,n21325);
xor (n21324,n21194,n20388);
or (n21325,n21326,n21330);
and (n21326,n21327,n21329);
xor (n21327,n21328,n9316);
and (n21328,n2565,n9765);
xor (n21329,n20408,n21220);
and (n21330,n21328,n9316);
and (n21331,n21324,n21325);
xor (n21332,n21191,n8886);
and (n21333,n21321,n21332);
or (n21334,n21335,n21348);
and (n21335,n21336,n1989);
xor (n21336,n21337,n21338);
xor (n21337,n21209,n9376);
or (n21338,n21339,n21347);
and (n21339,n21340,n9311);
xor (n21340,n21341,n21342);
xor (n21341,n21260,n8974);
or (n21342,n21343,n21346);
and (n21343,n21344,n8893);
xor (n21344,n8753,n21345);
xor (n21345,n21215,n21216);
and (n21346,n8753,n21345);
and (n21347,n21341,n21342);
and (n21348,n21337,n21338);
and (n21349,n21317,n21318);
and (n21350,n21303,n21304);
xor (n21351,n21180,n21228);
and (n21352,n21299,n21300);
xor (n21353,n21243,n21283);
and (n21354,n21295,n21296);
xor (n21355,n21240,n21286);
nand (n21356,n21357,n21463);
or (n21357,n21358,n21373);
nor (n21358,n21359,n21360);
xor (n21359,n21294,n21353);
or (n21360,n21361,n21372);
and (n21361,n21362,n21371);
xor (n21362,n21363,n21364);
xor (n21363,n21246,n21280);
or (n21364,n21365,n21370);
and (n21365,n21366,n21369);
xor (n21366,n21367,n21368);
xor (n21367,n21184,n9295);
xor (n21368,n21276,n1977);
xor (n21369,n21249,n21268);
and (n21370,n21367,n21368);
xor (n21371,n21298,n21351);
and (n21372,n21363,n21364);
and (n21373,n21374,n21462);
nand (n21374,n21375,n21390);
or (n21375,n21376,n21377);
xor (n21376,n21362,n21371);
or (n21377,n21378,n21389);
and (n21378,n21379,n21388);
xor (n21379,n21380,n21387);
or (n21380,n21381,n21386);
and (n21381,n21382,n21385);
xor (n21382,n21383,n21384);
xor (n21383,n21270,n1983);
xor (n21384,n21254,n8742);
xor (n21385,n21306,n9301);
and (n21386,n21383,n21384);
xor (n21387,n21302,n21314);
xor (n21388,n21366,n21369);
and (n21389,n21380,n21387);
nand (n21390,n21391,n21455);
nand (n21391,n21392,n21427,n21430);
or (n21392,n21393,n21426);
or (n21393,n21394,n21425);
and (n21394,n21395,n21424);
xor (n21395,n21396,n21413);
or (n21396,n21397,n21412);
and (n21397,n21398,n21411);
xor (n21398,n21399,n21400);
xor (n21399,n21320,n9307);
or (n21400,n21401,n21410);
and (n21401,n21402,n21409);
xor (n21402,n21403,n21404);
xor (n21403,n21323,n8750);
or (n21404,n21405,n21408);
and (n21405,n21406,n9318);
xor (n21406,n21407,n2000);
xor (n21407,n21327,n21329);
and (n21408,n21407,n2000);
xor (n21409,n21340,n9311);
and (n21410,n21403,n21404);
xor (n21411,n21336,n1989);
and (n21412,n21399,n21400);
or (n21413,n21414,n21423);
and (n21414,n21415,n21422);
xor (n21415,n21416,n21421);
or (n21416,n21417,n21420);
and (n21417,n21418,n1995);
xor (n21418,n9313,n21419);
xor (n21419,n21212,n8834);
and (n21420,n9313,n21419);
xor (n21421,n21257,n21263);
xor (n21422,n21310,n8746);
and (n21423,n21416,n21421);
xor (n21424,n21316,n21334);
and (n21425,n21396,n21413);
xor (n21426,n21379,n21388);
or (n21427,n21428,n21429);
xor (n21428,n21395,n21424);
xor (n21429,n21382,n21385);
nand (n21430,n21431,n21451);
or (n21431,n21432,n21435);
nor (n21432,n21433,n21434);
xor (n21433,n21398,n21411);
xor (n21434,n21415,n21422);
nand (n21435,n21436,n21439,n21442);
or (n21436,n21437,n21438);
xor (n21437,n21418,n1995);
xor (n21438,n21402,n21409);
or (n21439,n21440,n21441);
xor (n21440,n21344,n8893);
xor (n21441,n21406,n9318);
nand (n21442,n21443,n21446);
or (n21443,n21444,n21445);
not (n21444,n21440);
not (n21445,n21441);
nor (n21446,n21447,n21450);
and (n21447,n21448,n21449);
xor (n21448,n2565,n9765);
or (n21449,n2564,n9766);
and (n21450,n2564,n9766);
nor (n21451,n21452,n21454);
and (n21452,n21453,n21437,n21438);
not (n21453,n21432);
and (n21454,n21433,n21434);
nor (n21455,n21456,n21460);
and (n21456,n21426,n21457);
nand (n21457,n21458,n21459);
not (n21458,n21393);
nand (n21459,n21428,n21429);
and (n21460,n21461,n21393);
not (n21461,n21459);
nand (n21462,n21376,n21377);
nand (n21463,n21359,n21360);
and (n21464,n21292,n21355);
and (n21465,n21238,n21288);
and (n21466,n21151,n21152);
and (n21467,n21079,n21080);
and (n21468,n20700,n21019);
not (n21469,n21470);
or (n21470,n21471,n21474);
or (n21471,n21472,n21473);
and (n21472,n20701,n20968);
and (n21473,n20702,n20943);
nand (n21474,n21475,n21479);
not (n21475,n21476);
or (n21476,n21477,n21478);
and (n21477,n20969,n20981);
and (n21478,n20970,n20973);
nor (n21479,n21480,n21493);
not (n21480,n21481);
nor (n21481,n21482,n21490);
not (n21482,n21483);
nor (n21483,n21484,n21485);
and (n21484,n20980,n8713);
not (n21485,n21486);
nor (n21486,n21487,n21488);
and (n21487,n8851,n8712);
not (n21488,n21489);
xnor (n21489,n8708,n8848);
or (n21490,n21491,n21492);
and (n21491,n20974,n20979);
and (n21492,n20975,n20978);
and (n21493,n20944,n20965);
nor (n21494,n21495,n21499);
and (n21495,n21496,n21498);
not (n21496,n21497);
and (n21497,n17725,n19835);
not (n21498,n13872);
nand (n21499,n21500,n14125);
or (n21500,n21497,n19836);
endmodule
