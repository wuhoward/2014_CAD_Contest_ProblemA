module top (out,n3,n4,n5,n26,n28,n35,n36,n45,n52
        ,n54,n60,n66,n72,n80,n82,n92,n98,n111,n119
        ,n125,n136,n140,n145,n152,n160,n164,n168,n173,n183
        ,n189,n194,n202,n212);
output out;
input n3;
input n4;
input n5;
input n26;
input n28;
input n35;
input n36;
input n45;
input n52;
input n54;
input n60;
input n66;
input n72;
input n80;
input n82;
input n92;
input n98;
input n111;
input n119;
input n125;
input n136;
input n140;
input n145;
input n152;
input n160;
input n164;
input n168;
input n173;
input n183;
input n189;
input n194;
input n202;
input n212;
wire n0;
wire n1;
wire n2;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n24;
wire n25;
wire n27;
wire n29;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n53;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n81;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n137;
wire n138;
wire n139;
wire n141;
wire n142;
wire n143;
wire n144;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n161;
wire n162;
wire n163;
wire n165;
wire n166;
wire n167;
wire n169;
wire n170;
wire n171;
wire n172;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n190;
wire n191;
wire n192;
wire n193;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
xnor (out,n0,n811);
nor (n0,n1,n6);
and (n1,n2,n5);
nor (n2,n3,n4);
and (n6,n7,n808);
nand (n7,n8,n807);
or (n8,n9,n397);
not (n9,n10);
nand (n10,n11,n396);
nand (n11,n12,n363);
not (n12,n13);
xor (n13,n14,n310);
xor (n14,n15,n214);
xor (n15,n16,n177);
xor (n16,n17,n102);
or (n17,n18,n101);
and (n18,n19,n74);
xor (n19,n20,n47);
nand (n20,n21,n41);
or (n21,n22,n30);
not (n22,n23);
nor (n23,n24,n29);
and (n24,n25,n27);
not (n25,n26);
not (n27,n28);
and (n29,n26,n28);
nand (n30,n31,n38);
not (n31,n32);
nand (n32,n33,n37);
or (n33,n34,n36);
not (n34,n35);
nand (n37,n34,n36);
nand (n38,n39,n40);
or (n39,n28,n34);
nand (n40,n34,n28);
nand (n41,n42,n32);
nand (n42,n43,n46);
or (n43,n28,n44);
not (n44,n45);
or (n46,n27,n45);
nand (n47,n48,n68);
or (n48,n49,n57);
not (n49,n50);
nand (n50,n51,n55);
or (n51,n52,n53);
not (n53,n54);
or (n55,n56,n54);
not (n56,n52);
nand (n57,n58,n62);
nand (n58,n59,n61);
or (n59,n60,n56);
nand (n61,n56,n60);
not (n62,n63);
nand (n63,n64,n67);
or (n64,n65,n60);
not (n65,n66);
nand (n67,n60,n65);
nand (n68,n63,n69);
nand (n69,n70,n73);
or (n70,n52,n71);
not (n71,n72);
or (n73,n56,n72);
nand (n74,n75,n94);
or (n75,n76,n88);
not (n76,n77);
nor (n77,n78,n85);
nor (n78,n79,n83);
and (n79,n80,n81);
not (n81,n82);
and (n83,n82,n84);
not (n84,n80);
nand (n85,n86,n87);
or (n86,n56,n80);
nand (n87,n80,n56);
not (n88,n89);
nand (n89,n90,n93);
or (n90,n82,n91);
not (n91,n92);
or (n93,n81,n92);
or (n94,n95,n96);
not (n95,n85);
nor (n96,n97,n99);
and (n97,n81,n98);
and (n99,n82,n100);
not (n100,n98);
and (n101,n20,n47);
or (n102,n103,n176);
and (n103,n104,n154);
xor (n104,n105,n129);
nand (n105,n106,n122);
or (n106,n107,n117);
not (n107,n108);
nor (n108,n109,n113);
nand (n109,n110,n112);
or (n110,n27,n111);
nand (n112,n111,n27);
nor (n113,n114,n116);
and (n114,n115,n66);
not (n115,n111);
and (n116,n111,n65);
nor (n117,n118,n120);
and (n118,n65,n119);
and (n120,n66,n121);
not (n121,n119);
or (n122,n123,n128);
nor (n123,n124,n126);
and (n124,n65,n125);
and (n126,n66,n127);
not (n127,n125);
not (n128,n109);
nand (n129,n130,n148);
or (n130,n131,n143);
nand (n131,n132,n138);
not (n132,n133);
nand (n133,n134,n137);
or (n134,n135,n82);
not (n135,n136);
nand (n137,n82,n135);
nand (n138,n139,n141);
nand (n139,n135,n140);
nand (n141,n136,n142);
not (n142,n140);
nor (n143,n144,n146);
and (n144,n142,n145);
and (n146,n140,n147);
not (n147,n145);
or (n148,n149,n132);
nor (n149,n150,n153);
and (n150,n151,n140);
not (n151,n152);
and (n153,n152,n142);
nand (n154,n155,n170);
or (n155,n156,n165);
nand (n156,n157,n162);
nor (n157,n158,n161);
and (n158,n159,n140);
not (n159,n160);
and (n161,n160,n142);
xor (n162,n159,n163);
not (n163,n164);
nor (n165,n166,n169);
and (n166,n167,n164);
not (n167,n168);
and (n169,n168,n163);
or (n170,n171,n157);
nor (n171,n172,n174);
and (n172,n163,n173);
and (n174,n164,n175);
not (n175,n173);
and (n176,n105,n129);
xor (n177,n178,n204);
xor (n178,n179,n185);
nor (n179,n180,n167);
not (n180,n181);
nand (n181,n182,n184);
or (n182,n163,n183);
nand (n184,n163,n183);
nand (n185,n186,n197);
or (n186,n187,n190);
nand (n187,n188,n36);
not (n188,n189);
not (n190,n191);
nor (n191,n192,n196);
and (n192,n193,n195);
not (n193,n194);
not (n195,n36);
and (n196,n194,n36);
nand (n197,n198,n189);
not (n198,n199);
nor (n199,n200,n203);
and (n200,n201,n36);
not (n201,n202);
and (n203,n202,n195);
nand (n204,n205,n207);
or (n205,n30,n206);
not (n206,n42);
or (n207,n31,n208);
not (n208,n209);
nand (n209,n210,n213);
or (n210,n28,n211);
not (n211,n212);
or (n213,n27,n212);
xor (n214,n215,n264);
xor (n215,n216,n237);
xor (n216,n217,n231);
xor (n217,n218,n225);
nand (n218,n219,n221);
or (n219,n220,n57);
not (n220,n69);
nand (n221,n63,n222);
nor (n222,n223,n224);
and (n223,n121,n56);
and (n224,n119,n52);
nand (n225,n226,n227);
or (n226,n76,n96);
nand (n227,n85,n228);
nor (n228,n229,n230);
and (n229,n53,n81);
and (n230,n54,n82);
nand (n231,n232,n233);
or (n232,n107,n123);
or (n233,n234,n128);
nor (n234,n235,n236);
and (n235,n65,n26);
and (n236,n66,n25);
xor (n237,n238,n252);
xor (n238,n239,n246);
nand (n239,n240,n241);
or (n240,n149,n131);
nand (n241,n242,n133);
not (n242,n243);
nor (n243,n244,n245);
and (n244,n142,n92);
and (n245,n140,n91);
nand (n246,n247,n248);
or (n247,n171,n156);
or (n248,n157,n249);
nor (n249,n250,n251);
and (n250,n163,n145);
and (n251,n164,n147);
and (n252,n253,n258);
nor (n253,n254,n163);
nor (n254,n255,n257);
and (n255,n256,n142);
nand (n256,n168,n160);
and (n257,n167,n159);
nand (n258,n259,n260);
or (n259,n188,n190);
or (n260,n261,n187);
nor (n261,n262,n263);
and (n262,n211,n36);
and (n263,n212,n195);
or (n264,n265,n309);
and (n265,n266,n287);
xor (n266,n267,n268);
xor (n267,n253,n258);
or (n268,n269,n286);
and (n269,n270,n280);
xor (n270,n271,n273);
and (n271,n272,n168);
not (n272,n157);
nand (n273,n274,n279);
or (n274,n275,n30);
not (n275,n276);
nand (n276,n277,n278);
or (n277,n28,n127);
or (n278,n27,n125);
nand (n279,n32,n23);
nand (n280,n281,n282);
or (n281,n49,n62);
or (n282,n57,n283);
nor (n283,n284,n285);
and (n284,n100,n52);
and (n285,n98,n56);
and (n286,n271,n273);
or (n287,n288,n308);
and (n288,n289,n302);
xor (n289,n290,n296);
nand (n290,n291,n295);
or (n291,n292,n76);
nor (n292,n293,n294);
and (n293,n151,n82);
and (n294,n152,n81);
nand (n295,n89,n85);
nand (n296,n297,n301);
or (n297,n298,n187);
nor (n298,n299,n300);
and (n299,n195,n45);
and (n300,n36,n44);
or (n301,n261,n188);
nand (n302,n303,n307);
or (n303,n304,n131);
nor (n304,n305,n306);
and (n305,n142,n173);
and (n306,n140,n175);
or (n307,n143,n132);
and (n308,n290,n296);
and (n309,n267,n268);
or (n310,n311,n362);
and (n311,n312,n315);
xor (n312,n313,n314);
xor (n313,n104,n154);
xor (n314,n19,n74);
or (n315,n316,n361);
and (n316,n317,n339);
xor (n317,n318,n324);
nand (n318,n319,n323);
or (n319,n107,n320);
nor (n320,n321,n322);
and (n321,n65,n72);
and (n322,n66,n71);
or (n323,n117,n128);
and (n324,n325,n332);
nand (n325,n326,n331);
or (n326,n327,n30);
not (n327,n328);
nand (n328,n329,n330);
or (n329,n28,n121);
or (n330,n27,n119);
nand (n331,n32,n276);
not (n332,n333);
nand (n333,n334,n140);
nand (n334,n335,n336);
or (n335,n168,n136);
nand (n336,n337,n81);
not (n337,n338);
and (n338,n168,n136);
or (n339,n340,n360);
and (n340,n341,n354);
xor (n341,n342,n348);
nand (n342,n343,n347);
or (n343,n57,n344);
nor (n344,n345,n346);
and (n345,n92,n56);
and (n346,n91,n52);
or (n347,n283,n62);
nand (n348,n349,n353);
or (n349,n76,n350);
nor (n350,n351,n352);
and (n351,n145,n81);
and (n352,n147,n82);
or (n353,n95,n292);
nand (n354,n355,n359);
or (n355,n356,n187);
nor (n356,n357,n358);
and (n357,n195,n26);
and (n358,n36,n25);
or (n359,n298,n188);
and (n360,n342,n348);
and (n361,n318,n324);
and (n362,n313,n314);
not (n363,n364);
or (n364,n365,n395);
and (n365,n366,n394);
xor (n366,n367,n368);
xor (n367,n266,n287);
or (n368,n369,n393);
and (n369,n370,n373);
xor (n370,n371,n372);
xor (n371,n289,n302);
xor (n372,n270,n280);
or (n373,n374,n392);
and (n374,n375,n388);
xor (n375,n376,n382);
nand (n376,n377,n381);
or (n377,n131,n378);
nor (n378,n379,n380);
and (n379,n167,n140);
and (n380,n142,n168);
or (n381,n132,n304);
nand (n382,n383,n387);
or (n383,n107,n384);
nor (n384,n385,n386);
and (n385,n65,n54);
and (n386,n66,n53);
or (n387,n320,n128);
nand (n388,n389,n391);
or (n389,n332,n390);
not (n390,n325);
or (n391,n325,n333);
and (n392,n376,n382);
and (n393,n371,n372);
xor (n394,n312,n315);
and (n395,n367,n368);
nand (n396,n13,n364);
not (n397,n398);
nand (n398,n399,n802);
or (n399,n400,n504);
not (n400,n401);
nor (n401,n402,n455);
nor (n402,n403,n404);
xor (n403,n366,n394);
or (n404,n405,n454);
and (n405,n406,n453);
xor (n406,n407,n408);
xor (n407,n317,n339);
or (n408,n409,n452);
and (n409,n410,n451);
xor (n410,n411,n429);
or (n411,n412,n428);
and (n412,n413,n421);
xor (n413,n414,n415);
and (n414,n133,n168);
nand (n415,n416,n420);
or (n416,n417,n30);
nor (n417,n418,n419);
and (n418,n71,n28);
and (n419,n72,n27);
nand (n420,n32,n328);
nand (n421,n422,n427);
or (n422,n57,n423);
not (n423,n424);
nor (n424,n425,n426);
and (n425,n151,n56);
and (n426,n152,n52);
or (n427,n62,n344);
and (n428,n414,n415);
or (n429,n430,n450);
and (n430,n431,n444);
xor (n431,n432,n438);
nand (n432,n433,n437);
or (n433,n76,n434);
nor (n434,n435,n436);
and (n435,n175,n82);
and (n436,n173,n81);
or (n437,n95,n350);
nand (n438,n439,n443);
or (n439,n440,n187);
nor (n440,n441,n442);
and (n441,n195,n125);
and (n442,n36,n127);
or (n443,n356,n188);
nand (n444,n445,n449);
or (n445,n107,n446);
nor (n446,n447,n448);
and (n447,n65,n98);
and (n448,n66,n100);
or (n449,n384,n128);
and (n450,n432,n438);
xor (n451,n341,n354);
and (n452,n411,n429);
xor (n453,n370,n373);
and (n454,n407,n408);
nor (n455,n456,n503);
or (n456,n457,n502);
and (n457,n458,n461);
xor (n458,n459,n460);
xor (n459,n375,n388);
xor (n460,n410,n451);
or (n461,n462,n501);
and (n462,n463,n500);
xor (n463,n464,n477);
and (n464,n465,n471);
and (n465,n466,n82);
nand (n466,n467,n468);
or (n467,n168,n80);
nand (n468,n469,n56);
not (n469,n470);
and (n470,n168,n80);
nand (n471,n472,n476);
or (n472,n30,n473);
nor (n473,n474,n475);
and (n474,n27,n54);
and (n475,n28,n53);
or (n476,n31,n417);
or (n477,n478,n499);
and (n478,n479,n493);
xor (n479,n480,n487);
nand (n480,n481,n486);
or (n481,n482,n57);
not (n482,n483);
nor (n483,n484,n485);
and (n484,n145,n52);
and (n485,n147,n56);
nand (n486,n63,n424);
nand (n487,n488,n492);
or (n488,n76,n489);
nor (n489,n490,n491);
and (n490,n82,n167);
and (n491,n81,n168);
or (n492,n95,n434);
nand (n493,n494,n498);
or (n494,n187,n495);
nor (n495,n496,n497);
and (n496,n195,n119);
and (n497,n36,n121);
or (n498,n440,n188);
and (n499,n480,n487);
xor (n500,n413,n421);
and (n501,n464,n477);
and (n502,n459,n460);
xor (n503,n406,n453);
not (n504,n505);
nand (n505,n506,n791,n801);
nand (n506,n507,n546,n650);
nand (n507,n508,n510);
not (n508,n509);
xor (n509,n458,n461);
not (n510,n511);
or (n511,n512,n545);
and (n512,n513,n544);
xor (n513,n514,n515);
xor (n514,n431,n444);
or (n515,n516,n543);
and (n516,n517,n525);
xor (n517,n518,n524);
nand (n518,n519,n523);
or (n519,n107,n520);
nor (n520,n521,n522);
and (n521,n65,n92);
and (n522,n66,n91);
or (n523,n446,n128);
xor (n524,n465,n471);
or (n525,n526,n542);
and (n526,n527,n535);
xor (n527,n528,n529);
and (n528,n85,n168);
nand (n529,n530,n534);
or (n530,n531,n187);
nor (n531,n532,n533);
and (n532,n195,n72);
and (n533,n36,n71);
or (n534,n495,n188);
nand (n535,n536,n541);
or (n536,n57,n537);
not (n537,n538);
nand (n538,n539,n540);
or (n539,n52,n175);
or (n540,n56,n173);
or (n541,n62,n482);
and (n542,n528,n529);
and (n543,n518,n524);
xor (n544,n463,n500);
and (n545,n514,n515);
nor (n546,n547,n587);
not (n547,n548);
or (n548,n549,n550);
xor (n549,n513,n544);
or (n550,n551,n586);
and (n551,n552,n585);
xor (n552,n553,n554);
xor (n553,n479,n493);
or (n554,n555,n584);
and (n555,n556,n569);
xor (n556,n557,n563);
nand (n557,n558,n562);
or (n558,n30,n559);
nor (n559,n560,n561);
and (n560,n27,n98);
and (n561,n28,n100);
or (n562,n31,n473);
nand (n563,n564,n568);
or (n564,n107,n565);
nor (n565,n566,n567);
and (n566,n65,n152);
and (n567,n66,n151);
or (n568,n520,n128);
and (n569,n570,n577);
nor (n570,n571,n56);
nor (n571,n572,n575);
and (n572,n573,n65);
not (n573,n574);
and (n574,n168,n60);
and (n575,n167,n576);
not (n576,n60);
nand (n577,n578,n583);
or (n578,n187,n579);
not (n579,n580);
nor (n580,n581,n582);
and (n581,n54,n36);
and (n582,n53,n195);
or (n583,n531,n188);
and (n584,n557,n563);
xor (n585,n517,n525);
and (n586,n553,n554);
nand (n587,n588,n644);
not (n588,n589);
nor (n589,n590,n619);
xor (n590,n591,n618);
xor (n591,n592,n617);
or (n592,n593,n616);
and (n593,n594,n610);
xor (n594,n595,n602);
nand (n595,n596,n601);
or (n596,n597,n57);
not (n597,n598);
nand (n598,n599,n600);
or (n599,n56,n168);
or (n600,n52,n167);
nand (n601,n63,n538);
nand (n602,n603,n608);
or (n603,n604,n30);
not (n604,n605);
nand (n605,n606,n607);
or (n606,n28,n91);
or (n607,n27,n92);
nand (n608,n609,n32);
not (n609,n559);
nand (n610,n611,n615);
or (n611,n107,n612);
nor (n612,n613,n614);
and (n613,n65,n145);
and (n614,n66,n147);
or (n615,n565,n128);
and (n616,n595,n602);
xor (n617,n527,n535);
xor (n618,n556,n569);
or (n619,n620,n643);
and (n620,n621,n642);
xor (n621,n622,n623);
xor (n622,n570,n577);
or (n623,n624,n641);
and (n624,n625,n634);
xor (n625,n626,n627);
and (n626,n63,n168);
nand (n627,n628,n629);
or (n628,n188,n579);
or (n629,n630,n187);
not (n630,n631);
nand (n631,n632,n633);
or (n632,n98,n195);
nand (n633,n195,n98);
nand (n634,n635,n640);
or (n635,n636,n30);
not (n636,n637);
nand (n637,n638,n639);
or (n638,n28,n151);
or (n639,n27,n152);
nand (n640,n32,n605);
and (n641,n626,n627);
xor (n642,n594,n610);
and (n643,n622,n623);
not (n644,n645);
nor (n645,n646,n647);
xor (n646,n552,n585);
or (n647,n648,n649);
and (n648,n591,n618);
and (n649,n592,n617);
or (n650,n651,n790);
and (n651,n652,n679);
xor (n652,n653,n678);
or (n653,n654,n677);
and (n654,n655,n676);
xor (n655,n656,n662);
nand (n656,n657,n661);
or (n657,n107,n658);
nor (n658,n659,n660);
and (n659,n65,n173);
and (n660,n66,n175);
or (n661,n612,n128);
nor (n662,n663,n671);
not (n663,n664);
nand (n664,n665,n670);
or (n665,n187,n666);
not (n666,n667);
nor (n667,n668,n669);
and (n668,n92,n36);
and (n669,n91,n195);
nand (n670,n631,n189);
nand (n671,n672,n66);
nand (n672,n673,n675);
or (n673,n674,n28);
and (n674,n168,n111);
or (n675,n168,n111);
xor (n676,n625,n634);
and (n677,n656,n662);
xor (n678,n621,n642);
or (n679,n680,n789);
and (n680,n681,n705);
xor (n681,n682,n704);
or (n682,n683,n703);
and (n683,n684,n699);
xor (n684,n685,n692);
nand (n685,n686,n691);
or (n686,n687,n30);
not (n687,n688);
nor (n688,n689,n690);
and (n689,n147,n27);
and (n690,n145,n28);
nand (n691,n32,n637);
nand (n692,n693,n698);
or (n693,n694,n107);
not (n694,n695);
nand (n695,n696,n697);
or (n696,n65,n168);
or (n697,n167,n66);
or (n698,n658,n128);
nand (n699,n700,n702);
or (n700,n701,n663);
not (n701,n671);
or (n702,n664,n671);
and (n703,n685,n692);
xor (n704,n655,n676);
or (n705,n706,n788);
and (n706,n707,n728);
xor (n707,n708,n727);
or (n708,n709,n726);
and (n709,n710,n719);
xor (n710,n711,n712);
and (n711,n109,n168);
nand (n712,n713,n718);
or (n713,n714,n30);
not (n714,n715);
nor (n715,n716,n717);
and (n716,n175,n27);
and (n717,n173,n28);
nand (n718,n32,n688);
nand (n719,n720,n721);
or (n720,n188,n666);
or (n721,n187,n722);
not (n722,n723);
nor (n723,n724,n725);
and (n724,n151,n195);
and (n725,n152,n36);
and (n726,n711,n712);
xor (n727,n684,n699);
nand (n728,n729,n787);
or (n729,n730,n746);
nor (n730,n731,n732);
xor (n731,n710,n719);
and (n732,n733,n740);
nand (n733,n734,n735);
nand (n734,n723,n189);
nand (n735,n736,n739);
nor (n736,n737,n738);
and (n737,n147,n195);
and (n738,n145,n36);
not (n739,n187);
not (n740,n741);
nand (n741,n742,n28);
nand (n742,n743,n745);
or (n743,n744,n36);
and (n744,n168,n35);
or (n745,n168,n35);
nor (n746,n747,n786);
and (n747,n748,n760);
nand (n748,n749,n753);
nor (n749,n750,n752);
and (n750,n751,n740);
not (n751,n733);
and (n752,n733,n741);
nor (n753,n754,n755);
and (n754,n32,n715);
and (n755,n756,n757);
not (n756,n30);
nand (n757,n758,n759);
or (n758,n27,n168);
or (n759,n167,n28);
nand (n760,n761,n784);
or (n761,n762,n776);
not (n762,n763);
and (n763,n764,n774);
nand (n764,n765,n770);
or (n765,n188,n766);
not (n766,n767);
nor (n767,n768,n769);
and (n768,n175,n195);
and (n769,n173,n36);
nand (n770,n771,n739);
nand (n771,n772,n773);
or (n772,n195,n168);
or (n773,n36,n167);
nor (n774,n775,n195);
and (n775,n168,n189);
not (n776,n777);
nand (n777,n778,n783);
not (n778,n779);
nand (n779,n780,n782);
or (n780,n188,n781);
not (n781,n736);
nand (n782,n767,n739);
nand (n783,n32,n168);
nand (n784,n785,n779);
not (n785,n783);
nor (n786,n749,n753);
nand (n787,n731,n732);
and (n788,n708,n727);
and (n789,n682,n704);
and (n790,n653,n678);
nand (n791,n792,n507);
or (n792,n793,n795);
not (n793,n794);
nand (n794,n549,n550);
not (n795,n796);
nand (n796,n548,n797);
nand (n797,n798,n800);
or (n798,n645,n799);
nand (n799,n590,n619);
nand (n800,n646,n647);
nand (n801,n509,n511);
not (n802,n803);
nand (n803,n804,n806);
or (n804,n402,n805);
nand (n805,n456,n503);
nand (n806,n403,n404);
or (n807,n398,n10);
not (n808,n809);
nand (n809,n810,n3);
not (n810,n4);
wire s0n811,s1n811,notn811;
or (n811,s0n811,s1n811);
not(notn811,n4);
and (s0n811,notn811,n812);
and (s1n811,n4,1'b0);
wire s0n812,s1n812,notn812;
or (n812,s0n812,s1n812);
not(notn812,n3);
and (s0n812,notn812,n5);
and (s1n812,n3,n813);
xor (n813,n814,n1345);
xor (n814,n815,n1342);
xor (n815,n816,n1341);
xor (n816,n817,n1332);
xor (n817,n818,n1331);
xor (n818,n819,n1316);
xor (n819,n820,n1315);
xor (n820,n821,n1295);
xor (n821,n822,n1294);
xor (n822,n823,n1267);
xor (n823,n824,n1266);
xor (n824,n825,n1234);
xor (n825,n826,n1233);
xor (n826,n827,n1196);
xor (n827,n828,n1195);
xor (n828,n829,n1151);
xor (n829,n830,n1150);
xor (n830,n831,n1099);
xor (n831,n832,n1098);
xor (n832,n833,n1042);
xor (n833,n834,n1041);
xor (n834,n835,n981);
xor (n835,n836,n980);
xor (n836,n837,n912);
xor (n837,n838,n911);
xor (n838,n839,n841);
xor (n839,n840,n196);
and (n840,n202,n189);
or (n841,n842,n845);
and (n842,n843,n844);
and (n843,n194,n189);
and (n844,n212,n36);
and (n845,n846,n847);
xor (n846,n843,n844);
or (n847,n848,n851);
and (n848,n849,n850);
and (n849,n212,n189);
and (n850,n45,n36);
and (n851,n852,n853);
xor (n852,n849,n850);
or (n853,n854,n857);
and (n854,n855,n856);
and (n855,n45,n189);
and (n856,n26,n36);
and (n857,n858,n859);
xor (n858,n855,n856);
or (n859,n860,n863);
and (n860,n861,n862);
and (n861,n26,n189);
and (n862,n125,n36);
and (n863,n864,n865);
xor (n864,n861,n862);
or (n865,n866,n869);
and (n866,n867,n868);
and (n867,n125,n189);
and (n868,n119,n36);
and (n869,n870,n871);
xor (n870,n867,n868);
or (n871,n872,n875);
and (n872,n873,n874);
and (n873,n119,n189);
and (n874,n72,n36);
and (n875,n876,n877);
xor (n876,n873,n874);
or (n877,n878,n880);
and (n878,n879,n581);
and (n879,n72,n189);
and (n880,n881,n882);
xor (n881,n879,n581);
or (n882,n883,n886);
and (n883,n884,n885);
and (n884,n54,n189);
and (n885,n98,n36);
and (n886,n887,n888);
xor (n887,n884,n885);
or (n888,n889,n891);
and (n889,n890,n668);
and (n890,n98,n189);
and (n891,n892,n893);
xor (n892,n890,n668);
or (n893,n894,n896);
and (n894,n895,n725);
and (n895,n92,n189);
and (n896,n897,n898);
xor (n897,n895,n725);
or (n898,n899,n901);
and (n899,n900,n738);
and (n900,n152,n189);
and (n901,n902,n903);
xor (n902,n900,n738);
or (n903,n904,n906);
and (n904,n905,n769);
and (n905,n145,n189);
and (n906,n907,n908);
xor (n907,n905,n769);
and (n908,n909,n910);
and (n909,n173,n189);
and (n910,n168,n36);
and (n911,n212,n35);
or (n912,n913,n916);
and (n913,n914,n915);
xor (n914,n846,n847);
and (n915,n45,n35);
and (n916,n917,n918);
xor (n917,n914,n915);
or (n918,n919,n922);
and (n919,n920,n921);
xor (n920,n852,n853);
and (n921,n26,n35);
and (n922,n923,n924);
xor (n923,n920,n921);
or (n924,n925,n928);
and (n925,n926,n927);
xor (n926,n858,n859);
and (n927,n125,n35);
and (n928,n929,n930);
xor (n929,n926,n927);
or (n930,n931,n934);
and (n931,n932,n933);
xor (n932,n864,n865);
and (n933,n119,n35);
and (n934,n935,n936);
xor (n935,n932,n933);
or (n936,n937,n940);
and (n937,n938,n939);
xor (n938,n870,n871);
and (n939,n72,n35);
and (n940,n941,n942);
xor (n941,n938,n939);
or (n942,n943,n946);
and (n943,n944,n945);
xor (n944,n876,n877);
and (n945,n54,n35);
and (n946,n947,n948);
xor (n947,n944,n945);
or (n948,n949,n952);
and (n949,n950,n951);
xor (n950,n881,n882);
and (n951,n98,n35);
and (n952,n953,n954);
xor (n953,n950,n951);
or (n954,n955,n958);
and (n955,n956,n957);
xor (n956,n887,n888);
and (n957,n92,n35);
and (n958,n959,n960);
xor (n959,n956,n957);
or (n960,n961,n964);
and (n961,n962,n963);
xor (n962,n892,n893);
and (n963,n152,n35);
and (n964,n965,n966);
xor (n965,n962,n963);
or (n966,n967,n970);
and (n967,n968,n969);
xor (n968,n897,n898);
and (n969,n145,n35);
and (n970,n971,n972);
xor (n971,n968,n969);
or (n972,n973,n976);
and (n973,n974,n975);
xor (n974,n902,n903);
and (n975,n173,n35);
and (n976,n977,n978);
xor (n977,n974,n975);
and (n978,n979,n744);
xor (n979,n907,n908);
and (n980,n45,n28);
or (n981,n982,n984);
and (n982,n983,n29);
xor (n983,n917,n918);
and (n984,n985,n986);
xor (n985,n983,n29);
or (n986,n987,n990);
and (n987,n988,n989);
xor (n988,n923,n924);
and (n989,n125,n28);
and (n990,n991,n992);
xor (n991,n988,n989);
or (n992,n993,n996);
and (n993,n994,n995);
xor (n994,n929,n930);
and (n995,n119,n28);
and (n996,n997,n998);
xor (n997,n994,n995);
or (n998,n999,n1002);
and (n999,n1000,n1001);
xor (n1000,n935,n936);
and (n1001,n72,n28);
and (n1002,n1003,n1004);
xor (n1003,n1000,n1001);
or (n1004,n1005,n1008);
and (n1005,n1006,n1007);
xor (n1006,n941,n942);
and (n1007,n54,n28);
and (n1008,n1009,n1010);
xor (n1009,n1006,n1007);
or (n1010,n1011,n1014);
and (n1011,n1012,n1013);
xor (n1012,n947,n948);
and (n1013,n98,n28);
and (n1014,n1015,n1016);
xor (n1015,n1012,n1013);
or (n1016,n1017,n1020);
and (n1017,n1018,n1019);
xor (n1018,n953,n954);
and (n1019,n92,n28);
and (n1020,n1021,n1022);
xor (n1021,n1018,n1019);
or (n1022,n1023,n1026);
and (n1023,n1024,n1025);
xor (n1024,n959,n960);
and (n1025,n152,n28);
and (n1026,n1027,n1028);
xor (n1027,n1024,n1025);
or (n1028,n1029,n1031);
and (n1029,n1030,n690);
xor (n1030,n965,n966);
and (n1031,n1032,n1033);
xor (n1032,n1030,n690);
or (n1033,n1034,n1036);
and (n1034,n1035,n717);
xor (n1035,n971,n972);
and (n1036,n1037,n1038);
xor (n1037,n1035,n717);
and (n1038,n1039,n1040);
xor (n1039,n977,n978);
and (n1040,n168,n28);
and (n1041,n26,n111);
or (n1042,n1043,n1046);
and (n1043,n1044,n1045);
xor (n1044,n985,n986);
and (n1045,n125,n111);
and (n1046,n1047,n1048);
xor (n1047,n1044,n1045);
or (n1048,n1049,n1052);
and (n1049,n1050,n1051);
xor (n1050,n991,n992);
and (n1051,n119,n111);
and (n1052,n1053,n1054);
xor (n1053,n1050,n1051);
or (n1054,n1055,n1058);
and (n1055,n1056,n1057);
xor (n1056,n997,n998);
and (n1057,n72,n111);
and (n1058,n1059,n1060);
xor (n1059,n1056,n1057);
or (n1060,n1061,n1064);
and (n1061,n1062,n1063);
xor (n1062,n1003,n1004);
and (n1063,n54,n111);
and (n1064,n1065,n1066);
xor (n1065,n1062,n1063);
or (n1066,n1067,n1070);
and (n1067,n1068,n1069);
xor (n1068,n1009,n1010);
and (n1069,n98,n111);
and (n1070,n1071,n1072);
xor (n1071,n1068,n1069);
or (n1072,n1073,n1076);
and (n1073,n1074,n1075);
xor (n1074,n1015,n1016);
and (n1075,n92,n111);
and (n1076,n1077,n1078);
xor (n1077,n1074,n1075);
or (n1078,n1079,n1082);
and (n1079,n1080,n1081);
xor (n1080,n1021,n1022);
and (n1081,n152,n111);
and (n1082,n1083,n1084);
xor (n1083,n1080,n1081);
or (n1084,n1085,n1088);
and (n1085,n1086,n1087);
xor (n1086,n1027,n1028);
and (n1087,n145,n111);
and (n1088,n1089,n1090);
xor (n1089,n1086,n1087);
or (n1090,n1091,n1094);
and (n1091,n1092,n1093);
xor (n1092,n1032,n1033);
and (n1093,n173,n111);
and (n1094,n1095,n1096);
xor (n1095,n1092,n1093);
and (n1096,n1097,n674);
xor (n1097,n1037,n1038);
and (n1098,n125,n66);
or (n1099,n1100,n1103);
and (n1100,n1101,n1102);
xor (n1101,n1047,n1048);
and (n1102,n119,n66);
and (n1103,n1104,n1105);
xor (n1104,n1101,n1102);
or (n1105,n1106,n1109);
and (n1106,n1107,n1108);
xor (n1107,n1053,n1054);
and (n1108,n72,n66);
and (n1109,n1110,n1111);
xor (n1110,n1107,n1108);
or (n1111,n1112,n1115);
and (n1112,n1113,n1114);
xor (n1113,n1059,n1060);
and (n1114,n54,n66);
and (n1115,n1116,n1117);
xor (n1116,n1113,n1114);
or (n1117,n1118,n1121);
and (n1118,n1119,n1120);
xor (n1119,n1065,n1066);
and (n1120,n98,n66);
and (n1121,n1122,n1123);
xor (n1122,n1119,n1120);
or (n1123,n1124,n1127);
and (n1124,n1125,n1126);
xor (n1125,n1071,n1072);
and (n1126,n92,n66);
and (n1127,n1128,n1129);
xor (n1128,n1125,n1126);
or (n1129,n1130,n1133);
and (n1130,n1131,n1132);
xor (n1131,n1077,n1078);
and (n1132,n152,n66);
and (n1133,n1134,n1135);
xor (n1134,n1131,n1132);
or (n1135,n1136,n1139);
and (n1136,n1137,n1138);
xor (n1137,n1083,n1084);
and (n1138,n145,n66);
and (n1139,n1140,n1141);
xor (n1140,n1137,n1138);
or (n1141,n1142,n1145);
and (n1142,n1143,n1144);
xor (n1143,n1089,n1090);
and (n1144,n173,n66);
and (n1145,n1146,n1147);
xor (n1146,n1143,n1144);
and (n1147,n1148,n1149);
xor (n1148,n1095,n1096);
and (n1149,n168,n66);
and (n1150,n119,n60);
or (n1151,n1152,n1155);
and (n1152,n1153,n1154);
xor (n1153,n1104,n1105);
and (n1154,n72,n60);
and (n1155,n1156,n1157);
xor (n1156,n1153,n1154);
or (n1157,n1158,n1161);
and (n1158,n1159,n1160);
xor (n1159,n1110,n1111);
and (n1160,n54,n60);
and (n1161,n1162,n1163);
xor (n1162,n1159,n1160);
or (n1163,n1164,n1167);
and (n1164,n1165,n1166);
xor (n1165,n1116,n1117);
and (n1166,n98,n60);
and (n1167,n1168,n1169);
xor (n1168,n1165,n1166);
or (n1169,n1170,n1173);
and (n1170,n1171,n1172);
xor (n1171,n1122,n1123);
and (n1172,n92,n60);
and (n1173,n1174,n1175);
xor (n1174,n1171,n1172);
or (n1175,n1176,n1179);
and (n1176,n1177,n1178);
xor (n1177,n1128,n1129);
and (n1178,n152,n60);
and (n1179,n1180,n1181);
xor (n1180,n1177,n1178);
or (n1181,n1182,n1185);
and (n1182,n1183,n1184);
xor (n1183,n1134,n1135);
and (n1184,n145,n60);
and (n1185,n1186,n1187);
xor (n1186,n1183,n1184);
or (n1187,n1188,n1191);
and (n1188,n1189,n1190);
xor (n1189,n1140,n1141);
and (n1190,n173,n60);
and (n1191,n1192,n1193);
xor (n1192,n1189,n1190);
and (n1193,n1194,n574);
xor (n1194,n1146,n1147);
and (n1195,n72,n52);
or (n1196,n1197,n1200);
and (n1197,n1198,n1199);
xor (n1198,n1156,n1157);
and (n1199,n54,n52);
and (n1200,n1201,n1202);
xor (n1201,n1198,n1199);
or (n1202,n1203,n1206);
and (n1203,n1204,n1205);
xor (n1204,n1162,n1163);
and (n1205,n98,n52);
and (n1206,n1207,n1208);
xor (n1207,n1204,n1205);
or (n1208,n1209,n1212);
and (n1209,n1210,n1211);
xor (n1210,n1168,n1169);
and (n1211,n92,n52);
and (n1212,n1213,n1214);
xor (n1213,n1210,n1211);
or (n1214,n1215,n1217);
and (n1215,n1216,n426);
xor (n1216,n1174,n1175);
and (n1217,n1218,n1219);
xor (n1218,n1216,n426);
or (n1219,n1220,n1222);
and (n1220,n1221,n484);
xor (n1221,n1180,n1181);
and (n1222,n1223,n1224);
xor (n1223,n1221,n484);
or (n1224,n1225,n1228);
and (n1225,n1226,n1227);
xor (n1226,n1186,n1187);
and (n1227,n173,n52);
and (n1228,n1229,n1230);
xor (n1229,n1226,n1227);
and (n1230,n1231,n1232);
xor (n1231,n1192,n1193);
and (n1232,n168,n52);
and (n1233,n54,n80);
or (n1234,n1235,n1238);
and (n1235,n1236,n1237);
xor (n1236,n1201,n1202);
and (n1237,n98,n80);
and (n1238,n1239,n1240);
xor (n1239,n1236,n1237);
or (n1240,n1241,n1244);
and (n1241,n1242,n1243);
xor (n1242,n1207,n1208);
and (n1243,n92,n80);
and (n1244,n1245,n1246);
xor (n1245,n1242,n1243);
or (n1246,n1247,n1250);
and (n1247,n1248,n1249);
xor (n1248,n1213,n1214);
and (n1249,n152,n80);
and (n1250,n1251,n1252);
xor (n1251,n1248,n1249);
or (n1252,n1253,n1256);
and (n1253,n1254,n1255);
xor (n1254,n1218,n1219);
and (n1255,n145,n80);
and (n1256,n1257,n1258);
xor (n1257,n1254,n1255);
or (n1258,n1259,n1262);
and (n1259,n1260,n1261);
xor (n1260,n1223,n1224);
and (n1261,n173,n80);
and (n1262,n1263,n1264);
xor (n1263,n1260,n1261);
and (n1264,n1265,n470);
xor (n1265,n1229,n1230);
and (n1266,n98,n82);
or (n1267,n1268,n1271);
and (n1268,n1269,n1270);
xor (n1269,n1239,n1240);
and (n1270,n92,n82);
and (n1271,n1272,n1273);
xor (n1272,n1269,n1270);
or (n1273,n1274,n1277);
and (n1274,n1275,n1276);
xor (n1275,n1245,n1246);
and (n1276,n152,n82);
and (n1277,n1278,n1279);
xor (n1278,n1275,n1276);
or (n1279,n1280,n1283);
and (n1280,n1281,n1282);
xor (n1281,n1251,n1252);
and (n1282,n145,n82);
and (n1283,n1284,n1285);
xor (n1284,n1281,n1282);
or (n1285,n1286,n1289);
and (n1286,n1287,n1288);
xor (n1287,n1257,n1258);
and (n1288,n173,n82);
and (n1289,n1290,n1291);
xor (n1290,n1287,n1288);
and (n1291,n1292,n1293);
xor (n1292,n1263,n1264);
and (n1293,n168,n82);
and (n1294,n92,n136);
or (n1295,n1296,n1299);
and (n1296,n1297,n1298);
xor (n1297,n1272,n1273);
and (n1298,n152,n136);
and (n1299,n1300,n1301);
xor (n1300,n1297,n1298);
or (n1301,n1302,n1305);
and (n1302,n1303,n1304);
xor (n1303,n1278,n1279);
and (n1304,n145,n136);
and (n1305,n1306,n1307);
xor (n1306,n1303,n1304);
or (n1307,n1308,n1311);
and (n1308,n1309,n1310);
xor (n1309,n1284,n1285);
and (n1310,n173,n136);
and (n1311,n1312,n1313);
xor (n1312,n1309,n1310);
and (n1313,n1314,n338);
xor (n1314,n1290,n1291);
and (n1315,n152,n140);
or (n1316,n1317,n1320);
and (n1317,n1318,n1319);
xor (n1318,n1300,n1301);
and (n1319,n145,n140);
and (n1320,n1321,n1322);
xor (n1321,n1318,n1319);
or (n1322,n1323,n1326);
and (n1323,n1324,n1325);
xor (n1324,n1306,n1307);
and (n1325,n173,n140);
and (n1326,n1327,n1328);
xor (n1327,n1324,n1325);
and (n1328,n1329,n1330);
xor (n1329,n1312,n1313);
and (n1330,n168,n140);
and (n1331,n145,n160);
or (n1332,n1333,n1336);
and (n1333,n1334,n1335);
xor (n1334,n1321,n1322);
and (n1335,n173,n160);
and (n1336,n1337,n1338);
xor (n1337,n1334,n1335);
and (n1338,n1339,n1340);
xor (n1339,n1327,n1328);
not (n1340,n256);
and (n1341,n173,n164);
and (n1342,n1343,n1344);
xor (n1343,n1337,n1338);
and (n1344,n168,n164);
not (n1345,n1346);
nand (n1346,n168,n183);
endmodule
