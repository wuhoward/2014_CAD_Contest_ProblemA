module top (out,n4,n12,n14,n15,n17,n19,n20,n25,n31
        ,n34,n35,n41,n42,n57,n59,n60,n69,n70,n72
        ,n73,n83,n92,n105,n106,n113,n119,n132,n138,n157
        ,n163,n517);
output out;
input n4;
input n12;
input n14;
input n15;
input n17;
input n19;
input n20;
input n25;
input n31;
input n34;
input n35;
input n41;
input n42;
input n57;
input n59;
input n60;
input n69;
input n70;
input n72;
input n73;
input n83;
input n92;
input n105;
input n106;
input n113;
input n119;
input n132;
input n138;
input n157;
input n163;
input n517;
wire n0;
wire n1;
wire n2;
wire n3;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n13;
wire n16;
wire n18;
wire n21;
wire n22;
wire n23;
wire n24;
wire n26;
wire n27;
wire n28;
wire n29;
wire n30;
wire n32;
wire n33;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n58;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n71;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n91;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
xnor (out,n0,n518);
nand (n0,n1,n517);
nand (n1,n2,n43);
or (n2,n3,n5);
not (n3,n4);
not (n5,n6);
xor (n6,n7,n39);
xor (n7,n8,n36);
xor (n8,n9,n32);
xor (n9,n10,n21);
xor (n10,n11,n16);
and (n11,n12,n13);
wire s0n13,s1n13,notn13;
or (n13,s0n13,s1n13);
not(notn13,n4);
and (s0n13,notn13,n14);
and (s1n13,n4,n15);
and (n16,n17,n18);
wire s0n18,s1n18,notn18;
or (n18,s0n18,s1n18);
not(notn18,n4);
and (s0n18,notn18,n19);
and (s1n18,n4,n20);
or (n21,n22,n26);
and (n22,n23,n24);
and (n23,n17,n13);
and (n24,n25,n18);
and (n26,n27,n28);
xor (n27,n23,n24);
and (n28,n29,n30);
and (n29,n25,n13);
and (n30,n31,n18);
and (n32,n25,n33);
wire s0n33,s1n33,notn33;
or (n33,s0n33,s1n33);
not(notn33,n4);
and (s0n33,notn33,n34);
and (s1n33,n4,n35);
and (n36,n37,n38);
xor (n37,n27,n28);
and (n38,n31,n33);
and (n39,n31,n40);
wire s0n40,s1n40,notn40;
or (n40,s0n40,s1n40);
not(notn40,n4);
and (s0n40,notn40,n41);
and (s1n40,n4,n42);
nand (n43,n44,n3);
xnor (n44,n45,n266);
nand (n45,n46,n265);
nand (n46,n47,n224);
not (n47,n48);
xor (n48,n49,n201);
xor (n49,n50,n122);
xor (n50,n51,n97);
xor (n51,n52,n86);
nand (n52,n53,n79);
or (n53,n54,n64);
not (n54,n55);
nor (n55,n56,n61);
and (n56,n57,n58);
wire s0n58,s1n58,notn58;
or (n58,s0n58,s1n58);
not(notn58,n4);
and (s0n58,notn58,n59);
and (s1n58,n4,n60);
and (n61,n62,n63);
not (n62,n57);
not (n63,n58);
nand (n64,n65,n76);
nor (n65,n66,n74);
and (n66,n67,n71);
not (n67,n68);
wire s0n68,s1n68,notn68;
or (n68,s0n68,s1n68);
not(notn68,n4);
and (s0n68,notn68,n69);
and (s1n68,n4,n70);
wire s0n71,s1n71,notn71;
or (n71,s0n71,s1n71);
not(notn71,n4);
and (s0n71,notn71,n72);
and (s1n71,n4,n73);
and (n74,n68,n75);
not (n75,n71);
nand (n76,n77,n78);
or (n77,n67,n58);
nand (n78,n58,n67);
nand (n79,n80,n81);
not (n80,n65);
nor (n81,n82,n84);
and (n82,n83,n58);
and (n84,n85,n63);
not (n85,n83);
nor (n86,n87,n93);
nand (n87,n58,n88);
not (n88,n89);
wire s0n89,s1n89,notn89;
or (n89,s0n89,s1n89);
not(notn89,n4);
and (s0n89,notn89,1'b0);
and (s1n89,n4,n91);
and (n91,n92,n60);
nor (n93,n94,n96);
and (n94,n89,n95);
not (n95,n12);
and (n96,n88,n12);
nand (n97,n98,n116);
or (n98,n99,n111);
nand (n99,n100,n108);
not (n100,n101);
nand (n101,n102,n107);
or (n102,n103,n40);
not (n103,n104);
wire s0n104,s1n104,notn104;
or (n104,s0n104,s1n104);
not(notn104,n4);
and (s0n104,notn104,n105);
and (s1n104,n4,n106);
nand (n107,n40,n103);
nand (n108,n109,n110);
or (n109,n103,n71);
nand (n110,n71,n103);
nor (n111,n112,n114);
and (n112,n75,n113);
and (n114,n71,n115);
not (n115,n113);
or (n116,n100,n117);
nor (n117,n118,n120);
and (n118,n75,n119);
and (n120,n71,n121);
not (n121,n119);
xor (n122,n123,n179);
xor (n123,n124,n166);
xor (n124,n125,n142);
nand (n125,n126,n135);
or (n126,n127,n130);
not (n127,n128);
nor (n128,n129,n13);
not (n129,n18);
nor (n130,n131,n133);
and (n131,n129,n132);
and (n133,n18,n134);
not (n134,n132);
or (n135,n136,n141);
nor (n136,n137,n139);
and (n137,n129,n138);
and (n139,n18,n140);
not (n140,n138);
not (n141,n13);
nand (n142,n143,n160);
or (n143,n144,n154);
not (n144,n145);
and (n145,n146,n150);
nand (n146,n147,n149);
or (n147,n148,n40);
not (n148,n33);
nand (n149,n40,n148);
not (n150,n151);
nand (n151,n152,n153);
or (n152,n148,n18);
nand (n153,n18,n148);
nor (n154,n155,n158);
and (n155,n156,n157);
not (n156,n40);
and (n158,n40,n159);
not (n159,n157);
or (n160,n150,n161);
nor (n161,n162,n164);
and (n162,n156,n163);
and (n164,n40,n165);
not (n165,n163);
and (n166,n167,n173);
nand (n167,n168,n172);
or (n168,n127,n169);
nor (n169,n170,n171);
and (n170,n129,n163);
and (n171,n18,n165);
or (n172,n130,n141);
nand (n173,n174,n178);
or (n174,n144,n175);
nor (n175,n176,n177);
and (n176,n156,n119);
and (n177,n40,n121);
or (n178,n154,n150);
or (n179,n180,n200);
and (n180,n181,n194);
xor (n181,n182,n189);
nand (n182,n183,n188);
or (n183,n184,n64);
not (n184,n185);
nor (n185,n186,n187);
and (n186,n12,n58);
and (n187,n95,n63);
nand (n188,n80,n55);
nor (n189,n87,n190);
nor (n190,n191,n193);
and (n191,n89,n192);
not (n192,n17);
and (n193,n88,n17);
nand (n194,n195,n199);
or (n195,n99,n196);
nor (n196,n197,n198);
and (n197,n75,n83);
and (n198,n71,n85);
or (n199,n100,n111);
and (n200,n182,n189);
and (n201,n202,n203);
xor (n202,n167,n173);
or (n203,n204,n223);
and (n204,n205,n217);
xor (n205,n206,n212);
nand (n206,n207,n211);
or (n207,n208,n64);
nor (n208,n209,n210);
and (n209,n17,n63);
and (n210,n192,n58);
nand (n211,n185,n80);
nor (n212,n87,n213);
nor (n213,n214,n216);
and (n214,n89,n215);
not (n215,n25);
and (n216,n88,n25);
nand (n217,n218,n222);
or (n218,n127,n219);
nor (n219,n220,n221);
and (n220,n129,n157);
and (n221,n18,n159);
or (n222,n169,n141);
and (n223,n206,n212);
not (n224,n225);
or (n225,n226,n264);
and (n226,n227,n230);
xor (n227,n228,n229);
xor (n228,n181,n194);
xor (n229,n202,n203);
or (n230,n231,n263);
and (n231,n232,n245);
xor (n232,n233,n239);
nand (n233,n234,n238);
or (n234,n99,n235);
nor (n235,n236,n237);
and (n236,n75,n57);
and (n237,n71,n62);
or (n238,n100,n196);
nand (n239,n240,n244);
or (n240,n144,n241);
nor (n241,n242,n243);
and (n242,n156,n113);
and (n243,n40,n115);
or (n244,n175,n150);
or (n245,n246,n262);
and (n246,n247,n256);
xor (n247,n248,n250);
and (n248,n249,n31);
not (n249,n87);
nand (n250,n251,n255);
or (n251,n127,n252);
nor (n252,n253,n254);
and (n253,n121,n18);
and (n254,n119,n129);
or (n255,n219,n141);
nand (n256,n257,n261);
or (n257,n64,n258);
nor (n258,n259,n260);
and (n259,n25,n63);
and (n260,n215,n58);
or (n261,n65,n208);
and (n262,n248,n250);
and (n263,n233,n239);
and (n264,n228,n229);
nand (n265,n48,n225);
nand (n266,n267,n516);
or (n267,n268,n308);
nor (n268,n269,n270);
xor (n269,n227,n230);
or (n270,n271,n307);
and (n271,n272,n306);
xor (n272,n273,n274);
xor (n273,n205,n217);
or (n274,n275,n305);
and (n275,n276,n290);
xor (n276,n277,n284);
nand (n277,n278,n283);
or (n278,n144,n279);
not (n279,n280);
nor (n280,n281,n282);
and (n281,n83,n40);
and (n282,n85,n156);
or (n283,n150,n241);
nand (n284,n285,n289);
or (n285,n99,n286);
nor (n286,n287,n288);
and (n287,n75,n12);
and (n288,n71,n95);
or (n289,n100,n235);
and (n290,n291,n297);
nor (n291,n292,n63);
nor (n292,n293,n295);
and (n293,n75,n294);
nand (n294,n68,n31);
and (n295,n67,n296);
not (n296,n31);
nand (n297,n298,n303);
or (n298,n299,n127);
not (n299,n300);
nor (n300,n301,n302);
and (n301,n113,n18);
and (n302,n115,n129);
nand (n303,n304,n13);
not (n304,n252);
and (n305,n277,n284);
xor (n306,n232,n245);
and (n307,n273,n274);
not (n308,n309);
nand (n309,n310,n511);
not (n310,n311);
nor (n311,n312,n492);
nor (n312,n313,n490);
and (n313,n314,n464);
or (n314,n315,n463);
and (n315,n316,n380);
xor (n316,n317,n357);
or (n317,n318,n356);
and (n318,n319,n341);
xor (n319,n320,n330);
nand (n320,n321,n326);
or (n321,n322,n144);
not (n322,n323);
nor (n323,n324,n325);
and (n324,n192,n156);
and (n325,n17,n40);
nand (n326,n151,n327);
nor (n327,n328,n329);
and (n328,n12,n40);
and (n329,n156,n95);
nand (n330,n331,n336);
or (n331,n332,n100);
not (n332,n333);
nor (n333,n334,n335);
and (n334,n25,n71);
and (n335,n215,n75);
nand (n336,n337,n338);
not (n337,n99);
nand (n338,n339,n340);
or (n339,n75,n31);
or (n340,n71,n296);
xor (n341,n342,n347);
and (n342,n343,n71);
nand (n343,n344,n346);
or (n344,n40,n345);
and (n345,n31,n104);
or (n346,n104,n31);
nand (n347,n348,n352);
or (n348,n127,n349);
nor (n349,n350,n351);
and (n350,n129,n57);
and (n351,n18,n62);
or (n352,n353,n141);
nor (n353,n354,n355);
and (n354,n83,n129);
and (n355,n85,n18);
and (n356,n320,n330);
xor (n357,n358,n366);
xor (n358,n359,n365);
nand (n359,n360,n361);
or (n360,n332,n99);
or (n361,n100,n362);
nor (n362,n363,n364);
and (n363,n75,n17);
and (n364,n71,n192);
and (n365,n342,n347);
xor (n366,n367,n373);
xor (n367,n368,n369);
and (n368,n80,n31);
nand (n369,n370,n371);
or (n370,n141,n299);
nand (n371,n372,n128);
not (n372,n353);
nand (n373,n374,n376);
or (n374,n375,n144);
not (n375,n327);
nand (n376,n151,n377);
nand (n377,n378,n379);
or (n378,n40,n62);
or (n379,n156,n57);
or (n380,n381,n462);
and (n381,n382,n403);
xor (n382,n383,n402);
or (n383,n384,n401);
and (n384,n385,n394);
xor (n385,n386,n387);
and (n386,n101,n31);
nand (n387,n388,n393);
or (n388,n389,n144);
not (n389,n390);
nor (n390,n391,n392);
and (n391,n25,n40);
and (n392,n215,n156);
nand (n393,n323,n151);
nand (n394,n395,n400);
or (n395,n127,n396);
not (n396,n397);
nor (n397,n398,n399);
and (n398,n95,n129);
and (n399,n12,n18);
or (n400,n349,n141);
and (n401,n386,n387);
xor (n402,n319,n341);
or (n403,n404,n461);
and (n404,n405,n460);
xor (n405,n406,n419);
nor (n406,n407,n415);
not (n407,n408);
nand (n408,n409,n414);
or (n409,n410,n127);
not (n410,n411);
nand (n411,n412,n413);
or (n412,n192,n18);
nand (n413,n18,n192);
nand (n414,n397,n13);
nand (n415,n416,n40);
nand (n416,n417,n418);
or (n417,n18,n38);
or (n418,n33,n31);
nand (n419,n420,n458);
or (n420,n421,n444);
not (n421,n422);
nand (n422,n423,n443);
or (n423,n424,n433);
nor (n424,n425,n432);
nand (n425,n426,n431);
or (n426,n427,n127);
not (n427,n428);
nand (n428,n429,n430);
or (n429,n215,n18);
nand (n430,n18,n215);
nand (n431,n411,n13);
nor (n432,n150,n296);
nand (n433,n434,n441);
nand (n434,n435,n440);
or (n435,n436,n127);
not (n436,n437);
nand (n437,n438,n439);
or (n438,n129,n31);
or (n439,n18,n296);
nand (n440,n428,n13);
nor (n441,n442,n129);
and (n442,n31,n13);
nand (n443,n425,n432);
not (n444,n445);
nand (n445,n446,n454);
not (n446,n447);
nand (n447,n448,n453);
or (n448,n449,n144);
not (n449,n450);
nand (n450,n451,n452);
or (n451,n156,n31);
or (n452,n40,n296);
nand (n453,n151,n390);
nor (n454,n455,n457);
and (n455,n407,n456);
not (n456,n415);
and (n457,n408,n415);
nand (n458,n459,n447);
not (n459,n454);
xor (n460,n385,n394);
and (n461,n406,n419);
and (n462,n383,n402);
and (n463,n317,n357);
or (n464,n465,n487);
xor (n465,n466,n471);
xor (n466,n467,n468);
xor (n467,n291,n297);
or (n468,n469,n470);
and (n469,n367,n373);
and (n470,n368,n369);
xor (n471,n472,n484);
xor (n472,n473,n480);
nand (n473,n474,n479);
or (n474,n475,n64);
not (n475,n476);
nand (n476,n477,n478);
or (n477,n63,n31);
or (n478,n58,n296);
or (n479,n65,n258);
nand (n480,n481,n483);
or (n481,n482,n144);
not (n482,n377);
nand (n483,n151,n280);
nand (n484,n485,n486);
or (n485,n99,n362);
or (n486,n100,n286);
or (n487,n488,n489);
and (n488,n358,n366);
and (n489,n359,n365);
not (n490,n491);
nand (n491,n465,n487);
nand (n492,n493,n505);
not (n493,n494);
nor (n494,n495,n502);
xor (n495,n496,n501);
xor (n496,n497,n500);
or (n497,n498,n499);
and (n498,n472,n484);
and (n499,n473,n480);
xor (n500,n247,n256);
xor (n501,n276,n290);
or (n502,n503,n504);
and (n503,n466,n471);
and (n504,n467,n468);
not (n505,n506);
nor (n506,n507,n510);
or (n507,n508,n509);
and (n508,n496,n501);
and (n509,n497,n500);
xor (n510,n272,n306);
nor (n511,n512,n515);
and (n512,n505,n513);
not (n513,n514);
nand (n514,n495,n502);
and (n515,n507,n510);
nand (n516,n269,n270);
and (n518,n517,n519);
wire s0n519,s1n519,notn519;
or (n519,s0n519,s1n519);
not(notn519,n4);
and (s0n519,notn519,n520);
and (s1n519,n4,n6);
xor (n520,n521,n807);
xor (n521,n522,n815);
xor (n522,n523,n802);
xor (n523,n524,n808);
xor (n524,n525,n796);
xor (n525,n526,n793);
xor (n526,n527,n792);
xor (n527,n528,n772);
xor (n528,n529,n56);
xor (n529,n530,n745);
xor (n530,n531,n744);
xor (n531,n532,n712);
xor (n532,n533,n711);
xor (n533,n534,n673);
xor (n534,n535,n672);
xor (n535,n536,n633);
xor (n536,n537,n632);
xor (n537,n538,n587);
xor (n538,n539,n586);
xor (n539,n540,n543);
xor (n540,n541,n542);
and (n541,n138,n13);
and (n542,n132,n18);
or (n543,n544,n547);
and (n544,n545,n546);
and (n545,n132,n13);
and (n546,n163,n18);
and (n547,n548,n549);
xor (n548,n545,n546);
or (n549,n550,n553);
and (n550,n551,n552);
and (n551,n163,n13);
and (n552,n157,n18);
and (n553,n554,n555);
xor (n554,n551,n552);
or (n555,n556,n559);
and (n556,n557,n558);
and (n557,n157,n13);
and (n558,n119,n18);
and (n559,n560,n561);
xor (n560,n557,n558);
or (n561,n562,n564);
and (n562,n563,n301);
and (n563,n119,n13);
and (n564,n565,n566);
xor (n565,n563,n301);
or (n566,n567,n570);
and (n567,n568,n569);
and (n568,n113,n13);
and (n569,n83,n18);
and (n570,n571,n572);
xor (n571,n568,n569);
or (n572,n573,n576);
and (n573,n574,n575);
and (n574,n83,n13);
and (n575,n57,n18);
and (n576,n577,n578);
xor (n577,n574,n575);
or (n578,n579,n581);
and (n579,n580,n399);
and (n580,n57,n13);
and (n581,n582,n583);
xor (n582,n580,n399);
or (n583,n584,n585);
and (n584,n11,n16);
and (n585,n10,n21);
and (n586,n163,n33);
or (n587,n588,n591);
and (n588,n589,n590);
xor (n589,n548,n549);
and (n590,n157,n33);
and (n591,n592,n593);
xor (n592,n589,n590);
or (n593,n594,n597);
and (n594,n595,n596);
xor (n595,n554,n555);
and (n596,n119,n33);
and (n597,n598,n599);
xor (n598,n595,n596);
or (n599,n600,n603);
and (n600,n601,n602);
xor (n601,n560,n561);
and (n602,n113,n33);
and (n603,n604,n605);
xor (n604,n601,n602);
or (n605,n606,n609);
and (n606,n607,n608);
xor (n607,n565,n566);
and (n608,n83,n33);
and (n609,n610,n611);
xor (n610,n607,n608);
or (n611,n612,n615);
and (n612,n613,n614);
xor (n613,n571,n572);
and (n614,n57,n33);
and (n615,n616,n617);
xor (n616,n613,n614);
or (n617,n618,n621);
and (n618,n619,n620);
xor (n619,n577,n578);
and (n620,n12,n33);
and (n621,n622,n623);
xor (n622,n619,n620);
or (n623,n624,n627);
and (n624,n625,n626);
xor (n625,n582,n583);
and (n626,n17,n33);
and (n627,n628,n629);
xor (n628,n625,n626);
or (n629,n630,n631);
and (n630,n9,n32);
and (n631,n8,n36);
and (n632,n157,n40);
or (n633,n634,n637);
and (n634,n635,n636);
xor (n635,n592,n593);
and (n636,n119,n40);
and (n637,n638,n639);
xor (n638,n635,n636);
or (n639,n640,n643);
and (n640,n641,n642);
xor (n641,n598,n599);
and (n642,n113,n40);
and (n643,n644,n645);
xor (n644,n641,n642);
or (n645,n646,n648);
and (n646,n647,n281);
xor (n647,n604,n605);
and (n648,n649,n650);
xor (n649,n647,n281);
or (n650,n651,n654);
and (n651,n652,n653);
xor (n652,n610,n611);
and (n653,n57,n40);
and (n654,n655,n656);
xor (n655,n652,n653);
or (n656,n657,n659);
and (n657,n658,n328);
xor (n658,n616,n617);
and (n659,n660,n661);
xor (n660,n658,n328);
or (n661,n662,n664);
and (n662,n663,n325);
xor (n663,n622,n623);
and (n664,n665,n666);
xor (n665,n663,n325);
or (n666,n667,n669);
and (n667,n668,n391);
xor (n668,n628,n629);
and (n669,n670,n671);
xor (n670,n668,n391);
and (n671,n7,n39);
and (n672,n119,n104);
or (n673,n674,n677);
and (n674,n675,n676);
xor (n675,n638,n639);
and (n676,n113,n104);
and (n677,n678,n679);
xor (n678,n675,n676);
or (n679,n680,n683);
and (n680,n681,n682);
xor (n681,n644,n645);
and (n682,n83,n104);
and (n683,n684,n685);
xor (n684,n681,n682);
or (n685,n686,n689);
and (n686,n687,n688);
xor (n687,n649,n650);
and (n688,n57,n104);
and (n689,n690,n691);
xor (n690,n687,n688);
or (n691,n692,n695);
and (n692,n693,n694);
xor (n693,n655,n656);
and (n694,n12,n104);
and (n695,n696,n697);
xor (n696,n693,n694);
or (n697,n698,n701);
and (n698,n699,n700);
xor (n699,n660,n661);
and (n700,n17,n104);
and (n701,n702,n703);
xor (n702,n699,n700);
or (n703,n704,n707);
and (n704,n705,n706);
xor (n705,n665,n666);
and (n706,n25,n104);
and (n707,n708,n709);
xor (n708,n705,n706);
and (n709,n710,n345);
xor (n710,n670,n671);
and (n711,n113,n71);
or (n712,n713,n716);
and (n713,n714,n715);
xor (n714,n678,n679);
and (n715,n83,n71);
and (n716,n717,n718);
xor (n717,n714,n715);
or (n718,n719,n722);
and (n719,n720,n721);
xor (n720,n684,n685);
and (n721,n57,n71);
and (n722,n723,n724);
xor (n723,n720,n721);
or (n724,n725,n728);
and (n725,n726,n727);
xor (n726,n690,n691);
and (n727,n12,n71);
and (n728,n729,n730);
xor (n729,n726,n727);
or (n730,n731,n734);
and (n731,n732,n733);
xor (n732,n696,n697);
and (n733,n17,n71);
and (n734,n735,n736);
xor (n735,n732,n733);
or (n736,n737,n739);
and (n737,n738,n334);
xor (n738,n702,n703);
and (n739,n740,n741);
xor (n740,n738,n334);
and (n741,n742,n743);
xor (n742,n708,n709);
and (n743,n31,n71);
and (n744,n83,n68);
or (n745,n746,n749);
and (n746,n747,n748);
xor (n747,n717,n718);
and (n748,n57,n68);
and (n749,n750,n751);
xor (n750,n747,n748);
or (n751,n752,n755);
and (n752,n753,n754);
xor (n753,n723,n724);
and (n754,n12,n68);
and (n755,n756,n757);
xor (n756,n753,n754);
or (n757,n758,n761);
and (n758,n759,n760);
xor (n759,n729,n730);
and (n760,n17,n68);
and (n761,n762,n763);
xor (n762,n759,n760);
or (n763,n764,n767);
and (n764,n765,n766);
xor (n765,n735,n736);
and (n766,n25,n68);
and (n767,n768,n769);
xor (n768,n765,n766);
and (n769,n770,n771);
xor (n770,n740,n741);
not (n771,n294);
or (n772,n773,n775);
and (n773,n774,n186);
xor (n774,n750,n751);
and (n775,n776,n777);
xor (n776,n774,n186);
or (n777,n778,n781);
and (n778,n779,n780);
xor (n779,n756,n757);
and (n780,n17,n58);
and (n781,n782,n783);
xor (n782,n779,n780);
or (n783,n784,n787);
and (n784,n785,n786);
xor (n785,n762,n763);
and (n786,n25,n58);
and (n787,n788,n789);
xor (n788,n785,n786);
and (n789,n790,n791);
xor (n790,n768,n769);
and (n791,n31,n58);
and (n792,n12,n89);
or (n793,n794,n797);
and (n794,n795,n796);
xor (n795,n776,n777);
and (n796,n17,n89);
and (n797,n798,n799);
xor (n798,n795,n796);
or (n799,n800,n803);
and (n800,n801,n802);
xor (n801,n782,n783);
and (n802,n25,n89);
and (n803,n804,n805);
xor (n804,n801,n802);
and (n805,n806,n807);
xor (n806,n788,n789);
and (n807,n31,n89);
or (n808,n809,n811);
and (n809,n810,n802);
xor (n810,n798,n799);
and (n811,n812,n813);
xor (n812,n810,n802);
and (n813,n814,n807);
xor (n814,n804,n805);
and (n815,n816,n807);
xor (n816,n812,n813);
endmodule
