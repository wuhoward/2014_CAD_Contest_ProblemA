module top (out,n3,n4,n5,n23,n24,n28,n34,n39,n49
        ,n50,n55,n60,n67,n85,n92,n93,n102,n124,n126
        ,n132,n141,n158,n168,n178,n182,n189,n215,n297,n311);
output out;
input n3;
input n4;
input n5;
input n23;
input n24;
input n28;
input n34;
input n39;
input n49;
input n50;
input n55;
input n60;
input n67;
input n85;
input n92;
input n93;
input n102;
input n124;
input n126;
input n132;
input n141;
input n158;
input n168;
input n178;
input n182;
input n189;
input n215;
input n297;
input n311;
wire n0;
wire n1;
wire n2;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n25;
wire n26;
wire n27;
wire n29;
wire n30;
wire n31;
wire n32;
wire n33;
wire n35;
wire n36;
wire n37;
wire n38;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n51;
wire n52;
wire n53;
wire n54;
wire n56;
wire n57;
wire n58;
wire n59;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n125;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n179;
wire n180;
wire n181;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
xnor (out,n0,n628);
nor (n0,n1,n6);
and (n1,n2,n5);
nor (n2,n3,n4);
and (n6,n7,n625);
nor (n7,n8,n623);
and (n8,n9,n331);
nand (n9,n10,n330);
or (n10,n11,n262);
or (n11,n12,n261);
and (n12,n13,n218);
xor (n13,n14,n106);
xor (n14,n15,n70);
xor (n15,n16,n42);
nand (n16,n17,n36);
or (n17,n18,n31);
nand (n18,n19,n26);
not (n19,n20);
nand (n20,n21,n25);
or (n21,n22,n24);
not (n22,n23);
nand (n25,n24,n22);
nand (n26,n27,n29);
nand (n27,n22,n28);
nand (n29,n23,n30);
not (n30,n28);
nor (n31,n32,n35);
and (n32,n33,n28);
not (n33,n34);
and (n35,n34,n30);
or (n36,n19,n37);
nor (n37,n38,n40);
and (n38,n30,n39);
and (n40,n28,n41);
not (n41,n39);
nand (n42,n43,n63);
or (n43,n44,n58);
not (n44,n45);
nor (n45,n46,n52);
nand (n46,n47,n51);
or (n47,n48,n50);
not (n48,n49);
nand (n51,n50,n48);
nor (n52,n53,n56);
and (n53,n54,n55);
not (n54,n50);
and (n56,n50,n57);
not (n57,n55);
nor (n58,n59,n61);
and (n59,n57,n60);
and (n61,n55,n62);
not (n62,n60);
or (n63,n64,n65);
not (n64,n46);
nor (n65,n66,n68);
and (n66,n57,n67);
and (n68,n55,n69);
not (n69,n67);
nand (n70,n71,n105);
or (n71,n72,n80);
not (n72,n73);
nand (n73,n74,n28);
nand (n74,n75,n76);
or (n75,n34,n23);
nand (n76,n77,n79);
not (n77,n78);
and (n78,n34,n23);
not (n79,n24);
not (n80,n81);
nand (n81,n82,n95);
or (n82,n83,n88);
nor (n83,n84,n86);
and (n84,n85,n48);
and (n86,n87,n49);
not (n87,n85);
not (n88,n89);
nand (n89,n90,n94);
or (n90,n91,n93);
not (n91,n92);
nand (n94,n91,n93);
or (n95,n96,n100);
nand (n96,n88,n97);
nand (n97,n98,n99);
or (n98,n49,n91);
nand (n99,n91,n49);
nor (n100,n101,n103);
and (n101,n102,n48);
and (n103,n104,n49);
not (n104,n102);
or (n105,n81,n73);
xor (n106,n107,n194);
xor (n107,n108,n145);
or (n108,n109,n144);
and (n109,n110,n119);
xor (n110,n111,n112);
nor (n111,n19,n33);
nand (n112,n113,n117);
or (n113,n114,n96);
nor (n114,n115,n116);
and (n115,n48,n67);
and (n116,n49,n69);
nand (n117,n118,n89);
not (n118,n100);
nand (n119,n120,n134);
or (n120,n121,n129);
not (n121,n122);
nand (n122,n123,n127);
or (n123,n124,n125);
not (n125,n126);
or (n127,n128,n126);
not (n128,n124);
not (n129,n130);
nand (n130,n131,n133);
or (n131,n57,n132);
nand (n133,n132,n57);
or (n134,n135,n139);
nand (n135,n136,n129);
nand (n136,n137,n138);
or (n137,n132,n128);
nand (n138,n128,n132);
nor (n139,n140,n142);
and (n140,n128,n141);
and (n142,n124,n143);
not (n143,n141);
and (n144,n111,n112);
or (n145,n146,n193);
and (n146,n147,n185);
xor (n147,n148,n170);
nand (n148,n149,n164);
or (n149,n150,n154);
not (n150,n151);
nand (n151,n152,n153);
or (n152,n24,n41);
or (n153,n79,n39);
not (n154,n155);
nor (n155,n156,n161);
nor (n156,n157,n159);
and (n157,n158,n79);
and (n159,n24,n160);
not (n160,n158);
nand (n161,n162,n163);
or (n162,n128,n158);
nand (n163,n158,n128);
nand (n164,n161,n165);
nand (n165,n166,n169);
or (n166,n24,n167);
not (n167,n168);
or (n169,n79,n168);
nand (n170,n171,n179);
or (n171,n172,n176);
nor (n172,n173,n175);
and (n173,n174,n85);
not (n174,n93);
and (n175,n93,n87);
nand (n176,n177,n93);
not (n177,n178);
or (n179,n180,n177);
nor (n180,n181,n183);
and (n181,n174,n182);
and (n183,n93,n184);
not (n184,n182);
nand (n185,n186,n192);
or (n186,n44,n187);
nor (n187,n188,n190);
and (n188,n57,n189);
and (n190,n55,n191);
not (n191,n189);
or (n192,n64,n58);
and (n193,n148,n170);
xor (n194,n195,n209);
xor (n195,n196,n202);
nand (n196,n197,n198);
or (n197,n121,n135);
nand (n198,n130,n199);
nor (n199,n200,n201);
and (n200,n191,n128);
and (n201,n189,n124);
nand (n202,n203,n205);
or (n203,n204,n154);
not (n204,n165);
nand (n205,n161,n206);
nand (n206,n207,n208);
or (n207,n24,n143);
or (n208,n141,n79);
nand (n209,n210,n217);
or (n210,n177,n211);
not (n211,n212);
nor (n212,n213,n216);
and (n213,n214,n174);
not (n214,n215);
and (n216,n215,n93);
or (n217,n180,n176);
or (n218,n219,n260);
and (n219,n220,n259);
xor (n220,n221,n234);
and (n221,n222,n228);
and (n222,n223,n24);
nand (n223,n224,n225);
or (n224,n34,n158);
nand (n225,n226,n128);
not (n226,n227);
and (n227,n34,n158);
nand (n228,n229,n233);
or (n229,n96,n230);
nor (n230,n231,n232);
and (n231,n48,n60);
and (n232,n49,n62);
or (n233,n88,n114);
or (n234,n235,n258);
and (n235,n236,n252);
xor (n236,n237,n244);
nand (n237,n238,n242);
or (n238,n239,n135);
nor (n239,n240,n241);
and (n240,n128,n168);
and (n241,n124,n167);
nand (n242,n243,n130);
not (n243,n139);
nand (n244,n245,n247);
or (n245,n150,n246);
not (n246,n161);
nand (n247,n248,n155);
not (n248,n249);
nor (n249,n250,n251);
and (n250,n33,n24);
and (n251,n79,n34);
nand (n252,n253,n257);
or (n253,n176,n254);
nor (n254,n255,n256);
and (n255,n174,n102);
and (n256,n93,n104);
or (n257,n172,n177);
and (n258,n237,n244);
xor (n259,n110,n119);
and (n260,n221,n234);
and (n261,n14,n106);
xor (n262,n263,n279);
xor (n263,n264,n276);
xor (n264,n265,n273);
xor (n265,n266,n272);
nand (n266,n267,n268);
or (n267,n44,n65);
or (n268,n64,n269);
nor (n269,n270,n271);
and (n270,n57,n102);
and (n271,n55,n104);
and (n272,n81,n72);
or (n273,n274,n275);
and (n274,n195,n209);
and (n275,n196,n202);
or (n276,n277,n278);
and (n277,n107,n194);
and (n278,n108,n145);
xor (n279,n280,n327);
xor (n280,n281,n305);
xor (n281,n282,n299);
xor (n282,n283,n291);
nand (n283,n284,n286);
or (n284,n285,n154);
not (n285,n206);
nand (n286,n287,n161);
not (n287,n288);
nor (n288,n289,n290);
and (n289,n79,n126);
and (n290,n125,n24);
nand (n291,n292,n293);
or (n292,n176,n211);
nand (n293,n294,n178);
nor (n294,n295,n298);
and (n295,n296,n174);
not (n296,n297);
and (n298,n297,n93);
nand (n299,n300,n301);
or (n300,n18,n37);
or (n301,n19,n302);
nor (n302,n303,n304);
and (n303,n30,n168);
and (n304,n28,n167);
xor (n305,n306,n320);
xor (n306,n307,n313);
nor (n307,n308,n33);
nor (n308,n309,n312);
and (n309,n310,n28);
not (n310,n311);
and (n312,n311,n30);
nand (n313,n314,n315);
or (n314,n96,n83);
nand (n315,n316,n89);
not (n316,n317);
nor (n317,n318,n319);
and (n318,n182,n48);
and (n319,n184,n49);
nand (n320,n321,n323);
or (n321,n135,n322);
not (n322,n199);
or (n323,n129,n324);
nor (n324,n325,n326);
and (n325,n62,n124);
and (n326,n60,n128);
or (n327,n328,n329);
and (n328,n15,n70);
and (n329,n16,n42);
nand (n330,n11,n262);
not (n331,n332);
nand (n332,n333,n622);
or (n333,n334,n371);
not (n334,n335);
or (n335,n336,n337);
xor (n336,n13,n218);
or (n337,n338,n370);
and (n338,n339,n369);
xor (n339,n340,n341);
xor (n340,n147,n185);
or (n341,n342,n368);
and (n342,n343,n351);
xor (n343,n344,n350);
nand (n344,n345,n349);
or (n345,n44,n346);
nor (n346,n347,n348);
and (n347,n57,n126);
and (n348,n55,n125);
or (n349,n64,n187);
xor (n350,n222,n228);
or (n351,n352,n367);
and (n352,n353,n361);
xor (n353,n354,n355);
nor (n354,n246,n33);
nand (n355,n356,n360);
or (n356,n357,n176);
nor (n357,n358,n359);
and (n358,n69,n93);
and (n359,n67,n174);
or (n360,n254,n177);
nand (n361,n362,n366);
or (n362,n135,n363);
nor (n363,n364,n365);
and (n364,n128,n39);
and (n365,n124,n41);
or (n366,n129,n239);
and (n367,n354,n355);
and (n368,n344,n350);
xor (n369,n220,n259);
and (n370,n340,n341);
not (n371,n372);
or (n372,n373,n621);
and (n373,n374,n414);
xor (n374,n375,n413);
or (n375,n376,n412);
and (n376,n377,n411);
xor (n377,n378,n379);
xor (n378,n236,n252);
or (n379,n380,n410);
and (n380,n381,n396);
xor (n381,n382,n390);
nand (n382,n383,n388);
or (n383,n384,n96);
not (n384,n385);
nand (n385,n386,n387);
or (n386,n49,n191);
or (n387,n48,n189);
nand (n388,n389,n89);
not (n389,n230);
nand (n390,n391,n395);
or (n391,n44,n392);
nor (n392,n393,n394);
and (n393,n57,n141);
and (n394,n55,n143);
or (n395,n64,n346);
and (n396,n397,n403);
nor (n397,n398,n128);
nor (n398,n399,n401);
and (n399,n33,n400);
not (n400,n132);
nor (n401,n402,n55);
and (n402,n34,n132);
nand (n403,n404,n409);
or (n404,n176,n405);
not (n405,n406);
nor (n406,n407,n408);
and (n407,n62,n174);
and (n408,n60,n93);
or (n409,n357,n177);
and (n410,n382,n390);
xor (n411,n343,n351);
and (n412,n378,n379);
xor (n413,n339,n369);
nand (n414,n415,n618,n620);
nand (n415,n416,n451,n611);
nand (n416,n417,n419);
not (n417,n418);
xor (n418,n377,n411);
not (n419,n420);
or (n420,n421,n450);
and (n421,n422,n449);
xor (n422,n423,n448);
or (n423,n424,n447);
and (n424,n425,n441);
xor (n425,n426,n434);
nand (n426,n427,n432);
or (n427,n428,n135);
not (n428,n429);
nand (n429,n430,n431);
or (n430,n128,n34);
or (n431,n33,n124);
nand (n432,n433,n130);
not (n433,n363);
nand (n434,n435,n440);
or (n435,n436,n96);
not (n436,n437);
nand (n437,n438,n439);
or (n438,n49,n125);
or (n439,n48,n126);
nand (n440,n89,n385);
nand (n441,n442,n446);
or (n442,n44,n443);
nor (n443,n444,n445);
and (n444,n57,n168);
and (n445,n55,n167);
or (n446,n64,n392);
and (n447,n426,n434);
xor (n448,n353,n361);
xor (n449,n381,n396);
and (n450,n423,n448);
nand (n451,n452,n610);
or (n452,n453,n503);
not (n453,n454);
nand (n454,n455,n479);
not (n455,n456);
xor (n456,n457,n478);
xor (n457,n458,n459);
xor (n458,n397,n403);
or (n459,n460,n477);
and (n460,n461,n470);
xor (n461,n462,n463);
and (n462,n130,n34);
nand (n463,n464,n469);
or (n464,n176,n465);
not (n465,n466);
nor (n466,n467,n468);
and (n467,n191,n174);
and (n468,n189,n93);
nand (n469,n406,n178);
nand (n470,n471,n476);
or (n471,n472,n96);
not (n472,n473);
nor (n473,n474,n475);
and (n474,n143,n48);
and (n475,n141,n49);
nand (n476,n89,n437);
and (n477,n462,n463);
xor (n478,n425,n441);
not (n479,n480);
or (n480,n481,n502);
and (n481,n482,n501);
xor (n482,n483,n489);
nand (n483,n484,n488);
or (n484,n44,n485);
nor (n485,n486,n487);
and (n486,n41,n55);
and (n487,n39,n57);
or (n488,n64,n443);
and (n489,n490,n495);
and (n490,n491,n55);
nand (n491,n492,n494);
or (n492,n493,n49);
and (n493,n34,n50);
or (n494,n34,n50);
nand (n495,n496,n497);
or (n496,n177,n465);
or (n497,n498,n176);
nor (n498,n499,n500);
and (n499,n174,n126);
and (n500,n93,n125);
xor (n501,n461,n470);
and (n502,n483,n489);
not (n503,n504);
nand (n504,n505,n609);
or (n505,n506,n529);
not (n506,n507);
nand (n507,n508,n510);
not (n508,n509);
xor (n509,n482,n501);
not (n510,n511);
or (n511,n512,n528);
and (n512,n513,n527);
xor (n513,n514,n521);
nand (n514,n515,n520);
or (n515,n516,n96);
not (n516,n517);
nor (n517,n518,n519);
and (n518,n167,n48);
and (n519,n168,n49);
nand (n520,n473,n89);
nand (n521,n522,n523);
or (n522,n64,n485);
nand (n523,n45,n524);
nand (n524,n525,n526);
or (n525,n34,n57);
or (n526,n33,n55);
xor (n527,n490,n495);
and (n528,n514,n521);
not (n529,n530);
or (n530,n531,n608);
and (n531,n532,n553);
xor (n532,n533,n552);
or (n533,n534,n551);
and (n534,n535,n544);
xor (n535,n536,n537);
and (n536,n46,n34);
nand (n537,n538,n543);
or (n538,n539,n96);
not (n539,n540);
nor (n540,n541,n542);
and (n541,n41,n48);
and (n542,n39,n49);
nand (n543,n517,n89);
nand (n544,n545,n550);
or (n545,n176,n546);
not (n546,n547);
nor (n547,n548,n549);
and (n548,n143,n174);
and (n549,n141,n93);
or (n550,n498,n177);
and (n551,n536,n537);
xor (n552,n513,n527);
nand (n553,n554,n607);
or (n554,n555,n571);
nor (n555,n556,n557);
xor (n556,n535,n544);
nor (n557,n558,n566);
not (n558,n559);
nand (n559,n560,n561);
or (n560,n177,n546);
nand (n561,n562,n565);
nand (n562,n563,n564);
or (n563,n168,n174);
nand (n564,n174,n168);
not (n565,n176);
nand (n566,n567,n49);
nand (n567,n568,n570);
or (n568,n569,n93);
and (n569,n34,n92);
or (n570,n34,n92);
nor (n571,n572,n606);
and (n572,n573,n585);
nand (n573,n574,n581);
not (n574,n575);
nand (n575,n576,n580);
or (n576,n96,n577);
nor (n577,n578,n579);
and (n578,n49,n33);
and (n579,n34,n48);
or (n580,n88,n539);
nor (n581,n582,n583);
and (n582,n566,n559);
and (n583,n584,n558);
not (n584,n566);
or (n585,n586,n605);
and (n586,n587,n596);
xor (n587,n588,n589);
nor (n588,n88,n33);
nand (n589,n590,n595);
or (n590,n176,n591);
not (n591,n592);
nand (n592,n593,n594);
or (n593,n41,n93);
nand (n594,n93,n41);
nand (n595,n562,n178);
nor (n596,n597,n603);
nor (n597,n598,n599);
and (n598,n592,n178);
nor (n599,n600,n176);
nor (n600,n601,n602);
and (n601,n33,n93);
and (n602,n34,n174);
or (n603,n604,n174);
and (n604,n34,n178);
and (n605,n588,n589);
nor (n606,n574,n581);
nand (n607,n556,n557);
and (n608,n533,n552);
nand (n609,n509,n511);
nand (n610,n456,n480);
nand (n611,n612,n616);
not (n612,n613);
or (n613,n614,n615);
and (n614,n457,n478);
and (n615,n458,n459);
not (n616,n617);
xor (n617,n422,n449);
nand (n618,n416,n619);
and (n619,n617,n613);
nand (n620,n420,n418);
and (n621,n375,n413);
nand (n622,n336,n337);
and (n623,n624,n332);
not (n624,n9);
not (n625,n626);
nand (n626,n627,n3);
not (n627,n4);
wire s0n628,s1n628,notn628;
or (n628,s0n628,s1n628);
not(notn628,n4);
and (s0n628,notn628,n629);
and (s1n628,n4,1'b0);
wire s0n629,s1n629,notn629;
or (n629,s0n629,s1n629);
not(notn629,n3);
and (s0n629,notn629,n5);
and (s1n629,n3,n630);
xor (n630,n631,n1015);
xor (n631,n632,n1012);
xor (n632,n633,n1011);
xor (n633,n634,n1003);
xor (n634,n635,n1002);
xor (n635,n636,n987);
xor (n636,n637,n986);
xor (n637,n638,n966);
xor (n638,n639,n965);
xor (n639,n640,n938);
xor (n640,n641,n201);
xor (n641,n642,n906);
xor (n642,n643,n905);
xor (n643,n644,n866);
xor (n644,n645,n865);
xor (n645,n646,n821);
xor (n646,n647,n820);
xor (n647,n648,n772);
xor (n648,n649,n771);
xor (n649,n650,n715);
xor (n650,n651,n714);
xor (n651,n652,n654);
xor (n652,n653,n216);
and (n653,n297,n178);
or (n654,n655,n658);
and (n655,n656,n657);
and (n656,n215,n178);
and (n657,n182,n93);
and (n658,n659,n660);
xor (n659,n656,n657);
or (n660,n661,n664);
and (n661,n662,n663);
and (n662,n182,n178);
and (n663,n85,n93);
and (n664,n665,n666);
xor (n665,n662,n663);
or (n666,n667,n670);
and (n667,n668,n669);
and (n668,n85,n178);
and (n669,n102,n93);
and (n670,n671,n672);
xor (n671,n668,n669);
or (n672,n673,n676);
and (n673,n674,n675);
and (n674,n102,n178);
and (n675,n67,n93);
and (n676,n677,n678);
xor (n677,n674,n675);
or (n678,n679,n681);
and (n679,n680,n408);
and (n680,n67,n178);
and (n681,n682,n683);
xor (n682,n680,n408);
or (n683,n684,n686);
and (n684,n685,n468);
and (n685,n60,n178);
and (n686,n687,n688);
xor (n687,n685,n468);
or (n688,n689,n692);
and (n689,n690,n691);
and (n690,n189,n178);
and (n691,n126,n93);
and (n692,n693,n694);
xor (n693,n690,n691);
or (n694,n695,n697);
and (n695,n696,n549);
and (n696,n126,n178);
and (n697,n698,n699);
xor (n698,n696,n549);
or (n699,n700,n703);
and (n700,n701,n702);
and (n701,n141,n178);
and (n702,n168,n93);
and (n703,n704,n705);
xor (n704,n701,n702);
or (n705,n706,n709);
and (n706,n707,n708);
and (n707,n168,n178);
and (n708,n39,n93);
and (n709,n710,n711);
xor (n710,n707,n708);
and (n711,n712,n713);
and (n712,n39,n178);
and (n713,n34,n93);
and (n714,n182,n92);
or (n715,n716,n719);
and (n716,n717,n718);
xor (n717,n659,n660);
and (n718,n85,n92);
and (n719,n720,n721);
xor (n720,n717,n718);
or (n721,n722,n725);
and (n722,n723,n724);
xor (n723,n665,n666);
and (n724,n102,n92);
and (n725,n726,n727);
xor (n726,n723,n724);
or (n727,n728,n731);
and (n728,n729,n730);
xor (n729,n671,n672);
and (n730,n67,n92);
and (n731,n732,n733);
xor (n732,n729,n730);
or (n733,n734,n737);
and (n734,n735,n736);
xor (n735,n677,n678);
and (n736,n60,n92);
and (n737,n738,n739);
xor (n738,n735,n736);
or (n739,n740,n743);
and (n740,n741,n742);
xor (n741,n682,n683);
and (n742,n189,n92);
and (n743,n744,n745);
xor (n744,n741,n742);
or (n745,n746,n749);
and (n746,n747,n748);
xor (n747,n687,n688);
and (n748,n126,n92);
and (n749,n750,n751);
xor (n750,n747,n748);
or (n751,n752,n755);
and (n752,n753,n754);
xor (n753,n693,n694);
and (n754,n141,n92);
and (n755,n756,n757);
xor (n756,n753,n754);
or (n757,n758,n761);
and (n758,n759,n760);
xor (n759,n698,n699);
and (n760,n168,n92);
and (n761,n762,n763);
xor (n762,n759,n760);
or (n763,n764,n767);
and (n764,n765,n766);
xor (n765,n704,n705);
and (n766,n39,n92);
and (n767,n768,n769);
xor (n768,n765,n766);
and (n769,n770,n569);
xor (n770,n710,n711);
and (n771,n85,n49);
or (n772,n773,n776);
and (n773,n774,n775);
xor (n774,n720,n721);
and (n775,n102,n49);
and (n776,n777,n778);
xor (n777,n774,n775);
or (n778,n779,n782);
and (n779,n780,n781);
xor (n780,n726,n727);
and (n781,n67,n49);
and (n782,n783,n784);
xor (n783,n780,n781);
or (n784,n785,n788);
and (n785,n786,n787);
xor (n786,n732,n733);
and (n787,n60,n49);
and (n788,n789,n790);
xor (n789,n786,n787);
or (n790,n791,n794);
and (n791,n792,n793);
xor (n792,n738,n739);
and (n793,n189,n49);
and (n794,n795,n796);
xor (n795,n792,n793);
or (n796,n797,n800);
and (n797,n798,n799);
xor (n798,n744,n745);
and (n799,n126,n49);
and (n800,n801,n802);
xor (n801,n798,n799);
or (n802,n803,n805);
and (n803,n804,n475);
xor (n804,n750,n751);
and (n805,n806,n807);
xor (n806,n804,n475);
or (n807,n808,n810);
and (n808,n809,n519);
xor (n809,n756,n757);
and (n810,n811,n812);
xor (n811,n809,n519);
or (n812,n813,n815);
and (n813,n814,n542);
xor (n814,n762,n763);
and (n815,n816,n817);
xor (n816,n814,n542);
and (n817,n818,n819);
xor (n818,n768,n769);
and (n819,n34,n49);
and (n820,n102,n50);
or (n821,n822,n825);
and (n822,n823,n824);
xor (n823,n777,n778);
and (n824,n67,n50);
and (n825,n826,n827);
xor (n826,n823,n824);
or (n827,n828,n831);
and (n828,n829,n830);
xor (n829,n783,n784);
and (n830,n60,n50);
and (n831,n832,n833);
xor (n832,n829,n830);
or (n833,n834,n837);
and (n834,n835,n836);
xor (n835,n789,n790);
and (n836,n189,n50);
and (n837,n838,n839);
xor (n838,n835,n836);
or (n839,n840,n843);
and (n840,n841,n842);
xor (n841,n795,n796);
and (n842,n126,n50);
and (n843,n844,n845);
xor (n844,n841,n842);
or (n845,n846,n849);
and (n846,n847,n848);
xor (n847,n801,n802);
and (n848,n141,n50);
and (n849,n850,n851);
xor (n850,n847,n848);
or (n851,n852,n855);
and (n852,n853,n854);
xor (n853,n806,n807);
and (n854,n168,n50);
and (n855,n856,n857);
xor (n856,n853,n854);
or (n857,n858,n861);
and (n858,n859,n860);
xor (n859,n811,n812);
and (n860,n39,n50);
and (n861,n862,n863);
xor (n862,n859,n860);
and (n863,n864,n493);
xor (n864,n816,n817);
and (n865,n67,n55);
or (n866,n867,n870);
and (n867,n868,n869);
xor (n868,n826,n827);
and (n869,n60,n55);
and (n870,n871,n872);
xor (n871,n868,n869);
or (n872,n873,n876);
and (n873,n874,n875);
xor (n874,n832,n833);
and (n875,n189,n55);
and (n876,n877,n878);
xor (n877,n874,n875);
or (n878,n879,n882);
and (n879,n880,n881);
xor (n880,n838,n839);
and (n881,n126,n55);
and (n882,n883,n884);
xor (n883,n880,n881);
or (n884,n885,n888);
and (n885,n886,n887);
xor (n886,n844,n845);
and (n887,n141,n55);
and (n888,n889,n890);
xor (n889,n886,n887);
or (n890,n891,n894);
and (n891,n892,n893);
xor (n892,n850,n851);
and (n893,n168,n55);
and (n894,n895,n896);
xor (n895,n892,n893);
or (n896,n897,n900);
and (n897,n898,n899);
xor (n898,n856,n857);
and (n899,n39,n55);
and (n900,n901,n902);
xor (n901,n898,n899);
and (n902,n903,n904);
xor (n903,n862,n863);
and (n904,n34,n55);
and (n905,n60,n132);
or (n906,n907,n910);
and (n907,n908,n909);
xor (n908,n871,n872);
and (n909,n189,n132);
and (n910,n911,n912);
xor (n911,n908,n909);
or (n912,n913,n916);
and (n913,n914,n915);
xor (n914,n877,n878);
and (n915,n126,n132);
and (n916,n917,n918);
xor (n917,n914,n915);
or (n918,n919,n922);
and (n919,n920,n921);
xor (n920,n883,n884);
and (n921,n141,n132);
and (n922,n923,n924);
xor (n923,n920,n921);
or (n924,n925,n928);
and (n925,n926,n927);
xor (n926,n889,n890);
and (n927,n168,n132);
and (n928,n929,n930);
xor (n929,n926,n927);
or (n930,n931,n934);
and (n931,n932,n933);
xor (n932,n895,n896);
and (n933,n39,n132);
and (n934,n935,n936);
xor (n935,n932,n933);
and (n936,n937,n402);
xor (n937,n901,n902);
or (n938,n939,n942);
and (n939,n940,n941);
xor (n940,n911,n912);
and (n941,n126,n124);
and (n942,n943,n944);
xor (n943,n940,n941);
or (n944,n945,n948);
and (n945,n946,n947);
xor (n946,n917,n918);
and (n947,n141,n124);
and (n948,n949,n950);
xor (n949,n946,n947);
or (n950,n951,n954);
and (n951,n952,n953);
xor (n952,n923,n924);
and (n953,n168,n124);
and (n954,n955,n956);
xor (n955,n952,n953);
or (n956,n957,n960);
and (n957,n958,n959);
xor (n958,n929,n930);
and (n959,n39,n124);
and (n960,n961,n962);
xor (n961,n958,n959);
and (n962,n963,n964);
xor (n963,n935,n936);
and (n964,n34,n124);
and (n965,n126,n158);
or (n966,n967,n970);
and (n967,n968,n969);
xor (n968,n943,n944);
and (n969,n141,n158);
and (n970,n971,n972);
xor (n971,n968,n969);
or (n972,n973,n976);
and (n973,n974,n975);
xor (n974,n949,n950);
and (n975,n168,n158);
and (n976,n977,n978);
xor (n977,n974,n975);
or (n978,n979,n982);
and (n979,n980,n981);
xor (n980,n955,n956);
and (n981,n39,n158);
and (n982,n983,n984);
xor (n983,n980,n981);
and (n984,n985,n227);
xor (n985,n961,n962);
and (n986,n141,n24);
or (n987,n988,n991);
and (n988,n989,n990);
xor (n989,n971,n972);
and (n990,n168,n24);
and (n991,n992,n993);
xor (n992,n989,n990);
or (n993,n994,n997);
and (n994,n995,n996);
xor (n995,n977,n978);
and (n996,n39,n24);
and (n997,n998,n999);
xor (n998,n995,n996);
and (n999,n1000,n1001);
xor (n1000,n983,n984);
and (n1001,n34,n24);
and (n1002,n168,n23);
or (n1003,n1004,n1007);
and (n1004,n1005,n1006);
xor (n1005,n992,n993);
and (n1006,n39,n23);
and (n1007,n1008,n1009);
xor (n1008,n1005,n1006);
and (n1009,n1010,n78);
xor (n1010,n998,n999);
and (n1011,n39,n28);
and (n1012,n1013,n1014);
xor (n1013,n1008,n1009);
and (n1014,n34,n28);
not (n1015,n1016);
nand (n1016,n34,n311);
endmodule
