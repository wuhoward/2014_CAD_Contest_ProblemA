module top (out,n23,n24,n28,n30,n37,n44,n51,n58,n65
        ,n72,n79,n86,n93,n99,n101,n168,n235,n302,n369
        ,n436,n503,n570,n637,n704,n790,n791,n795,n797,n804
        ,n811,n818,n825,n832,n839,n846,n853,n860,n866,n868
        ,n935,n1002,n1069,n1136,n1203,n1270,n1337,n1404,n1471,n1535);
output out;
input n23;
input n24;
input n28;
input n30;
input n37;
input n44;
input n51;
input n58;
input n65;
input n72;
input n79;
input n86;
input n93;
input n99;
input n101;
input n168;
input n235;
input n302;
input n369;
input n436;
input n503;
input n570;
input n637;
input n704;
input n790;
input n791;
input n795;
input n797;
input n804;
input n811;
input n818;
input n825;
input n832;
input n839;
input n846;
input n853;
input n860;
input n866;
input n868;
input n935;
input n1002;
input n1069;
input n1136;
input n1203;
input n1270;
input n1337;
input n1404;
input n1471;
input n1535;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n25;
wire n26;
wire n27;
wire n29;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n100;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n792;
wire n793;
wire n794;
wire n796;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n867;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
xor (out,n0,n1536);
wire s0n0,s1n0,notn0;
or (n0,s0n0,s1n0);
not(notn0,n1535);
and (s0n0,notn0,n1);
and (s1n0,n1535,n768);
xor (n1,n2,n705);
xor (n2,n3,n703);
or (n3,n4,n638);
and (n4,n5,n636);
or (n5,n6,n571);
and (n6,n7,n569);
or (n7,n8,n504);
and (n8,n9,n502);
or (n9,n10,n437);
and (n10,n11,n435);
or (n11,n12,n370);
and (n12,n13,n368);
or (n13,n14,n303);
and (n14,n15,n301);
or (n15,n16,n236);
and (n16,n17,n234);
or (n17,n18,n169);
and (n18,n19,n167);
or (n19,n20,n102);
and (n20,n21,n100);
and (n21,n22,n25);
and (n22,n23,n24);
or (n25,n26,n31);
and (n26,n27,n29);
and (n27,n23,n28);
and (n29,n30,n24);
and (n31,n32,n33);
xor (n32,n27,n29);
or (n33,n34,n38);
and (n34,n35,n36);
and (n35,n30,n28);
and (n36,n37,n24);
and (n38,n39,n40);
xor (n39,n35,n36);
or (n40,n41,n45);
and (n41,n42,n43);
and (n42,n37,n28);
and (n43,n44,n24);
and (n45,n46,n47);
xor (n46,n42,n43);
or (n47,n48,n52);
and (n48,n49,n50);
and (n49,n44,n28);
and (n50,n51,n24);
and (n52,n53,n54);
xor (n53,n49,n50);
or (n54,n55,n59);
and (n55,n56,n57);
and (n56,n51,n28);
and (n57,n58,n24);
and (n59,n60,n61);
xor (n60,n56,n57);
or (n61,n62,n66);
and (n62,n63,n64);
and (n63,n58,n28);
and (n64,n65,n24);
and (n66,n67,n68);
xor (n67,n63,n64);
or (n68,n69,n73);
and (n69,n70,n71);
and (n70,n65,n28);
and (n71,n72,n24);
and (n73,n74,n75);
xor (n74,n70,n71);
or (n75,n76,n80);
and (n76,n77,n78);
and (n77,n72,n28);
and (n78,n79,n24);
and (n80,n81,n82);
xor (n81,n77,n78);
or (n82,n83,n87);
and (n83,n84,n85);
and (n84,n79,n28);
and (n85,n86,n24);
and (n87,n88,n89);
xor (n88,n84,n85);
or (n89,n90,n94);
and (n90,n91,n92);
and (n91,n86,n28);
and (n92,n93,n24);
and (n94,n95,n96);
xor (n95,n91,n92);
and (n96,n97,n98);
and (n97,n93,n28);
and (n98,n99,n24);
and (n100,n23,n101);
and (n102,n103,n104);
xor (n103,n21,n100);
or (n104,n105,n108);
and (n105,n106,n107);
xor (n106,n22,n25);
and (n107,n30,n101);
and (n108,n109,n110);
xor (n109,n106,n107);
or (n110,n111,n114);
and (n111,n112,n113);
xor (n112,n32,n33);
and (n113,n37,n101);
and (n114,n115,n116);
xor (n115,n112,n113);
or (n116,n117,n120);
and (n117,n118,n119);
xor (n118,n39,n40);
and (n119,n44,n101);
and (n120,n121,n122);
xor (n121,n118,n119);
or (n122,n123,n126);
and (n123,n124,n125);
xor (n124,n46,n47);
and (n125,n51,n101);
and (n126,n127,n128);
xor (n127,n124,n125);
or (n128,n129,n132);
and (n129,n130,n131);
xor (n130,n53,n54);
and (n131,n58,n101);
and (n132,n133,n134);
xor (n133,n130,n131);
or (n134,n135,n138);
and (n135,n136,n137);
xor (n136,n60,n61);
and (n137,n65,n101);
and (n138,n139,n140);
xor (n139,n136,n137);
or (n140,n141,n144);
and (n141,n142,n143);
xor (n142,n67,n68);
and (n143,n72,n101);
and (n144,n145,n146);
xor (n145,n142,n143);
or (n146,n147,n150);
and (n147,n148,n149);
xor (n148,n74,n75);
and (n149,n79,n101);
and (n150,n151,n152);
xor (n151,n148,n149);
or (n152,n153,n156);
and (n153,n154,n155);
xor (n154,n81,n82);
and (n155,n86,n101);
and (n156,n157,n158);
xor (n157,n154,n155);
or (n158,n159,n162);
and (n159,n160,n161);
xor (n160,n88,n89);
and (n161,n93,n101);
and (n162,n163,n164);
xor (n163,n160,n161);
and (n164,n165,n166);
xor (n165,n95,n96);
and (n166,n99,n101);
and (n167,n23,n168);
and (n169,n170,n171);
xor (n170,n19,n167);
or (n171,n172,n175);
and (n172,n173,n174);
xor (n173,n103,n104);
and (n174,n30,n168);
and (n175,n176,n177);
xor (n176,n173,n174);
or (n177,n178,n181);
and (n178,n179,n180);
xor (n179,n109,n110);
and (n180,n37,n168);
and (n181,n182,n183);
xor (n182,n179,n180);
or (n183,n184,n187);
and (n184,n185,n186);
xor (n185,n115,n116);
and (n186,n44,n168);
and (n187,n188,n189);
xor (n188,n185,n186);
or (n189,n190,n193);
and (n190,n191,n192);
xor (n191,n121,n122);
and (n192,n51,n168);
and (n193,n194,n195);
xor (n194,n191,n192);
or (n195,n196,n199);
and (n196,n197,n198);
xor (n197,n127,n128);
and (n198,n58,n168);
and (n199,n200,n201);
xor (n200,n197,n198);
or (n201,n202,n205);
and (n202,n203,n204);
xor (n203,n133,n134);
and (n204,n65,n168);
and (n205,n206,n207);
xor (n206,n203,n204);
or (n207,n208,n211);
and (n208,n209,n210);
xor (n209,n139,n140);
and (n210,n72,n168);
and (n211,n212,n213);
xor (n212,n209,n210);
or (n213,n214,n217);
and (n214,n215,n216);
xor (n215,n145,n146);
and (n216,n79,n168);
and (n217,n218,n219);
xor (n218,n215,n216);
or (n219,n220,n223);
and (n220,n221,n222);
xor (n221,n151,n152);
and (n222,n86,n168);
and (n223,n224,n225);
xor (n224,n221,n222);
or (n225,n226,n229);
and (n226,n227,n228);
xor (n227,n157,n158);
and (n228,n93,n168);
and (n229,n230,n231);
xor (n230,n227,n228);
and (n231,n232,n233);
xor (n232,n163,n164);
and (n233,n99,n168);
and (n234,n23,n235);
and (n236,n237,n238);
xor (n237,n17,n234);
or (n238,n239,n242);
and (n239,n240,n241);
xor (n240,n170,n171);
and (n241,n30,n235);
and (n242,n243,n244);
xor (n243,n240,n241);
or (n244,n245,n248);
and (n245,n246,n247);
xor (n246,n176,n177);
and (n247,n37,n235);
and (n248,n249,n250);
xor (n249,n246,n247);
or (n250,n251,n254);
and (n251,n252,n253);
xor (n252,n182,n183);
and (n253,n44,n235);
and (n254,n255,n256);
xor (n255,n252,n253);
or (n256,n257,n260);
and (n257,n258,n259);
xor (n258,n188,n189);
and (n259,n51,n235);
and (n260,n261,n262);
xor (n261,n258,n259);
or (n262,n263,n266);
and (n263,n264,n265);
xor (n264,n194,n195);
and (n265,n58,n235);
and (n266,n267,n268);
xor (n267,n264,n265);
or (n268,n269,n272);
and (n269,n270,n271);
xor (n270,n200,n201);
and (n271,n65,n235);
and (n272,n273,n274);
xor (n273,n270,n271);
or (n274,n275,n278);
and (n275,n276,n277);
xor (n276,n206,n207);
and (n277,n72,n235);
and (n278,n279,n280);
xor (n279,n276,n277);
or (n280,n281,n284);
and (n281,n282,n283);
xor (n282,n212,n213);
and (n283,n79,n235);
and (n284,n285,n286);
xor (n285,n282,n283);
or (n286,n287,n290);
and (n287,n288,n289);
xor (n288,n218,n219);
and (n289,n86,n235);
and (n290,n291,n292);
xor (n291,n288,n289);
or (n292,n293,n296);
and (n293,n294,n295);
xor (n294,n224,n225);
and (n295,n93,n235);
and (n296,n297,n298);
xor (n297,n294,n295);
and (n298,n299,n300);
xor (n299,n230,n231);
and (n300,n99,n235);
and (n301,n23,n302);
and (n303,n304,n305);
xor (n304,n15,n301);
or (n305,n306,n309);
and (n306,n307,n308);
xor (n307,n237,n238);
and (n308,n30,n302);
and (n309,n310,n311);
xor (n310,n307,n308);
or (n311,n312,n315);
and (n312,n313,n314);
xor (n313,n243,n244);
and (n314,n37,n302);
and (n315,n316,n317);
xor (n316,n313,n314);
or (n317,n318,n321);
and (n318,n319,n320);
xor (n319,n249,n250);
and (n320,n44,n302);
and (n321,n322,n323);
xor (n322,n319,n320);
or (n323,n324,n327);
and (n324,n325,n326);
xor (n325,n255,n256);
and (n326,n51,n302);
and (n327,n328,n329);
xor (n328,n325,n326);
or (n329,n330,n333);
and (n330,n331,n332);
xor (n331,n261,n262);
and (n332,n58,n302);
and (n333,n334,n335);
xor (n334,n331,n332);
or (n335,n336,n339);
and (n336,n337,n338);
xor (n337,n267,n268);
and (n338,n65,n302);
and (n339,n340,n341);
xor (n340,n337,n338);
or (n341,n342,n345);
and (n342,n343,n344);
xor (n343,n273,n274);
and (n344,n72,n302);
and (n345,n346,n347);
xor (n346,n343,n344);
or (n347,n348,n351);
and (n348,n349,n350);
xor (n349,n279,n280);
and (n350,n79,n302);
and (n351,n352,n353);
xor (n352,n349,n350);
or (n353,n354,n357);
and (n354,n355,n356);
xor (n355,n285,n286);
and (n356,n86,n302);
and (n357,n358,n359);
xor (n358,n355,n356);
or (n359,n360,n363);
and (n360,n361,n362);
xor (n361,n291,n292);
and (n362,n93,n302);
and (n363,n364,n365);
xor (n364,n361,n362);
and (n365,n366,n367);
xor (n366,n297,n298);
and (n367,n99,n302);
and (n368,n23,n369);
and (n370,n371,n372);
xor (n371,n13,n368);
or (n372,n373,n376);
and (n373,n374,n375);
xor (n374,n304,n305);
and (n375,n30,n369);
and (n376,n377,n378);
xor (n377,n374,n375);
or (n378,n379,n382);
and (n379,n380,n381);
xor (n380,n310,n311);
and (n381,n37,n369);
and (n382,n383,n384);
xor (n383,n380,n381);
or (n384,n385,n388);
and (n385,n386,n387);
xor (n386,n316,n317);
and (n387,n44,n369);
and (n388,n389,n390);
xor (n389,n386,n387);
or (n390,n391,n394);
and (n391,n392,n393);
xor (n392,n322,n323);
and (n393,n51,n369);
and (n394,n395,n396);
xor (n395,n392,n393);
or (n396,n397,n400);
and (n397,n398,n399);
xor (n398,n328,n329);
and (n399,n58,n369);
and (n400,n401,n402);
xor (n401,n398,n399);
or (n402,n403,n406);
and (n403,n404,n405);
xor (n404,n334,n335);
and (n405,n65,n369);
and (n406,n407,n408);
xor (n407,n404,n405);
or (n408,n409,n412);
and (n409,n410,n411);
xor (n410,n340,n341);
and (n411,n72,n369);
and (n412,n413,n414);
xor (n413,n410,n411);
or (n414,n415,n418);
and (n415,n416,n417);
xor (n416,n346,n347);
and (n417,n79,n369);
and (n418,n419,n420);
xor (n419,n416,n417);
or (n420,n421,n424);
and (n421,n422,n423);
xor (n422,n352,n353);
and (n423,n86,n369);
and (n424,n425,n426);
xor (n425,n422,n423);
or (n426,n427,n430);
and (n427,n428,n429);
xor (n428,n358,n359);
and (n429,n93,n369);
and (n430,n431,n432);
xor (n431,n428,n429);
and (n432,n433,n434);
xor (n433,n364,n365);
and (n434,n99,n369);
and (n435,n23,n436);
and (n437,n438,n439);
xor (n438,n11,n435);
or (n439,n440,n443);
and (n440,n441,n442);
xor (n441,n371,n372);
and (n442,n30,n436);
and (n443,n444,n445);
xor (n444,n441,n442);
or (n445,n446,n449);
and (n446,n447,n448);
xor (n447,n377,n378);
and (n448,n37,n436);
and (n449,n450,n451);
xor (n450,n447,n448);
or (n451,n452,n455);
and (n452,n453,n454);
xor (n453,n383,n384);
and (n454,n44,n436);
and (n455,n456,n457);
xor (n456,n453,n454);
or (n457,n458,n461);
and (n458,n459,n460);
xor (n459,n389,n390);
and (n460,n51,n436);
and (n461,n462,n463);
xor (n462,n459,n460);
or (n463,n464,n467);
and (n464,n465,n466);
xor (n465,n395,n396);
and (n466,n58,n436);
and (n467,n468,n469);
xor (n468,n465,n466);
or (n469,n470,n473);
and (n470,n471,n472);
xor (n471,n401,n402);
and (n472,n65,n436);
and (n473,n474,n475);
xor (n474,n471,n472);
or (n475,n476,n479);
and (n476,n477,n478);
xor (n477,n407,n408);
and (n478,n72,n436);
and (n479,n480,n481);
xor (n480,n477,n478);
or (n481,n482,n485);
and (n482,n483,n484);
xor (n483,n413,n414);
and (n484,n79,n436);
and (n485,n486,n487);
xor (n486,n483,n484);
or (n487,n488,n491);
and (n488,n489,n490);
xor (n489,n419,n420);
and (n490,n86,n436);
and (n491,n492,n493);
xor (n492,n489,n490);
or (n493,n494,n497);
and (n494,n495,n496);
xor (n495,n425,n426);
and (n496,n93,n436);
and (n497,n498,n499);
xor (n498,n495,n496);
and (n499,n500,n501);
xor (n500,n431,n432);
and (n501,n99,n436);
and (n502,n23,n503);
and (n504,n505,n506);
xor (n505,n9,n502);
or (n506,n507,n510);
and (n507,n508,n509);
xor (n508,n438,n439);
and (n509,n30,n503);
and (n510,n511,n512);
xor (n511,n508,n509);
or (n512,n513,n516);
and (n513,n514,n515);
xor (n514,n444,n445);
and (n515,n37,n503);
and (n516,n517,n518);
xor (n517,n514,n515);
or (n518,n519,n522);
and (n519,n520,n521);
xor (n520,n450,n451);
and (n521,n44,n503);
and (n522,n523,n524);
xor (n523,n520,n521);
or (n524,n525,n528);
and (n525,n526,n527);
xor (n526,n456,n457);
and (n527,n51,n503);
and (n528,n529,n530);
xor (n529,n526,n527);
or (n530,n531,n534);
and (n531,n532,n533);
xor (n532,n462,n463);
and (n533,n58,n503);
and (n534,n535,n536);
xor (n535,n532,n533);
or (n536,n537,n540);
and (n537,n538,n539);
xor (n538,n468,n469);
and (n539,n65,n503);
and (n540,n541,n542);
xor (n541,n538,n539);
or (n542,n543,n546);
and (n543,n544,n545);
xor (n544,n474,n475);
and (n545,n72,n503);
and (n546,n547,n548);
xor (n547,n544,n545);
or (n548,n549,n552);
and (n549,n550,n551);
xor (n550,n480,n481);
and (n551,n79,n503);
and (n552,n553,n554);
xor (n553,n550,n551);
or (n554,n555,n558);
and (n555,n556,n557);
xor (n556,n486,n487);
and (n557,n86,n503);
and (n558,n559,n560);
xor (n559,n556,n557);
or (n560,n561,n564);
and (n561,n562,n563);
xor (n562,n492,n493);
and (n563,n93,n503);
and (n564,n565,n566);
xor (n565,n562,n563);
and (n566,n567,n568);
xor (n567,n498,n499);
and (n568,n99,n503);
and (n569,n23,n570);
and (n571,n572,n573);
xor (n572,n7,n569);
or (n573,n574,n577);
and (n574,n575,n576);
xor (n575,n505,n506);
and (n576,n30,n570);
and (n577,n578,n579);
xor (n578,n575,n576);
or (n579,n580,n583);
and (n580,n581,n582);
xor (n581,n511,n512);
and (n582,n37,n570);
and (n583,n584,n585);
xor (n584,n581,n582);
or (n585,n586,n589);
and (n586,n587,n588);
xor (n587,n517,n518);
and (n588,n44,n570);
and (n589,n590,n591);
xor (n590,n587,n588);
or (n591,n592,n595);
and (n592,n593,n594);
xor (n593,n523,n524);
and (n594,n51,n570);
and (n595,n596,n597);
xor (n596,n593,n594);
or (n597,n598,n601);
and (n598,n599,n600);
xor (n599,n529,n530);
and (n600,n58,n570);
and (n601,n602,n603);
xor (n602,n599,n600);
or (n603,n604,n607);
and (n604,n605,n606);
xor (n605,n535,n536);
and (n606,n65,n570);
and (n607,n608,n609);
xor (n608,n605,n606);
or (n609,n610,n613);
and (n610,n611,n612);
xor (n611,n541,n542);
and (n612,n72,n570);
and (n613,n614,n615);
xor (n614,n611,n612);
or (n615,n616,n619);
and (n616,n617,n618);
xor (n617,n547,n548);
and (n618,n79,n570);
and (n619,n620,n621);
xor (n620,n617,n618);
or (n621,n622,n625);
and (n622,n623,n624);
xor (n623,n553,n554);
and (n624,n86,n570);
and (n625,n626,n627);
xor (n626,n623,n624);
or (n627,n628,n631);
and (n628,n629,n630);
xor (n629,n559,n560);
and (n630,n93,n570);
and (n631,n632,n633);
xor (n632,n629,n630);
and (n633,n634,n635);
xor (n634,n565,n566);
and (n635,n99,n570);
and (n636,n23,n637);
and (n638,n639,n640);
xor (n639,n5,n636);
or (n640,n641,n644);
and (n641,n642,n643);
xor (n642,n572,n573);
and (n643,n30,n637);
and (n644,n645,n646);
xor (n645,n642,n643);
or (n646,n647,n650);
and (n647,n648,n649);
xor (n648,n578,n579);
and (n649,n37,n637);
and (n650,n651,n652);
xor (n651,n648,n649);
or (n652,n653,n656);
and (n653,n654,n655);
xor (n654,n584,n585);
and (n655,n44,n637);
and (n656,n657,n658);
xor (n657,n654,n655);
or (n658,n659,n662);
and (n659,n660,n661);
xor (n660,n590,n591);
and (n661,n51,n637);
and (n662,n663,n664);
xor (n663,n660,n661);
or (n664,n665,n668);
and (n665,n666,n667);
xor (n666,n596,n597);
and (n667,n58,n637);
and (n668,n669,n670);
xor (n669,n666,n667);
or (n670,n671,n674);
and (n671,n672,n673);
xor (n672,n602,n603);
and (n673,n65,n637);
and (n674,n675,n676);
xor (n675,n672,n673);
or (n676,n677,n680);
and (n677,n678,n679);
xor (n678,n608,n609);
and (n679,n72,n637);
and (n680,n681,n682);
xor (n681,n678,n679);
or (n682,n683,n686);
and (n683,n684,n685);
xor (n684,n614,n615);
and (n685,n79,n637);
and (n686,n687,n688);
xor (n687,n684,n685);
or (n688,n689,n692);
and (n689,n690,n691);
xor (n690,n620,n621);
and (n691,n86,n637);
and (n692,n693,n694);
xor (n693,n690,n691);
or (n694,n695,n698);
and (n695,n696,n697);
xor (n696,n626,n627);
and (n697,n93,n637);
and (n698,n699,n700);
xor (n699,n696,n697);
and (n700,n701,n702);
xor (n701,n632,n633);
and (n702,n99,n637);
and (n703,n23,n704);
or (n705,n706,n709);
and (n706,n707,n708);
xor (n707,n639,n640);
and (n708,n30,n704);
and (n709,n710,n711);
xor (n710,n707,n708);
or (n711,n712,n715);
and (n712,n713,n714);
xor (n713,n645,n646);
and (n714,n37,n704);
and (n715,n716,n717);
xor (n716,n713,n714);
or (n717,n718,n721);
and (n718,n719,n720);
xor (n719,n651,n652);
and (n720,n44,n704);
and (n721,n722,n723);
xor (n722,n719,n720);
or (n723,n724,n727);
and (n724,n725,n726);
xor (n725,n657,n658);
and (n726,n51,n704);
and (n727,n728,n729);
xor (n728,n725,n726);
or (n729,n730,n733);
and (n730,n731,n732);
xor (n731,n663,n664);
and (n732,n58,n704);
and (n733,n734,n735);
xor (n734,n731,n732);
or (n735,n736,n739);
and (n736,n737,n738);
xor (n737,n669,n670);
and (n738,n65,n704);
and (n739,n740,n741);
xor (n740,n737,n738);
or (n741,n742,n745);
and (n742,n743,n744);
xor (n743,n675,n676);
and (n744,n72,n704);
and (n745,n746,n747);
xor (n746,n743,n744);
or (n747,n748,n751);
and (n748,n749,n750);
xor (n749,n681,n682);
and (n750,n79,n704);
and (n751,n752,n753);
xor (n752,n749,n750);
or (n753,n754,n757);
and (n754,n755,n756);
xor (n755,n687,n688);
and (n756,n86,n704);
and (n757,n758,n759);
xor (n758,n755,n756);
or (n759,n760,n763);
and (n760,n761,n762);
xor (n761,n693,n694);
and (n762,n93,n704);
and (n763,n764,n765);
xor (n764,n761,n762);
and (n765,n766,n767);
xor (n766,n699,n700);
and (n767,n99,n704);
xor (n768,n769,n1472);
xor (n769,n770,n1470);
or (n770,n771,n1405);
and (n771,n772,n1403);
or (n772,n773,n1338);
and (n773,n774,n1336);
or (n774,n775,n1271);
and (n775,n776,n1269);
or (n776,n777,n1204);
and (n777,n778,n1202);
or (n778,n779,n1137);
and (n779,n780,n1135);
or (n780,n781,n1070);
and (n781,n782,n1068);
or (n782,n783,n1003);
and (n783,n784,n1001);
or (n784,n785,n936);
and (n785,n786,n934);
or (n786,n787,n869);
and (n787,n788,n867);
and (n788,n789,n792);
and (n789,n790,n791);
or (n792,n793,n798);
and (n793,n794,n796);
and (n794,n790,n795);
and (n796,n797,n791);
and (n798,n799,n800);
xor (n799,n794,n796);
or (n800,n801,n805);
and (n801,n802,n803);
and (n802,n797,n795);
and (n803,n804,n791);
and (n805,n806,n807);
xor (n806,n802,n803);
or (n807,n808,n812);
and (n808,n809,n810);
and (n809,n804,n795);
and (n810,n811,n791);
and (n812,n813,n814);
xor (n813,n809,n810);
or (n814,n815,n819);
and (n815,n816,n817);
and (n816,n811,n795);
and (n817,n818,n791);
and (n819,n820,n821);
xor (n820,n816,n817);
or (n821,n822,n826);
and (n822,n823,n824);
and (n823,n818,n795);
and (n824,n825,n791);
and (n826,n827,n828);
xor (n827,n823,n824);
or (n828,n829,n833);
and (n829,n830,n831);
and (n830,n825,n795);
and (n831,n832,n791);
and (n833,n834,n835);
xor (n834,n830,n831);
or (n835,n836,n840);
and (n836,n837,n838);
and (n837,n832,n795);
and (n838,n839,n791);
and (n840,n841,n842);
xor (n841,n837,n838);
or (n842,n843,n847);
and (n843,n844,n845);
and (n844,n839,n795);
and (n845,n846,n791);
and (n847,n848,n849);
xor (n848,n844,n845);
or (n849,n850,n854);
and (n850,n851,n852);
and (n851,n846,n795);
and (n852,n853,n791);
and (n854,n855,n856);
xor (n855,n851,n852);
or (n856,n857,n861);
and (n857,n858,n859);
and (n858,n853,n795);
and (n859,n860,n791);
and (n861,n862,n863);
xor (n862,n858,n859);
and (n863,n864,n865);
and (n864,n860,n795);
and (n865,n866,n791);
and (n867,n790,n868);
and (n869,n870,n871);
xor (n870,n788,n867);
or (n871,n872,n875);
and (n872,n873,n874);
xor (n873,n789,n792);
and (n874,n797,n868);
and (n875,n876,n877);
xor (n876,n873,n874);
or (n877,n878,n881);
and (n878,n879,n880);
xor (n879,n799,n800);
and (n880,n804,n868);
and (n881,n882,n883);
xor (n882,n879,n880);
or (n883,n884,n887);
and (n884,n885,n886);
xor (n885,n806,n807);
and (n886,n811,n868);
and (n887,n888,n889);
xor (n888,n885,n886);
or (n889,n890,n893);
and (n890,n891,n892);
xor (n891,n813,n814);
and (n892,n818,n868);
and (n893,n894,n895);
xor (n894,n891,n892);
or (n895,n896,n899);
and (n896,n897,n898);
xor (n897,n820,n821);
and (n898,n825,n868);
and (n899,n900,n901);
xor (n900,n897,n898);
or (n901,n902,n905);
and (n902,n903,n904);
xor (n903,n827,n828);
and (n904,n832,n868);
and (n905,n906,n907);
xor (n906,n903,n904);
or (n907,n908,n911);
and (n908,n909,n910);
xor (n909,n834,n835);
and (n910,n839,n868);
and (n911,n912,n913);
xor (n912,n909,n910);
or (n913,n914,n917);
and (n914,n915,n916);
xor (n915,n841,n842);
and (n916,n846,n868);
and (n917,n918,n919);
xor (n918,n915,n916);
or (n919,n920,n923);
and (n920,n921,n922);
xor (n921,n848,n849);
and (n922,n853,n868);
and (n923,n924,n925);
xor (n924,n921,n922);
or (n925,n926,n929);
and (n926,n927,n928);
xor (n927,n855,n856);
and (n928,n860,n868);
and (n929,n930,n931);
xor (n930,n927,n928);
and (n931,n932,n933);
xor (n932,n862,n863);
and (n933,n866,n868);
and (n934,n790,n935);
and (n936,n937,n938);
xor (n937,n786,n934);
or (n938,n939,n942);
and (n939,n940,n941);
xor (n940,n870,n871);
and (n941,n797,n935);
and (n942,n943,n944);
xor (n943,n940,n941);
or (n944,n945,n948);
and (n945,n946,n947);
xor (n946,n876,n877);
and (n947,n804,n935);
and (n948,n949,n950);
xor (n949,n946,n947);
or (n950,n951,n954);
and (n951,n952,n953);
xor (n952,n882,n883);
and (n953,n811,n935);
and (n954,n955,n956);
xor (n955,n952,n953);
or (n956,n957,n960);
and (n957,n958,n959);
xor (n958,n888,n889);
and (n959,n818,n935);
and (n960,n961,n962);
xor (n961,n958,n959);
or (n962,n963,n966);
and (n963,n964,n965);
xor (n964,n894,n895);
and (n965,n825,n935);
and (n966,n967,n968);
xor (n967,n964,n965);
or (n968,n969,n972);
and (n969,n970,n971);
xor (n970,n900,n901);
and (n971,n832,n935);
and (n972,n973,n974);
xor (n973,n970,n971);
or (n974,n975,n978);
and (n975,n976,n977);
xor (n976,n906,n907);
and (n977,n839,n935);
and (n978,n979,n980);
xor (n979,n976,n977);
or (n980,n981,n984);
and (n981,n982,n983);
xor (n982,n912,n913);
and (n983,n846,n935);
and (n984,n985,n986);
xor (n985,n982,n983);
or (n986,n987,n990);
and (n987,n988,n989);
xor (n988,n918,n919);
and (n989,n853,n935);
and (n990,n991,n992);
xor (n991,n988,n989);
or (n992,n993,n996);
and (n993,n994,n995);
xor (n994,n924,n925);
and (n995,n860,n935);
and (n996,n997,n998);
xor (n997,n994,n995);
and (n998,n999,n1000);
xor (n999,n930,n931);
and (n1000,n866,n935);
and (n1001,n790,n1002);
and (n1003,n1004,n1005);
xor (n1004,n784,n1001);
or (n1005,n1006,n1009);
and (n1006,n1007,n1008);
xor (n1007,n937,n938);
and (n1008,n797,n1002);
and (n1009,n1010,n1011);
xor (n1010,n1007,n1008);
or (n1011,n1012,n1015);
and (n1012,n1013,n1014);
xor (n1013,n943,n944);
and (n1014,n804,n1002);
and (n1015,n1016,n1017);
xor (n1016,n1013,n1014);
or (n1017,n1018,n1021);
and (n1018,n1019,n1020);
xor (n1019,n949,n950);
and (n1020,n811,n1002);
and (n1021,n1022,n1023);
xor (n1022,n1019,n1020);
or (n1023,n1024,n1027);
and (n1024,n1025,n1026);
xor (n1025,n955,n956);
and (n1026,n818,n1002);
and (n1027,n1028,n1029);
xor (n1028,n1025,n1026);
or (n1029,n1030,n1033);
and (n1030,n1031,n1032);
xor (n1031,n961,n962);
and (n1032,n825,n1002);
and (n1033,n1034,n1035);
xor (n1034,n1031,n1032);
or (n1035,n1036,n1039);
and (n1036,n1037,n1038);
xor (n1037,n967,n968);
and (n1038,n832,n1002);
and (n1039,n1040,n1041);
xor (n1040,n1037,n1038);
or (n1041,n1042,n1045);
and (n1042,n1043,n1044);
xor (n1043,n973,n974);
and (n1044,n839,n1002);
and (n1045,n1046,n1047);
xor (n1046,n1043,n1044);
or (n1047,n1048,n1051);
and (n1048,n1049,n1050);
xor (n1049,n979,n980);
and (n1050,n846,n1002);
and (n1051,n1052,n1053);
xor (n1052,n1049,n1050);
or (n1053,n1054,n1057);
and (n1054,n1055,n1056);
xor (n1055,n985,n986);
and (n1056,n853,n1002);
and (n1057,n1058,n1059);
xor (n1058,n1055,n1056);
or (n1059,n1060,n1063);
and (n1060,n1061,n1062);
xor (n1061,n991,n992);
and (n1062,n860,n1002);
and (n1063,n1064,n1065);
xor (n1064,n1061,n1062);
and (n1065,n1066,n1067);
xor (n1066,n997,n998);
and (n1067,n866,n1002);
and (n1068,n790,n1069);
and (n1070,n1071,n1072);
xor (n1071,n782,n1068);
or (n1072,n1073,n1076);
and (n1073,n1074,n1075);
xor (n1074,n1004,n1005);
and (n1075,n797,n1069);
and (n1076,n1077,n1078);
xor (n1077,n1074,n1075);
or (n1078,n1079,n1082);
and (n1079,n1080,n1081);
xor (n1080,n1010,n1011);
and (n1081,n804,n1069);
and (n1082,n1083,n1084);
xor (n1083,n1080,n1081);
or (n1084,n1085,n1088);
and (n1085,n1086,n1087);
xor (n1086,n1016,n1017);
and (n1087,n811,n1069);
and (n1088,n1089,n1090);
xor (n1089,n1086,n1087);
or (n1090,n1091,n1094);
and (n1091,n1092,n1093);
xor (n1092,n1022,n1023);
and (n1093,n818,n1069);
and (n1094,n1095,n1096);
xor (n1095,n1092,n1093);
or (n1096,n1097,n1100);
and (n1097,n1098,n1099);
xor (n1098,n1028,n1029);
and (n1099,n825,n1069);
and (n1100,n1101,n1102);
xor (n1101,n1098,n1099);
or (n1102,n1103,n1106);
and (n1103,n1104,n1105);
xor (n1104,n1034,n1035);
and (n1105,n832,n1069);
and (n1106,n1107,n1108);
xor (n1107,n1104,n1105);
or (n1108,n1109,n1112);
and (n1109,n1110,n1111);
xor (n1110,n1040,n1041);
and (n1111,n839,n1069);
and (n1112,n1113,n1114);
xor (n1113,n1110,n1111);
or (n1114,n1115,n1118);
and (n1115,n1116,n1117);
xor (n1116,n1046,n1047);
and (n1117,n846,n1069);
and (n1118,n1119,n1120);
xor (n1119,n1116,n1117);
or (n1120,n1121,n1124);
and (n1121,n1122,n1123);
xor (n1122,n1052,n1053);
and (n1123,n853,n1069);
and (n1124,n1125,n1126);
xor (n1125,n1122,n1123);
or (n1126,n1127,n1130);
and (n1127,n1128,n1129);
xor (n1128,n1058,n1059);
and (n1129,n860,n1069);
and (n1130,n1131,n1132);
xor (n1131,n1128,n1129);
and (n1132,n1133,n1134);
xor (n1133,n1064,n1065);
and (n1134,n866,n1069);
and (n1135,n790,n1136);
and (n1137,n1138,n1139);
xor (n1138,n780,n1135);
or (n1139,n1140,n1143);
and (n1140,n1141,n1142);
xor (n1141,n1071,n1072);
and (n1142,n797,n1136);
and (n1143,n1144,n1145);
xor (n1144,n1141,n1142);
or (n1145,n1146,n1149);
and (n1146,n1147,n1148);
xor (n1147,n1077,n1078);
and (n1148,n804,n1136);
and (n1149,n1150,n1151);
xor (n1150,n1147,n1148);
or (n1151,n1152,n1155);
and (n1152,n1153,n1154);
xor (n1153,n1083,n1084);
and (n1154,n811,n1136);
and (n1155,n1156,n1157);
xor (n1156,n1153,n1154);
or (n1157,n1158,n1161);
and (n1158,n1159,n1160);
xor (n1159,n1089,n1090);
and (n1160,n818,n1136);
and (n1161,n1162,n1163);
xor (n1162,n1159,n1160);
or (n1163,n1164,n1167);
and (n1164,n1165,n1166);
xor (n1165,n1095,n1096);
and (n1166,n825,n1136);
and (n1167,n1168,n1169);
xor (n1168,n1165,n1166);
or (n1169,n1170,n1173);
and (n1170,n1171,n1172);
xor (n1171,n1101,n1102);
and (n1172,n832,n1136);
and (n1173,n1174,n1175);
xor (n1174,n1171,n1172);
or (n1175,n1176,n1179);
and (n1176,n1177,n1178);
xor (n1177,n1107,n1108);
and (n1178,n839,n1136);
and (n1179,n1180,n1181);
xor (n1180,n1177,n1178);
or (n1181,n1182,n1185);
and (n1182,n1183,n1184);
xor (n1183,n1113,n1114);
and (n1184,n846,n1136);
and (n1185,n1186,n1187);
xor (n1186,n1183,n1184);
or (n1187,n1188,n1191);
and (n1188,n1189,n1190);
xor (n1189,n1119,n1120);
and (n1190,n853,n1136);
and (n1191,n1192,n1193);
xor (n1192,n1189,n1190);
or (n1193,n1194,n1197);
and (n1194,n1195,n1196);
xor (n1195,n1125,n1126);
and (n1196,n860,n1136);
and (n1197,n1198,n1199);
xor (n1198,n1195,n1196);
and (n1199,n1200,n1201);
xor (n1200,n1131,n1132);
and (n1201,n866,n1136);
and (n1202,n790,n1203);
and (n1204,n1205,n1206);
xor (n1205,n778,n1202);
or (n1206,n1207,n1210);
and (n1207,n1208,n1209);
xor (n1208,n1138,n1139);
and (n1209,n797,n1203);
and (n1210,n1211,n1212);
xor (n1211,n1208,n1209);
or (n1212,n1213,n1216);
and (n1213,n1214,n1215);
xor (n1214,n1144,n1145);
and (n1215,n804,n1203);
and (n1216,n1217,n1218);
xor (n1217,n1214,n1215);
or (n1218,n1219,n1222);
and (n1219,n1220,n1221);
xor (n1220,n1150,n1151);
and (n1221,n811,n1203);
and (n1222,n1223,n1224);
xor (n1223,n1220,n1221);
or (n1224,n1225,n1228);
and (n1225,n1226,n1227);
xor (n1226,n1156,n1157);
and (n1227,n818,n1203);
and (n1228,n1229,n1230);
xor (n1229,n1226,n1227);
or (n1230,n1231,n1234);
and (n1231,n1232,n1233);
xor (n1232,n1162,n1163);
and (n1233,n825,n1203);
and (n1234,n1235,n1236);
xor (n1235,n1232,n1233);
or (n1236,n1237,n1240);
and (n1237,n1238,n1239);
xor (n1238,n1168,n1169);
and (n1239,n832,n1203);
and (n1240,n1241,n1242);
xor (n1241,n1238,n1239);
or (n1242,n1243,n1246);
and (n1243,n1244,n1245);
xor (n1244,n1174,n1175);
and (n1245,n839,n1203);
and (n1246,n1247,n1248);
xor (n1247,n1244,n1245);
or (n1248,n1249,n1252);
and (n1249,n1250,n1251);
xor (n1250,n1180,n1181);
and (n1251,n846,n1203);
and (n1252,n1253,n1254);
xor (n1253,n1250,n1251);
or (n1254,n1255,n1258);
and (n1255,n1256,n1257);
xor (n1256,n1186,n1187);
and (n1257,n853,n1203);
and (n1258,n1259,n1260);
xor (n1259,n1256,n1257);
or (n1260,n1261,n1264);
and (n1261,n1262,n1263);
xor (n1262,n1192,n1193);
and (n1263,n860,n1203);
and (n1264,n1265,n1266);
xor (n1265,n1262,n1263);
and (n1266,n1267,n1268);
xor (n1267,n1198,n1199);
and (n1268,n866,n1203);
and (n1269,n790,n1270);
and (n1271,n1272,n1273);
xor (n1272,n776,n1269);
or (n1273,n1274,n1277);
and (n1274,n1275,n1276);
xor (n1275,n1205,n1206);
and (n1276,n797,n1270);
and (n1277,n1278,n1279);
xor (n1278,n1275,n1276);
or (n1279,n1280,n1283);
and (n1280,n1281,n1282);
xor (n1281,n1211,n1212);
and (n1282,n804,n1270);
and (n1283,n1284,n1285);
xor (n1284,n1281,n1282);
or (n1285,n1286,n1289);
and (n1286,n1287,n1288);
xor (n1287,n1217,n1218);
and (n1288,n811,n1270);
and (n1289,n1290,n1291);
xor (n1290,n1287,n1288);
or (n1291,n1292,n1295);
and (n1292,n1293,n1294);
xor (n1293,n1223,n1224);
and (n1294,n818,n1270);
and (n1295,n1296,n1297);
xor (n1296,n1293,n1294);
or (n1297,n1298,n1301);
and (n1298,n1299,n1300);
xor (n1299,n1229,n1230);
and (n1300,n825,n1270);
and (n1301,n1302,n1303);
xor (n1302,n1299,n1300);
or (n1303,n1304,n1307);
and (n1304,n1305,n1306);
xor (n1305,n1235,n1236);
and (n1306,n832,n1270);
and (n1307,n1308,n1309);
xor (n1308,n1305,n1306);
or (n1309,n1310,n1313);
and (n1310,n1311,n1312);
xor (n1311,n1241,n1242);
and (n1312,n839,n1270);
and (n1313,n1314,n1315);
xor (n1314,n1311,n1312);
or (n1315,n1316,n1319);
and (n1316,n1317,n1318);
xor (n1317,n1247,n1248);
and (n1318,n846,n1270);
and (n1319,n1320,n1321);
xor (n1320,n1317,n1318);
or (n1321,n1322,n1325);
and (n1322,n1323,n1324);
xor (n1323,n1253,n1254);
and (n1324,n853,n1270);
and (n1325,n1326,n1327);
xor (n1326,n1323,n1324);
or (n1327,n1328,n1331);
and (n1328,n1329,n1330);
xor (n1329,n1259,n1260);
and (n1330,n860,n1270);
and (n1331,n1332,n1333);
xor (n1332,n1329,n1330);
and (n1333,n1334,n1335);
xor (n1334,n1265,n1266);
and (n1335,n866,n1270);
and (n1336,n790,n1337);
and (n1338,n1339,n1340);
xor (n1339,n774,n1336);
or (n1340,n1341,n1344);
and (n1341,n1342,n1343);
xor (n1342,n1272,n1273);
and (n1343,n797,n1337);
and (n1344,n1345,n1346);
xor (n1345,n1342,n1343);
or (n1346,n1347,n1350);
and (n1347,n1348,n1349);
xor (n1348,n1278,n1279);
and (n1349,n804,n1337);
and (n1350,n1351,n1352);
xor (n1351,n1348,n1349);
or (n1352,n1353,n1356);
and (n1353,n1354,n1355);
xor (n1354,n1284,n1285);
and (n1355,n811,n1337);
and (n1356,n1357,n1358);
xor (n1357,n1354,n1355);
or (n1358,n1359,n1362);
and (n1359,n1360,n1361);
xor (n1360,n1290,n1291);
and (n1361,n818,n1337);
and (n1362,n1363,n1364);
xor (n1363,n1360,n1361);
or (n1364,n1365,n1368);
and (n1365,n1366,n1367);
xor (n1366,n1296,n1297);
and (n1367,n825,n1337);
and (n1368,n1369,n1370);
xor (n1369,n1366,n1367);
or (n1370,n1371,n1374);
and (n1371,n1372,n1373);
xor (n1372,n1302,n1303);
and (n1373,n832,n1337);
and (n1374,n1375,n1376);
xor (n1375,n1372,n1373);
or (n1376,n1377,n1380);
and (n1377,n1378,n1379);
xor (n1378,n1308,n1309);
and (n1379,n839,n1337);
and (n1380,n1381,n1382);
xor (n1381,n1378,n1379);
or (n1382,n1383,n1386);
and (n1383,n1384,n1385);
xor (n1384,n1314,n1315);
and (n1385,n846,n1337);
and (n1386,n1387,n1388);
xor (n1387,n1384,n1385);
or (n1388,n1389,n1392);
and (n1389,n1390,n1391);
xor (n1390,n1320,n1321);
and (n1391,n853,n1337);
and (n1392,n1393,n1394);
xor (n1393,n1390,n1391);
or (n1394,n1395,n1398);
and (n1395,n1396,n1397);
xor (n1396,n1326,n1327);
and (n1397,n860,n1337);
and (n1398,n1399,n1400);
xor (n1399,n1396,n1397);
and (n1400,n1401,n1402);
xor (n1401,n1332,n1333);
and (n1402,n866,n1337);
and (n1403,n790,n1404);
and (n1405,n1406,n1407);
xor (n1406,n772,n1403);
or (n1407,n1408,n1411);
and (n1408,n1409,n1410);
xor (n1409,n1339,n1340);
and (n1410,n797,n1404);
and (n1411,n1412,n1413);
xor (n1412,n1409,n1410);
or (n1413,n1414,n1417);
and (n1414,n1415,n1416);
xor (n1415,n1345,n1346);
and (n1416,n804,n1404);
and (n1417,n1418,n1419);
xor (n1418,n1415,n1416);
or (n1419,n1420,n1423);
and (n1420,n1421,n1422);
xor (n1421,n1351,n1352);
and (n1422,n811,n1404);
and (n1423,n1424,n1425);
xor (n1424,n1421,n1422);
or (n1425,n1426,n1429);
and (n1426,n1427,n1428);
xor (n1427,n1357,n1358);
and (n1428,n818,n1404);
and (n1429,n1430,n1431);
xor (n1430,n1427,n1428);
or (n1431,n1432,n1435);
and (n1432,n1433,n1434);
xor (n1433,n1363,n1364);
and (n1434,n825,n1404);
and (n1435,n1436,n1437);
xor (n1436,n1433,n1434);
or (n1437,n1438,n1441);
and (n1438,n1439,n1440);
xor (n1439,n1369,n1370);
and (n1440,n832,n1404);
and (n1441,n1442,n1443);
xor (n1442,n1439,n1440);
or (n1443,n1444,n1447);
and (n1444,n1445,n1446);
xor (n1445,n1375,n1376);
and (n1446,n839,n1404);
and (n1447,n1448,n1449);
xor (n1448,n1445,n1446);
or (n1449,n1450,n1453);
and (n1450,n1451,n1452);
xor (n1451,n1381,n1382);
and (n1452,n846,n1404);
and (n1453,n1454,n1455);
xor (n1454,n1451,n1452);
or (n1455,n1456,n1459);
and (n1456,n1457,n1458);
xor (n1457,n1387,n1388);
and (n1458,n853,n1404);
and (n1459,n1460,n1461);
xor (n1460,n1457,n1458);
or (n1461,n1462,n1465);
and (n1462,n1463,n1464);
xor (n1463,n1393,n1394);
and (n1464,n860,n1404);
and (n1465,n1466,n1467);
xor (n1466,n1463,n1464);
and (n1467,n1468,n1469);
xor (n1468,n1399,n1400);
and (n1469,n866,n1404);
and (n1470,n790,n1471);
or (n1472,n1473,n1476);
and (n1473,n1474,n1475);
xor (n1474,n1406,n1407);
and (n1475,n797,n1471);
and (n1476,n1477,n1478);
xor (n1477,n1474,n1475);
or (n1478,n1479,n1482);
and (n1479,n1480,n1481);
xor (n1480,n1412,n1413);
and (n1481,n804,n1471);
and (n1482,n1483,n1484);
xor (n1483,n1480,n1481);
or (n1484,n1485,n1488);
and (n1485,n1486,n1487);
xor (n1486,n1418,n1419);
and (n1487,n811,n1471);
and (n1488,n1489,n1490);
xor (n1489,n1486,n1487);
or (n1490,n1491,n1494);
and (n1491,n1492,n1493);
xor (n1492,n1424,n1425);
and (n1493,n818,n1471);
and (n1494,n1495,n1496);
xor (n1495,n1492,n1493);
or (n1496,n1497,n1500);
and (n1497,n1498,n1499);
xor (n1498,n1430,n1431);
and (n1499,n825,n1471);
and (n1500,n1501,n1502);
xor (n1501,n1498,n1499);
or (n1502,n1503,n1506);
and (n1503,n1504,n1505);
xor (n1504,n1436,n1437);
and (n1505,n832,n1471);
and (n1506,n1507,n1508);
xor (n1507,n1504,n1505);
or (n1508,n1509,n1512);
and (n1509,n1510,n1511);
xor (n1510,n1442,n1443);
and (n1511,n839,n1471);
and (n1512,n1513,n1514);
xor (n1513,n1510,n1511);
or (n1514,n1515,n1518);
and (n1515,n1516,n1517);
xor (n1516,n1448,n1449);
and (n1517,n846,n1471);
and (n1518,n1519,n1520);
xor (n1519,n1516,n1517);
or (n1520,n1521,n1524);
and (n1521,n1522,n1523);
xor (n1522,n1454,n1455);
and (n1523,n853,n1471);
and (n1524,n1525,n1526);
xor (n1525,n1522,n1523);
or (n1526,n1527,n1530);
and (n1527,n1528,n1529);
xor (n1528,n1460,n1461);
and (n1529,n860,n1471);
and (n1530,n1531,n1532);
xor (n1531,n1528,n1529);
and (n1532,n1533,n1534);
xor (n1533,n1466,n1467);
and (n1534,n866,n1471);
xor (n1536,n1537,n2240);
xor (n1537,n1538,n2238);
or (n1538,n1539,n2173);
and (n1539,n1540,n2171);
or (n1540,n1541,n2106);
and (n1541,n1542,n2104);
or (n1542,n1543,n2039);
and (n1543,n1544,n2037);
or (n1544,n1545,n1972);
and (n1545,n1546,n1970);
or (n1546,n1547,n1905);
and (n1547,n1548,n1903);
or (n1548,n1549,n1838);
and (n1549,n1550,n1836);
or (n1550,n1551,n1771);
and (n1551,n1552,n1769);
or (n1552,n1553,n1704);
and (n1553,n1554,n1702);
or (n1554,n1555,n1637);
and (n1555,n1556,n1635);
and (n1556,n1557,n1560);
and (n1557,n1558,n1559);
wire s0n1558,s1n1558,notn1558;
or (n1558,s0n1558,s1n1558);
not(notn1558,n1535);
and (s0n1558,notn1558,n23);
and (s1n1558,n1535,n790);
wire s0n1559,s1n1559,notn1559;
or (n1559,s0n1559,s1n1559);
not(notn1559,n1535);
and (s0n1559,notn1559,n24);
and (s1n1559,n1535,n791);
or (n1560,n1561,n1566);
and (n1561,n1562,n1564);
and (n1562,n1558,n1563);
wire s0n1563,s1n1563,notn1563;
or (n1563,s0n1563,s1n1563);
not(notn1563,n1535);
and (s0n1563,notn1563,n28);
and (s1n1563,n1535,n795);
and (n1564,n1565,n1559);
wire s0n1565,s1n1565,notn1565;
or (n1565,s0n1565,s1n1565);
not(notn1565,n1535);
and (s0n1565,notn1565,n30);
and (s1n1565,n1535,n797);
and (n1566,n1567,n1568);
xor (n1567,n1562,n1564);
or (n1568,n1569,n1573);
and (n1569,n1570,n1571);
and (n1570,n1565,n1563);
and (n1571,n1572,n1559);
wire s0n1572,s1n1572,notn1572;
or (n1572,s0n1572,s1n1572);
not(notn1572,n1535);
and (s0n1572,notn1572,n37);
and (s1n1572,n1535,n804);
and (n1573,n1574,n1575);
xor (n1574,n1570,n1571);
or (n1575,n1576,n1580);
and (n1576,n1577,n1578);
and (n1577,n1572,n1563);
and (n1578,n1579,n1559);
wire s0n1579,s1n1579,notn1579;
or (n1579,s0n1579,s1n1579);
not(notn1579,n1535);
and (s0n1579,notn1579,n44);
and (s1n1579,n1535,n811);
and (n1580,n1581,n1582);
xor (n1581,n1577,n1578);
or (n1582,n1583,n1587);
and (n1583,n1584,n1585);
and (n1584,n1579,n1563);
and (n1585,n1586,n1559);
wire s0n1586,s1n1586,notn1586;
or (n1586,s0n1586,s1n1586);
not(notn1586,n1535);
and (s0n1586,notn1586,n51);
and (s1n1586,n1535,n818);
and (n1587,n1588,n1589);
xor (n1588,n1584,n1585);
or (n1589,n1590,n1594);
and (n1590,n1591,n1592);
and (n1591,n1586,n1563);
and (n1592,n1593,n1559);
wire s0n1593,s1n1593,notn1593;
or (n1593,s0n1593,s1n1593);
not(notn1593,n1535);
and (s0n1593,notn1593,n58);
and (s1n1593,n1535,n825);
and (n1594,n1595,n1596);
xor (n1595,n1591,n1592);
or (n1596,n1597,n1601);
and (n1597,n1598,n1599);
and (n1598,n1593,n1563);
and (n1599,n1600,n1559);
wire s0n1600,s1n1600,notn1600;
or (n1600,s0n1600,s1n1600);
not(notn1600,n1535);
and (s0n1600,notn1600,n65);
and (s1n1600,n1535,n832);
and (n1601,n1602,n1603);
xor (n1602,n1598,n1599);
or (n1603,n1604,n1608);
and (n1604,n1605,n1606);
and (n1605,n1600,n1563);
and (n1606,n1607,n1559);
wire s0n1607,s1n1607,notn1607;
or (n1607,s0n1607,s1n1607);
not(notn1607,n1535);
and (s0n1607,notn1607,n72);
and (s1n1607,n1535,n839);
and (n1608,n1609,n1610);
xor (n1609,n1605,n1606);
or (n1610,n1611,n1615);
and (n1611,n1612,n1613);
and (n1612,n1607,n1563);
and (n1613,n1614,n1559);
wire s0n1614,s1n1614,notn1614;
or (n1614,s0n1614,s1n1614);
not(notn1614,n1535);
and (s0n1614,notn1614,n79);
and (s1n1614,n1535,n846);
and (n1615,n1616,n1617);
xor (n1616,n1612,n1613);
or (n1617,n1618,n1622);
and (n1618,n1619,n1620);
and (n1619,n1614,n1563);
and (n1620,n1621,n1559);
wire s0n1621,s1n1621,notn1621;
or (n1621,s0n1621,s1n1621);
not(notn1621,n1535);
and (s0n1621,notn1621,n86);
and (s1n1621,n1535,n853);
and (n1622,n1623,n1624);
xor (n1623,n1619,n1620);
or (n1624,n1625,n1629);
and (n1625,n1626,n1627);
and (n1626,n1621,n1563);
and (n1627,n1628,n1559);
wire s0n1628,s1n1628,notn1628;
or (n1628,s0n1628,s1n1628);
not(notn1628,n1535);
and (s0n1628,notn1628,n93);
and (s1n1628,n1535,n860);
and (n1629,n1630,n1631);
xor (n1630,n1626,n1627);
and (n1631,n1632,n1633);
and (n1632,n1628,n1563);
and (n1633,n1634,n1559);
wire s0n1634,s1n1634,notn1634;
or (n1634,s0n1634,s1n1634);
not(notn1634,n1535);
and (s0n1634,notn1634,n99);
and (s1n1634,n1535,n866);
and (n1635,n1558,n1636);
wire s0n1636,s1n1636,notn1636;
or (n1636,s0n1636,s1n1636);
not(notn1636,n1535);
and (s0n1636,notn1636,n101);
and (s1n1636,n1535,n868);
and (n1637,n1638,n1639);
xor (n1638,n1556,n1635);
or (n1639,n1640,n1643);
and (n1640,n1641,n1642);
xor (n1641,n1557,n1560);
and (n1642,n1565,n1636);
and (n1643,n1644,n1645);
xor (n1644,n1641,n1642);
or (n1645,n1646,n1649);
and (n1646,n1647,n1648);
xor (n1647,n1567,n1568);
and (n1648,n1572,n1636);
and (n1649,n1650,n1651);
xor (n1650,n1647,n1648);
or (n1651,n1652,n1655);
and (n1652,n1653,n1654);
xor (n1653,n1574,n1575);
and (n1654,n1579,n1636);
and (n1655,n1656,n1657);
xor (n1656,n1653,n1654);
or (n1657,n1658,n1661);
and (n1658,n1659,n1660);
xor (n1659,n1581,n1582);
and (n1660,n1586,n1636);
and (n1661,n1662,n1663);
xor (n1662,n1659,n1660);
or (n1663,n1664,n1667);
and (n1664,n1665,n1666);
xor (n1665,n1588,n1589);
and (n1666,n1593,n1636);
and (n1667,n1668,n1669);
xor (n1668,n1665,n1666);
or (n1669,n1670,n1673);
and (n1670,n1671,n1672);
xor (n1671,n1595,n1596);
and (n1672,n1600,n1636);
and (n1673,n1674,n1675);
xor (n1674,n1671,n1672);
or (n1675,n1676,n1679);
and (n1676,n1677,n1678);
xor (n1677,n1602,n1603);
and (n1678,n1607,n1636);
and (n1679,n1680,n1681);
xor (n1680,n1677,n1678);
or (n1681,n1682,n1685);
and (n1682,n1683,n1684);
xor (n1683,n1609,n1610);
and (n1684,n1614,n1636);
and (n1685,n1686,n1687);
xor (n1686,n1683,n1684);
or (n1687,n1688,n1691);
and (n1688,n1689,n1690);
xor (n1689,n1616,n1617);
and (n1690,n1621,n1636);
and (n1691,n1692,n1693);
xor (n1692,n1689,n1690);
or (n1693,n1694,n1697);
and (n1694,n1695,n1696);
xor (n1695,n1623,n1624);
and (n1696,n1628,n1636);
and (n1697,n1698,n1699);
xor (n1698,n1695,n1696);
and (n1699,n1700,n1701);
xor (n1700,n1630,n1631);
and (n1701,n1634,n1636);
and (n1702,n1558,n1703);
wire s0n1703,s1n1703,notn1703;
or (n1703,s0n1703,s1n1703);
not(notn1703,n1535);
and (s0n1703,notn1703,n168);
and (s1n1703,n1535,n935);
and (n1704,n1705,n1706);
xor (n1705,n1554,n1702);
or (n1706,n1707,n1710);
and (n1707,n1708,n1709);
xor (n1708,n1638,n1639);
and (n1709,n1565,n1703);
and (n1710,n1711,n1712);
xor (n1711,n1708,n1709);
or (n1712,n1713,n1716);
and (n1713,n1714,n1715);
xor (n1714,n1644,n1645);
and (n1715,n1572,n1703);
and (n1716,n1717,n1718);
xor (n1717,n1714,n1715);
or (n1718,n1719,n1722);
and (n1719,n1720,n1721);
xor (n1720,n1650,n1651);
and (n1721,n1579,n1703);
and (n1722,n1723,n1724);
xor (n1723,n1720,n1721);
or (n1724,n1725,n1728);
and (n1725,n1726,n1727);
xor (n1726,n1656,n1657);
and (n1727,n1586,n1703);
and (n1728,n1729,n1730);
xor (n1729,n1726,n1727);
or (n1730,n1731,n1734);
and (n1731,n1732,n1733);
xor (n1732,n1662,n1663);
and (n1733,n1593,n1703);
and (n1734,n1735,n1736);
xor (n1735,n1732,n1733);
or (n1736,n1737,n1740);
and (n1737,n1738,n1739);
xor (n1738,n1668,n1669);
and (n1739,n1600,n1703);
and (n1740,n1741,n1742);
xor (n1741,n1738,n1739);
or (n1742,n1743,n1746);
and (n1743,n1744,n1745);
xor (n1744,n1674,n1675);
and (n1745,n1607,n1703);
and (n1746,n1747,n1748);
xor (n1747,n1744,n1745);
or (n1748,n1749,n1752);
and (n1749,n1750,n1751);
xor (n1750,n1680,n1681);
and (n1751,n1614,n1703);
and (n1752,n1753,n1754);
xor (n1753,n1750,n1751);
or (n1754,n1755,n1758);
and (n1755,n1756,n1757);
xor (n1756,n1686,n1687);
and (n1757,n1621,n1703);
and (n1758,n1759,n1760);
xor (n1759,n1756,n1757);
or (n1760,n1761,n1764);
and (n1761,n1762,n1763);
xor (n1762,n1692,n1693);
and (n1763,n1628,n1703);
and (n1764,n1765,n1766);
xor (n1765,n1762,n1763);
and (n1766,n1767,n1768);
xor (n1767,n1698,n1699);
and (n1768,n1634,n1703);
and (n1769,n1558,n1770);
wire s0n1770,s1n1770,notn1770;
or (n1770,s0n1770,s1n1770);
not(notn1770,n1535);
and (s0n1770,notn1770,n235);
and (s1n1770,n1535,n1002);
and (n1771,n1772,n1773);
xor (n1772,n1552,n1769);
or (n1773,n1774,n1777);
and (n1774,n1775,n1776);
xor (n1775,n1705,n1706);
and (n1776,n1565,n1770);
and (n1777,n1778,n1779);
xor (n1778,n1775,n1776);
or (n1779,n1780,n1783);
and (n1780,n1781,n1782);
xor (n1781,n1711,n1712);
and (n1782,n1572,n1770);
and (n1783,n1784,n1785);
xor (n1784,n1781,n1782);
or (n1785,n1786,n1789);
and (n1786,n1787,n1788);
xor (n1787,n1717,n1718);
and (n1788,n1579,n1770);
and (n1789,n1790,n1791);
xor (n1790,n1787,n1788);
or (n1791,n1792,n1795);
and (n1792,n1793,n1794);
xor (n1793,n1723,n1724);
and (n1794,n1586,n1770);
and (n1795,n1796,n1797);
xor (n1796,n1793,n1794);
or (n1797,n1798,n1801);
and (n1798,n1799,n1800);
xor (n1799,n1729,n1730);
and (n1800,n1593,n1770);
and (n1801,n1802,n1803);
xor (n1802,n1799,n1800);
or (n1803,n1804,n1807);
and (n1804,n1805,n1806);
xor (n1805,n1735,n1736);
and (n1806,n1600,n1770);
and (n1807,n1808,n1809);
xor (n1808,n1805,n1806);
or (n1809,n1810,n1813);
and (n1810,n1811,n1812);
xor (n1811,n1741,n1742);
and (n1812,n1607,n1770);
and (n1813,n1814,n1815);
xor (n1814,n1811,n1812);
or (n1815,n1816,n1819);
and (n1816,n1817,n1818);
xor (n1817,n1747,n1748);
and (n1818,n1614,n1770);
and (n1819,n1820,n1821);
xor (n1820,n1817,n1818);
or (n1821,n1822,n1825);
and (n1822,n1823,n1824);
xor (n1823,n1753,n1754);
and (n1824,n1621,n1770);
and (n1825,n1826,n1827);
xor (n1826,n1823,n1824);
or (n1827,n1828,n1831);
and (n1828,n1829,n1830);
xor (n1829,n1759,n1760);
and (n1830,n1628,n1770);
and (n1831,n1832,n1833);
xor (n1832,n1829,n1830);
and (n1833,n1834,n1835);
xor (n1834,n1765,n1766);
and (n1835,n1634,n1770);
and (n1836,n1558,n1837);
wire s0n1837,s1n1837,notn1837;
or (n1837,s0n1837,s1n1837);
not(notn1837,n1535);
and (s0n1837,notn1837,n302);
and (s1n1837,n1535,n1069);
and (n1838,n1839,n1840);
xor (n1839,n1550,n1836);
or (n1840,n1841,n1844);
and (n1841,n1842,n1843);
xor (n1842,n1772,n1773);
and (n1843,n1565,n1837);
and (n1844,n1845,n1846);
xor (n1845,n1842,n1843);
or (n1846,n1847,n1850);
and (n1847,n1848,n1849);
xor (n1848,n1778,n1779);
and (n1849,n1572,n1837);
and (n1850,n1851,n1852);
xor (n1851,n1848,n1849);
or (n1852,n1853,n1856);
and (n1853,n1854,n1855);
xor (n1854,n1784,n1785);
and (n1855,n1579,n1837);
and (n1856,n1857,n1858);
xor (n1857,n1854,n1855);
or (n1858,n1859,n1862);
and (n1859,n1860,n1861);
xor (n1860,n1790,n1791);
and (n1861,n1586,n1837);
and (n1862,n1863,n1864);
xor (n1863,n1860,n1861);
or (n1864,n1865,n1868);
and (n1865,n1866,n1867);
xor (n1866,n1796,n1797);
and (n1867,n1593,n1837);
and (n1868,n1869,n1870);
xor (n1869,n1866,n1867);
or (n1870,n1871,n1874);
and (n1871,n1872,n1873);
xor (n1872,n1802,n1803);
and (n1873,n1600,n1837);
and (n1874,n1875,n1876);
xor (n1875,n1872,n1873);
or (n1876,n1877,n1880);
and (n1877,n1878,n1879);
xor (n1878,n1808,n1809);
and (n1879,n1607,n1837);
and (n1880,n1881,n1882);
xor (n1881,n1878,n1879);
or (n1882,n1883,n1886);
and (n1883,n1884,n1885);
xor (n1884,n1814,n1815);
and (n1885,n1614,n1837);
and (n1886,n1887,n1888);
xor (n1887,n1884,n1885);
or (n1888,n1889,n1892);
and (n1889,n1890,n1891);
xor (n1890,n1820,n1821);
and (n1891,n1621,n1837);
and (n1892,n1893,n1894);
xor (n1893,n1890,n1891);
or (n1894,n1895,n1898);
and (n1895,n1896,n1897);
xor (n1896,n1826,n1827);
and (n1897,n1628,n1837);
and (n1898,n1899,n1900);
xor (n1899,n1896,n1897);
and (n1900,n1901,n1902);
xor (n1901,n1832,n1833);
and (n1902,n1634,n1837);
and (n1903,n1558,n1904);
wire s0n1904,s1n1904,notn1904;
or (n1904,s0n1904,s1n1904);
not(notn1904,n1535);
and (s0n1904,notn1904,n369);
and (s1n1904,n1535,n1136);
and (n1905,n1906,n1907);
xor (n1906,n1548,n1903);
or (n1907,n1908,n1911);
and (n1908,n1909,n1910);
xor (n1909,n1839,n1840);
and (n1910,n1565,n1904);
and (n1911,n1912,n1913);
xor (n1912,n1909,n1910);
or (n1913,n1914,n1917);
and (n1914,n1915,n1916);
xor (n1915,n1845,n1846);
and (n1916,n1572,n1904);
and (n1917,n1918,n1919);
xor (n1918,n1915,n1916);
or (n1919,n1920,n1923);
and (n1920,n1921,n1922);
xor (n1921,n1851,n1852);
and (n1922,n1579,n1904);
and (n1923,n1924,n1925);
xor (n1924,n1921,n1922);
or (n1925,n1926,n1929);
and (n1926,n1927,n1928);
xor (n1927,n1857,n1858);
and (n1928,n1586,n1904);
and (n1929,n1930,n1931);
xor (n1930,n1927,n1928);
or (n1931,n1932,n1935);
and (n1932,n1933,n1934);
xor (n1933,n1863,n1864);
and (n1934,n1593,n1904);
and (n1935,n1936,n1937);
xor (n1936,n1933,n1934);
or (n1937,n1938,n1941);
and (n1938,n1939,n1940);
xor (n1939,n1869,n1870);
and (n1940,n1600,n1904);
and (n1941,n1942,n1943);
xor (n1942,n1939,n1940);
or (n1943,n1944,n1947);
and (n1944,n1945,n1946);
xor (n1945,n1875,n1876);
and (n1946,n1607,n1904);
and (n1947,n1948,n1949);
xor (n1948,n1945,n1946);
or (n1949,n1950,n1953);
and (n1950,n1951,n1952);
xor (n1951,n1881,n1882);
and (n1952,n1614,n1904);
and (n1953,n1954,n1955);
xor (n1954,n1951,n1952);
or (n1955,n1956,n1959);
and (n1956,n1957,n1958);
xor (n1957,n1887,n1888);
and (n1958,n1621,n1904);
and (n1959,n1960,n1961);
xor (n1960,n1957,n1958);
or (n1961,n1962,n1965);
and (n1962,n1963,n1964);
xor (n1963,n1893,n1894);
and (n1964,n1628,n1904);
and (n1965,n1966,n1967);
xor (n1966,n1963,n1964);
and (n1967,n1968,n1969);
xor (n1968,n1899,n1900);
and (n1969,n1634,n1904);
and (n1970,n1558,n1971);
wire s0n1971,s1n1971,notn1971;
or (n1971,s0n1971,s1n1971);
not(notn1971,n1535);
and (s0n1971,notn1971,n436);
and (s1n1971,n1535,n1203);
and (n1972,n1973,n1974);
xor (n1973,n1546,n1970);
or (n1974,n1975,n1978);
and (n1975,n1976,n1977);
xor (n1976,n1906,n1907);
and (n1977,n1565,n1971);
and (n1978,n1979,n1980);
xor (n1979,n1976,n1977);
or (n1980,n1981,n1984);
and (n1981,n1982,n1983);
xor (n1982,n1912,n1913);
and (n1983,n1572,n1971);
and (n1984,n1985,n1986);
xor (n1985,n1982,n1983);
or (n1986,n1987,n1990);
and (n1987,n1988,n1989);
xor (n1988,n1918,n1919);
and (n1989,n1579,n1971);
and (n1990,n1991,n1992);
xor (n1991,n1988,n1989);
or (n1992,n1993,n1996);
and (n1993,n1994,n1995);
xor (n1994,n1924,n1925);
and (n1995,n1586,n1971);
and (n1996,n1997,n1998);
xor (n1997,n1994,n1995);
or (n1998,n1999,n2002);
and (n1999,n2000,n2001);
xor (n2000,n1930,n1931);
and (n2001,n1593,n1971);
and (n2002,n2003,n2004);
xor (n2003,n2000,n2001);
or (n2004,n2005,n2008);
and (n2005,n2006,n2007);
xor (n2006,n1936,n1937);
and (n2007,n1600,n1971);
and (n2008,n2009,n2010);
xor (n2009,n2006,n2007);
or (n2010,n2011,n2014);
and (n2011,n2012,n2013);
xor (n2012,n1942,n1943);
and (n2013,n1607,n1971);
and (n2014,n2015,n2016);
xor (n2015,n2012,n2013);
or (n2016,n2017,n2020);
and (n2017,n2018,n2019);
xor (n2018,n1948,n1949);
and (n2019,n1614,n1971);
and (n2020,n2021,n2022);
xor (n2021,n2018,n2019);
or (n2022,n2023,n2026);
and (n2023,n2024,n2025);
xor (n2024,n1954,n1955);
and (n2025,n1621,n1971);
and (n2026,n2027,n2028);
xor (n2027,n2024,n2025);
or (n2028,n2029,n2032);
and (n2029,n2030,n2031);
xor (n2030,n1960,n1961);
and (n2031,n1628,n1971);
and (n2032,n2033,n2034);
xor (n2033,n2030,n2031);
and (n2034,n2035,n2036);
xor (n2035,n1966,n1967);
and (n2036,n1634,n1971);
and (n2037,n1558,n2038);
wire s0n2038,s1n2038,notn2038;
or (n2038,s0n2038,s1n2038);
not(notn2038,n1535);
and (s0n2038,notn2038,n503);
and (s1n2038,n1535,n1270);
and (n2039,n2040,n2041);
xor (n2040,n1544,n2037);
or (n2041,n2042,n2045);
and (n2042,n2043,n2044);
xor (n2043,n1973,n1974);
and (n2044,n1565,n2038);
and (n2045,n2046,n2047);
xor (n2046,n2043,n2044);
or (n2047,n2048,n2051);
and (n2048,n2049,n2050);
xor (n2049,n1979,n1980);
and (n2050,n1572,n2038);
and (n2051,n2052,n2053);
xor (n2052,n2049,n2050);
or (n2053,n2054,n2057);
and (n2054,n2055,n2056);
xor (n2055,n1985,n1986);
and (n2056,n1579,n2038);
and (n2057,n2058,n2059);
xor (n2058,n2055,n2056);
or (n2059,n2060,n2063);
and (n2060,n2061,n2062);
xor (n2061,n1991,n1992);
and (n2062,n1586,n2038);
and (n2063,n2064,n2065);
xor (n2064,n2061,n2062);
or (n2065,n2066,n2069);
and (n2066,n2067,n2068);
xor (n2067,n1997,n1998);
and (n2068,n1593,n2038);
and (n2069,n2070,n2071);
xor (n2070,n2067,n2068);
or (n2071,n2072,n2075);
and (n2072,n2073,n2074);
xor (n2073,n2003,n2004);
and (n2074,n1600,n2038);
and (n2075,n2076,n2077);
xor (n2076,n2073,n2074);
or (n2077,n2078,n2081);
and (n2078,n2079,n2080);
xor (n2079,n2009,n2010);
and (n2080,n1607,n2038);
and (n2081,n2082,n2083);
xor (n2082,n2079,n2080);
or (n2083,n2084,n2087);
and (n2084,n2085,n2086);
xor (n2085,n2015,n2016);
and (n2086,n1614,n2038);
and (n2087,n2088,n2089);
xor (n2088,n2085,n2086);
or (n2089,n2090,n2093);
and (n2090,n2091,n2092);
xor (n2091,n2021,n2022);
and (n2092,n1621,n2038);
and (n2093,n2094,n2095);
xor (n2094,n2091,n2092);
or (n2095,n2096,n2099);
and (n2096,n2097,n2098);
xor (n2097,n2027,n2028);
and (n2098,n1628,n2038);
and (n2099,n2100,n2101);
xor (n2100,n2097,n2098);
and (n2101,n2102,n2103);
xor (n2102,n2033,n2034);
and (n2103,n1634,n2038);
and (n2104,n1558,n2105);
wire s0n2105,s1n2105,notn2105;
or (n2105,s0n2105,s1n2105);
not(notn2105,n1535);
and (s0n2105,notn2105,n570);
and (s1n2105,n1535,n1337);
and (n2106,n2107,n2108);
xor (n2107,n1542,n2104);
or (n2108,n2109,n2112);
and (n2109,n2110,n2111);
xor (n2110,n2040,n2041);
and (n2111,n1565,n2105);
and (n2112,n2113,n2114);
xor (n2113,n2110,n2111);
or (n2114,n2115,n2118);
and (n2115,n2116,n2117);
xor (n2116,n2046,n2047);
and (n2117,n1572,n2105);
and (n2118,n2119,n2120);
xor (n2119,n2116,n2117);
or (n2120,n2121,n2124);
and (n2121,n2122,n2123);
xor (n2122,n2052,n2053);
and (n2123,n1579,n2105);
and (n2124,n2125,n2126);
xor (n2125,n2122,n2123);
or (n2126,n2127,n2130);
and (n2127,n2128,n2129);
xor (n2128,n2058,n2059);
and (n2129,n1586,n2105);
and (n2130,n2131,n2132);
xor (n2131,n2128,n2129);
or (n2132,n2133,n2136);
and (n2133,n2134,n2135);
xor (n2134,n2064,n2065);
and (n2135,n1593,n2105);
and (n2136,n2137,n2138);
xor (n2137,n2134,n2135);
or (n2138,n2139,n2142);
and (n2139,n2140,n2141);
xor (n2140,n2070,n2071);
and (n2141,n1600,n2105);
and (n2142,n2143,n2144);
xor (n2143,n2140,n2141);
or (n2144,n2145,n2148);
and (n2145,n2146,n2147);
xor (n2146,n2076,n2077);
and (n2147,n1607,n2105);
and (n2148,n2149,n2150);
xor (n2149,n2146,n2147);
or (n2150,n2151,n2154);
and (n2151,n2152,n2153);
xor (n2152,n2082,n2083);
and (n2153,n1614,n2105);
and (n2154,n2155,n2156);
xor (n2155,n2152,n2153);
or (n2156,n2157,n2160);
and (n2157,n2158,n2159);
xor (n2158,n2088,n2089);
and (n2159,n1621,n2105);
and (n2160,n2161,n2162);
xor (n2161,n2158,n2159);
or (n2162,n2163,n2166);
and (n2163,n2164,n2165);
xor (n2164,n2094,n2095);
and (n2165,n1628,n2105);
and (n2166,n2167,n2168);
xor (n2167,n2164,n2165);
and (n2168,n2169,n2170);
xor (n2169,n2100,n2101);
and (n2170,n1634,n2105);
and (n2171,n1558,n2172);
wire s0n2172,s1n2172,notn2172;
or (n2172,s0n2172,s1n2172);
not(notn2172,n1535);
and (s0n2172,notn2172,n637);
and (s1n2172,n1535,n1404);
and (n2173,n2174,n2175);
xor (n2174,n1540,n2171);
or (n2175,n2176,n2179);
and (n2176,n2177,n2178);
xor (n2177,n2107,n2108);
and (n2178,n1565,n2172);
and (n2179,n2180,n2181);
xor (n2180,n2177,n2178);
or (n2181,n2182,n2185);
and (n2182,n2183,n2184);
xor (n2183,n2113,n2114);
and (n2184,n1572,n2172);
and (n2185,n2186,n2187);
xor (n2186,n2183,n2184);
or (n2187,n2188,n2191);
and (n2188,n2189,n2190);
xor (n2189,n2119,n2120);
and (n2190,n1579,n2172);
and (n2191,n2192,n2193);
xor (n2192,n2189,n2190);
or (n2193,n2194,n2197);
and (n2194,n2195,n2196);
xor (n2195,n2125,n2126);
and (n2196,n1586,n2172);
and (n2197,n2198,n2199);
xor (n2198,n2195,n2196);
or (n2199,n2200,n2203);
and (n2200,n2201,n2202);
xor (n2201,n2131,n2132);
and (n2202,n1593,n2172);
and (n2203,n2204,n2205);
xor (n2204,n2201,n2202);
or (n2205,n2206,n2209);
and (n2206,n2207,n2208);
xor (n2207,n2137,n2138);
and (n2208,n1600,n2172);
and (n2209,n2210,n2211);
xor (n2210,n2207,n2208);
or (n2211,n2212,n2215);
and (n2212,n2213,n2214);
xor (n2213,n2143,n2144);
and (n2214,n1607,n2172);
and (n2215,n2216,n2217);
xor (n2216,n2213,n2214);
or (n2217,n2218,n2221);
and (n2218,n2219,n2220);
xor (n2219,n2149,n2150);
and (n2220,n1614,n2172);
and (n2221,n2222,n2223);
xor (n2222,n2219,n2220);
or (n2223,n2224,n2227);
and (n2224,n2225,n2226);
xor (n2225,n2155,n2156);
and (n2226,n1621,n2172);
and (n2227,n2228,n2229);
xor (n2228,n2225,n2226);
or (n2229,n2230,n2233);
and (n2230,n2231,n2232);
xor (n2231,n2161,n2162);
and (n2232,n1628,n2172);
and (n2233,n2234,n2235);
xor (n2234,n2231,n2232);
and (n2235,n2236,n2237);
xor (n2236,n2167,n2168);
and (n2237,n1634,n2172);
and (n2238,n1558,n2239);
wire s0n2239,s1n2239,notn2239;
or (n2239,s0n2239,s1n2239);
not(notn2239,n1535);
and (s0n2239,notn2239,n704);
and (s1n2239,n1535,n1471);
or (n2240,n2241,n2244);
and (n2241,n2242,n2243);
xor (n2242,n2174,n2175);
and (n2243,n1565,n2239);
and (n2244,n2245,n2246);
xor (n2245,n2242,n2243);
or (n2246,n2247,n2250);
and (n2247,n2248,n2249);
xor (n2248,n2180,n2181);
and (n2249,n1572,n2239);
and (n2250,n2251,n2252);
xor (n2251,n2248,n2249);
or (n2252,n2253,n2256);
and (n2253,n2254,n2255);
xor (n2254,n2186,n2187);
and (n2255,n1579,n2239);
and (n2256,n2257,n2258);
xor (n2257,n2254,n2255);
or (n2258,n2259,n2262);
and (n2259,n2260,n2261);
xor (n2260,n2192,n2193);
and (n2261,n1586,n2239);
and (n2262,n2263,n2264);
xor (n2263,n2260,n2261);
or (n2264,n2265,n2268);
and (n2265,n2266,n2267);
xor (n2266,n2198,n2199);
and (n2267,n1593,n2239);
and (n2268,n2269,n2270);
xor (n2269,n2266,n2267);
or (n2270,n2271,n2274);
and (n2271,n2272,n2273);
xor (n2272,n2204,n2205);
and (n2273,n1600,n2239);
and (n2274,n2275,n2276);
xor (n2275,n2272,n2273);
or (n2276,n2277,n2280);
and (n2277,n2278,n2279);
xor (n2278,n2210,n2211);
and (n2279,n1607,n2239);
and (n2280,n2281,n2282);
xor (n2281,n2278,n2279);
or (n2282,n2283,n2286);
and (n2283,n2284,n2285);
xor (n2284,n2216,n2217);
and (n2285,n1614,n2239);
and (n2286,n2287,n2288);
xor (n2287,n2284,n2285);
or (n2288,n2289,n2292);
and (n2289,n2290,n2291);
xor (n2290,n2222,n2223);
and (n2291,n1621,n2239);
and (n2292,n2293,n2294);
xor (n2293,n2290,n2291);
or (n2294,n2295,n2298);
and (n2295,n2296,n2297);
xor (n2296,n2228,n2229);
and (n2297,n1628,n2239);
and (n2298,n2299,n2300);
xor (n2299,n2296,n2297);
and (n2300,n2301,n2302);
xor (n2301,n2234,n2235);
and (n2302,n1634,n2239);
endmodule
