module top (out,n3,n18,n20,n21,n30,n31,n33,n34,n44
        ,n53,n57,n67,n68,n70,n71,n78,n84,n96,n97
        ,n99,n100,n103,n109,n121,n122,n131,n137,n167,n191
        ,n226,n511,n517,n535,n541);
output out;
input n3;
input n18;
input n20;
input n21;
input n30;
input n31;
input n33;
input n34;
input n44;
input n53;
input n57;
input n67;
input n68;
input n70;
input n71;
input n78;
input n84;
input n96;
input n97;
input n99;
input n100;
input n103;
input n109;
input n121;
input n122;
input n131;
input n137;
input n167;
input n191;
input n226;
input n511;
input n517;
input n535;
input n541;
wire n0;
wire n1;
wire n2;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n19;
wire n22;
wire n23;
wire n24;
wire n25;
wire n26;
wire n27;
wire n28;
wire n29;
wire n32;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n52;
wire n54;
wire n55;
wire n56;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n69;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n98;
wire n101;
wire n102;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
xor (out,n0,n913);
nand (n0,n1,n495);
or (n1,n2,n4);
not (n2,n3);
not (n4,n5);
xnor (n5,n6,n243);
nand (n6,n7,n242);
nand (n7,n8,n200);
not (n8,n9);
xor (n9,n10,n176);
xor (n10,n11,n87);
xor (n11,n12,n59);
xor (n12,n13,n47);
nand (n13,n14,n40);
or (n14,n15,n25);
not (n15,n16);
nor (n16,n17,n22);
and (n17,n18,n19);
wire s0n19,s1n19,notn19;
or (n19,s0n19,s1n19);
not(notn19,n3);
and (s0n19,notn19,n20);
and (s1n19,n3,n21);
and (n22,n23,n24);
not (n23,n18);
not (n24,n19);
nand (n25,n26,n37);
nor (n26,n27,n35);
and (n27,n28,n32);
not (n28,n29);
wire s0n29,s1n29,notn29;
or (n29,s0n29,s1n29);
not(notn29,n3);
and (s0n29,notn29,n30);
and (s1n29,n3,n31);
wire s0n32,s1n32,notn32;
or (n32,s0n32,s1n32);
not(notn32,n3);
and (s0n32,notn32,n33);
and (s1n32,n3,n34);
and (n35,n29,n36);
not (n36,n32);
nand (n37,n38,n39);
or (n38,n28,n19);
nand (n39,n19,n28);
nand (n40,n41,n42);
not (n41,n26);
nor (n42,n43,n45);
and (n43,n44,n19);
and (n45,n46,n24);
not (n46,n44);
nor (n47,n48,n54);
nand (n48,n19,n49);
not (n49,n50);
wire s0n50,s1n50,notn50;
or (n50,s0n50,s1n50);
not(notn50,n3);
and (s0n50,notn50,1'b0);
and (s1n50,n3,n52);
and (n52,n53,n21);
nor (n54,n55,n58);
and (n55,n50,n56);
not (n56,n57);
and (n58,n49,n57);
nand (n59,n60,n81);
or (n60,n61,n76);
nand (n61,n62,n73);
not (n62,n63);
nand (n63,n64,n72);
or (n64,n65,n69);
not (n65,n66);
wire s0n66,s1n66,notn66;
or (n66,s0n66,s1n66);
not(notn66,n3);
and (s0n66,notn66,n67);
and (s1n66,n3,n68);
wire s0n69,s1n69,notn69;
or (n69,s0n69,s1n69);
not(notn69,n3);
and (s0n69,notn69,n70);
and (s1n69,n3,n71);
nand (n72,n69,n65);
nand (n73,n74,n75);
or (n74,n65,n32);
nand (n75,n32,n65);
nor (n76,n77,n79);
and (n77,n36,n78);
and (n79,n32,n80);
not (n80,n78);
or (n81,n62,n82);
nor (n82,n83,n85);
and (n83,n36,n84);
and (n85,n32,n86);
not (n86,n84);
xor (n87,n88,n153);
xor (n88,n89,n140);
xor (n89,n90,n113);
nand (n90,n91,n106);
or (n91,n92,n101);
not (n92,n93);
nor (n93,n94,n98);
not (n94,n95);
wire s0n95,s1n95,notn95;
or (n95,s0n95,s1n95);
not(notn95,n3);
and (s0n95,notn95,n96);
and (s1n95,n3,n97);
wire s0n98,s1n98,notn98;
or (n98,s0n98,s1n98);
not(notn98,n3);
and (s0n98,notn98,n99);
and (s1n98,n3,n100);
nor (n101,n102,n104);
and (n102,n94,n103);
and (n104,n95,n105);
not (n105,n103);
or (n106,n107,n112);
nor (n107,n108,n110);
and (n108,n94,n109);
and (n110,n95,n111);
not (n111,n109);
not (n112,n98);
nand (n113,n114,n134);
or (n114,n115,n128);
not (n115,n116);
and (n116,n117,n124);
nand (n117,n118,n123);
or (n118,n119,n69);
not (n119,n120);
wire s0n120,s1n120,notn120;
or (n120,s0n120,s1n120);
not(notn120,n3);
and (s0n120,notn120,n121);
and (s1n120,n3,n122);
nand (n123,n69,n119);
not (n124,n125);
nand (n125,n126,n127);
or (n126,n119,n95);
nand (n127,n95,n119);
nor (n128,n129,n132);
and (n129,n130,n131);
not (n130,n69);
and (n132,n69,n133);
not (n133,n131);
or (n134,n124,n135);
nor (n135,n136,n138);
and (n136,n130,n137);
and (n138,n69,n139);
not (n139,n137);
and (n140,n141,n147);
nand (n141,n142,n146);
or (n142,n92,n143);
nor (n143,n144,n145);
and (n144,n94,n137);
and (n145,n95,n139);
or (n146,n101,n112);
nand (n147,n148,n152);
or (n148,n115,n149);
nor (n149,n150,n151);
and (n150,n130,n84);
and (n151,n69,n86);
or (n152,n128,n124);
or (n153,n154,n175);
and (n154,n155,n169);
xor (n155,n156,n163);
nand (n156,n157,n162);
or (n157,n158,n25);
not (n158,n159);
nor (n159,n160,n161);
and (n160,n57,n19);
and (n161,n56,n24);
nand (n162,n41,n16);
nor (n163,n48,n164);
nor (n164,n165,n168);
and (n165,n50,n166);
not (n166,n167);
and (n168,n49,n167);
nand (n169,n170,n174);
or (n170,n61,n171);
nor (n171,n172,n173);
and (n172,n36,n44);
and (n173,n32,n46);
or (n174,n62,n76);
and (n175,n156,n163);
and (n176,n177,n178);
xor (n177,n141,n147);
or (n178,n179,n199);
and (n179,n180,n193);
xor (n180,n181,n187);
nand (n181,n182,n186);
or (n182,n183,n25);
nor (n183,n184,n185);
and (n184,n167,n24);
and (n185,n166,n19);
nand (n186,n159,n41);
nor (n187,n48,n188);
nor (n188,n189,n192);
and (n189,n50,n190);
not (n190,n191);
and (n192,n49,n191);
nand (n193,n194,n198);
or (n194,n92,n195);
nor (n195,n196,n197);
and (n196,n94,n131);
and (n197,n95,n133);
or (n198,n143,n112);
and (n199,n181,n187);
not (n200,n201);
or (n201,n202,n241);
and (n202,n203,n206);
xor (n203,n204,n205);
xor (n204,n155,n169);
xor (n205,n177,n178);
or (n206,n207,n240);
and (n207,n208,n221);
xor (n208,n209,n215);
nand (n209,n210,n214);
or (n210,n61,n211);
nor (n211,n212,n213);
and (n212,n36,n18);
and (n213,n32,n23);
or (n214,n62,n171);
nand (n215,n216,n220);
or (n216,n115,n217);
nor (n217,n218,n219);
and (n218,n130,n78);
and (n219,n69,n80);
or (n220,n149,n124);
or (n221,n222,n239);
and (n222,n223,n233);
xor (n223,n224,n227);
and (n224,n225,n226);
not (n225,n48);
nand (n227,n228,n232);
or (n228,n92,n229);
nor (n229,n230,n231);
and (n230,n86,n95);
and (n231,n84,n94);
or (n232,n195,n112);
nand (n233,n234,n238);
or (n234,n25,n235);
nor (n235,n236,n237);
and (n236,n191,n24);
and (n237,n190,n19);
or (n238,n26,n183);
and (n239,n224,n227);
and (n240,n209,n215);
and (n241,n204,n205);
nand (n242,n9,n201);
nand (n243,n244,n494);
or (n244,n245,n285);
nor (n245,n246,n247);
xor (n246,n203,n206);
or (n247,n248,n284);
and (n248,n249,n283);
xor (n249,n250,n251);
xor (n250,n180,n193);
or (n251,n252,n282);
and (n252,n253,n267);
xor (n253,n254,n261);
nand (n254,n255,n260);
or (n255,n115,n256);
not (n256,n257);
nor (n257,n258,n259);
and (n258,n44,n69);
and (n259,n46,n130);
or (n260,n124,n217);
nand (n261,n262,n266);
or (n262,n61,n263);
nor (n263,n264,n265);
and (n264,n36,n57);
and (n265,n32,n56);
or (n266,n62,n211);
and (n267,n268,n274);
nor (n268,n269,n24);
nor (n269,n270,n272);
and (n270,n36,n271);
nand (n271,n29,n226);
and (n272,n28,n273);
not (n273,n226);
nand (n274,n275,n280);
or (n275,n276,n92);
not (n276,n277);
nor (n277,n278,n279);
and (n278,n78,n95);
and (n279,n80,n94);
nand (n280,n281,n98);
not (n281,n229);
and (n282,n254,n261);
xor (n283,n208,n221);
and (n284,n250,n251);
not (n285,n286);
nand (n286,n287,n489);
not (n287,n288);
nor (n288,n289,n470);
nor (n289,n290,n468);
and (n290,n291,n442);
or (n291,n292,n441);
and (n292,n293,n357);
xor (n293,n294,n334);
or (n294,n295,n333);
and (n295,n296,n318);
xor (n296,n297,n307);
nand (n297,n298,n303);
or (n298,n299,n115);
not (n299,n300);
nor (n300,n301,n302);
and (n301,n166,n130);
and (n302,n167,n69);
nand (n303,n125,n304);
nor (n304,n305,n306);
and (n305,n57,n69);
and (n306,n130,n56);
nand (n307,n308,n313);
or (n308,n309,n62);
not (n309,n310);
nor (n310,n311,n312);
and (n311,n191,n32);
and (n312,n190,n36);
nand (n313,n314,n315);
not (n314,n61);
nand (n315,n316,n317);
or (n316,n36,n226);
or (n317,n32,n273);
xor (n318,n319,n324);
and (n319,n320,n32);
nand (n320,n321,n323);
or (n321,n69,n322);
and (n322,n226,n66);
or (n323,n66,n226);
nand (n324,n325,n329);
or (n325,n92,n326);
nor (n326,n327,n328);
and (n327,n94,n18);
and (n328,n95,n23);
or (n329,n330,n112);
nor (n330,n331,n332);
and (n331,n44,n94);
and (n332,n46,n95);
and (n333,n297,n307);
xor (n334,n335,n343);
xor (n335,n336,n342);
nand (n336,n337,n338);
or (n337,n309,n61);
or (n338,n62,n339);
nor (n339,n340,n341);
and (n340,n36,n167);
and (n341,n32,n166);
and (n342,n319,n324);
xor (n343,n344,n350);
xor (n344,n345,n346);
and (n345,n41,n226);
nand (n346,n347,n348);
or (n347,n112,n276);
nand (n348,n349,n93);
not (n349,n330);
nand (n350,n351,n353);
or (n351,n352,n115);
not (n352,n304);
nand (n353,n125,n354);
nand (n354,n355,n356);
or (n355,n69,n23);
or (n356,n130,n18);
or (n357,n358,n440);
and (n358,n359,n380);
xor (n359,n360,n379);
or (n360,n361,n378);
and (n361,n362,n371);
xor (n362,n363,n364);
and (n363,n63,n226);
nand (n364,n365,n370);
or (n365,n366,n115);
not (n366,n367);
nor (n367,n368,n369);
and (n368,n191,n69);
and (n369,n190,n130);
nand (n370,n300,n125);
nand (n371,n372,n377);
or (n372,n92,n373);
not (n373,n374);
nor (n374,n375,n376);
and (n375,n56,n94);
and (n376,n57,n95);
or (n377,n326,n112);
and (n378,n363,n364);
xor (n379,n296,n318);
or (n380,n381,n439);
and (n381,n382,n438);
xor (n382,n383,n397);
nor (n383,n384,n392);
not (n384,n385);
nand (n385,n386,n391);
or (n386,n387,n92);
not (n387,n388);
nand (n388,n389,n390);
or (n389,n166,n95);
nand (n390,n95,n166);
nand (n391,n374,n98);
nand (n392,n393,n69);
nand (n393,n394,n396);
or (n394,n95,n395);
and (n395,n226,n120);
or (n396,n120,n226);
nand (n397,n398,n436);
or (n398,n399,n422);
not (n399,n400);
nand (n400,n401,n421);
or (n401,n402,n411);
nor (n402,n403,n410);
nand (n403,n404,n409);
or (n404,n405,n92);
not (n405,n406);
nand (n406,n407,n408);
or (n407,n190,n95);
nand (n408,n95,n190);
nand (n409,n388,n98);
nor (n410,n124,n273);
nand (n411,n412,n419);
nand (n412,n413,n418);
or (n413,n414,n92);
not (n414,n415);
nand (n415,n416,n417);
or (n416,n94,n226);
or (n417,n95,n273);
nand (n418,n406,n98);
nor (n419,n420,n94);
and (n420,n226,n98);
nand (n421,n403,n410);
not (n422,n423);
nand (n423,n424,n432);
not (n424,n425);
nand (n425,n426,n431);
or (n426,n427,n115);
not (n427,n428);
nand (n428,n429,n430);
or (n429,n130,n226);
or (n430,n69,n273);
nand (n431,n125,n367);
nor (n432,n433,n435);
and (n433,n384,n434);
not (n434,n392);
and (n435,n385,n392);
nand (n436,n437,n425);
not (n437,n432);
xor (n438,n362,n371);
and (n439,n383,n397);
and (n440,n360,n379);
and (n441,n294,n334);
or (n442,n443,n465);
xor (n443,n444,n449);
xor (n444,n445,n446);
xor (n445,n268,n274);
or (n446,n447,n448);
and (n447,n344,n350);
and (n448,n345,n346);
xor (n449,n450,n462);
xor (n450,n451,n458);
nand (n451,n452,n457);
or (n452,n453,n25);
not (n453,n454);
nand (n454,n455,n456);
or (n455,n24,n226);
or (n456,n19,n273);
or (n457,n26,n235);
nand (n458,n459,n461);
or (n459,n460,n115);
not (n460,n354);
nand (n461,n125,n257);
nand (n462,n463,n464);
or (n463,n61,n339);
or (n464,n62,n263);
or (n465,n466,n467);
and (n466,n335,n343);
and (n467,n336,n342);
not (n468,n469);
nand (n469,n443,n465);
nand (n470,n471,n483);
not (n471,n472);
nor (n472,n473,n480);
xor (n473,n474,n479);
xor (n474,n475,n478);
or (n475,n476,n477);
and (n476,n450,n462);
and (n477,n451,n458);
xor (n478,n223,n233);
xor (n479,n253,n267);
or (n480,n481,n482);
and (n481,n444,n449);
and (n482,n445,n446);
not (n483,n484);
nor (n484,n485,n488);
or (n485,n486,n487);
and (n486,n474,n479);
and (n487,n475,n478);
xor (n488,n249,n283);
nor (n489,n490,n493);
and (n490,n483,n491);
not (n491,n492);
nand (n492,n473,n480);
and (n493,n485,n488);
nand (n494,n246,n247);
nand (n495,n496,n2);
nand (n496,n497,n912);
or (n497,n498,n659);
nand (n498,n499,n658);
nand (n499,n500,n611);
not (n500,n501);
xor (n501,n502,n572);
xor (n502,n503,n529);
xor (n503,n504,n525);
xor (n504,n505,n513);
nand (n505,n506,n507);
or (n506,n116,n125);
nand (n507,n508,n512);
or (n508,n69,n509);
not (n509,n510);
and (n510,n53,n511);
or (n512,n130,n510);
nand (n513,n514,n520);
or (n514,n61,n515);
nor (n515,n516,n518);
and (n516,n36,n517);
and (n518,n32,n519);
not (n519,n517);
or (n520,n62,n521);
nor (n521,n522,n523);
and (n522,n36,n511);
and (n523,n32,n524);
not (n524,n511);
nor (n525,n48,n526);
nor (n526,n527,n528);
and (n527,n50,n111);
and (n528,n49,n109);
xor (n529,n530,n552);
xor (n530,n531,n544);
nand (n531,n532,n538);
or (n532,n25,n533);
nor (n533,n534,n536);
and (n534,n24,n535);
and (n536,n19,n537);
not (n537,n535);
or (n538,n26,n539);
nor (n539,n540,n542);
and (n540,n24,n541);
and (n542,n19,n543);
not (n543,n541);
nand (n544,n545,n547);
or (n545,n546,n124);
not (n546,n507);
nand (n547,n548,n116);
not (n548,n549);
nor (n549,n550,n551);
and (n550,n130,n511);
and (n551,n69,n524);
or (n552,n553,n571);
and (n553,n554,n565);
xor (n554,n555,n559);
nor (n555,n48,n556);
nor (n556,n557,n558);
and (n557,n50,n105);
and (n558,n49,n103);
nand (n559,n560,n564);
or (n560,n61,n561);
nor (n561,n562,n563);
and (n562,n541,n36);
and (n563,n543,n32);
or (n564,n62,n515);
nand (n565,n566,n570);
or (n566,n25,n567);
nor (n567,n568,n569);
and (n568,n24,n109);
and (n569,n19,n111);
or (n570,n26,n533);
and (n571,n555,n559);
or (n572,n573,n610);
and (n573,n574,n590);
xor (n574,n575,n576);
not (n575,n544);
or (n576,n577,n583);
nand (n577,n578,n582);
or (n578,n25,n579);
nor (n579,n580,n581);
and (n580,n24,n103);
and (n581,n19,n105);
or (n582,n26,n567);
nand (n583,n584,n589);
or (n584,n115,n585);
not (n585,n586);
nand (n586,n587,n588);
or (n587,n69,n519);
or (n588,n130,n517);
or (n589,n124,n549);
or (n590,n591,n609);
and (n591,n592,n603);
xor (n592,n593,n597);
nor (n593,n48,n594);
nor (n594,n595,n596);
and (n595,n50,n139);
and (n596,n49,n137);
nand (n597,n598,n599);
or (n598,n98,n93);
not (n599,n600);
nor (n600,n601,n602);
and (n601,n94,n510);
and (n602,n95,n509);
nand (n603,n604,n605);
or (n604,n561,n62);
or (n605,n61,n606);
nor (n606,n607,n608);
and (n607,n36,n535);
and (n608,n32,n537);
and (n609,n593,n597);
and (n610,n575,n576);
not (n611,n612);
or (n612,n613,n657);
and (n613,n614,n617);
xor (n614,n615,n616);
xor (n615,n554,n565);
xor (n616,n574,n590);
or (n617,n618,n656);
and (n618,n619,n652);
xor (n619,n620,n631);
and (n620,n621,n627);
nand (n621,n622,n626);
or (n622,n92,n623);
nor (n623,n624,n625);
and (n624,n94,n511);
and (n625,n95,n524);
or (n626,n600,n112);
nand (n627,n628,n630);
or (n628,n629,n115);
xor (n629,n541,n130);
nand (n630,n125,n586);
or (n631,n632,n651);
and (n632,n633,n645);
xor (n633,n634,n641);
nand (n634,n635,n640);
or (n635,n636,n25);
not (n636,n637);
nor (n637,n638,n639);
and (n638,n137,n19);
and (n639,n139,n24);
or (n640,n26,n579);
nor (n641,n48,n642);
nor (n642,n643,n644);
and (n643,n50,n133);
and (n644,n49,n131);
nand (n645,n646,n650);
or (n646,n61,n647);
nor (n647,n648,n649);
and (n648,n36,n109);
and (n649,n32,n111);
or (n650,n62,n606);
and (n651,n634,n641);
nand (n652,n653,n576);
or (n653,n654,n655);
not (n654,n583);
not (n655,n577);
and (n656,n620,n631);
and (n657,n615,n616);
or (n658,n500,n611);
nand (n659,n660,n911);
or (n660,n661,n708);
nor (n661,n662,n663);
xor (n662,n614,n617);
or (n663,n664,n707);
and (n664,n665,n706);
xor (n665,n666,n667);
xor (n666,n592,n603);
or (n667,n668,n705);
and (n668,n669,n684);
xor (n669,n670,n671);
xor (n670,n621,n627);
and (n671,n672,n678);
nand (n672,n673,n677);
or (n673,n92,n674);
nor (n674,n675,n676);
and (n675,n94,n517);
and (n676,n95,n519);
or (n677,n623,n112);
nand (n678,n679,n683);
or (n679,n115,n680);
nor (n680,n681,n682);
and (n681,n130,n535);
and (n682,n69,n537);
or (n683,n629,n124);
or (n684,n685,n704);
and (n685,n686,n698);
xor (n686,n687,n694);
nand (n687,n688,n693);
or (n688,n689,n25);
not (n689,n690);
nor (n690,n691,n692);
and (n691,n131,n19);
and (n692,n133,n24);
nand (n693,n41,n637);
nor (n694,n48,n695);
nor (n695,n696,n697);
and (n696,n50,n86);
and (n697,n49,n84);
nand (n698,n699,n703);
or (n699,n61,n700);
nor (n700,n701,n702);
and (n701,n36,n103);
and (n702,n32,n105);
or (n703,n62,n647);
and (n704,n687,n694);
and (n705,n670,n671);
xor (n706,n619,n652);
and (n707,n666,n667);
not (n708,n709);
nand (n709,n710,n907);
or (n710,n711,n808);
not (n711,n712);
nor (n712,n713,n800);
nor (n713,n714,n793);
or (n714,n715,n792);
and (n715,n716,n754);
xor (n716,n717,n718);
xor (n717,n686,n698);
xor (n718,n719,n734);
xor (n719,n720,n721);
xor (n720,n672,n678);
and (n721,n722,n728);
nand (n722,n723,n727);
or (n723,n92,n724);
nor (n724,n725,n726);
and (n725,n94,n541);
and (n726,n95,n543);
or (n727,n674,n112);
nand (n728,n729,n733);
or (n729,n115,n730);
nor (n730,n731,n732);
and (n731,n130,n109);
and (n732,n69,n111);
or (n733,n124,n680);
or (n734,n735,n753);
and (n735,n736,n747);
xor (n736,n737,n743);
nand (n737,n738,n742);
or (n738,n739,n25);
nor (n739,n740,n741);
and (n740,n84,n24);
and (n741,n86,n19);
nand (n742,n41,n690);
nor (n743,n48,n744);
nor (n744,n745,n746);
and (n745,n50,n80);
and (n746,n49,n78);
nand (n747,n748,n752);
or (n748,n61,n749);
nor (n749,n750,n751);
and (n750,n36,n137);
and (n751,n32,n139);
or (n752,n62,n700);
and (n753,n737,n743);
or (n754,n755,n791);
and (n755,n756,n771);
xor (n756,n757,n758);
xor (n757,n722,n728);
and (n758,n759,n765);
nand (n759,n760,n764);
or (n760,n92,n761);
nor (n761,n762,n763);
and (n762,n94,n535);
and (n763,n95,n537);
or (n764,n724,n112);
nand (n765,n766,n770);
or (n766,n115,n767);
nor (n767,n768,n769);
and (n768,n130,n103);
and (n769,n69,n105);
or (n770,n730,n124);
or (n771,n772,n790);
and (n772,n773,n784);
xor (n773,n774,n780);
nand (n774,n775,n779);
or (n775,n25,n776);
nor (n776,n777,n778);
and (n777,n24,n78);
and (n778,n19,n80);
or (n779,n26,n739);
nor (n780,n48,n781);
nor (n781,n782,n783);
and (n782,n50,n46);
and (n783,n49,n44);
nand (n784,n785,n786);
or (n785,n749,n62);
or (n786,n61,n787);
nor (n787,n788,n789);
and (n788,n36,n131);
and (n789,n32,n133);
and (n790,n774,n780);
and (n791,n757,n758);
and (n792,n717,n718);
xor (n793,n794,n797);
xor (n794,n795,n796);
xor (n795,n633,n645);
xor (n796,n669,n684);
or (n797,n798,n799);
and (n798,n719,n734);
and (n799,n720,n721);
not (n800,n801);
nand (n801,n802,n804);
not (n802,n803);
xor (n803,n665,n706);
not (n804,n805);
or (n805,n806,n807);
and (n806,n794,n797);
and (n807,n795,n796);
not (n808,n809);
nand (n809,n810,n896,n906);
nand (n810,n811,n817);
nand (n811,n812,n815,n242);
nand (n812,n813,n7);
nand (n813,n814,n494);
or (n814,n489,n245);
nand (n815,n7,n288,n816);
not (n816,n245);
nor (n817,n818,n875);
nand (n818,n819,n868);
not (n819,n820);
nor (n820,n821,n859);
xor (n821,n822,n850);
xor (n822,n823,n824);
xor (n823,n773,n784);
xor (n824,n825,n834);
xor (n825,n826,n827);
xor (n826,n759,n765);
and (n827,n828,n831);
nand (n828,n829,n830);
or (n829,n92,n107);
or (n830,n761,n112);
nand (n831,n832,n833);
or (n832,n115,n135);
or (n833,n767,n124);
or (n834,n835,n849);
and (n835,n836,n846);
xor (n836,n837,n842);
nand (n837,n838,n840);
or (n838,n839,n25);
not (n839,n42);
nand (n840,n841,n41);
not (n841,n776);
nor (n842,n48,n843);
nor (n843,n844,n845);
and (n844,n50,n23);
and (n845,n49,n18);
nand (n846,n847,n848);
or (n847,n61,n82);
or (n848,n62,n787);
and (n849,n837,n842);
or (n850,n851,n858);
and (n851,n852,n855);
xor (n852,n853,n854);
xor (n853,n828,n831);
and (n854,n90,n113);
or (n855,n856,n857);
and (n856,n12,n59);
and (n857,n13,n47);
and (n858,n853,n854);
or (n859,n860,n867);
and (n860,n861,n864);
xor (n861,n862,n863);
xor (n862,n836,n846);
xor (n863,n852,n855);
or (n864,n865,n866);
and (n865,n88,n153);
and (n866,n89,n140);
and (n867,n862,n863);
nand (n868,n869,n871);
not (n869,n870);
xor (n870,n861,n864);
not (n871,n872);
or (n872,n873,n874);
and (n873,n10,n176);
and (n874,n11,n87);
nand (n875,n876,n889);
nand (n876,n877,n885);
not (n877,n878);
xor (n878,n879,n882);
xor (n879,n880,n881);
xor (n880,n736,n747);
xor (n881,n756,n771);
or (n882,n883,n884);
and (n883,n825,n834);
and (n884,n826,n827);
not (n885,n886);
or (n886,n887,n888);
and (n887,n822,n850);
and (n888,n823,n824);
nand (n889,n890,n892);
not (n890,n891);
xor (n891,n716,n754);
not (n892,n893);
or (n893,n894,n895);
and (n894,n879,n882);
and (n895,n880,n881);
nand (n896,n897,n889);
nand (n897,n898,n905);
or (n898,n899,n900);
not (n899,n876);
not (n900,n901);
nand (n901,n902,n904);
or (n902,n820,n903);
nand (n903,n870,n872);
nand (n904,n821,n859);
nand (n905,n878,n886);
nand (n906,n893,n891);
nor (n907,n908,n910);
and (n908,n909,n801);
and (n909,n714,n793);
nor (n910,n802,n804);
nand (n911,n662,n663);
nand (n912,n659,n498);
wire s0n913,s1n913,notn913;
or (n913,s0n913,s1n913);
not(notn913,n3);
and (s0n913,notn913,n914);
and (s1n913,n3,n1845);
xor (n914,n915,n1599);
xor (n915,n916,n1843);
xor (n916,n917,n1594);
xor (n917,n918,n1836);
xor (n918,n919,n1588);
xor (n919,n920,n1824);
xor (n920,n921,n1582);
xor (n921,n922,n1807);
xor (n922,n923,n1576);
xor (n923,n924,n1785);
xor (n924,n925,n1570);
xor (n925,n926,n1758);
xor (n926,n927,n1564);
xor (n927,n928,n1726);
xor (n928,n929,n1558);
xor (n929,n930,n1689);
xor (n930,n931,n1552);
xor (n931,n932,n1647);
xor (n932,n933,n1546);
xor (n933,n934,n1600);
xor (n934,n935,n1540);
xor (n935,n936,n1537);
xor (n936,n937,n1536);
xor (n937,n938,n1472);
xor (n938,n939,n1471);
xor (n939,n940,n1396);
xor (n940,n941,n1395);
xor (n941,n942,n1315);
xor (n942,n943,n1314);
xor (n943,n944,n1228);
xor (n944,n945,n1227);
xor (n945,n946,n957);
xor (n946,n947,n956);
xor (n947,n948,n955);
xor (n948,n949,n954);
xor (n949,n950,n953);
xor (n950,n951,n952);
and (n951,n510,n98);
and (n952,n510,n95);
and (n953,n951,n952);
and (n954,n510,n120);
and (n955,n949,n954);
and (n956,n510,n69);
or (n957,n958,n1142);
and (n958,n959,n1141);
xor (n959,n948,n960);
or (n960,n961,n1053);
and (n961,n962,n1052);
xor (n962,n950,n963);
or (n963,n953,n964);
and (n964,n965,n967);
xor (n965,n951,n966);
and (n966,n511,n95);
or (n967,n968,n971);
and (n968,n969,n970);
and (n969,n511,n98);
and (n970,n517,n95);
and (n971,n972,n973);
xor (n972,n969,n970);
or (n973,n974,n977);
and (n974,n975,n976);
and (n975,n517,n98);
and (n976,n541,n95);
and (n977,n978,n979);
xor (n978,n975,n976);
or (n979,n980,n983);
and (n980,n981,n982);
and (n981,n541,n98);
and (n982,n535,n95);
and (n983,n984,n985);
xor (n984,n981,n982);
or (n985,n986,n989);
and (n986,n987,n988);
and (n987,n535,n98);
and (n988,n109,n95);
and (n989,n990,n991);
xor (n990,n987,n988);
or (n991,n992,n995);
and (n992,n993,n994);
and (n993,n109,n98);
and (n994,n103,n95);
and (n995,n996,n997);
xor (n996,n993,n994);
or (n997,n998,n1001);
and (n998,n999,n1000);
and (n999,n103,n98);
and (n1000,n137,n95);
and (n1001,n1002,n1003);
xor (n1002,n999,n1000);
or (n1003,n1004,n1007);
and (n1004,n1005,n1006);
and (n1005,n137,n98);
and (n1006,n131,n95);
and (n1007,n1008,n1009);
xor (n1008,n1005,n1006);
or (n1009,n1010,n1013);
and (n1010,n1011,n1012);
and (n1011,n131,n98);
and (n1012,n84,n95);
and (n1013,n1014,n1015);
xor (n1014,n1011,n1012);
or (n1015,n1016,n1018);
and (n1016,n1017,n278);
and (n1017,n84,n98);
and (n1018,n1019,n1020);
xor (n1019,n1017,n278);
or (n1020,n1021,n1024);
and (n1021,n1022,n1023);
and (n1022,n78,n98);
and (n1023,n44,n95);
and (n1024,n1025,n1026);
xor (n1025,n1022,n1023);
or (n1026,n1027,n1030);
and (n1027,n1028,n1029);
and (n1028,n44,n98);
and (n1029,n18,n95);
and (n1030,n1031,n1032);
xor (n1031,n1028,n1029);
or (n1032,n1033,n1035);
and (n1033,n1034,n376);
and (n1034,n18,n98);
and (n1035,n1036,n1037);
xor (n1036,n1034,n376);
or (n1037,n1038,n1041);
and (n1038,n1039,n1040);
and (n1039,n57,n98);
and (n1040,n167,n95);
and (n1041,n1042,n1043);
xor (n1042,n1039,n1040);
or (n1043,n1044,n1047);
and (n1044,n1045,n1046);
and (n1045,n167,n98);
and (n1046,n191,n95);
and (n1047,n1048,n1049);
xor (n1048,n1045,n1046);
and (n1049,n1050,n1051);
and (n1050,n191,n98);
and (n1051,n226,n95);
and (n1052,n511,n120);
and (n1053,n1054,n1055);
xor (n1054,n962,n1052);
or (n1055,n1056,n1059);
and (n1056,n1057,n1058);
xor (n1057,n965,n967);
and (n1058,n517,n120);
and (n1059,n1060,n1061);
xor (n1060,n1057,n1058);
or (n1061,n1062,n1065);
and (n1062,n1063,n1064);
xor (n1063,n972,n973);
and (n1064,n541,n120);
and (n1065,n1066,n1067);
xor (n1066,n1063,n1064);
or (n1067,n1068,n1071);
and (n1068,n1069,n1070);
xor (n1069,n978,n979);
and (n1070,n535,n120);
and (n1071,n1072,n1073);
xor (n1072,n1069,n1070);
or (n1073,n1074,n1077);
and (n1074,n1075,n1076);
xor (n1075,n984,n985);
and (n1076,n109,n120);
and (n1077,n1078,n1079);
xor (n1078,n1075,n1076);
or (n1079,n1080,n1083);
and (n1080,n1081,n1082);
xor (n1081,n990,n991);
and (n1082,n103,n120);
and (n1083,n1084,n1085);
xor (n1084,n1081,n1082);
or (n1085,n1086,n1089);
and (n1086,n1087,n1088);
xor (n1087,n996,n997);
and (n1088,n137,n120);
and (n1089,n1090,n1091);
xor (n1090,n1087,n1088);
or (n1091,n1092,n1095);
and (n1092,n1093,n1094);
xor (n1093,n1002,n1003);
and (n1094,n131,n120);
and (n1095,n1096,n1097);
xor (n1096,n1093,n1094);
or (n1097,n1098,n1101);
and (n1098,n1099,n1100);
xor (n1099,n1008,n1009);
and (n1100,n84,n120);
and (n1101,n1102,n1103);
xor (n1102,n1099,n1100);
or (n1103,n1104,n1107);
and (n1104,n1105,n1106);
xor (n1105,n1014,n1015);
and (n1106,n78,n120);
and (n1107,n1108,n1109);
xor (n1108,n1105,n1106);
or (n1109,n1110,n1113);
and (n1110,n1111,n1112);
xor (n1111,n1019,n1020);
and (n1112,n44,n120);
and (n1113,n1114,n1115);
xor (n1114,n1111,n1112);
or (n1115,n1116,n1119);
and (n1116,n1117,n1118);
xor (n1117,n1025,n1026);
and (n1118,n18,n120);
and (n1119,n1120,n1121);
xor (n1120,n1117,n1118);
or (n1121,n1122,n1125);
and (n1122,n1123,n1124);
xor (n1123,n1031,n1032);
and (n1124,n57,n120);
and (n1125,n1126,n1127);
xor (n1126,n1123,n1124);
or (n1127,n1128,n1131);
and (n1128,n1129,n1130);
xor (n1129,n1036,n1037);
and (n1130,n167,n120);
and (n1131,n1132,n1133);
xor (n1132,n1129,n1130);
or (n1133,n1134,n1137);
and (n1134,n1135,n1136);
xor (n1135,n1042,n1043);
and (n1136,n191,n120);
and (n1137,n1138,n1139);
xor (n1138,n1135,n1136);
and (n1139,n1140,n395);
xor (n1140,n1048,n1049);
and (n1141,n511,n69);
and (n1142,n1143,n1144);
xor (n1143,n959,n1141);
or (n1144,n1145,n1148);
and (n1145,n1146,n1147);
xor (n1146,n1054,n1055);
and (n1147,n517,n69);
and (n1148,n1149,n1150);
xor (n1149,n1146,n1147);
or (n1150,n1151,n1154);
and (n1151,n1152,n1153);
xor (n1152,n1060,n1061);
and (n1153,n541,n69);
and (n1154,n1155,n1156);
xor (n1155,n1152,n1153);
or (n1156,n1157,n1160);
and (n1157,n1158,n1159);
xor (n1158,n1066,n1067);
and (n1159,n535,n69);
and (n1160,n1161,n1162);
xor (n1161,n1158,n1159);
or (n1162,n1163,n1166);
and (n1163,n1164,n1165);
xor (n1164,n1072,n1073);
and (n1165,n109,n69);
and (n1166,n1167,n1168);
xor (n1167,n1164,n1165);
or (n1168,n1169,n1172);
and (n1169,n1170,n1171);
xor (n1170,n1078,n1079);
and (n1171,n103,n69);
and (n1172,n1173,n1174);
xor (n1173,n1170,n1171);
or (n1174,n1175,n1178);
and (n1175,n1176,n1177);
xor (n1176,n1084,n1085);
and (n1177,n137,n69);
and (n1178,n1179,n1180);
xor (n1179,n1176,n1177);
or (n1180,n1181,n1184);
and (n1181,n1182,n1183);
xor (n1182,n1090,n1091);
and (n1183,n131,n69);
and (n1184,n1185,n1186);
xor (n1185,n1182,n1183);
or (n1186,n1187,n1190);
and (n1187,n1188,n1189);
xor (n1188,n1096,n1097);
and (n1189,n84,n69);
and (n1190,n1191,n1192);
xor (n1191,n1188,n1189);
or (n1192,n1193,n1196);
and (n1193,n1194,n1195);
xor (n1194,n1102,n1103);
and (n1195,n78,n69);
and (n1196,n1197,n1198);
xor (n1197,n1194,n1195);
or (n1198,n1199,n1201);
and (n1199,n1200,n258);
xor (n1200,n1108,n1109);
and (n1201,n1202,n1203);
xor (n1202,n1200,n258);
or (n1203,n1204,n1207);
and (n1204,n1205,n1206);
xor (n1205,n1114,n1115);
and (n1206,n18,n69);
and (n1207,n1208,n1209);
xor (n1208,n1205,n1206);
or (n1209,n1210,n1212);
and (n1210,n1211,n305);
xor (n1211,n1120,n1121);
and (n1212,n1213,n1214);
xor (n1213,n1211,n305);
or (n1214,n1215,n1217);
and (n1215,n1216,n302);
xor (n1216,n1126,n1127);
and (n1217,n1218,n1219);
xor (n1218,n1216,n302);
or (n1219,n1220,n1222);
and (n1220,n1221,n368);
xor (n1221,n1132,n1133);
and (n1222,n1223,n1224);
xor (n1223,n1221,n368);
and (n1224,n1225,n1226);
xor (n1225,n1138,n1139);
and (n1226,n226,n69);
and (n1227,n511,n66);
or (n1228,n1229,n1232);
and (n1229,n1230,n1231);
xor (n1230,n1143,n1144);
and (n1231,n517,n66);
and (n1232,n1233,n1234);
xor (n1233,n1230,n1231);
or (n1234,n1235,n1238);
and (n1235,n1236,n1237);
xor (n1236,n1149,n1150);
and (n1237,n541,n66);
and (n1238,n1239,n1240);
xor (n1239,n1236,n1237);
or (n1240,n1241,n1244);
and (n1241,n1242,n1243);
xor (n1242,n1155,n1156);
and (n1243,n535,n66);
and (n1244,n1245,n1246);
xor (n1245,n1242,n1243);
or (n1246,n1247,n1250);
and (n1247,n1248,n1249);
xor (n1248,n1161,n1162);
and (n1249,n109,n66);
and (n1250,n1251,n1252);
xor (n1251,n1248,n1249);
or (n1252,n1253,n1256);
and (n1253,n1254,n1255);
xor (n1254,n1167,n1168);
and (n1255,n103,n66);
and (n1256,n1257,n1258);
xor (n1257,n1254,n1255);
or (n1258,n1259,n1262);
and (n1259,n1260,n1261);
xor (n1260,n1173,n1174);
and (n1261,n137,n66);
and (n1262,n1263,n1264);
xor (n1263,n1260,n1261);
or (n1264,n1265,n1268);
and (n1265,n1266,n1267);
xor (n1266,n1179,n1180);
and (n1267,n131,n66);
and (n1268,n1269,n1270);
xor (n1269,n1266,n1267);
or (n1270,n1271,n1274);
and (n1271,n1272,n1273);
xor (n1272,n1185,n1186);
and (n1273,n84,n66);
and (n1274,n1275,n1276);
xor (n1275,n1272,n1273);
or (n1276,n1277,n1280);
and (n1277,n1278,n1279);
xor (n1278,n1191,n1192);
and (n1279,n78,n66);
and (n1280,n1281,n1282);
xor (n1281,n1278,n1279);
or (n1282,n1283,n1286);
and (n1283,n1284,n1285);
xor (n1284,n1197,n1198);
and (n1285,n44,n66);
and (n1286,n1287,n1288);
xor (n1287,n1284,n1285);
or (n1288,n1289,n1292);
and (n1289,n1290,n1291);
xor (n1290,n1202,n1203);
and (n1291,n18,n66);
and (n1292,n1293,n1294);
xor (n1293,n1290,n1291);
or (n1294,n1295,n1298);
and (n1295,n1296,n1297);
xor (n1296,n1208,n1209);
and (n1297,n57,n66);
and (n1298,n1299,n1300);
xor (n1299,n1296,n1297);
or (n1300,n1301,n1304);
and (n1301,n1302,n1303);
xor (n1302,n1213,n1214);
and (n1303,n167,n66);
and (n1304,n1305,n1306);
xor (n1305,n1302,n1303);
or (n1306,n1307,n1310);
and (n1307,n1308,n1309);
xor (n1308,n1218,n1219);
and (n1309,n191,n66);
and (n1310,n1311,n1312);
xor (n1311,n1308,n1309);
and (n1312,n1313,n322);
xor (n1313,n1223,n1224);
and (n1314,n517,n32);
or (n1315,n1316,n1319);
and (n1316,n1317,n1318);
xor (n1317,n1233,n1234);
and (n1318,n541,n32);
and (n1319,n1320,n1321);
xor (n1320,n1317,n1318);
or (n1321,n1322,n1325);
and (n1322,n1323,n1324);
xor (n1323,n1239,n1240);
and (n1324,n535,n32);
and (n1325,n1326,n1327);
xor (n1326,n1323,n1324);
or (n1327,n1328,n1331);
and (n1328,n1329,n1330);
xor (n1329,n1245,n1246);
and (n1330,n109,n32);
and (n1331,n1332,n1333);
xor (n1332,n1329,n1330);
or (n1333,n1334,n1337);
and (n1334,n1335,n1336);
xor (n1335,n1251,n1252);
and (n1336,n103,n32);
and (n1337,n1338,n1339);
xor (n1338,n1335,n1336);
or (n1339,n1340,n1343);
and (n1340,n1341,n1342);
xor (n1341,n1257,n1258);
and (n1342,n137,n32);
and (n1343,n1344,n1345);
xor (n1344,n1341,n1342);
or (n1345,n1346,n1349);
and (n1346,n1347,n1348);
xor (n1347,n1263,n1264);
and (n1348,n131,n32);
and (n1349,n1350,n1351);
xor (n1350,n1347,n1348);
or (n1351,n1352,n1355);
and (n1352,n1353,n1354);
xor (n1353,n1269,n1270);
and (n1354,n84,n32);
and (n1355,n1356,n1357);
xor (n1356,n1353,n1354);
or (n1357,n1358,n1361);
and (n1358,n1359,n1360);
xor (n1359,n1275,n1276);
and (n1360,n78,n32);
and (n1361,n1362,n1363);
xor (n1362,n1359,n1360);
or (n1363,n1364,n1367);
and (n1364,n1365,n1366);
xor (n1365,n1281,n1282);
and (n1366,n44,n32);
and (n1367,n1368,n1369);
xor (n1368,n1365,n1366);
or (n1369,n1370,n1373);
and (n1370,n1371,n1372);
xor (n1371,n1287,n1288);
and (n1372,n18,n32);
and (n1373,n1374,n1375);
xor (n1374,n1371,n1372);
or (n1375,n1376,n1379);
and (n1376,n1377,n1378);
xor (n1377,n1293,n1294);
and (n1378,n57,n32);
and (n1379,n1380,n1381);
xor (n1380,n1377,n1378);
or (n1381,n1382,n1385);
and (n1382,n1383,n1384);
xor (n1383,n1299,n1300);
and (n1384,n167,n32);
and (n1385,n1386,n1387);
xor (n1386,n1383,n1384);
or (n1387,n1388,n1390);
and (n1388,n1389,n311);
xor (n1389,n1305,n1306);
and (n1390,n1391,n1392);
xor (n1391,n1389,n311);
and (n1392,n1393,n1394);
xor (n1393,n1311,n1312);
and (n1394,n226,n32);
and (n1395,n541,n29);
or (n1396,n1397,n1400);
and (n1397,n1398,n1399);
xor (n1398,n1320,n1321);
and (n1399,n535,n29);
and (n1400,n1401,n1402);
xor (n1401,n1398,n1399);
or (n1402,n1403,n1406);
and (n1403,n1404,n1405);
xor (n1404,n1326,n1327);
and (n1405,n109,n29);
and (n1406,n1407,n1408);
xor (n1407,n1404,n1405);
or (n1408,n1409,n1412);
and (n1409,n1410,n1411);
xor (n1410,n1332,n1333);
and (n1411,n103,n29);
and (n1412,n1413,n1414);
xor (n1413,n1410,n1411);
or (n1414,n1415,n1418);
and (n1415,n1416,n1417);
xor (n1416,n1338,n1339);
and (n1417,n137,n29);
and (n1418,n1419,n1420);
xor (n1419,n1416,n1417);
or (n1420,n1421,n1424);
and (n1421,n1422,n1423);
xor (n1422,n1344,n1345);
and (n1423,n131,n29);
and (n1424,n1425,n1426);
xor (n1425,n1422,n1423);
or (n1426,n1427,n1430);
and (n1427,n1428,n1429);
xor (n1428,n1350,n1351);
and (n1429,n84,n29);
and (n1430,n1431,n1432);
xor (n1431,n1428,n1429);
or (n1432,n1433,n1436);
and (n1433,n1434,n1435);
xor (n1434,n1356,n1357);
and (n1435,n78,n29);
and (n1436,n1437,n1438);
xor (n1437,n1434,n1435);
or (n1438,n1439,n1442);
and (n1439,n1440,n1441);
xor (n1440,n1362,n1363);
and (n1441,n44,n29);
and (n1442,n1443,n1444);
xor (n1443,n1440,n1441);
or (n1444,n1445,n1448);
and (n1445,n1446,n1447);
xor (n1446,n1368,n1369);
and (n1447,n18,n29);
and (n1448,n1449,n1450);
xor (n1449,n1446,n1447);
or (n1450,n1451,n1454);
and (n1451,n1452,n1453);
xor (n1452,n1374,n1375);
and (n1453,n57,n29);
and (n1454,n1455,n1456);
xor (n1455,n1452,n1453);
or (n1456,n1457,n1460);
and (n1457,n1458,n1459);
xor (n1458,n1380,n1381);
and (n1459,n167,n29);
and (n1460,n1461,n1462);
xor (n1461,n1458,n1459);
or (n1462,n1463,n1466);
and (n1463,n1464,n1465);
xor (n1464,n1386,n1387);
and (n1465,n191,n29);
and (n1466,n1467,n1468);
xor (n1467,n1464,n1465);
and (n1468,n1469,n1470);
xor (n1469,n1391,n1392);
not (n1470,n271);
and (n1471,n535,n19);
or (n1472,n1473,n1476);
and (n1473,n1474,n1475);
xor (n1474,n1401,n1402);
and (n1475,n109,n19);
and (n1476,n1477,n1478);
xor (n1477,n1474,n1475);
or (n1478,n1479,n1482);
and (n1479,n1480,n1481);
xor (n1480,n1407,n1408);
and (n1481,n103,n19);
and (n1482,n1483,n1484);
xor (n1483,n1480,n1481);
or (n1484,n1485,n1487);
and (n1485,n1486,n638);
xor (n1486,n1413,n1414);
and (n1487,n1488,n1489);
xor (n1488,n1486,n638);
or (n1489,n1490,n1492);
and (n1490,n1491,n691);
xor (n1491,n1419,n1420);
and (n1492,n1493,n1494);
xor (n1493,n1491,n691);
or (n1494,n1495,n1498);
and (n1495,n1496,n1497);
xor (n1496,n1425,n1426);
and (n1497,n84,n19);
and (n1498,n1499,n1500);
xor (n1499,n1496,n1497);
or (n1500,n1501,n1504);
and (n1501,n1502,n1503);
xor (n1502,n1431,n1432);
and (n1503,n78,n19);
and (n1504,n1505,n1506);
xor (n1505,n1502,n1503);
or (n1506,n1507,n1509);
and (n1507,n1508,n43);
xor (n1508,n1437,n1438);
and (n1509,n1510,n1511);
xor (n1510,n1508,n43);
or (n1511,n1512,n1514);
and (n1512,n1513,n17);
xor (n1513,n1443,n1444);
and (n1514,n1515,n1516);
xor (n1515,n1513,n17);
or (n1516,n1517,n1519);
and (n1517,n1518,n160);
xor (n1518,n1449,n1450);
and (n1519,n1520,n1521);
xor (n1520,n1518,n160);
or (n1521,n1522,n1525);
and (n1522,n1523,n1524);
xor (n1523,n1455,n1456);
and (n1524,n167,n19);
and (n1525,n1526,n1527);
xor (n1526,n1523,n1524);
or (n1527,n1528,n1531);
and (n1528,n1529,n1530);
xor (n1529,n1461,n1462);
and (n1530,n191,n19);
and (n1531,n1532,n1533);
xor (n1532,n1529,n1530);
and (n1533,n1534,n1535);
xor (n1534,n1467,n1468);
and (n1535,n226,n19);
and (n1536,n109,n50);
or (n1537,n1538,n1541);
and (n1538,n1539,n1540);
xor (n1539,n1477,n1478);
and (n1540,n103,n50);
and (n1541,n1542,n1543);
xor (n1542,n1539,n1540);
or (n1543,n1544,n1547);
and (n1544,n1545,n1546);
xor (n1545,n1483,n1484);
and (n1546,n137,n50);
and (n1547,n1548,n1549);
xor (n1548,n1545,n1546);
or (n1549,n1550,n1553);
and (n1550,n1551,n1552);
xor (n1551,n1488,n1489);
and (n1552,n131,n50);
and (n1553,n1554,n1555);
xor (n1554,n1551,n1552);
or (n1555,n1556,n1559);
and (n1556,n1557,n1558);
xor (n1557,n1493,n1494);
and (n1558,n84,n50);
and (n1559,n1560,n1561);
xor (n1560,n1557,n1558);
or (n1561,n1562,n1565);
and (n1562,n1563,n1564);
xor (n1563,n1499,n1500);
and (n1564,n78,n50);
and (n1565,n1566,n1567);
xor (n1566,n1563,n1564);
or (n1567,n1568,n1571);
and (n1568,n1569,n1570);
xor (n1569,n1505,n1506);
and (n1570,n44,n50);
and (n1571,n1572,n1573);
xor (n1572,n1569,n1570);
or (n1573,n1574,n1577);
and (n1574,n1575,n1576);
xor (n1575,n1510,n1511);
and (n1576,n18,n50);
and (n1577,n1578,n1579);
xor (n1578,n1575,n1576);
or (n1579,n1580,n1583);
and (n1580,n1581,n1582);
xor (n1581,n1515,n1516);
and (n1582,n57,n50);
and (n1583,n1584,n1585);
xor (n1584,n1581,n1582);
or (n1585,n1586,n1589);
and (n1586,n1587,n1588);
xor (n1587,n1520,n1521);
and (n1588,n167,n50);
and (n1589,n1590,n1591);
xor (n1590,n1587,n1588);
or (n1591,n1592,n1595);
and (n1592,n1593,n1594);
xor (n1593,n1526,n1527);
and (n1594,n191,n50);
and (n1595,n1596,n1597);
xor (n1596,n1593,n1594);
and (n1597,n1598,n1599);
xor (n1598,n1532,n1533);
and (n1599,n226,n50);
or (n1600,n1601,n1603);
and (n1601,n1602,n1546);
xor (n1602,n1542,n1543);
and (n1603,n1604,n1605);
xor (n1604,n1602,n1546);
or (n1605,n1606,n1608);
and (n1606,n1607,n1552);
xor (n1607,n1548,n1549);
and (n1608,n1609,n1610);
xor (n1609,n1607,n1552);
or (n1610,n1611,n1613);
and (n1611,n1612,n1558);
xor (n1612,n1554,n1555);
and (n1613,n1614,n1615);
xor (n1614,n1612,n1558);
or (n1615,n1616,n1618);
and (n1616,n1617,n1564);
xor (n1617,n1560,n1561);
and (n1618,n1619,n1620);
xor (n1619,n1617,n1564);
or (n1620,n1621,n1623);
and (n1621,n1622,n1570);
xor (n1622,n1566,n1567);
and (n1623,n1624,n1625);
xor (n1624,n1622,n1570);
or (n1625,n1626,n1628);
and (n1626,n1627,n1576);
xor (n1627,n1572,n1573);
and (n1628,n1629,n1630);
xor (n1629,n1627,n1576);
or (n1630,n1631,n1633);
and (n1631,n1632,n1582);
xor (n1632,n1578,n1579);
and (n1633,n1634,n1635);
xor (n1634,n1632,n1582);
or (n1635,n1636,n1638);
and (n1636,n1637,n1588);
xor (n1637,n1584,n1585);
and (n1638,n1639,n1640);
xor (n1639,n1637,n1588);
or (n1640,n1641,n1643);
and (n1641,n1642,n1594);
xor (n1642,n1590,n1591);
and (n1643,n1644,n1645);
xor (n1644,n1642,n1594);
and (n1645,n1646,n1599);
xor (n1646,n1596,n1597);
or (n1647,n1648,n1650);
and (n1648,n1649,n1552);
xor (n1649,n1604,n1605);
and (n1650,n1651,n1652);
xor (n1651,n1649,n1552);
or (n1652,n1653,n1655);
and (n1653,n1654,n1558);
xor (n1654,n1609,n1610);
and (n1655,n1656,n1657);
xor (n1656,n1654,n1558);
or (n1657,n1658,n1660);
and (n1658,n1659,n1564);
xor (n1659,n1614,n1615);
and (n1660,n1661,n1662);
xor (n1661,n1659,n1564);
or (n1662,n1663,n1665);
and (n1663,n1664,n1570);
xor (n1664,n1619,n1620);
and (n1665,n1666,n1667);
xor (n1666,n1664,n1570);
or (n1667,n1668,n1670);
and (n1668,n1669,n1576);
xor (n1669,n1624,n1625);
and (n1670,n1671,n1672);
xor (n1671,n1669,n1576);
or (n1672,n1673,n1675);
and (n1673,n1674,n1582);
xor (n1674,n1629,n1630);
and (n1675,n1676,n1677);
xor (n1676,n1674,n1582);
or (n1677,n1678,n1680);
and (n1678,n1679,n1588);
xor (n1679,n1634,n1635);
and (n1680,n1681,n1682);
xor (n1681,n1679,n1588);
or (n1682,n1683,n1685);
and (n1683,n1684,n1594);
xor (n1684,n1639,n1640);
and (n1685,n1686,n1687);
xor (n1686,n1684,n1594);
and (n1687,n1688,n1599);
xor (n1688,n1644,n1645);
or (n1689,n1690,n1692);
and (n1690,n1691,n1558);
xor (n1691,n1651,n1652);
and (n1692,n1693,n1694);
xor (n1693,n1691,n1558);
or (n1694,n1695,n1697);
and (n1695,n1696,n1564);
xor (n1696,n1656,n1657);
and (n1697,n1698,n1699);
xor (n1698,n1696,n1564);
or (n1699,n1700,n1702);
and (n1700,n1701,n1570);
xor (n1701,n1661,n1662);
and (n1702,n1703,n1704);
xor (n1703,n1701,n1570);
or (n1704,n1705,n1707);
and (n1705,n1706,n1576);
xor (n1706,n1666,n1667);
and (n1707,n1708,n1709);
xor (n1708,n1706,n1576);
or (n1709,n1710,n1712);
and (n1710,n1711,n1582);
xor (n1711,n1671,n1672);
and (n1712,n1713,n1714);
xor (n1713,n1711,n1582);
or (n1714,n1715,n1717);
and (n1715,n1716,n1588);
xor (n1716,n1676,n1677);
and (n1717,n1718,n1719);
xor (n1718,n1716,n1588);
or (n1719,n1720,n1722);
and (n1720,n1721,n1594);
xor (n1721,n1681,n1682);
and (n1722,n1723,n1724);
xor (n1723,n1721,n1594);
and (n1724,n1725,n1599);
xor (n1725,n1686,n1687);
or (n1726,n1727,n1729);
and (n1727,n1728,n1564);
xor (n1728,n1693,n1694);
and (n1729,n1730,n1731);
xor (n1730,n1728,n1564);
or (n1731,n1732,n1734);
and (n1732,n1733,n1570);
xor (n1733,n1698,n1699);
and (n1734,n1735,n1736);
xor (n1735,n1733,n1570);
or (n1736,n1737,n1739);
and (n1737,n1738,n1576);
xor (n1738,n1703,n1704);
and (n1739,n1740,n1741);
xor (n1740,n1738,n1576);
or (n1741,n1742,n1744);
and (n1742,n1743,n1582);
xor (n1743,n1708,n1709);
and (n1744,n1745,n1746);
xor (n1745,n1743,n1582);
or (n1746,n1747,n1749);
and (n1747,n1748,n1588);
xor (n1748,n1713,n1714);
and (n1749,n1750,n1751);
xor (n1750,n1748,n1588);
or (n1751,n1752,n1754);
and (n1752,n1753,n1594);
xor (n1753,n1718,n1719);
and (n1754,n1755,n1756);
xor (n1755,n1753,n1594);
and (n1756,n1757,n1599);
xor (n1757,n1723,n1724);
or (n1758,n1759,n1761);
and (n1759,n1760,n1570);
xor (n1760,n1730,n1731);
and (n1761,n1762,n1763);
xor (n1762,n1760,n1570);
or (n1763,n1764,n1766);
and (n1764,n1765,n1576);
xor (n1765,n1735,n1736);
and (n1766,n1767,n1768);
xor (n1767,n1765,n1576);
or (n1768,n1769,n1771);
and (n1769,n1770,n1582);
xor (n1770,n1740,n1741);
and (n1771,n1772,n1773);
xor (n1772,n1770,n1582);
or (n1773,n1774,n1776);
and (n1774,n1775,n1588);
xor (n1775,n1745,n1746);
and (n1776,n1777,n1778);
xor (n1777,n1775,n1588);
or (n1778,n1779,n1781);
and (n1779,n1780,n1594);
xor (n1780,n1750,n1751);
and (n1781,n1782,n1783);
xor (n1782,n1780,n1594);
and (n1783,n1784,n1599);
xor (n1784,n1755,n1756);
or (n1785,n1786,n1788);
and (n1786,n1787,n1576);
xor (n1787,n1762,n1763);
and (n1788,n1789,n1790);
xor (n1789,n1787,n1576);
or (n1790,n1791,n1793);
and (n1791,n1792,n1582);
xor (n1792,n1767,n1768);
and (n1793,n1794,n1795);
xor (n1794,n1792,n1582);
or (n1795,n1796,n1798);
and (n1796,n1797,n1588);
xor (n1797,n1772,n1773);
and (n1798,n1799,n1800);
xor (n1799,n1797,n1588);
or (n1800,n1801,n1803);
and (n1801,n1802,n1594);
xor (n1802,n1777,n1778);
and (n1803,n1804,n1805);
xor (n1804,n1802,n1594);
and (n1805,n1806,n1599);
xor (n1806,n1782,n1783);
or (n1807,n1808,n1810);
and (n1808,n1809,n1582);
xor (n1809,n1789,n1790);
and (n1810,n1811,n1812);
xor (n1811,n1809,n1582);
or (n1812,n1813,n1815);
and (n1813,n1814,n1588);
xor (n1814,n1794,n1795);
and (n1815,n1816,n1817);
xor (n1816,n1814,n1588);
or (n1817,n1818,n1820);
and (n1818,n1819,n1594);
xor (n1819,n1799,n1800);
and (n1820,n1821,n1822);
xor (n1821,n1819,n1594);
and (n1822,n1823,n1599);
xor (n1823,n1804,n1805);
or (n1824,n1825,n1827);
and (n1825,n1826,n1588);
xor (n1826,n1811,n1812);
and (n1827,n1828,n1829);
xor (n1828,n1826,n1588);
or (n1829,n1830,n1832);
and (n1830,n1831,n1594);
xor (n1831,n1816,n1817);
and (n1832,n1833,n1834);
xor (n1833,n1831,n1594);
and (n1834,n1835,n1599);
xor (n1835,n1821,n1822);
or (n1836,n1837,n1839);
and (n1837,n1838,n1594);
xor (n1838,n1828,n1829);
and (n1839,n1840,n1841);
xor (n1840,n1838,n1594);
and (n1841,n1842,n1599);
xor (n1842,n1833,n1834);
and (n1843,n1844,n1599);
xor (n1844,n1840,n1841);
xor (n1845,n1725,n1599);
endmodule
