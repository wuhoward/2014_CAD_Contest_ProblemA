module top (out,n12,n15,n17,n18,n21,n22,n36,n46,n52
        ,n61,n96,n100,n148,n178,n231,n340,n343,n346,n360
        ,n369,n418,n493,n545);
output out;
input n12;
input n15;
input n17;
input n18;
input n21;
input n22;
input n36;
input n46;
input n52;
input n61;
input n96;
input n100;
input n148;
input n178;
input n231;
input n340;
input n343;
input n346;
input n360;
input n369;
input n418;
input n493;
input n545;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n13;
wire n14;
wire n16;
wire n19;
wire n20;
wire n23;
wire n24;
wire n25;
wire n26;
wire n27;
wire n28;
wire n29;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n97;
wire n98;
wire n99;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n341;
wire n342;
wire n344;
wire n345;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
xor (out,n0,n717);
xor (n0,n1,n644);
xor (n1,n2,n330);
xor (n2,n3,n80);
xor (n3,n4,n38);
xor (n4,n5,n33);
xor (n5,n6,n30);
or (n6,n7,n27,n29);
and (n7,n8,n24);
or (n8,n9,n19,n23);
and (n9,n10,n16);
nor (n10,n11,n13);
not (n11,n12);
and (n13,n14,n12);
not (n14,n15);
and (n16,n17,n18);
and (n19,n16,n20);
and (n20,n21,n22);
and (n23,n10,n20);
nor (n24,n25,n26);
not (n25,n17);
and (n26,n14,n17);
and (n27,n24,n28);
and (n28,n21,n18);
and (n29,n8,n28);
nor (n30,n31,n32);
not (n31,n21);
and (n32,n14,n21);
nor (n33,n34,n37);
and (n34,n35,n18);
not (n35,n36);
not (n37,n18);
or (n38,n39,n76,n79);
and (n39,n40,n73);
or (n40,n41,n69,n72);
and (n41,n42,n55);
or (n42,n43,n49,n54);
and (n43,n44,n48);
nor (n44,n45,n47);
not (n45,n46);
and (n47,n14,n46);
and (n48,n12,n18);
and (n49,n48,n50);
nor (n50,n51,n53);
and (n51,n35,n52);
not (n53,n52);
and (n54,n44,n50);
or (n55,n56,n66,n68);
and (n56,n57,n65);
or (n57,n58,n62,n64);
and (n58,n59,n60);
and (n59,n12,n22);
and (n60,n17,n61);
and (n62,n60,n63);
and (n63,n21,n52);
and (n64,n59,n63);
and (n65,n17,n22);
and (n66,n65,n67);
and (n67,n21,n61);
and (n68,n57,n67);
and (n69,n55,n70);
xor (n70,n71,n20);
xor (n71,n10,n16);
and (n72,n42,n70);
nor (n73,n74,n75);
and (n74,n35,n22);
not (n75,n22);
and (n76,n73,n77);
xor (n77,n78,n28);
xor (n78,n8,n24);
and (n79,n40,n77);
or (n80,n81,n119);
and (n81,n82,n84);
xor (n82,n83,n77);
xor (n83,n40,n73);
or (n84,n85,n115,n118);
and (n85,n86,n112);
or (n86,n87,n108,n111);
and (n87,n88,n106);
or (n88,n89,n102,n105);
and (n89,n90,n98);
or (n90,n91,n94,n97);
and (n91,n92,n93);
and (n92,n12,n61);
and (n93,n17,n52);
and (n94,n93,n95);
and (n95,n21,n96);
and (n97,n92,n95);
and (n98,n99,n101);
and (n99,n100,n18);
and (n101,n46,n22);
and (n102,n98,n103);
xor (n103,n104,n63);
xor (n104,n59,n60);
and (n105,n90,n103);
xor (n106,n107,n50);
xor (n107,n44,n48);
and (n108,n106,n109);
xor (n109,n110,n67);
xor (n110,n57,n65);
and (n111,n88,n109);
nor (n112,n113,n114);
and (n113,n35,n61);
not (n114,n61);
and (n115,n112,n116);
xor (n116,n117,n70);
xor (n117,n42,n55);
and (n118,n86,n116);
and (n119,n120,n121);
xor (n120,n82,n84);
or (n121,n122,n165);
and (n122,n123,n125);
xor (n123,n124,n116);
xor (n124,n86,n112);
or (n125,n126,n161,n164);
and (n126,n127,n138);
or (n127,n128,n133,n137);
and (n128,n129,n132);
nor (n129,n130,n131);
not (n130,n100);
and (n131,n14,n100);
and (n132,n46,n18);
and (n133,n132,n134);
nor (n134,n135,n136);
and (n135,n35,n96);
not (n136,n96);
and (n137,n129,n134);
or (n138,n139,n157,n160);
and (n139,n140,n155);
or (n140,n141,n152,n154);
and (n141,n142,n150);
or (n142,n143,n146,n149);
and (n143,n144,n145);
and (n144,n12,n52);
and (n145,n17,n96);
and (n146,n145,n147);
and (n147,n21,n148);
and (n149,n144,n147);
xor (n150,n151,n95);
xor (n151,n92,n93);
and (n152,n150,n153);
xor (n153,n99,n101);
and (n154,n142,n153);
xor (n155,n156,n134);
xor (n156,n129,n132);
and (n157,n155,n158);
xor (n158,n159,n103);
xor (n159,n90,n98);
and (n160,n140,n158);
and (n161,n138,n162);
xor (n162,n163,n109);
xor (n163,n88,n106);
and (n164,n127,n162);
and (n165,n166,n167);
xor (n166,n123,n125);
or (n167,n168,n214);
and (n168,n169,n171);
xor (n169,n170,n162);
xor (n170,n127,n138);
or (n171,n172,n210,n213);
and (n172,n173,n191);
or (n173,n174,n186,n190);
and (n174,n175,n183);
or (n175,n176,n180,n182);
and (n176,n177,n179);
and (n177,n178,n18);
and (n179,n100,n22);
and (n180,n179,n181);
and (n181,n46,n61);
and (n182,n177,n181);
nor (n183,n184,n185);
not (n184,n178);
and (n185,n14,n178);
and (n186,n183,n187);
nor (n187,n188,n189);
and (n188,n35,n148);
not (n189,n148);
and (n190,n175,n187);
or (n191,n192,n206,n209);
and (n192,n193,n204);
or (n193,n194,n200,n203);
and (n194,n195,n198);
and (n195,n196,n197);
and (n196,n12,n96);
and (n197,n17,n148);
xor (n198,n199,n181);
xor (n199,n177,n179);
and (n200,n198,n201);
xor (n201,n202,n147);
xor (n202,n144,n145);
and (n203,n195,n201);
xor (n204,n205,n187);
xor (n205,n175,n183);
and (n206,n204,n207);
xor (n207,n208,n153);
xor (n208,n142,n150);
and (n209,n193,n207);
and (n210,n191,n211);
xor (n211,n212,n158);
xor (n212,n140,n155);
and (n213,n173,n211);
and (n214,n215,n216);
xor (n215,n169,n171);
or (n216,n217,n236);
and (n217,n218,n220);
xor (n218,n219,n211);
xor (n219,n173,n191);
and (n220,n221,n234);
or (n221,n222,n228,n233);
and (n222,n223,n226);
and (n223,n224,n225);
and (n224,n46,n52);
xor (n225,n196,n197);
xor (n226,n227,n201);
xor (n227,n195,n198);
and (n228,n226,n229);
nor (n229,n230,n232);
not (n230,n231);
and (n232,n14,n231);
and (n233,n223,n229);
xor (n234,n235,n207);
xor (n235,n193,n204);
and (n236,n237,n238);
xor (n237,n218,n220);
or (n238,n239,n269);
and (n239,n240,n241);
xor (n240,n221,n234);
or (n241,n242,n265,n268);
and (n242,n243,n250);
or (n243,n244,n247,n249);
and (n244,n245,n246);
and (n245,n231,n18);
and (n246,n178,n22);
and (n247,n246,n248);
and (n248,n100,n61);
and (n249,n245,n248);
or (n250,n251,n262,n264);
and (n251,n252,n260);
or (n252,n253,n256,n259);
and (n253,n254,n255);
and (n254,n100,n96);
and (n255,n46,n148);
and (n256,n257,n258);
and (n257,n46,n96);
and (n258,n12,n148);
and (n259,n253,n258);
xor (n260,n261,n248);
xor (n261,n245,n246);
and (n262,n260,n263);
xor (n263,n224,n225);
and (n264,n252,n263);
and (n265,n250,n266);
xor (n266,n267,n229);
xor (n267,n223,n226);
and (n268,n243,n266);
and (n269,n270,n271);
xor (n270,n240,n241);
or (n271,n272,n300);
and (n272,n273,n275);
xor (n273,n274,n266);
xor (n274,n243,n250);
or (n275,n276,n296,n299);
and (n276,n277,n280);
and (n277,n278,n279);
and (n278,n178,n61);
and (n279,n100,n52);
or (n280,n281,n292,n295);
and (n281,n282,n291);
or (n282,n283,n288,n290);
and (n283,n284,n287);
and (n284,n285,n286);
and (n285,n178,n96);
and (n286,n100,n148);
and (n287,n178,n52);
and (n288,n287,n289);
xor (n289,n254,n255);
and (n290,n284,n289);
xor (n291,n278,n279);
and (n292,n291,n293);
xor (n293,n294,n258);
xor (n294,n253,n257);
and (n295,n282,n293);
and (n296,n280,n297);
xor (n297,n298,n263);
xor (n298,n252,n260);
and (n299,n277,n297);
and (n300,n301,n302);
xor (n301,n273,n275);
or (n302,n303,n325);
and (n303,n304,n306);
xor (n304,n305,n297);
xor (n305,n277,n280);
and (n306,n307,n323);
or (n307,n308,n319,n322);
and (n308,n309,n318);
or (n309,n310,n315,n317);
and (n310,n311,n314);
and (n311,n312,n313);
and (n312,n231,n96);
and (n313,n178,n148);
and (n314,n231,n52);
and (n315,n314,n316);
xor (n316,n285,n286);
and (n317,n311,n316);
and (n318,n231,n61);
and (n319,n318,n320);
xor (n320,n321,n289);
xor (n321,n284,n287);
and (n322,n309,n320);
xor (n323,n324,n293);
xor (n324,n282,n291);
and (n325,n326,n327);
xor (n326,n304,n306);
and (n327,n328,n329);
and (n328,n231,n22);
xor (n329,n307,n323);
xor (n330,n331,n399);
xor (n331,n332,n361);
xor (n332,n333,n357);
xor (n333,n334,n354);
or (n334,n335,n351,n353);
and (n335,n336,n348);
or (n336,n337,n344,n347);
and (n337,n338,n342);
nor (n338,n339,n341);
not (n339,n340);
and (n341,n14,n340);
and (n342,n343,n18);
and (n344,n342,n345);
and (n345,n346,n22);
and (n347,n338,n345);
nor (n348,n349,n350);
not (n349,n343);
and (n350,n14,n343);
and (n351,n348,n352);
and (n352,n346,n18);
and (n353,n336,n352);
nor (n354,n355,n356);
not (n355,n346);
and (n356,n14,n346);
nor (n357,n358,n37);
and (n358,n359,n18);
not (n359,n360);
or (n361,n362,n395,n398);
and (n362,n363,n393);
or (n363,n364,n389,n392);
and (n364,n365,n376);
or (n365,n366,n372,n375);
and (n366,n367,n371);
nor (n367,n368,n370);
not (n368,n369);
and (n370,n14,n369);
and (n371,n340,n18);
and (n372,n371,n373);
nor (n373,n374,n53);
and (n374,n359,n52);
and (n375,n367,n373);
or (n376,n377,n386,n388);
and (n377,n378,n385);
or (n378,n379,n382,n384);
and (n379,n380,n381);
and (n380,n340,n22);
and (n381,n343,n61);
and (n382,n381,n383);
and (n383,n346,n52);
and (n384,n380,n383);
and (n385,n343,n22);
and (n386,n385,n387);
and (n387,n346,n61);
and (n388,n378,n387);
and (n389,n376,n390);
xor (n390,n391,n345);
xor (n391,n338,n342);
and (n392,n365,n390);
nor (n393,n394,n75);
and (n394,n359,n22);
and (n395,n393,n396);
xor (n396,n397,n352);
xor (n397,n336,n348);
and (n398,n363,n396);
or (n399,n400,n436);
and (n400,n401,n403);
xor (n401,n402,n396);
xor (n402,n363,n393);
or (n403,n404,n432,n435);
and (n404,n405,n430);
or (n405,n406,n426,n429);
and (n406,n407,n424);
or (n407,n408,n420,n423);
and (n408,n409,n416);
or (n409,n410,n413,n415);
and (n410,n411,n412);
and (n411,n340,n61);
and (n412,n343,n52);
and (n413,n412,n414);
and (n414,n346,n96);
and (n415,n411,n414);
and (n416,n417,n419);
and (n417,n418,n18);
and (n419,n369,n22);
and (n420,n416,n421);
xor (n421,n422,n383);
xor (n422,n380,n381);
and (n423,n409,n421);
xor (n424,n425,n373);
xor (n425,n367,n371);
and (n426,n424,n427);
xor (n427,n428,n387);
xor (n428,n378,n385);
and (n429,n407,n427);
nor (n430,n431,n114);
and (n431,n359,n61);
and (n432,n430,n433);
xor (n433,n434,n390);
xor (n434,n365,n376);
and (n435,n405,n433);
and (n436,n437,n438);
xor (n437,n401,n403);
or (n438,n439,n480);
and (n439,n440,n442);
xor (n440,n441,n433);
xor (n441,n405,n430);
or (n442,n443,n476,n479);
and (n443,n444,n454);
or (n444,n445,n450,n453);
and (n445,n446,n449);
nor (n446,n447,n448);
not (n447,n418);
and (n448,n14,n418);
and (n449,n369,n18);
and (n450,n449,n451);
nor (n451,n452,n136);
and (n452,n359,n96);
and (n453,n446,n451);
or (n454,n455,n472,n475);
and (n455,n456,n470);
or (n456,n457,n467,n469);
and (n457,n458,n465);
or (n458,n459,n462,n464);
and (n459,n460,n461);
and (n460,n340,n52);
and (n461,n343,n96);
and (n462,n461,n463);
and (n463,n346,n148);
and (n464,n460,n463);
xor (n465,n466,n414);
xor (n466,n411,n412);
and (n467,n465,n468);
xor (n468,n417,n419);
and (n469,n458,n468);
xor (n470,n471,n451);
xor (n471,n446,n449);
and (n472,n470,n473);
xor (n473,n474,n421);
xor (n474,n409,n416);
and (n475,n456,n473);
and (n476,n454,n477);
xor (n477,n478,n427);
xor (n478,n407,n424);
and (n479,n444,n477);
and (n480,n481,n482);
xor (n481,n440,n442);
or (n482,n483,n528);
and (n483,n484,n486);
xor (n484,n485,n477);
xor (n485,n444,n454);
or (n486,n487,n524,n527);
and (n487,n488,n505);
or (n488,n489,n501,n504);
and (n489,n490,n498);
or (n490,n491,n495,n497);
and (n491,n492,n494);
and (n492,n493,n18);
and (n494,n418,n22);
and (n495,n494,n496);
and (n496,n369,n61);
and (n497,n492,n496);
nor (n498,n499,n500);
not (n499,n493);
and (n500,n14,n493);
and (n501,n498,n502);
nor (n502,n503,n189);
and (n503,n359,n148);
and (n504,n490,n502);
or (n505,n506,n520,n523);
and (n506,n507,n518);
or (n507,n508,n514,n517);
and (n508,n509,n512);
and (n509,n510,n511);
and (n510,n340,n96);
and (n511,n343,n148);
xor (n512,n513,n496);
xor (n513,n492,n494);
and (n514,n512,n515);
xor (n515,n516,n463);
xor (n516,n460,n461);
and (n517,n509,n515);
xor (n518,n519,n502);
xor (n519,n490,n498);
and (n520,n518,n521);
xor (n521,n522,n468);
xor (n522,n458,n465);
and (n523,n507,n521);
and (n524,n505,n525);
xor (n525,n526,n473);
xor (n526,n456,n470);
and (n527,n488,n525);
and (n528,n529,n530);
xor (n529,n484,n486);
or (n530,n531,n550);
and (n531,n532,n534);
xor (n532,n533,n525);
xor (n533,n488,n505);
and (n534,n535,n548);
or (n535,n536,n542,n547);
and (n536,n537,n540);
and (n537,n538,n539);
and (n538,n369,n52);
xor (n539,n510,n511);
xor (n540,n541,n515);
xor (n541,n509,n512);
and (n542,n540,n543);
nor (n543,n544,n546);
not (n544,n545);
and (n546,n14,n545);
and (n547,n537,n543);
xor (n548,n549,n521);
xor (n549,n507,n518);
and (n550,n551,n552);
xor (n551,n532,n534);
or (n552,n553,n583);
and (n553,n554,n555);
xor (n554,n535,n548);
or (n555,n556,n579,n582);
and (n556,n557,n564);
or (n557,n558,n561,n563);
and (n558,n559,n560);
and (n559,n545,n18);
and (n560,n493,n22);
and (n561,n560,n562);
and (n562,n418,n61);
and (n563,n559,n562);
or (n564,n565,n576,n578);
and (n565,n566,n574);
or (n566,n567,n570,n573);
and (n567,n568,n569);
and (n568,n418,n96);
and (n569,n369,n148);
and (n570,n571,n572);
and (n571,n369,n96);
and (n572,n340,n148);
and (n573,n567,n572);
xor (n574,n575,n562);
xor (n575,n559,n560);
and (n576,n574,n577);
xor (n577,n538,n539);
and (n578,n566,n577);
and (n579,n564,n580);
xor (n580,n581,n543);
xor (n581,n537,n540);
and (n582,n557,n580);
and (n583,n584,n585);
xor (n584,n554,n555);
or (n585,n586,n614);
and (n586,n587,n589);
xor (n587,n588,n580);
xor (n588,n557,n564);
or (n589,n590,n610,n613);
and (n590,n591,n594);
and (n591,n592,n593);
and (n592,n493,n61);
and (n593,n418,n52);
or (n594,n595,n606,n609);
and (n595,n596,n605);
or (n596,n597,n602,n604);
and (n597,n598,n601);
and (n598,n599,n600);
and (n599,n493,n96);
and (n600,n418,n148);
and (n601,n493,n52);
and (n602,n601,n603);
xor (n603,n568,n569);
and (n604,n598,n603);
xor (n605,n592,n593);
and (n606,n605,n607);
xor (n607,n608,n572);
xor (n608,n567,n571);
and (n609,n596,n607);
and (n610,n594,n611);
xor (n611,n612,n577);
xor (n612,n566,n574);
and (n613,n591,n611);
and (n614,n615,n616);
xor (n615,n587,n589);
or (n616,n617,n639);
and (n617,n618,n620);
xor (n618,n619,n611);
xor (n619,n591,n594);
and (n620,n621,n637);
or (n621,n622,n633,n636);
and (n622,n623,n632);
or (n623,n624,n629,n631);
and (n624,n625,n628);
and (n625,n626,n627);
and (n626,n545,n96);
and (n627,n493,n148);
and (n628,n545,n52);
and (n629,n628,n630);
xor (n630,n599,n600);
and (n631,n625,n630);
and (n632,n545,n61);
and (n633,n632,n634);
xor (n634,n635,n603);
xor (n635,n598,n601);
and (n636,n623,n634);
xor (n637,n638,n607);
xor (n638,n596,n605);
and (n639,n640,n641);
xor (n640,n618,n620);
and (n641,n642,n643);
and (n642,n545,n22);
xor (n643,n621,n637);
or (n644,n645,n648,n716);
and (n645,n646,n647);
xor (n646,n120,n121);
xor (n647,n437,n438);
and (n648,n647,n649);
or (n649,n650,n653,n715);
and (n650,n651,n652);
xor (n651,n166,n167);
xor (n652,n481,n482);
and (n653,n652,n654);
or (n654,n655,n658,n714);
and (n655,n656,n657);
xor (n656,n215,n216);
xor (n657,n529,n530);
and (n658,n657,n659);
or (n659,n660,n663,n713);
and (n660,n661,n662);
xor (n661,n237,n238);
xor (n662,n551,n552);
and (n663,n662,n664);
or (n664,n665,n668,n712);
and (n665,n666,n667);
xor (n666,n270,n271);
xor (n667,n584,n585);
and (n668,n667,n669);
or (n669,n670,n673,n711);
and (n670,n671,n672);
xor (n671,n301,n302);
xor (n672,n615,n616);
and (n673,n672,n674);
or (n674,n675,n678,n710);
and (n675,n676,n677);
xor (n676,n326,n327);
xor (n677,n640,n641);
and (n678,n677,n679);
or (n679,n680,n683,n709);
and (n680,n681,n682);
xor (n681,n328,n329);
xor (n682,n642,n643);
and (n683,n682,n684);
or (n684,n685,n690,n708);
and (n685,n686,n688);
xor (n686,n687,n320);
xor (n687,n309,n318);
xor (n688,n689,n634);
xor (n689,n623,n632);
and (n690,n688,n691);
or (n691,n692,n697,n707);
and (n692,n693,n695);
xor (n693,n694,n316);
xor (n694,n311,n314);
xor (n695,n696,n630);
xor (n696,n625,n628);
and (n697,n695,n698);
or (n698,n699,n702,n706);
and (n699,n700,n701);
xor (n700,n312,n313);
xor (n701,n626,n627);
and (n702,n701,n703);
and (n703,n704,n705);
and (n704,n231,n148);
and (n705,n545,n148);
and (n706,n700,n703);
and (n707,n693,n698);
and (n708,n686,n691);
and (n709,n681,n684);
and (n710,n676,n679);
and (n711,n671,n674);
and (n712,n666,n669);
and (n713,n661,n664);
and (n714,n656,n659);
and (n715,n651,n654);
and (n716,n646,n649);
xor (n717,n718,n847);
xor (n718,n719,n805);
xor (n719,n720,n795);
xor (n720,n721,n793);
or (n721,n722,n784,n792);
and (n722,n723,n767);
or (n723,n724,n750,n766);
and (n724,n725,n743);
nor (n725,n726,n742);
not (n726,n727);
xor (n727,n728,n729);
xor (n728,n12,n340);
or (n729,n730,n731,n741);
and (n730,n46,n369);
and (n731,n369,n732);
or (n732,n733,n734,n740);
and (n733,n100,n418);
and (n734,n418,n735);
or (n735,n736,n737,n739);
and (n736,n178,n493);
and (n737,n493,n738);
and (n738,n231,n545);
and (n739,n178,n738);
and (n740,n100,n735);
and (n741,n46,n732);
and (n742,n14,n727);
and (n743,n744,n18);
xor (n744,n745,n746);
xor (n745,n17,n343);
or (n746,n747,n748,n749);
and (n747,n12,n340);
and (n748,n340,n729);
and (n749,n12,n729);
and (n750,n743,n751);
nor (n751,n752,n53);
and (n752,n753,n52);
not (n753,n754);
or (n754,n755,n756,n765);
and (n755,n36,n360);
and (n756,n360,n757);
or (n757,n758,n759,n764);
and (n758,n21,n346);
and (n759,n346,n760);
or (n760,n761,n762,n763);
and (n761,n17,n343);
and (n762,n343,n746);
and (n763,n17,n746);
and (n764,n21,n760);
and (n765,n36,n757);
and (n766,n725,n751);
or (n767,n768,n781,n783);
and (n768,n769,n780);
or (n769,n770,n775,n779);
and (n770,n771,n772);
and (n771,n744,n22);
and (n772,n773,n61);
xor (n773,n774,n760);
xor (n774,n21,n346);
and (n775,n772,n776);
and (n776,n777,n52);
xor (n777,n778,n757);
xor (n778,n36,n360);
and (n779,n771,n776);
and (n780,n773,n22);
and (n781,n780,n782);
and (n782,n777,n61);
and (n783,n769,n782);
and (n784,n767,n785);
xor (n785,n786,n791);
xor (n786,n787,n790);
nor (n787,n788,n789);
not (n788,n744);
and (n789,n14,n744);
and (n790,n773,n18);
and (n791,n777,n22);
and (n792,n723,n785);
nor (n793,n794,n75);
and (n794,n753,n22);
xor (n795,n796,n804);
xor (n796,n797,n801);
or (n797,n798,n799,n800);
and (n798,n787,n790);
and (n799,n790,n791);
and (n800,n787,n791);
nor (n801,n802,n803);
not (n802,n773);
and (n803,n14,n773);
and (n804,n777,n18);
or (n805,n806,n843,n846);
and (n806,n807,n841);
or (n807,n808,n837,n840);
and (n808,n809,n835);
or (n809,n810,n831,n834);
and (n810,n811,n818);
or (n811,n812,n815,n817);
and (n812,n813,n814);
and (n813,n744,n61);
and (n814,n773,n52);
and (n815,n814,n816);
and (n816,n777,n96);
and (n817,n813,n816);
or (n818,n819,n828,n830);
and (n819,n820,n825);
nor (n820,n821,n824);
not (n821,n822);
xor (n822,n823,n735);
xor (n823,n100,n418);
and (n824,n14,n822);
and (n825,n826,n18);
xor (n826,n827,n732);
xor (n827,n46,n369);
and (n828,n825,n829);
and (n829,n727,n22);
and (n830,n820,n829);
and (n831,n818,n832);
xor (n832,n833,n776);
xor (n833,n771,n772);
and (n834,n811,n832);
xor (n835,n836,n751);
xor (n836,n725,n743);
and (n837,n835,n838);
xor (n838,n839,n782);
xor (n839,n769,n780);
and (n840,n809,n838);
nor (n841,n842,n114);
and (n842,n753,n61);
and (n843,n841,n844);
xor (n844,n845,n785);
xor (n845,n723,n767);
and (n846,n807,n844);
or (n847,n848,n890);
and (n848,n849,n851);
xor (n849,n850,n844);
xor (n850,n807,n841);
or (n851,n852,n886,n889);
and (n852,n853,n863);
or (n853,n854,n859,n862);
and (n854,n855,n858);
nor (n855,n856,n857);
not (n856,n826);
and (n857,n14,n826);
and (n858,n727,n18);
and (n859,n858,n860);
nor (n860,n861,n136);
and (n861,n753,n96);
and (n862,n855,n860);
or (n863,n864,n882,n885);
and (n864,n865,n880);
or (n865,n866,n876,n879);
and (n866,n867,n874);
or (n867,n868,n871,n873);
and (n868,n869,n870);
and (n869,n744,n52);
and (n870,n773,n96);
and (n871,n870,n872);
and (n872,n777,n148);
and (n873,n869,n872);
xor (n874,n875,n816);
xor (n875,n813,n814);
and (n876,n874,n877);
xor (n877,n878,n829);
xor (n878,n820,n825);
and (n879,n867,n877);
xor (n880,n881,n860);
xor (n881,n855,n858);
and (n882,n880,n883);
xor (n883,n884,n832);
xor (n884,n811,n818);
and (n885,n865,n883);
and (n886,n863,n887);
xor (n887,n888,n838);
xor (n888,n809,n835);
and (n889,n853,n887);
and (n890,n891,n892);
xor (n891,n849,n851);
or (n892,n893,n932);
and (n893,n894,n896);
xor (n894,n895,n887);
xor (n895,n853,n863);
or (n896,n897,n928,n931);
and (n897,n898,n908);
and (n898,n899,n906);
or (n899,n900,n903,n905);
and (n900,n901,n902);
and (n901,n822,n18);
and (n902,n826,n22);
and (n903,n902,n904);
and (n904,n727,n61);
and (n905,n901,n904);
nor (n906,n907,n189);
and (n907,n753,n148);
or (n908,n909,n925,n927);
and (n909,n910,n923);
or (n910,n911,n919,n922);
and (n911,n912,n917);
nor (n912,n913,n916);
not (n913,n914);
xor (n914,n915,n738);
xor (n915,n178,n493);
and (n916,n14,n914);
xor (n917,n918,n872);
xor (n918,n869,n870);
and (n919,n917,n920);
xor (n920,n921,n904);
xor (n921,n901,n902);
and (n922,n912,n920);
xor (n923,n924,n877);
xor (n924,n867,n874);
and (n925,n923,n926);
xor (n926,n899,n906);
and (n927,n910,n926);
and (n928,n908,n929);
xor (n929,n930,n883);
xor (n930,n865,n880);
and (n931,n898,n929);
and (n932,n933,n934);
xor (n933,n894,n896);
or (n934,n935,n972);
and (n935,n936,n938);
xor (n936,n937,n929);
xor (n937,n898,n908);
or (n938,n939,n968,n971);
and (n939,n940,n951);
and (n940,n941,n948);
or (n941,n942,n945,n947);
and (n942,n943,n944);
and (n943,n822,n22);
and (n944,n826,n61);
and (n945,n944,n946);
and (n946,n727,n52);
and (n947,n943,n946);
and (n948,n949,n950);
and (n949,n744,n96);
and (n950,n773,n148);
or (n951,n952,n964,n967);
and (n952,n953,n963);
or (n953,n954,n960,n962);
and (n954,n955,n958);
and (n955,n956,n957);
and (n956,n727,n96);
and (n957,n744,n148);
xor (n958,n959,n946);
xor (n959,n943,n944);
and (n960,n958,n961);
xor (n961,n949,n950);
and (n962,n955,n961);
xor (n963,n941,n948);
and (n964,n963,n965);
xor (n965,n966,n920);
xor (n966,n912,n917);
and (n967,n953,n965);
and (n968,n951,n969);
xor (n969,n970,n926);
xor (n970,n910,n923);
and (n971,n940,n969);
and (n972,n973,n974);
xor (n973,n936,n938);
or (n974,n975,n1000);
and (n975,n976,n978);
xor (n976,n977,n969);
xor (n977,n940,n951);
or (n978,n979,n996,n999);
and (n979,n980,n986);
and (n980,n981,n985);
nor (n981,n982,n984);
not (n982,n983);
xor (n983,n231,n545);
and (n984,n14,n983);
and (n985,n914,n18);
or (n986,n987,n993,n995);
and (n987,n988,n991);
and (n988,n989,n990);
and (n989,n826,n52);
xor (n990,n956,n957);
xor (n991,n992,n961);
xor (n992,n955,n958);
and (n993,n991,n994);
xor (n994,n981,n985);
and (n995,n988,n994);
and (n996,n986,n997);
xor (n997,n998,n965);
xor (n998,n953,n963);
and (n999,n980,n997);
and (n1000,n1001,n1002);
xor (n1001,n976,n978);
or (n1002,n1003,n1034);
and (n1003,n1004,n1006);
xor (n1004,n1005,n997);
xor (n1005,n980,n986);
or (n1006,n1007,n1030,n1033);
and (n1007,n1008,n1015);
or (n1008,n1009,n1012,n1014);
and (n1009,n1010,n1011);
and (n1010,n983,n18);
and (n1011,n914,n22);
and (n1012,n1011,n1013);
and (n1013,n822,n61);
and (n1014,n1010,n1013);
or (n1015,n1016,n1027,n1029);
and (n1016,n1017,n1025);
or (n1017,n1018,n1021,n1024);
and (n1018,n1019,n1020);
and (n1019,n822,n96);
and (n1020,n826,n148);
and (n1021,n1022,n1023);
and (n1022,n826,n96);
and (n1023,n727,n148);
and (n1024,n1018,n1023);
xor (n1025,n1026,n1013);
xor (n1026,n1010,n1011);
and (n1027,n1025,n1028);
xor (n1028,n989,n990);
and (n1029,n1017,n1028);
and (n1030,n1015,n1031);
xor (n1031,n1032,n994);
xor (n1032,n988,n991);
and (n1033,n1008,n1031);
and (n1034,n1035,n1036);
xor (n1035,n1004,n1006);
or (n1036,n1037,n1065);
and (n1037,n1038,n1040);
xor (n1038,n1039,n1031);
xor (n1039,n1008,n1015);
or (n1040,n1041,n1061,n1064);
and (n1041,n1042,n1045);
and (n1042,n1043,n1044);
and (n1043,n914,n61);
and (n1044,n822,n52);
or (n1045,n1046,n1057,n1060);
and (n1046,n1047,n1056);
or (n1047,n1048,n1053,n1055);
and (n1048,n1049,n1052);
and (n1049,n1050,n1051);
and (n1050,n914,n96);
and (n1051,n822,n148);
and (n1052,n914,n52);
and (n1053,n1052,n1054);
xor (n1054,n1019,n1020);
and (n1055,n1049,n1054);
xor (n1056,n1043,n1044);
and (n1057,n1056,n1058);
xor (n1058,n1059,n1023);
xor (n1059,n1018,n1022);
and (n1060,n1047,n1058);
and (n1061,n1045,n1062);
xor (n1062,n1063,n1028);
xor (n1063,n1017,n1025);
and (n1064,n1042,n1062);
and (n1065,n1066,n1067);
xor (n1066,n1038,n1040);
or (n1067,n1068,n1090);
and (n1068,n1069,n1071);
xor (n1069,n1070,n1062);
xor (n1070,n1042,n1045);
and (n1071,n1072,n1088);
or (n1072,n1073,n1084,n1087);
and (n1073,n1074,n1083);
or (n1074,n1075,n1080,n1082);
and (n1075,n1076,n1079);
and (n1076,n1077,n1078);
and (n1077,n983,n96);
and (n1078,n914,n148);
and (n1079,n983,n52);
and (n1080,n1079,n1081);
xor (n1081,n1050,n1051);
and (n1082,n1076,n1081);
and (n1083,n983,n61);
and (n1084,n1083,n1085);
xor (n1085,n1086,n1054);
xor (n1086,n1049,n1052);
and (n1087,n1074,n1085);
xor (n1088,n1089,n1058);
xor (n1089,n1047,n1056);
and (n1090,n1091,n1092);
xor (n1091,n1069,n1071);
and (n1092,n1093,n1094);
and (n1093,n983,n22);
xor (n1094,n1072,n1088);
endmodule
