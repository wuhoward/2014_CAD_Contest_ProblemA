module top (out,n18,n19,n25,n29,n35,n42,n43,n47,n48
        ,n55,n65,n77,n84,n85,n95,n103,n105,n113,n121
        ,n130,n137,n143,n185,n188,n194,n203,n219,n808);
output out;
input n18;
input n19;
input n25;
input n29;
input n35;
input n42;
input n43;
input n47;
input n48;
input n55;
input n65;
input n77;
input n84;
input n85;
input n95;
input n103;
input n105;
input n113;
input n121;
input n130;
input n137;
input n143;
input n185;
input n188;
input n194;
input n203;
input n219;
input n808;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n20;
wire n21;
wire n22;
wire n23;
wire n24;
wire n26;
wire n27;
wire n28;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n44;
wire n45;
wire n46;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n104;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n186;
wire n187;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
xor (out,n0,n834);
nand (n0,n1,n833);
or (n1,n2,n758);
nand (n2,n3,n754);
or (n3,n4,n345);
nor (n4,n5,n313);
xor (n5,n6,n260);
xor (n6,n7,n149);
nand (n7,n8,n147);
or (n8,n9,n67);
or (n9,n10,n66);
and (n10,n11,n64);
xor (n11,n12,n38);
nand (n12,n13,n32);
or (n13,n14,n27);
nand (n14,n15,n22);
nor (n15,n16,n20);
and (n16,n17,n19);
not (n17,n18);
and (n20,n18,n21);
not (n21,n19);
nand (n22,n23,n26);
or (n23,n19,n24);
not (n24,n25);
nand (n26,n24,n19);
nor (n27,n28,n30);
and (n28,n24,n29);
and (n30,n25,n31);
not (n31,n29);
or (n32,n33,n15);
nor (n33,n34,n36);
and (n34,n35,n24);
and (n36,n25,n37);
not (n37,n35);
nand (n38,n39,n51);
or (n39,n40,n44);
not (n40,n41);
xor (n41,n42,n43);
nor (n44,n45,n49);
and (n45,n46,n48);
not (n46,n47);
and (n49,n47,n50);
not (n50,n48);
nand (n51,n52,n59);
not (n52,n53);
nor (n53,n54,n57);
and (n54,n55,n56);
not (n56,n43);
and (n57,n58,n43);
not (n58,n55);
not (n59,n60);
nand (n60,n44,n61);
nand (n61,n62,n63);
or (n62,n50,n43);
nand (n63,n50,n43);
and (n64,n43,n65);
and (n66,n12,n38);
not (n67,n68);
or (n68,n69,n146);
and (n69,n70,n123);
xor (n70,n71,n98);
nand (n71,n72,n91);
or (n72,n73,n79);
not (n73,n74);
nand (n74,n75,n78);
or (n75,n18,n76);
not (n76,n77);
or (n78,n17,n77);
not (n79,n80);
nor (n80,n81,n87);
nand (n81,n82,n86);
or (n82,n83,n85);
not (n83,n84);
nand (n86,n83,n85);
nor (n87,n88,n89);
and (n88,n17,n85);
and (n89,n18,n90);
not (n90,n85);
nand (n91,n92,n81);
not (n92,n93);
nor (n93,n94,n96);
and (n94,n17,n95);
and (n96,n18,n97);
not (n97,n95);
nand (n98,n99,n116);
or (n99,n100,n111);
nand (n100,n101,n107);
nand (n101,n102,n106);
or (n102,n103,n104);
not (n104,n105);
nand (n106,n104,n103);
not (n107,n108);
nand (n108,n109,n110);
or (n109,n24,n103);
nand (n110,n24,n103);
nor (n111,n112,n114);
and (n112,n104,n113);
and (n114,n105,n115);
not (n115,n113);
or (n116,n107,n117);
not (n117,n118);
nor (n118,n119,n122);
and (n119,n120,n104);
not (n120,n121);
and (n122,n105,n121);
nand (n123,n124,n140);
or (n124,n125,n135);
not (n125,n126);
and (n126,n127,n132);
not (n127,n128);
nand (n128,n129,n131);
or (n129,n130,n104);
nand (n131,n130,n104);
nand (n132,n133,n134);
or (n133,n130,n46);
nand (n134,n46,n130);
nor (n135,n136,n138);
and (n136,n46,n137);
and (n138,n47,n139);
not (n139,n137);
or (n140,n127,n141);
nor (n141,n142,n144);
and (n142,n46,n143);
and (n144,n47,n145);
not (n145,n143);
and (n146,n71,n98);
or (n147,n68,n148);
not (n148,n9);
xor (n149,n150,n206);
xor (n150,n151,n171);
xor (n151,n152,n165);
xor (n152,n153,n159);
nand (n153,n154,n155);
or (n154,n117,n100);
nand (n155,n108,n156);
nor (n156,n157,n158);
and (n157,n31,n104);
and (n158,n105,n29);
nand (n159,n160,n161);
or (n160,n125,n141);
nand (n161,n128,n162);
nand (n162,n163,n164);
or (n163,n47,n115);
or (n164,n46,n113);
nand (n165,n166,n167);
or (n166,n14,n33);
or (n167,n15,n168);
nor (n168,n169,n170);
and (n169,n77,n24);
and (n170,n25,n76);
xor (n171,n172,n180);
xor (n172,n173,n179);
nand (n173,n174,n175);
or (n174,n40,n60);
or (n175,n44,n176);
nor (n176,n177,n178);
and (n177,n137,n56);
and (n178,n43,n139);
and (n179,n43,n55);
xor (n180,n181,n197);
nand (n181,n182,n191);
or (n182,n183,n186);
nand (n183,n84,n184);
not (n184,n185);
nor (n186,n187,n189);
and (n187,n83,n188);
and (n189,n84,n190);
not (n190,n188);
or (n191,n192,n184);
nor (n192,n193,n195);
and (n193,n83,n194);
and (n195,n84,n196);
not (n196,n194);
nand (n197,n198,n199);
or (n198,n79,n93);
or (n199,n200,n201);
not (n200,n81);
nor (n201,n202,n204);
and (n202,n17,n203);
and (n204,n18,n205);
not (n205,n203);
or (n206,n207,n259);
and (n207,n208,n233);
xor (n208,n209,n215);
nand (n209,n210,n214);
or (n210,n183,n211);
nor (n211,n212,n213);
and (n212,n83,n203);
and (n213,n84,n205);
or (n214,n186,n184);
or (n215,n216,n232);
and (n216,n217,n226);
xor (n217,n218,n220);
and (n218,n43,n219);
nand (n220,n221,n222);
or (n221,n200,n73);
nand (n222,n80,n223);
nand (n223,n224,n225);
or (n224,n18,n37);
or (n225,n17,n35);
nand (n226,n227,n231);
or (n227,n100,n228);
nor (n228,n229,n230);
and (n229,n104,n143);
and (n230,n105,n145);
or (n231,n111,n107);
and (n232,n218,n220);
or (n233,n234,n258);
and (n234,n235,n251);
xor (n235,n236,n245);
nand (n236,n237,n243);
or (n237,n238,n125);
not (n238,n239);
nor (n239,n240,n242);
and (n240,n241,n46);
not (n241,n42);
and (n242,n47,n42);
nand (n243,n244,n128);
not (n244,n135);
nand (n245,n246,n250);
or (n246,n247,n183);
nor (n247,n248,n249);
and (n248,n83,n95);
and (n249,n84,n97);
or (n250,n211,n184);
nand (n251,n252,n257);
or (n252,n60,n253);
nor (n253,n254,n255);
and (n254,n56,n65);
and (n255,n43,n256);
not (n256,n65);
or (n257,n44,n53);
and (n258,n236,n245);
and (n259,n209,n215);
or (n260,n261,n312);
and (n261,n262,n265);
xor (n262,n263,n264);
xor (n263,n11,n64);
xor (n264,n70,n123);
or (n265,n266,n311);
and (n266,n267,n289);
xor (n267,n268,n274);
nand (n268,n269,n273);
or (n269,n14,n270);
nor (n270,n271,n272);
and (n271,n24,n121);
and (n272,n25,n120);
or (n273,n15,n27);
nor (n274,n275,n283);
not (n275,n276);
nand (n276,n277,n282);
or (n277,n278,n79);
not (n278,n279);
nand (n279,n280,n281);
or (n280,n18,n31);
or (n281,n17,n29);
nand (n282,n81,n223);
nand (n283,n284,n43);
nand (n284,n285,n286);
or (n285,n47,n48);
nand (n286,n287,n288);
or (n287,n50,n46);
not (n288,n219);
or (n289,n290,n310);
and (n290,n291,n304);
xor (n291,n292,n298);
nand (n292,n293,n297);
or (n293,n100,n294);
nor (n294,n295,n296);
and (n295,n104,n137);
and (n296,n105,n139);
or (n297,n107,n228);
nand (n298,n299,n303);
or (n299,n125,n300);
nor (n300,n301,n302);
and (n301,n46,n55);
and (n302,n47,n58);
or (n303,n127,n238);
nand (n304,n305,n309);
or (n305,n306,n183);
nor (n306,n307,n308);
and (n307,n83,n77);
and (n308,n84,n76);
or (n309,n247,n184);
and (n310,n292,n298);
and (n311,n268,n274);
and (n312,n263,n264);
or (n313,n314,n344);
and (n314,n315,n343);
xor (n315,n316,n317);
xor (n316,n208,n233);
or (n317,n318,n342);
and (n318,n319,n322);
xor (n319,n320,n321);
xor (n320,n235,n251);
xor (n321,n217,n226);
or (n322,n323,n341);
and (n323,n324,n337);
xor (n324,n325,n331);
nand (n325,n326,n330);
or (n326,n60,n327);
nor (n327,n328,n329);
and (n328,n219,n56);
and (n329,n288,n43);
or (n330,n44,n253);
nand (n331,n332,n336);
or (n332,n14,n333);
nor (n333,n334,n335);
and (n334,n24,n113);
and (n335,n25,n115);
or (n336,n15,n270);
nand (n337,n338,n340);
or (n338,n339,n275);
not (n339,n283);
or (n340,n276,n283);
and (n341,n325,n331);
and (n342,n320,n321);
xor (n343,n262,n265);
and (n344,n316,n317);
not (n345,n346);
nand (n346,n347,n749);
or (n347,n348,n458);
not (n348,n349);
nor (n349,n350,n453);
not (n350,n351);
or (n351,n352,n446);
or (n352,n353,n445);
and (n353,n354,n402);
xor (n354,n355,n356);
xor (n355,n324,n337);
xor (n356,n357,n401);
xor (n357,n358,n377);
or (n358,n359,n376);
and (n359,n360,n368);
xor (n360,n361,n362);
nor (n361,n44,n288);
nand (n362,n363,n367);
or (n363,n364,n79);
nor (n364,n365,n366);
and (n365,n120,n18);
and (n366,n121,n17);
nand (n367,n279,n81);
nand (n368,n369,n374);
or (n369,n370,n100);
not (n370,n371);
nand (n371,n372,n373);
or (n372,n105,n241);
or (n373,n104,n42);
nand (n374,n375,n108);
not (n375,n294);
and (n376,n361,n362);
or (n377,n378,n400);
and (n378,n379,n394);
xor (n379,n380,n388);
nand (n380,n381,n386);
or (n381,n382,n125);
not (n382,n383);
nand (n383,n384,n385);
or (n384,n47,n256);
or (n385,n46,n65);
nand (n386,n387,n128);
not (n387,n300);
nand (n388,n389,n393);
or (n389,n390,n183);
nor (n390,n391,n392);
and (n391,n83,n35);
and (n392,n84,n37);
or (n393,n306,n184);
nand (n394,n395,n399);
or (n395,n14,n396);
nor (n396,n397,n398);
and (n397,n24,n143);
and (n398,n25,n145);
or (n399,n15,n333);
and (n400,n380,n388);
xor (n401,n291,n304);
or (n402,n403,n444);
and (n403,n404,n443);
xor (n404,n405,n419);
and (n405,n406,n412);
and (n406,n407,n47);
nand (n407,n408,n409);
or (n408,n105,n130);
nand (n409,n410,n288);
or (n410,n411,n104);
not (n411,n130);
nand (n412,n413,n418);
or (n413,n414,n79);
not (n414,n415);
nand (n415,n416,n417);
or (n416,n18,n115);
or (n417,n17,n113);
or (n418,n200,n364);
or (n419,n420,n442);
and (n420,n421,n435);
xor (n421,n422,n428);
nand (n422,n423,n424);
or (n423,n107,n370);
or (n424,n425,n100);
nor (n425,n426,n427);
and (n426,n58,n105);
and (n427,n55,n104);
nand (n428,n429,n434);
or (n429,n430,n125);
not (n430,n431);
nand (n431,n432,n433);
or (n432,n47,n288);
or (n433,n46,n219);
nand (n434,n383,n128);
nand (n435,n436,n441);
or (n436,n437,n183);
not (n437,n438);
nor (n438,n439,n440);
and (n439,n31,n83);
and (n440,n84,n29);
or (n441,n390,n184);
and (n442,n422,n428);
xor (n443,n360,n368);
and (n444,n405,n419);
and (n445,n355,n356);
xor (n446,n447,n452);
xor (n447,n448,n449);
xor (n448,n267,n289);
or (n449,n450,n451);
and (n450,n357,n401);
and (n451,n358,n377);
xor (n452,n319,n322);
nor (n453,n454,n455);
xor (n454,n315,n343);
or (n455,n456,n457);
and (n456,n447,n452);
and (n457,n448,n449);
not (n458,n459);
nand (n459,n460,n737,n748);
nand (n460,n461,n499,n598);
nand (n461,n462,n464);
not (n462,n463);
xor (n463,n354,n402);
not (n464,n465);
or (n465,n466,n498);
and (n466,n467,n497);
xor (n467,n468,n469);
xor (n468,n379,n394);
or (n469,n470,n496);
and (n470,n471,n479);
xor (n471,n472,n478);
nand (n472,n473,n477);
or (n473,n14,n474);
nor (n474,n475,n476);
and (n475,n24,n137);
and (n476,n25,n139);
or (n477,n396,n15);
xor (n478,n406,n412);
or (n479,n480,n495);
and (n480,n481,n489);
xor (n481,n482,n483);
and (n482,n128,n219);
nand (n483,n484,n485);
or (n484,n184,n437);
or (n485,n486,n183);
nor (n486,n487,n488);
and (n487,n83,n121);
and (n488,n84,n120);
nand (n489,n490,n494);
or (n490,n100,n491);
nor (n491,n492,n493);
and (n492,n104,n65);
and (n493,n105,n256);
or (n494,n107,n425);
and (n495,n482,n483);
and (n496,n472,n478);
xor (n497,n404,n443);
and (n498,n468,n469);
nor (n499,n500,n593);
not (n500,n501);
nor (n501,n502,n566);
nor (n502,n503,n538);
xor (n503,n504,n537);
xor (n504,n505,n506);
xor (n505,n421,n435);
or (n506,n507,n536);
and (n507,n508,n522);
xor (n508,n509,n516);
nand (n509,n510,n515);
or (n510,n511,n79);
not (n511,n512);
nand (n512,n513,n514);
or (n513,n18,n145);
or (n514,n17,n143);
nand (n515,n81,n415);
nand (n516,n517,n521);
or (n517,n14,n518);
nor (n518,n519,n520);
and (n519,n42,n24);
and (n520,n25,n241);
or (n521,n15,n474);
and (n522,n523,n529);
nor (n523,n524,n104);
nor (n524,n525,n527);
and (n525,n526,n288);
nand (n526,n25,n103);
and (n527,n24,n528);
not (n528,n103);
nand (n529,n530,n535);
or (n530,n183,n531);
not (n531,n532);
nor (n532,n533,n534);
and (n533,n84,n113);
and (n534,n115,n83);
or (n535,n486,n184);
and (n536,n509,n516);
xor (n537,n471,n479);
or (n538,n539,n565);
and (n539,n540,n564);
xor (n540,n541,n563);
or (n541,n542,n562);
and (n542,n543,n556);
xor (n543,n544,n550);
nand (n544,n545,n549);
or (n545,n100,n546);
nor (n546,n547,n548);
and (n547,n104,n219);
and (n548,n105,n288);
or (n549,n491,n107);
nand (n550,n551,n552);
or (n551,n511,n200);
nand (n552,n80,n553);
nand (n553,n554,n555);
or (n554,n18,n139);
or (n555,n17,n137);
nand (n556,n557,n561);
or (n557,n14,n558);
nor (n558,n559,n560);
and (n559,n24,n55);
and (n560,n25,n58);
or (n561,n15,n518);
and (n562,n544,n550);
xor (n563,n481,n489);
xor (n564,n508,n522);
and (n565,n541,n563);
nor (n566,n567,n568);
xor (n567,n540,n564);
or (n568,n569,n592);
and (n569,n570,n591);
xor (n570,n571,n572);
xor (n571,n523,n529);
or (n572,n573,n590);
and (n573,n574,n583);
xor (n574,n575,n576);
and (n575,n108,n219);
nand (n576,n577,n578);
or (n577,n184,n531);
or (n578,n579,n183);
not (n579,n580);
nand (n580,n581,n582);
or (n581,n143,n83);
nand (n582,n83,n143);
nand (n583,n584,n589);
or (n584,n585,n79);
not (n585,n586);
nor (n586,n587,n588);
and (n587,n18,n42);
and (n588,n241,n17);
nand (n589,n81,n553);
and (n590,n575,n576);
xor (n591,n543,n556);
and (n592,n571,n572);
nor (n593,n594,n595);
xor (n594,n467,n497);
or (n595,n596,n597);
and (n596,n504,n537);
and (n597,n505,n506);
or (n598,n599,n736);
and (n599,n600,n627);
xor (n600,n601,n626);
or (n601,n602,n625);
and (n602,n603,n624);
xor (n603,n604,n610);
nand (n604,n605,n609);
or (n605,n14,n606);
nor (n606,n607,n608);
and (n607,n24,n65);
and (n608,n25,n256);
or (n609,n15,n558);
and (n610,n611,n618);
nand (n611,n612,n617);
or (n612,n183,n613);
not (n613,n614);
nor (n614,n615,n616);
and (n615,n84,n137);
and (n616,n139,n83);
nand (n617,n580,n185);
not (n618,n619);
nand (n619,n620,n25);
nand (n620,n621,n622);
or (n621,n18,n19);
nand (n622,n623,n288);
or (n623,n21,n17);
xor (n624,n574,n583);
and (n625,n604,n610);
xor (n626,n570,n591);
or (n627,n628,n735);
and (n628,n629,n653);
xor (n629,n630,n652);
or (n630,n631,n651);
and (n631,n632,n647);
xor (n632,n633,n640);
nand (n633,n634,n639);
or (n634,n635,n79);
not (n635,n636);
nand (n636,n637,n638);
or (n637,n18,n58);
or (n638,n17,n55);
nand (n639,n81,n586);
nand (n640,n641,n646);
or (n641,n642,n14);
not (n642,n643);
nand (n643,n644,n645);
or (n644,n288,n25);
or (n645,n24,n219);
or (n646,n15,n606);
nand (n647,n648,n650);
or (n648,n618,n649);
not (n649,n611);
or (n650,n611,n619);
and (n651,n633,n640);
xor (n652,n603,n624);
or (n653,n654,n734);
and (n654,n655,n676);
xor (n655,n656,n675);
or (n656,n657,n674);
and (n657,n658,n667);
xor (n658,n659,n660);
nor (n659,n15,n288);
nand (n660,n661,n666);
or (n661,n662,n79);
not (n662,n663);
nor (n663,n664,n665);
and (n664,n256,n17);
and (n665,n18,n65);
nand (n666,n81,n636);
nand (n667,n668,n673);
or (n668,n183,n669);
not (n669,n670);
nor (n670,n671,n672);
and (n671,n241,n83);
and (n672,n84,n42);
or (n673,n613,n184);
and (n674,n659,n660);
xor (n675,n632,n647);
or (n676,n677,n733);
and (n677,n678,n732);
xor (n678,n679,n693);
nor (n679,n680,n688);
not (n680,n681);
nand (n681,n682,n683);
or (n682,n184,n669);
nand (n683,n684,n687);
nor (n684,n685,n686);
and (n685,n58,n83);
and (n686,n84,n55);
not (n687,n183);
nand (n688,n689,n18);
nand (n689,n690,n691);
or (n690,n85,n84);
or (n691,n692,n219);
and (n692,n84,n85);
nand (n693,n694,n731);
or (n694,n695,n719);
not (n695,n696);
nand (n696,n697,n718);
or (n697,n698,n707);
nor (n698,n699,n700);
and (n699,n81,n219);
nand (n700,n701,n703);
or (n701,n184,n702);
not (n702,n684);
nand (n703,n704,n687);
nand (n704,n705,n706);
or (n705,n256,n84);
or (n706,n83,n65);
nand (n707,n708,n711);
not (n708,n709);
nand (n709,n710,n84);
nand (n710,n219,n185);
nand (n711,n712,n714);
or (n712,n184,n713);
not (n713,n704);
nand (n714,n715,n687);
nor (n715,n716,n717);
and (n716,n288,n83);
and (n717,n84,n219);
nand (n718,n699,n700);
not (n719,n720);
nand (n720,n721,n725);
nor (n721,n722,n723);
and (n722,n688,n681);
and (n723,n724,n680);
not (n724,n688);
nor (n725,n726,n730);
and (n726,n80,n727);
nand (n727,n728,n729);
or (n728,n18,n288);
or (n729,n17,n219);
and (n730,n81,n663);
or (n731,n721,n725);
xor (n732,n658,n667);
and (n733,n679,n693);
and (n734,n656,n675);
and (n735,n630,n652);
and (n736,n601,n626);
nand (n737,n738,n461);
nand (n738,n739,n747);
or (n739,n593,n740);
nand (n740,n741,n746);
or (n741,n742,n744);
not (n742,n743);
nand (n743,n567,n568);
not (n744,n745);
nand (n745,n503,n538);
not (n746,n502);
nand (n747,n594,n595);
nand (n748,n463,n465);
not (n749,n750);
nand (n750,n751,n753);
or (n751,n453,n752);
nand (n752,n446,n352);
nand (n753,n454,n455);
not (n754,n755);
nor (n755,n756,n757);
not (n756,n5);
not (n757,n313);
nand (n758,n759,n831);
not (n759,n760);
and (n760,n761,n828);
xor (n761,n762,n825);
xor (n762,n763,n791);
xor (n763,n764,n769);
xor (n764,n765,n766);
and (n765,n181,n197);
or (n766,n767,n768);
and (n767,n152,n165);
and (n768,n153,n159);
xor (n769,n770,n785);
xor (n770,n771,n778);
nand (n771,n772,n774);
or (n772,n773,n100);
not (n773,n156);
nand (n774,n775,n108);
nor (n775,n776,n777);
and (n776,n37,n104);
and (n777,n35,n105);
nand (n778,n779,n781);
or (n779,n780,n125);
not (n780,n162);
nand (n781,n128,n782);
nor (n782,n783,n784);
and (n783,n120,n46);
and (n784,n121,n47);
nand (n785,n786,n787);
or (n786,n14,n168);
or (n787,n788,n15);
nor (n788,n789,n790);
and (n789,n24,n95);
and (n790,n25,n97);
xor (n791,n792,n824);
xor (n792,n793,n821);
xor (n793,n794,n802);
xor (n794,n795,n801);
nand (n795,n796,n797);
or (n796,n60,n176);
or (n797,n798,n44);
nor (n798,n799,n800);
and (n799,n143,n56);
and (n800,n43,n145);
and (n801,n43,n42);
xor (n802,n803,n813);
nand (n803,n804,n811);
or (n804,n184,n805);
not (n805,n806);
nor (n806,n807,n809);
and (n807,n808,n84);
and (n809,n810,n83);
not (n810,n808);
nand (n811,n812,n687);
not (n812,n192);
nand (n813,n814,n819);
or (n814,n200,n815);
not (n815,n816);
nand (n816,n817,n818);
or (n817,n18,n190);
or (n818,n17,n188);
nand (n819,n820,n80);
not (n820,n201);
or (n821,n822,n823);
and (n822,n172,n180);
and (n823,n173,n179);
and (n824,n68,n9);
or (n825,n826,n827);
and (n826,n150,n206);
and (n827,n151,n171);
or (n828,n829,n830);
and (n829,n6,n260);
and (n830,n7,n149);
not (n831,n832);
nor (n832,n761,n828);
nand (n833,n2,n758);
xor (n834,n835,n1417);
xor (n835,n836,n1414);
xor (n836,n837,n1413);
xor (n837,n838,n1404);
xor (n838,n839,n1403);
xor (n839,n840,n1388);
xor (n840,n841,n1387);
xor (n841,n842,n1366);
xor (n842,n843,n1365);
xor (n843,n844,n1338);
xor (n844,n845,n1337);
xor (n845,n846,n1304);
xor (n846,n847,n1303);
xor (n847,n848,n1265);
xor (n848,n849,n158);
xor (n849,n850,n1221);
xor (n850,n851,n1220);
xor (n851,n852,n1170);
xor (n852,n853,n1169);
xor (n853,n854,n1112);
xor (n854,n855,n1111);
xor (n855,n856,n1049);
xor (n856,n857,n1048);
or (n857,n858,n986);
and (n858,n859,n801);
or (n859,n860,n922);
and (n860,n861,n179);
and (n861,n64,n862);
or (n862,n863,n865);
and (n863,n218,n864);
and (n864,n48,n65);
and (n865,n866,n867);
xor (n866,n218,n864);
or (n867,n868,n871);
and (n868,n869,n870);
and (n869,n48,n219);
and (n870,n47,n65);
and (n871,n872,n873);
xor (n872,n869,n870);
or (n873,n874,n877);
and (n874,n875,n876);
and (n875,n47,n219);
and (n876,n130,n65);
and (n877,n878,n879);
xor (n878,n875,n876);
or (n879,n880,n883);
and (n880,n881,n882);
and (n881,n130,n219);
and (n882,n105,n65);
and (n883,n884,n885);
xor (n884,n881,n882);
or (n885,n886,n889);
and (n886,n887,n888);
and (n887,n105,n219);
and (n888,n103,n65);
and (n889,n890,n891);
xor (n890,n887,n888);
or (n891,n892,n895);
and (n892,n893,n894);
and (n893,n103,n219);
and (n894,n25,n65);
and (n895,n896,n897);
xor (n896,n893,n894);
or (n897,n898,n901);
and (n898,n899,n900);
and (n899,n25,n219);
and (n900,n19,n65);
and (n901,n902,n903);
xor (n902,n899,n900);
or (n903,n904,n906);
and (n904,n905,n665);
and (n905,n19,n219);
and (n906,n907,n908);
xor (n907,n905,n665);
or (n908,n909,n912);
and (n909,n910,n911);
and (n910,n18,n219);
and (n911,n85,n65);
and (n912,n913,n914);
xor (n913,n910,n911);
or (n914,n915,n918);
and (n915,n916,n917);
and (n916,n85,n219);
and (n917,n84,n65);
and (n918,n919,n920);
xor (n919,n916,n917);
and (n920,n717,n921);
and (n921,n185,n65);
and (n922,n923,n924);
xor (n923,n861,n179);
or (n924,n925,n928);
and (n925,n926,n927);
xor (n926,n64,n862);
and (n927,n48,n55);
and (n928,n929,n930);
xor (n929,n926,n927);
or (n930,n931,n934);
and (n931,n932,n933);
xor (n932,n866,n867);
and (n933,n47,n55);
and (n934,n935,n936);
xor (n935,n932,n933);
or (n936,n937,n940);
and (n937,n938,n939);
xor (n938,n872,n873);
and (n939,n130,n55);
and (n940,n941,n942);
xor (n941,n938,n939);
or (n942,n943,n946);
and (n943,n944,n945);
xor (n944,n878,n879);
and (n945,n105,n55);
and (n946,n947,n948);
xor (n947,n944,n945);
or (n948,n949,n952);
and (n949,n950,n951);
xor (n950,n884,n885);
and (n951,n103,n55);
and (n952,n953,n954);
xor (n953,n950,n951);
or (n954,n955,n958);
and (n955,n956,n957);
xor (n956,n890,n891);
and (n957,n25,n55);
and (n958,n959,n960);
xor (n959,n956,n957);
or (n960,n961,n964);
and (n961,n962,n963);
xor (n962,n896,n897);
and (n963,n19,n55);
and (n964,n965,n966);
xor (n965,n962,n963);
or (n966,n967,n970);
and (n967,n968,n969);
xor (n968,n902,n903);
and (n969,n18,n55);
and (n970,n971,n972);
xor (n971,n968,n969);
or (n972,n973,n976);
and (n973,n974,n975);
xor (n974,n907,n908);
and (n975,n85,n55);
and (n976,n977,n978);
xor (n977,n974,n975);
or (n978,n979,n981);
and (n979,n980,n686);
xor (n980,n913,n914);
and (n981,n982,n983);
xor (n982,n980,n686);
and (n983,n984,n985);
xor (n984,n919,n920);
and (n985,n185,n55);
and (n986,n987,n988);
xor (n987,n859,n801);
or (n988,n989,n992);
and (n989,n990,n991);
xor (n990,n923,n924);
and (n991,n48,n42);
and (n992,n993,n994);
xor (n993,n990,n991);
or (n994,n995,n997);
and (n995,n996,n242);
xor (n996,n929,n930);
and (n997,n998,n999);
xor (n998,n996,n242);
or (n999,n1000,n1003);
and (n1000,n1001,n1002);
xor (n1001,n935,n936);
and (n1002,n130,n42);
and (n1003,n1004,n1005);
xor (n1004,n1001,n1002);
or (n1005,n1006,n1009);
and (n1006,n1007,n1008);
xor (n1007,n941,n942);
and (n1008,n105,n42);
and (n1009,n1010,n1011);
xor (n1010,n1007,n1008);
or (n1011,n1012,n1015);
and (n1012,n1013,n1014);
xor (n1013,n947,n948);
and (n1014,n103,n42);
and (n1015,n1016,n1017);
xor (n1016,n1013,n1014);
or (n1017,n1018,n1021);
and (n1018,n1019,n1020);
xor (n1019,n953,n954);
and (n1020,n25,n42);
and (n1021,n1022,n1023);
xor (n1022,n1019,n1020);
or (n1023,n1024,n1027);
and (n1024,n1025,n1026);
xor (n1025,n959,n960);
and (n1026,n19,n42);
and (n1027,n1028,n1029);
xor (n1028,n1025,n1026);
or (n1029,n1030,n1032);
and (n1030,n1031,n587);
xor (n1031,n965,n966);
and (n1032,n1033,n1034);
xor (n1033,n1031,n587);
or (n1034,n1035,n1038);
and (n1035,n1036,n1037);
xor (n1036,n971,n972);
and (n1037,n85,n42);
and (n1038,n1039,n1040);
xor (n1039,n1036,n1037);
or (n1040,n1041,n1043);
and (n1041,n1042,n672);
xor (n1042,n977,n978);
and (n1043,n1044,n1045);
xor (n1044,n1042,n672);
and (n1045,n1046,n1047);
xor (n1046,n982,n983);
and (n1047,n185,n42);
and (n1048,n43,n137);
or (n1049,n1050,n1053);
and (n1050,n1051,n1052);
xor (n1051,n987,n988);
and (n1052,n48,n137);
and (n1053,n1054,n1055);
xor (n1054,n1051,n1052);
or (n1055,n1056,n1059);
and (n1056,n1057,n1058);
xor (n1057,n993,n994);
and (n1058,n47,n137);
and (n1059,n1060,n1061);
xor (n1060,n1057,n1058);
or (n1061,n1062,n1065);
and (n1062,n1063,n1064);
xor (n1063,n998,n999);
and (n1064,n130,n137);
and (n1065,n1066,n1067);
xor (n1066,n1063,n1064);
or (n1067,n1068,n1071);
and (n1068,n1069,n1070);
xor (n1069,n1004,n1005);
and (n1070,n105,n137);
and (n1071,n1072,n1073);
xor (n1072,n1069,n1070);
or (n1073,n1074,n1077);
and (n1074,n1075,n1076);
xor (n1075,n1010,n1011);
and (n1076,n103,n137);
and (n1077,n1078,n1079);
xor (n1078,n1075,n1076);
or (n1079,n1080,n1083);
and (n1080,n1081,n1082);
xor (n1081,n1016,n1017);
and (n1082,n25,n137);
and (n1083,n1084,n1085);
xor (n1084,n1081,n1082);
or (n1085,n1086,n1089);
and (n1086,n1087,n1088);
xor (n1087,n1022,n1023);
and (n1088,n19,n137);
and (n1089,n1090,n1091);
xor (n1090,n1087,n1088);
or (n1091,n1092,n1095);
and (n1092,n1093,n1094);
xor (n1093,n1028,n1029);
and (n1094,n18,n137);
and (n1095,n1096,n1097);
xor (n1096,n1093,n1094);
or (n1097,n1098,n1101);
and (n1098,n1099,n1100);
xor (n1099,n1033,n1034);
and (n1100,n85,n137);
and (n1101,n1102,n1103);
xor (n1102,n1099,n1100);
or (n1103,n1104,n1106);
and (n1104,n1105,n615);
xor (n1105,n1039,n1040);
and (n1106,n1107,n1108);
xor (n1107,n1105,n615);
and (n1108,n1109,n1110);
xor (n1109,n1044,n1045);
and (n1110,n185,n137);
and (n1111,n48,n143);
or (n1112,n1113,n1116);
and (n1113,n1114,n1115);
xor (n1114,n1054,n1055);
and (n1115,n47,n143);
and (n1116,n1117,n1118);
xor (n1117,n1114,n1115);
or (n1118,n1119,n1122);
and (n1119,n1120,n1121);
xor (n1120,n1060,n1061);
and (n1121,n130,n143);
and (n1122,n1123,n1124);
xor (n1123,n1120,n1121);
or (n1124,n1125,n1128);
and (n1125,n1126,n1127);
xor (n1126,n1066,n1067);
and (n1127,n105,n143);
and (n1128,n1129,n1130);
xor (n1129,n1126,n1127);
or (n1130,n1131,n1134);
and (n1131,n1132,n1133);
xor (n1132,n1072,n1073);
and (n1133,n103,n143);
and (n1134,n1135,n1136);
xor (n1135,n1132,n1133);
or (n1136,n1137,n1140);
and (n1137,n1138,n1139);
xor (n1138,n1078,n1079);
and (n1139,n25,n143);
and (n1140,n1141,n1142);
xor (n1141,n1138,n1139);
or (n1142,n1143,n1146);
and (n1143,n1144,n1145);
xor (n1144,n1084,n1085);
and (n1145,n19,n143);
and (n1146,n1147,n1148);
xor (n1147,n1144,n1145);
or (n1148,n1149,n1152);
and (n1149,n1150,n1151);
xor (n1150,n1090,n1091);
and (n1151,n18,n143);
and (n1152,n1153,n1154);
xor (n1153,n1150,n1151);
or (n1154,n1155,n1158);
and (n1155,n1156,n1157);
xor (n1156,n1096,n1097);
and (n1157,n85,n143);
and (n1158,n1159,n1160);
xor (n1159,n1156,n1157);
or (n1160,n1161,n1164);
and (n1161,n1162,n1163);
xor (n1162,n1102,n1103);
and (n1163,n84,n143);
and (n1164,n1165,n1166);
xor (n1165,n1162,n1163);
and (n1166,n1167,n1168);
xor (n1167,n1107,n1108);
and (n1168,n185,n143);
and (n1169,n47,n113);
or (n1170,n1171,n1174);
and (n1171,n1172,n1173);
xor (n1172,n1117,n1118);
and (n1173,n130,n113);
and (n1174,n1175,n1176);
xor (n1175,n1172,n1173);
or (n1176,n1177,n1180);
and (n1177,n1178,n1179);
xor (n1178,n1123,n1124);
and (n1179,n105,n113);
and (n1180,n1181,n1182);
xor (n1181,n1178,n1179);
or (n1182,n1183,n1186);
and (n1183,n1184,n1185);
xor (n1184,n1129,n1130);
and (n1185,n103,n113);
and (n1186,n1187,n1188);
xor (n1187,n1184,n1185);
or (n1188,n1189,n1192);
and (n1189,n1190,n1191);
xor (n1190,n1135,n1136);
and (n1191,n25,n113);
and (n1192,n1193,n1194);
xor (n1193,n1190,n1191);
or (n1194,n1195,n1198);
and (n1195,n1196,n1197);
xor (n1196,n1141,n1142);
and (n1197,n19,n113);
and (n1198,n1199,n1200);
xor (n1199,n1196,n1197);
or (n1200,n1201,n1204);
and (n1201,n1202,n1203);
xor (n1202,n1147,n1148);
and (n1203,n18,n113);
and (n1204,n1205,n1206);
xor (n1205,n1202,n1203);
or (n1206,n1207,n1210);
and (n1207,n1208,n1209);
xor (n1208,n1153,n1154);
and (n1209,n85,n113);
and (n1210,n1211,n1212);
xor (n1211,n1208,n1209);
or (n1212,n1213,n1215);
and (n1213,n1214,n533);
xor (n1214,n1159,n1160);
and (n1215,n1216,n1217);
xor (n1216,n1214,n533);
and (n1217,n1218,n1219);
xor (n1218,n1165,n1166);
and (n1219,n185,n113);
and (n1220,n130,n121);
or (n1221,n1222,n1224);
and (n1222,n1223,n122);
xor (n1223,n1175,n1176);
and (n1224,n1225,n1226);
xor (n1225,n1223,n122);
or (n1226,n1227,n1230);
and (n1227,n1228,n1229);
xor (n1228,n1181,n1182);
and (n1229,n103,n121);
and (n1230,n1231,n1232);
xor (n1231,n1228,n1229);
or (n1232,n1233,n1236);
and (n1233,n1234,n1235);
xor (n1234,n1187,n1188);
and (n1235,n25,n121);
and (n1236,n1237,n1238);
xor (n1237,n1234,n1235);
or (n1238,n1239,n1242);
and (n1239,n1240,n1241);
xor (n1240,n1193,n1194);
and (n1241,n19,n121);
and (n1242,n1243,n1244);
xor (n1243,n1240,n1241);
or (n1244,n1245,n1248);
and (n1245,n1246,n1247);
xor (n1246,n1199,n1200);
and (n1247,n18,n121);
and (n1248,n1249,n1250);
xor (n1249,n1246,n1247);
or (n1250,n1251,n1254);
and (n1251,n1252,n1253);
xor (n1252,n1205,n1206);
and (n1253,n85,n121);
and (n1254,n1255,n1256);
xor (n1255,n1252,n1253);
or (n1256,n1257,n1260);
and (n1257,n1258,n1259);
xor (n1258,n1211,n1212);
and (n1259,n84,n121);
and (n1260,n1261,n1262);
xor (n1261,n1258,n1259);
and (n1262,n1263,n1264);
xor (n1263,n1216,n1217);
and (n1264,n185,n121);
or (n1265,n1266,n1269);
and (n1266,n1267,n1268);
xor (n1267,n1225,n1226);
and (n1268,n103,n29);
and (n1269,n1270,n1271);
xor (n1270,n1267,n1268);
or (n1271,n1272,n1275);
and (n1272,n1273,n1274);
xor (n1273,n1231,n1232);
and (n1274,n25,n29);
and (n1275,n1276,n1277);
xor (n1276,n1273,n1274);
or (n1277,n1278,n1281);
and (n1278,n1279,n1280);
xor (n1279,n1237,n1238);
and (n1280,n19,n29);
and (n1281,n1282,n1283);
xor (n1282,n1279,n1280);
or (n1283,n1284,n1287);
and (n1284,n1285,n1286);
xor (n1285,n1243,n1244);
and (n1286,n18,n29);
and (n1287,n1288,n1289);
xor (n1288,n1285,n1286);
or (n1289,n1290,n1293);
and (n1290,n1291,n1292);
xor (n1291,n1249,n1250);
and (n1292,n85,n29);
and (n1293,n1294,n1295);
xor (n1294,n1291,n1292);
or (n1295,n1296,n1298);
and (n1296,n1297,n440);
xor (n1297,n1255,n1256);
and (n1298,n1299,n1300);
xor (n1299,n1297,n440);
and (n1300,n1301,n1302);
xor (n1301,n1261,n1262);
and (n1302,n185,n29);
and (n1303,n103,n35);
or (n1304,n1305,n1308);
and (n1305,n1306,n1307);
xor (n1306,n1270,n1271);
and (n1307,n25,n35);
and (n1308,n1309,n1310);
xor (n1309,n1306,n1307);
or (n1310,n1311,n1314);
and (n1311,n1312,n1313);
xor (n1312,n1276,n1277);
and (n1313,n19,n35);
and (n1314,n1315,n1316);
xor (n1315,n1312,n1313);
or (n1316,n1317,n1320);
and (n1317,n1318,n1319);
xor (n1318,n1282,n1283);
and (n1319,n18,n35);
and (n1320,n1321,n1322);
xor (n1321,n1318,n1319);
or (n1322,n1323,n1326);
and (n1323,n1324,n1325);
xor (n1324,n1288,n1289);
and (n1325,n85,n35);
and (n1326,n1327,n1328);
xor (n1327,n1324,n1325);
or (n1328,n1329,n1332);
and (n1329,n1330,n1331);
xor (n1330,n1294,n1295);
and (n1331,n84,n35);
and (n1332,n1333,n1334);
xor (n1333,n1330,n1331);
and (n1334,n1335,n1336);
xor (n1335,n1299,n1300);
and (n1336,n185,n35);
and (n1337,n25,n77);
or (n1338,n1339,n1342);
and (n1339,n1340,n1341);
xor (n1340,n1309,n1310);
and (n1341,n19,n77);
and (n1342,n1343,n1344);
xor (n1343,n1340,n1341);
or (n1344,n1345,n1348);
and (n1345,n1346,n1347);
xor (n1346,n1315,n1316);
and (n1347,n18,n77);
and (n1348,n1349,n1350);
xor (n1349,n1346,n1347);
or (n1350,n1351,n1354);
and (n1351,n1352,n1353);
xor (n1352,n1321,n1322);
and (n1353,n85,n77);
and (n1354,n1355,n1356);
xor (n1355,n1352,n1353);
or (n1356,n1357,n1360);
and (n1357,n1358,n1359);
xor (n1358,n1327,n1328);
and (n1359,n84,n77);
and (n1360,n1361,n1362);
xor (n1361,n1358,n1359);
and (n1362,n1363,n1364);
xor (n1363,n1333,n1334);
and (n1364,n185,n77);
and (n1365,n19,n95);
or (n1366,n1367,n1370);
and (n1367,n1368,n1369);
xor (n1368,n1343,n1344);
and (n1369,n18,n95);
and (n1370,n1371,n1372);
xor (n1371,n1368,n1369);
or (n1372,n1373,n1376);
and (n1373,n1374,n1375);
xor (n1374,n1349,n1350);
and (n1375,n85,n95);
and (n1376,n1377,n1378);
xor (n1377,n1374,n1375);
or (n1378,n1379,n1382);
and (n1379,n1380,n1381);
xor (n1380,n1355,n1356);
and (n1381,n84,n95);
and (n1382,n1383,n1384);
xor (n1383,n1380,n1381);
and (n1384,n1385,n1386);
xor (n1385,n1361,n1362);
and (n1386,n185,n95);
and (n1387,n18,n203);
or (n1388,n1389,n1392);
and (n1389,n1390,n1391);
xor (n1390,n1371,n1372);
and (n1391,n85,n203);
and (n1392,n1393,n1394);
xor (n1393,n1390,n1391);
or (n1394,n1395,n1398);
and (n1395,n1396,n1397);
xor (n1396,n1377,n1378);
and (n1397,n84,n203);
and (n1398,n1399,n1400);
xor (n1399,n1396,n1397);
and (n1400,n1401,n1402);
xor (n1401,n1383,n1384);
and (n1402,n185,n203);
and (n1403,n85,n188);
or (n1404,n1405,n1408);
and (n1405,n1406,n1407);
xor (n1406,n1393,n1394);
and (n1407,n84,n188);
and (n1408,n1409,n1410);
xor (n1409,n1406,n1407);
and (n1410,n1411,n1412);
xor (n1411,n1399,n1400);
and (n1412,n185,n188);
and (n1413,n84,n194);
and (n1414,n1415,n1416);
xor (n1415,n1409,n1410);
and (n1416,n185,n194);
and (n1417,n185,n808);
endmodule
