module top (out,n18,n28,n30,n31,n33,n38,n41,n43,n48
        ,n52,n60,n64,n65,n66,n78,n82,n83,n84,n99
        ,n100,n101,n102,n103,n107,n108,n109,n114,n116,n118
        ,n155,n157,n158,n159,n170,n171,n172,n173,n185,n186
        ,n187,n188,n202,n208,n210,n211,n215,n216,n219,n221
        ,n222,n223,n296,n351,n354,n356,n444,n446,n447,n562
        ,n563,n564,n565,n572,n574,n578,n589,n592,n594,n595
        ,n597,n601,n607,n610,n612,n614,n618,n621,n623,n625
        ,n629,n632,n634,n636,n638,n644,n647,n649,n651,n655
        ,n658,n660,n662,n666,n669,n671,n673,n677,n680,n682
        ,n684,n691,n694,n696,n698,n702,n705,n707,n709,n713
        ,n716,n718,n720,n724,n727,n729,n731,n740,n744,n746
        ,n748,n770,n774,n776,n778,n788,n792,n794,n796,n806
        ,n810,n812,n814,n826,n828,n830,n832,n845,n847,n849
        ,n851,n860,n864,n866,n868,n939,n942,n944,n946,n950
        ,n953,n955,n957,n961,n964,n966,n968,n972,n975,n977
        ,n979,n991,n993,n995,n997,n1009,n1011,n1013,n1015,n1027
        ,n1029,n1031,n1033,n1045,n1047,n1049,n1051,n1063,n1065,n1067
        ,n1069,n1079,n1083,n1085,n1087,n1099,n1101,n1103,n1105,n1116
        ,n1118,n1120,n1122,n1188,n1192,n1194,n1196,n1205,n1209,n1211
        ,n1213,n1229,n1233,n1235,n1237,n1247,n1251,n1253,n1255,n1265
        ,n1269,n1271,n1273,n1283,n1287,n1289,n1291,n1301,n1305,n1307
        ,n1309,n1320,n1322,n1324,n1326,n1401,n1404,n1406,n1408,n1412
        ,n1415,n1417,n1419,n1423,n1426,n1428,n1430,n1434,n1437,n1439
        ,n1441,n1449,n1452,n1454,n1456,n1460,n1463,n1465,n1467,n1471
        ,n1474,n1476,n1478,n1482,n1485,n1487,n1489,n1502,n1506,n1508
        ,n1510,n1520,n1524,n1526,n1528,n1540,n1542,n1544,n1546,n1558
        ,n1560,n1562,n1564,n1574,n1578,n1580,n1582,n1594,n1596,n1598
        ,n1600,n1610,n1614,n1616,n1618,n1627,n1631,n1633,n1635);
output out;
input n18;
input n28;
input n30;
input n31;
input n33;
input n38;
input n41;
input n43;
input n48;
input n52;
input n60;
input n64;
input n65;
input n66;
input n78;
input n82;
input n83;
input n84;
input n99;
input n100;
input n101;
input n102;
input n103;
input n107;
input n108;
input n109;
input n114;
input n116;
input n118;
input n155;
input n157;
input n158;
input n159;
input n170;
input n171;
input n172;
input n173;
input n185;
input n186;
input n187;
input n188;
input n202;
input n208;
input n210;
input n211;
input n215;
input n216;
input n219;
input n221;
input n222;
input n223;
input n296;
input n351;
input n354;
input n356;
input n444;
input n446;
input n447;
input n562;
input n563;
input n564;
input n565;
input n572;
input n574;
input n578;
input n589;
input n592;
input n594;
input n595;
input n597;
input n601;
input n607;
input n610;
input n612;
input n614;
input n618;
input n621;
input n623;
input n625;
input n629;
input n632;
input n634;
input n636;
input n638;
input n644;
input n647;
input n649;
input n651;
input n655;
input n658;
input n660;
input n662;
input n666;
input n669;
input n671;
input n673;
input n677;
input n680;
input n682;
input n684;
input n691;
input n694;
input n696;
input n698;
input n702;
input n705;
input n707;
input n709;
input n713;
input n716;
input n718;
input n720;
input n724;
input n727;
input n729;
input n731;
input n740;
input n744;
input n746;
input n748;
input n770;
input n774;
input n776;
input n778;
input n788;
input n792;
input n794;
input n796;
input n806;
input n810;
input n812;
input n814;
input n826;
input n828;
input n830;
input n832;
input n845;
input n847;
input n849;
input n851;
input n860;
input n864;
input n866;
input n868;
input n939;
input n942;
input n944;
input n946;
input n950;
input n953;
input n955;
input n957;
input n961;
input n964;
input n966;
input n968;
input n972;
input n975;
input n977;
input n979;
input n991;
input n993;
input n995;
input n997;
input n1009;
input n1011;
input n1013;
input n1015;
input n1027;
input n1029;
input n1031;
input n1033;
input n1045;
input n1047;
input n1049;
input n1051;
input n1063;
input n1065;
input n1067;
input n1069;
input n1079;
input n1083;
input n1085;
input n1087;
input n1099;
input n1101;
input n1103;
input n1105;
input n1116;
input n1118;
input n1120;
input n1122;
input n1188;
input n1192;
input n1194;
input n1196;
input n1205;
input n1209;
input n1211;
input n1213;
input n1229;
input n1233;
input n1235;
input n1237;
input n1247;
input n1251;
input n1253;
input n1255;
input n1265;
input n1269;
input n1271;
input n1273;
input n1283;
input n1287;
input n1289;
input n1291;
input n1301;
input n1305;
input n1307;
input n1309;
input n1320;
input n1322;
input n1324;
input n1326;
input n1401;
input n1404;
input n1406;
input n1408;
input n1412;
input n1415;
input n1417;
input n1419;
input n1423;
input n1426;
input n1428;
input n1430;
input n1434;
input n1437;
input n1439;
input n1441;
input n1449;
input n1452;
input n1454;
input n1456;
input n1460;
input n1463;
input n1465;
input n1467;
input n1471;
input n1474;
input n1476;
input n1478;
input n1482;
input n1485;
input n1487;
input n1489;
input n1502;
input n1506;
input n1508;
input n1510;
input n1520;
input n1524;
input n1526;
input n1528;
input n1540;
input n1542;
input n1544;
input n1546;
input n1558;
input n1560;
input n1562;
input n1564;
input n1574;
input n1578;
input n1580;
input n1582;
input n1594;
input n1596;
input n1598;
input n1600;
input n1610;
input n1614;
input n1616;
input n1618;
input n1627;
input n1631;
input n1633;
input n1635;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n24;
wire n25;
wire n26;
wire n27;
wire n29;
wire n32;
wire n34;
wire n35;
wire n36;
wire n37;
wire n39;
wire n40;
wire n42;
wire n44;
wire n45;
wire n46;
wire n47;
wire n49;
wire n50;
wire n51;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n61;
wire n62;
wire n63;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n79;
wire n80;
wire n81;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n104;
wire n105;
wire n106;
wire n110;
wire n111;
wire n112;
wire n113;
wire n115;
wire n117;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n156;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n209;
wire n212;
wire n213;
wire n214;
wire n217;
wire n218;
wire n220;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n352;
wire n353;
wire n355;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n445;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n573;
wire n575;
wire n576;
wire n577;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n590;
wire n591;
wire n593;
wire n596;
wire n598;
wire n599;
wire n600;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n608;
wire n609;
wire n611;
wire n613;
wire n615;
wire n616;
wire n617;
wire n619;
wire n620;
wire n622;
wire n624;
wire n626;
wire n627;
wire n628;
wire n630;
wire n631;
wire n633;
wire n635;
wire n637;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n645;
wire n646;
wire n648;
wire n650;
wire n652;
wire n653;
wire n654;
wire n656;
wire n657;
wire n659;
wire n661;
wire n663;
wire n664;
wire n665;
wire n667;
wire n668;
wire n670;
wire n672;
wire n674;
wire n675;
wire n676;
wire n678;
wire n679;
wire n681;
wire n683;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n692;
wire n693;
wire n695;
wire n697;
wire n699;
wire n700;
wire n701;
wire n703;
wire n704;
wire n706;
wire n708;
wire n710;
wire n711;
wire n712;
wire n714;
wire n715;
wire n717;
wire n719;
wire n721;
wire n722;
wire n723;
wire n725;
wire n726;
wire n728;
wire n730;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n741;
wire n742;
wire n743;
wire n745;
wire n747;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n771;
wire n772;
wire n773;
wire n775;
wire n777;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n789;
wire n790;
wire n791;
wire n793;
wire n795;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n807;
wire n808;
wire n809;
wire n811;
wire n813;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n827;
wire n829;
wire n831;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n846;
wire n848;
wire n850;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n861;
wire n862;
wire n863;
wire n865;
wire n867;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n940;
wire n941;
wire n943;
wire n945;
wire n947;
wire n948;
wire n949;
wire n951;
wire n952;
wire n954;
wire n956;
wire n958;
wire n959;
wire n960;
wire n962;
wire n963;
wire n965;
wire n967;
wire n969;
wire n970;
wire n971;
wire n973;
wire n974;
wire n976;
wire n978;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n992;
wire n994;
wire n996;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1010;
wire n1012;
wire n1014;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1028;
wire n1030;
wire n1032;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1046;
wire n1048;
wire n1050;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1064;
wire n1066;
wire n1068;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1080;
wire n1081;
wire n1082;
wire n1084;
wire n1086;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1100;
wire n1102;
wire n1104;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1117;
wire n1119;
wire n1121;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1189;
wire n1190;
wire n1191;
wire n1193;
wire n1195;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1206;
wire n1207;
wire n1208;
wire n1210;
wire n1212;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1230;
wire n1231;
wire n1232;
wire n1234;
wire n1236;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1248;
wire n1249;
wire n1250;
wire n1252;
wire n1254;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1266;
wire n1267;
wire n1268;
wire n1270;
wire n1272;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1284;
wire n1285;
wire n1286;
wire n1288;
wire n1290;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1302;
wire n1303;
wire n1304;
wire n1306;
wire n1308;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1321;
wire n1323;
wire n1325;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1402;
wire n1403;
wire n1405;
wire n1407;
wire n1409;
wire n1410;
wire n1411;
wire n1413;
wire n1414;
wire n1416;
wire n1418;
wire n1420;
wire n1421;
wire n1422;
wire n1424;
wire n1425;
wire n1427;
wire n1429;
wire n1431;
wire n1432;
wire n1433;
wire n1435;
wire n1436;
wire n1438;
wire n1440;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1450;
wire n1451;
wire n1453;
wire n1455;
wire n1457;
wire n1458;
wire n1459;
wire n1461;
wire n1462;
wire n1464;
wire n1466;
wire n1468;
wire n1469;
wire n1470;
wire n1472;
wire n1473;
wire n1475;
wire n1477;
wire n1479;
wire n1480;
wire n1481;
wire n1483;
wire n1484;
wire n1486;
wire n1488;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1503;
wire n1504;
wire n1505;
wire n1507;
wire n1509;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1521;
wire n1522;
wire n1523;
wire n1525;
wire n1527;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1541;
wire n1543;
wire n1545;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1559;
wire n1561;
wire n1563;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1575;
wire n1576;
wire n1577;
wire n1579;
wire n1581;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1595;
wire n1597;
wire n1599;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1611;
wire n1612;
wire n1613;
wire n1615;
wire n1617;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1628;
wire n1629;
wire n1630;
wire n1632;
wire n1634;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
xor (out,n0,n2252);
nor (n0,n1,n2096);
not (n1,n2);
nor (n2,n3,n1946);
not (n3,n4);
nor (n4,n5,n1769);
not (n5,n6);
nor (n6,n7,n1706);
not (n7,n8);
nor (n8,n9,n1491);
and (n9,n10,n1182);
xor (n10,n11,n981);
wire s0n11,s1n11,notn11;
or (n11,s0n11,s1n11);
not(notn11,n934);
and (s0n11,notn11,1'b0);
and (s1n11,n934,n13);
xor (n13,n14,n733);
wire s0n14,s1n14,notn14;
or (n14,s0n14,s1n14);
not(notn14,n583);
and (s0n14,notn14,1'b0);
and (s1n14,n583,n15);
nand (n15,n16,n568);
or (n16,n17,n19);
not (n17,n18);
not (n19,n20);
and (n20,n21,n566);
nor (n21,n22,n559);
not (n22,n23);
nor (n23,n24,n57);
nor (n24,n25,n44);
and (n25,n26,n43);
or (n26,n27,n32,n37,n40);
and (n27,n28,n29);
and (n29,n30,n31);
and (n32,n33,n34);
not (n34,n35);
nand (n35,n36,n31);
not (n36,n30);
and (n37,n38,n39);
nor (n39,n36,n31);
and (n40,n41,n42);
nor (n42,n30,n31);
nor (n44,n45,n53,n43);
and (n45,n46,n51);
nand (n46,n47,n49);
or (n47,n48,n41);
or (n49,n50,n33);
not (n50,n48);
not (n51,n52);
and (n53,n54,n52);
nand (n54,n55,n56);
or (n55,n48,n38);
or (n56,n50,n28);
nand (n57,n58,n67);
or (n58,n59,n61);
not (n59,n60);
not (n61,n62);
nand (n62,n63,n66);
nor (n63,n64,n65);
nand (n67,n68,n523);
nand (n68,n69,n515);
or (n69,n70,n439);
not (n70,n71);
or (n71,1'b0,n72,n359,n437);
and (n72,n73,n358);
wire s0n73,s1n73,notn73;
or (n73,s0n73,s1n73);
not(notn73,n349);
and (s0n73,notn73,n74);
and (s1n73,n349,1'b0);
wire s0n74,s1n74,notn74;
or (n74,s0n74,s1n74);
not(notn74,n285);
and (s0n74,notn74,1'b0);
and (s1n74,n285,n75);
or (n75,n76,n259,n265,n271,n276,1'b0,1'b0,1'b0);
and (n76,n77,n85);
xnor (n77,n78,n79);
not (n79,n80);
nor (n80,n81,n84);
or (n81,n82,n83);
and (n85,n86,n228,n247,n255);
wire s0n86,s1n86,notn86;
or (n86,s0n86,s1n86);
not(notn86,n119);
and (s0n86,notn86,n87);
and (s1n86,n119,1'b0);
wire s0n87,s1n87,notn87;
or (n87,s0n87,s1n87);
not(notn87,n117);
and (s0n87,notn87,n88);
and (s1n87,n117,n115);
wire s0n88,s1n88,notn88;
or (n88,s0n88,s1n88);
not(notn88,n110);
and (s0n88,notn88,n89);
and (s1n88,n110,n104);
wire s0n89,s1n89,notn89;
or (n89,s0n89,s1n89);
not(notn89,n103);
and (s0n89,notn89,n90);
and (s1n89,n103,1'b0);
wire s0n90,s1n90,notn90;
or (n90,s0n90,s1n90);
not(notn90,n102);
and (s0n90,notn90,n91);
and (s1n90,n102,1'b1);
wire s0n91,s1n91,notn91;
or (n91,s0n91,s1n91);
not(notn91,n101);
and (s0n91,notn91,n92);
and (s1n91,n101,1'b0);
wire s0n92,s1n92,notn92;
or (n92,s0n92,s1n92);
not(notn92,n100);
and (s0n92,notn92,n93);
and (s1n92,n100,1'b1);
wire s0n93,s1n93,notn93;
or (n93,s0n93,s1n93);
not(notn93,n99);
and (s0n93,notn93,n94);
and (s1n93,n99,1'b0);
wire s0n94,s1n94,notn94;
or (n94,s0n94,s1n94);
not(notn94,n78);
and (s0n94,notn94,n95);
and (s1n94,n78,1'b1);
wire s0n95,s1n95,notn95;
or (n95,s0n95,s1n95);
not(notn95,n84);
and (s0n95,notn95,n96);
and (s1n95,n84,1'b0);
wire s0n96,s1n96,notn96;
or (n96,s0n96,s1n96);
not(notn96,n82);
and (s0n96,notn96,n97);
and (s1n96,n82,1'b1);
not (n97,n83);
wire s0n104,s1n104,notn104;
or (n104,s0n104,s1n104);
not(notn104,n109);
and (s0n104,notn104,n105);
and (s1n104,n109,1'b0);
wire s0n105,s1n105,notn105;
or (n105,s0n105,s1n105);
not(notn105,n108);
and (s0n105,notn105,n106);
and (s1n105,n108,1'b1);
not (n106,n107);
or (n110,n111,n114);
or (n111,n109,n112);
not (n112,n113);
nor (n113,n108,n107);
not (n115,n116);
or (n117,n116,n118);
not (n119,n120);
or (n120,n121,n226);
or (n121,n122,n224);
or (n122,n123,n218);
or (n123,n124,n217);
or (n124,n125,n213);
or (n125,n126,n212);
or (n126,n127,n207);
or (n127,n128,n206);
or (n128,n129,n205);
or (n129,n130,n203);
or (n130,n131,n200);
or (n131,n132,n199);
or (n132,n133,n198);
or (n133,n134,n197);
or (n134,n135,n196);
or (n135,n136,n194);
or (n136,n137,n192);
or (n137,n138,n191);
or (n138,n139,n189);
or (n139,n140,n183);
or (n140,n141,n182);
or (n141,n142,n181);
or (n142,n143,n180);
or (n143,n144,n179);
or (n144,n145,n178);
or (n145,n146,n176);
or (n146,n147,n174);
or (n147,n148,n168);
or (n148,n149,n167);
or (n149,n150,n166);
or (n150,n151,n165);
or (n151,n152,n164);
or (n152,n153,n162);
or (n153,n154,n160);
nor (n154,n155,n156,n158,n159);
not (n156,n157);
nor (n160,n155,n156,n161,n159);
not (n161,n158);
and (n162,n155,n157,n158,n163);
not (n163,n159);
and (n164,n155,n156,n158,n163);
nor (n165,n155,n157,n161,n159);
and (n166,n155,n156,n158,n159);
and (n167,n155,n157,n158,n159);
nor (n168,n169,n171,n172,n173);
not (n169,n170);
nor (n174,n169,n175,n172,n173);
not (n175,n171);
and (n176,n169,n171,n172,n177);
not (n177,n173);
and (n178,n170,n171,n172,n177);
and (n179,n170,n175,n172,n177);
and (n180,n169,n175,n172,n173);
and (n181,n170,n175,n172,n173);
and (n182,n170,n171,n172,n173);
nor (n183,n184,n186,n187,n188);
not (n184,n185);
nor (n189,n184,n190,n187,n188);
not (n190,n186);
nor (n191,n185,n190,n187,n188);
nor (n192,n184,n190,n193,n188);
not (n193,n187);
nor (n194,n185,n186,n193,n195);
not (n195,n188);
and (n196,n184,n186,n187,n188);
and (n197,n184,n186,n193,n188);
and (n198,n185,n186,n193,n188);
and (n199,n185,n190,n193,n188);
nor (n200,n201,n66,n64,n65);
not (n201,n202);
nor (n203,n202,n204,n64,n65);
not (n204,n66);
and (n205,n201,n204,n64,n65);
and (n206,n202,n204,n64,n65);
nor (n207,n208,n209,n211);
not (n209,n210);
and (n212,n208,n210,n211);
nor (n213,n214,n216);
not (n214,n215);
and (n217,n214,n216);
nor (n218,n219,n220,n222,n223);
not (n220,n221);
and (n224,n219,n221,n222,n225);
not (n225,n223);
and (n226,n227,n220,n222,n225);
not (n227,n219);
not (n228,n229);
or (n229,n119,n230);
nand (n230,n231,n246);
or (n231,n232,n245);
nor (n232,n233,n243);
nor (n233,n234,n240);
and (n234,n235,n239);
nand (n235,n236,n237);
or (n236,n82,n84);
wire s0n237,s1n237,notn237;
or (n237,s0n237,s1n237);
not(notn237,n99);
and (s0n237,notn237,n238);
and (s1n237,n99,1'b0);
not (n238,n78);
nor (n239,n100,n101);
not (n240,n241);
wire s0n241,s1n241,notn241;
or (n241,s0n241,s1n241);
not(notn241,n103);
and (s0n241,notn241,n242);
and (s1n241,n103,1'b0);
not (n242,n102);
nand (n243,n244,n106);
not (n244,n114);
or (n245,n109,n108);
not (n246,n117);
wire s0n247,s1n247,notn247;
or (n247,s0n247,s1n247);
not(notn247,n119);
and (s0n247,notn247,n248);
and (s1n247,n119,1'b0);
wire s0n248,s1n248,notn248;
or (n248,s0n248,s1n248);
not(notn248,n117);
and (s0n248,notn248,n249);
and (s1n248,n117,1'b0);
wire s0n249,s1n249,notn249;
or (n249,s0n249,s1n249);
not(notn249,n110);
and (s0n249,notn249,n250);
and (s1n249,n110,n254);
wire s0n250,s1n250,notn250;
or (n250,s0n250,s1n250);
not(notn250,n103);
and (s0n250,notn250,n251);
and (s1n250,n103,1'b1);
wire s0n251,s1n251,notn251;
or (n251,s0n251,s1n251);
not(notn251,n102);
and (s0n251,notn251,n252);
and (s1n251,n102,1'b1);
wire s0n252,s1n252,notn252;
or (n252,s0n252,s1n252);
not(notn252,n101);
and (s0n252,notn252,n253);
and (s1n252,n101,1'b0);
wire s0n253,s1n253,notn253;
or (n253,s0n253,s1n253);
not(notn253,n100);
and (s0n253,notn253,n237);
and (s1n253,n100,1'b0);
not (n254,n245);
not (n255,n256);
wire s0n256,s1n256,notn256;
or (n256,s0n256,s1n256);
not(notn256,n119);
and (s0n256,notn256,n257);
and (s1n256,n119,1'b0);
wire s0n257,s1n257,notn257;
or (n257,s0n257,s1n257);
not(notn257,n117);
and (s0n257,notn257,n258);
and (s1n257,n117,1'b0);
wire s0n258,s1n258,notn258;
or (n258,s0n258,s1n258);
not(notn258,n110);
and (s0n258,notn258,n241);
and (s1n258,n110,1'b0);
and (n259,n260,n263);
xnor (n260,n100,n261);
or (n261,n99,n262);
or (n262,n78,n84);
and (n263,n264,n228,n247,n255);
not (n264,n86);
and (n265,n266,n270);
xnor (n266,n102,n267);
not (n267,n268);
nor (n268,n269,n101);
or (n269,n100,n99);
and (n270,n86,n229,n247,n255);
and (n271,n272,n275);
xnor (n272,n114,n273);
or (n273,n103,n274);
or (n274,n102,n101);
and (n275,n264,n229,n247,n255);
and (n276,n277,n280);
not (n277,n278);
nand (n278,n279,n255,n86,n228);
not (n279,n247);
not (n280,n281);
nand (n281,n282,n108);
or (n282,n107,n283);
not (n283,n284);
nor (n284,n103,n114);
or (n285,n286,n332);
or (n286,n287,n308,n316,n322);
nand (n287,n288,n299);
or (n288,n289,n208);
nand (n289,n290,n297,n210);
nor (n290,n291,n65);
not (n291,n292);
and (n292,n293,n294,n195);
nor (n293,n187,n186);
nor (n294,n295,n185);
not (n295,n296);
nor (n297,n298,n202);
nand (n298,n204,n64);
nor (n299,n300,n302);
and (n300,n290,n301,n215);
nor (n301,n201,n298);
nand (n302,n303,n307);
or (n303,n304,n306);
nor (n304,n305,n293);
and (n305,n186,n195);
nand (n306,n185,n296);
nand (n307,n193,n294,n186);
nor (n308,n309,n314,n173);
nand (n309,n290,n310);
and (n310,n311,n313,n204);
not (n311,n312);
or (n312,n155,n157,n158,n159);
nor (n313,n64,n202);
nor (n314,n315,n170);
and (n315,n172,n171);
nor (n316,n317,n318,n319,n311);
not (n317,n313);
not (n318,n290);
nor (n319,n320,n321);
and (n320,n158,n155);
nor (n321,n155,n159);
nor (n322,n323,n330);
nor (n323,n324,n297);
and (n324,n325,n329);
not (n325,n326);
nor (n326,n327,n328);
and (n327,n313,n66);
and (n328,n202,n204);
not (n329,n65);
nand (n330,n331,n292);
or (n331,n298,n65);
wire s0n332,s1n332,notn332;
or (n332,s0n332,s1n332);
not(notn332,n295);
and (s0n332,notn332,n333);
and (s1n332,n295,1'b0);
wire s0n333,s1n333,notn333;
or (n333,s0n333,s1n333);
not(notn333,n348);
and (s0n333,notn333,n334);
and (s1n333,n348,n347);
wire s0n334,s1n334,notn334;
or (n334,s0n334,s1n334);
not(notn334,n346);
and (s0n334,notn334,n335);
and (s1n334,n346,n338);
wire s0n335,s1n335,notn335;
or (n335,s0n335,s1n335);
not(notn335,n312);
and (s0n335,notn335,n336);
and (s1n335,n312,1'b0);
or (n336,n337,n182);
or (n337,n180,n181);
or (n338,1'b0,n206,n339,n344,1'b0);
and (n339,n340,n343);
or (n340,1'b0,n212,n341,1'b0);
and (n341,n342,n210,n211);
not (n342,n208);
and (n343,n201,n204,n64,n329);
and (n344,n216,n345);
and (n345,n202,n204,n64,n329);
or (n346,n202,n66,n64,n65);
or (n347,n196,n198);
or (n348,n185,n186,n187,n188);
nor (n349,n350,n352,n355);
not (n350,n351);
not (n352,n353);
xor (n353,n354,n351);
xor (n355,n356,n357);
and (n357,n354,n351);
and (n358,n286,n332);
and (n359,n360,n435);
wire s0n360,s1n360,notn360;
or (n360,s0n360,s1n360);
not(notn360,n420);
and (s0n360,notn360,n361);
and (s1n360,n420,n416);
xor (n361,n362,n378);
not (n362,n363);
wire s0n363,s1n363,notn363;
or (n363,s0n363,s1n363);
not(notn363,n285);
and (s0n363,notn363,1'b0);
and (s1n363,n285,n364);
or (n364,n365,n368,n371,n375,1'b0,1'b0,1'b0,1'b0);
and (n365,n366,n85);
xnor (n366,n99,n367);
or (n367,n81,n262);
and (n368,n369,n263);
xnor (n369,n101,n370);
or (n370,n100,n261);
and (n371,n372,n270);
xnor (n372,n103,n373);
not (n373,n374);
and (n374,n268,n242);
and (n375,n376,n275);
xnor (n376,n107,n377);
or (n377,n114,n273);
and (n378,n379,n380);
not (n379,n74);
and (n380,n381,n398);
not (n381,n382);
wire s0n382,s1n382,notn382;
or (n382,s0n382,s1n382);
not(notn382,n285);
and (s0n382,notn382,1'b0);
and (s1n382,n285,n383);
or (n383,n384,n386,n388,n390,n392,n395,1'b0,1'b0);
and (n384,n385,n85);
xnor (n385,n84,n81);
and (n386,n387,n263);
xnor (n387,n99,n262);
and (n388,n389,n270);
xnor (n389,n101,n269);
and (n390,n391,n275);
xnor (n391,n103,n274);
nor (n392,n393,n278);
not (n393,n394);
xnor (n394,n107,n283);
and (n395,n396,n397);
xnor (n396,n109,n112);
nor (n397,n86,n229,n247,n256);
not (n398,n399);
wire s0n399,s1n399,notn399;
or (n399,s0n399,s1n399);
not(notn399,n285);
and (s0n399,notn399,1'b0);
and (s1n399,n285,n400);
or (n400,n401,n403,n405,n407,n409,n411,n413,1'b0);
and (n401,n402,n85);
xnor (n402,n82,n83);
and (n403,n404,n263);
xnor (n404,n78,n84);
and (n405,n406,n270);
xnor (n406,n100,n99);
and (n407,n408,n275);
xnor (n408,n102,n101);
and (n409,n410,n277);
xnor (n410,n114,n103);
and (n411,n412,n397);
xnor (n412,n108,n107);
and (n413,n414,n415);
xnor (n414,n118,n109);
nor (n415,n264,n228,n247,n256);
xor (n416,n363,n417);
and (n417,n74,n418);
and (n418,n382,n419);
and (n419,n399,n420);
wire s0n420,s1n420,notn420;
or (n420,s0n420,s1n420);
not(notn420,n285);
and (s0n420,notn420,1'b0);
and (s1n420,n285,n421);
or (n421,n422,n423,n425,n427,n429,n432,n433,1'b0);
and (n422,n97,n85);
and (n423,n424,n263);
not (n424,n84);
and (n425,n426,n270);
not (n426,n99);
and (n427,n428,n275);
not (n428,n101);
not (n429,n430);
nand (n430,n277,n431);
not (n431,n103);
and (n432,n106,n397);
and (n433,n434,n415);
not (n434,n109);
nor (n435,n436,n286);
not (n436,n332);
and (n437,n74,n438);
and (n438,n286,n436);
not (n439,n440);
nand (n440,n441,n465);
or (n441,n442,n449);
or (n442,n443,n448);
nor (n443,n444,n445,n447);
not (n445,n446);
and (n448,n444,n446,n447);
not (n449,n450);
nand (n450,n451,n459);
or (n451,1'b0,n452,n454,n458);
and (n452,n453,n358);
wire s0n453,s1n453,notn453;
or (n453,s0n453,s1n453);
not(notn453,n349);
and (s0n453,notn453,n382);
and (s1n453,n349,1'b0);
and (n454,n455,n435);
wire s0n455,s1n455,notn455;
or (n455,s0n455,s1n455);
not(notn455,n420);
and (s0n455,notn455,n456);
and (s1n455,n420,n457);
xor (n456,n379,n380);
xor (n457,n74,n418);
and (n458,n382,n438);
or (n459,1'b0,n460,n462,n464);
and (n460,n461,n358);
wire s0n461,s1n461,notn461;
or (n461,s0n461,s1n461);
not(notn461,n349);
and (s0n461,notn461,n399);
and (s1n461,n349,1'b0);
and (n462,n463,n435);
xor (n463,n381,n398);
and (n464,n399,n438);
nor (n465,n466,n489);
not (n466,n467);
or (n467,1'b0,n468,n470,n488);
and (n468,n469,n358);
wire s0n469,s1n469,notn469;
or (n469,s0n469,s1n469);
not(notn469,n349);
and (s0n469,notn469,n363);
and (s1n469,n349,1'b0);
and (n470,n471,n435);
wire s0n471,s1n471,notn471;
or (n471,s0n471,s1n471);
not(notn471,n420);
and (s0n471,notn471,n472);
and (s1n471,n420,n486);
xor (n472,n473,n485);
not (n473,n474);
wire s0n474,s1n474,notn474;
or (n474,s0n474,s1n474);
not(notn474,n285);
and (s0n474,notn474,1'b0);
and (s1n474,n285,n475);
or (n475,n476,n479,n482,1'b0,1'b0,1'b0,1'b0,1'b0);
and (n476,n477,n85);
xnor (n477,n100,n478);
or (n478,n367,n99);
and (n479,n480,n263);
xnor (n480,n102,n481);
or (n481,n101,n370);
and (n482,n483,n270);
xnor (n483,n114,n484);
or (n484,n103,n373);
and (n485,n362,n378);
xor (n486,n474,n487);
and (n487,n363,n417);
and (n488,n363,n438);
nor (n489,n490,n493);
nand (n490,n491,n492);
not (n491,n451);
not (n492,n459);
or (n493,1'b0,n494,n512,n514);
and (n494,n495,n358);
wire s0n495,s1n495,notn495;
or (n495,s0n495,s1n495);
not(notn495,n349);
and (s0n495,notn495,n420);
and (s1n495,n349,n496);
not (n496,n497);
nor (n497,n420,n399,n382,n74,n363,n474,n498,n509);
wire s0n498,s1n498,notn498;
or (n498,s0n498,s1n498);
not(notn498,n285);
and (s0n498,notn498,1'b0);
and (s1n498,n285,n499);
or (n499,n500,n506,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0);
and (n500,n501,n85);
nand (n501,n502,n504);
or (n502,n503,n428);
nor (n503,n367,n269);
nand (n504,n505,n268);
not (n505,n367);
and (n506,n507,n263);
xnor (n507,n103,n508);
or (n508,n102,n481);
wire s0n509,s1n509,notn509;
or (n509,s0n509,s1n509);
not(notn509,n285);
and (s0n509,notn509,1'b0);
and (s1n509,n285,n510);
and (n510,n511,n85);
xnor (n511,n102,n504);
and (n512,n513,n435);
xor (n513,n399,n420);
and (n514,n420,n438);
nand (n515,n516,n70);
or (n516,n517,n519);
not (n517,n518);
nor (n518,n467,n442);
not (n519,n520);
nand (n520,n521,n451);
nand (n521,n522,n492);
not (n522,n493);
nor (n523,n524,n558);
nand (n524,n525,n540,n549);
not (n525,n526);
or (n526,1'b0,n527,n529,n539);
and (n527,n528,n358);
wire s0n528,s1n528,notn528;
or (n528,s0n528,s1n528);
not(notn528,n349);
and (s0n528,notn528,n498);
and (s1n528,n349,1'b0);
and (n529,n530,n435);
wire s0n530,s1n530,notn530;
or (n530,s0n530,s1n530);
not(notn530,n420);
and (s0n530,notn530,n531);
and (s1n530,n420,n536);
xor (n531,n532,n533);
not (n532,n509);
and (n533,n534,n535);
not (n534,n498);
and (n535,n473,n485);
xor (n536,n509,n537);
and (n537,n498,n538);
and (n538,n474,n487);
and (n539,n498,n438);
not (n540,n541);
or (n541,1'b0,n542,n544,n548);
and (n542,n543,n358);
wire s0n543,s1n543,notn543;
or (n543,s0n543,s1n543);
not(notn543,n349);
and (s0n543,notn543,n474);
and (s1n543,n349,1'b0);
and (n544,n545,n435);
wire s0n545,s1n545,notn545;
or (n545,s0n545,s1n545);
not(notn545,n420);
and (s0n545,notn545,n546);
and (s1n545,n420,n547);
xor (n546,n534,n535);
xor (n547,n498,n538);
and (n548,n474,n438);
not (n549,n550);
or (n550,1'b0,n551,n553,n557);
and (n551,n552,n358);
wire s0n552,s1n552,notn552;
or (n552,s0n552,s1n552);
not(notn552,n349);
and (s0n552,notn552,n509);
and (s1n552,n349,1'b0);
and (n553,n554,n435);
wire s0n554,s1n554,notn554;
or (n554,s0n554,s1n554);
not(notn554,n420);
and (s0n554,notn554,n555);
and (s1n554,n420,1'b0);
not (n555,n556);
and (n556,n532,n533);
and (n557,n509,n438);
not (n558,n203);
not (n559,n560);
nor (n560,n561,n563,n564,n565);
not (n561,n562);
and (n566,n567,n43);
not (n567,n57);
nand (n568,n569,n570);
and (n569,n22,n566);
or (n570,1'b0,n571,n573,n577,n580);
and (n571,n572,n560);
and (n573,n574,n575);
nor (n575,n562,n576,n564,n565);
not (n576,n563);
and (n577,n578,n579);
nor (n579,n561,n576,n564,n565);
and (n580,n18,n581);
nor (n581,n562,n563,n582,n565);
not (n582,n564);
nor (n583,n584,n639,n686);
wire s0n584,s1n584,notn584;
or (n584,s0n584,s1n584);
not(notn584,n566);
and (s0n584,notn584,1'b0);
and (s1n584,n566,n585);
wire s0n585,s1n585,notn585;
or (n585,s0n585,s1n585);
not(notn585,n638);
and (s0n585,notn585,n586);
and (s1n585,n638,n629);
or (n586,n587,n605,n616,n627);
and (n587,n588,n29);
wire s0n588,s1n588,notn588;
or (n588,s0n588,s1n588);
not(notn588,n23);
and (s0n588,notn588,n589);
and (s1n588,n23,n590);
or (n590,n591,n596,n600,n603);
and (n591,n592,n593);
nor (n593,n594,n595);
and (n596,n597,n598);
and (n598,n594,n599);
not (n599,n595);
and (n600,n601,n602);
nor (n602,n594,n599);
and (n603,n589,n604);
and (n604,n594,n595);
and (n605,n606,n34);
wire s0n606,s1n606,notn606;
or (n606,s0n606,s1n606);
not(notn606,n23);
and (s0n606,notn606,n607);
and (s1n606,n23,n608);
or (n608,n609,n611,n613,n615);
and (n609,n610,n593);
and (n611,n612,n598);
and (n613,n614,n602);
and (n615,n607,n604);
and (n616,n617,n39);
wire s0n617,s1n617,notn617;
or (n617,s0n617,s1n617);
not(notn617,n23);
and (s0n617,notn617,n618);
and (s1n617,n23,n619);
or (n619,n620,n622,n624,n626);
and (n620,n621,n593);
and (n622,n623,n598);
and (n624,n625,n602);
and (n626,n618,n604);
and (n627,n628,n42);
wire s0n628,s1n628,notn628;
or (n628,s0n628,s1n628);
not(notn628,n23);
and (s0n628,notn628,n629);
and (s1n628,n23,n630);
or (n630,n631,n633,n635,n637);
and (n631,n632,n593);
and (n633,n634,n598);
and (n635,n636,n602);
and (n637,n629,n604);
wire s0n639,s1n639,notn639;
or (n639,s0n639,s1n639);
not(notn639,n566);
and (s0n639,notn639,1'b0);
and (s1n639,n566,n640);
wire s0n640,s1n640,notn640;
or (n640,s0n640,s1n640);
not(notn640,n638);
and (s0n640,notn640,n641);
and (s1n640,n638,n677);
or (n641,n642,n653,n664,n675);
and (n642,n643,n29);
wire s0n643,s1n643,notn643;
or (n643,s0n643,s1n643);
not(notn643,n23);
and (s0n643,notn643,n644);
and (s1n643,n23,n645);
or (n645,n646,n648,n650,n652);
and (n646,n647,n593);
and (n648,n649,n598);
and (n650,n651,n602);
and (n652,n644,n604);
and (n653,n654,n34);
wire s0n654,s1n654,notn654;
or (n654,s0n654,s1n654);
not(notn654,n23);
and (s0n654,notn654,n655);
and (s1n654,n23,n656);
or (n656,n657,n659,n661,n663);
and (n657,n658,n593);
and (n659,n660,n598);
and (n661,n662,n602);
and (n663,n655,n604);
and (n664,n665,n39);
wire s0n665,s1n665,notn665;
or (n665,s0n665,s1n665);
not(notn665,n23);
and (s0n665,notn665,n666);
and (s1n665,n23,n667);
or (n667,n668,n670,n672,n674);
and (n668,n669,n593);
and (n670,n671,n598);
and (n672,n673,n602);
and (n674,n666,n604);
and (n675,n676,n42);
wire s0n676,s1n676,notn676;
or (n676,s0n676,s1n676);
not(notn676,n23);
and (s0n676,notn676,n677);
and (s1n676,n23,n678);
or (n678,n679,n681,n683,n685);
and (n679,n680,n593);
and (n681,n682,n598);
and (n683,n684,n602);
and (n685,n677,n604);
wire s0n686,s1n686,notn686;
or (n686,s0n686,s1n686);
not(notn686,n566);
and (s0n686,notn686,1'b0);
and (s1n686,n566,n687);
wire s0n687,s1n687,notn687;
or (n687,s0n687,s1n687);
not(notn687,n638);
and (s0n687,notn687,n688);
and (s1n687,n638,n724);
or (n688,n689,n700,n711,n722);
and (n689,n690,n29);
wire s0n690,s1n690,notn690;
or (n690,s0n690,s1n690);
not(notn690,n23);
and (s0n690,notn690,n691);
and (s1n690,n23,n692);
or (n692,n693,n695,n697,n699);
and (n693,n694,n593);
and (n695,n696,n598);
and (n697,n698,n602);
and (n699,n691,n604);
and (n700,n701,n34);
wire s0n701,s1n701,notn701;
or (n701,s0n701,s1n701);
not(notn701,n23);
and (s0n701,notn701,n702);
and (s1n701,n23,n703);
or (n703,n704,n706,n708,n710);
and (n704,n705,n593);
and (n706,n707,n598);
and (n708,n709,n602);
and (n710,n702,n604);
and (n711,n712,n39);
wire s0n712,s1n712,notn712;
or (n712,s0n712,s1n712);
not(notn712,n23);
and (s0n712,notn712,n713);
and (s1n712,n23,n714);
or (n714,n715,n717,n719,n721);
and (n715,n716,n593);
and (n717,n718,n598);
and (n719,n720,n602);
and (n721,n713,n604);
and (n722,n723,n42);
wire s0n723,s1n723,notn723;
or (n723,s0n723,s1n723);
not(notn723,n23);
and (s0n723,notn723,n724);
and (s1n723,n23,n725);
or (n725,n726,n728,n730,n732);
and (n726,n727,n593);
and (n728,n729,n598);
and (n730,n731,n602);
and (n732,n724,n604);
or (n733,n734,n875,n933);
and (n734,n735,n756);
xor (n735,n736,n750);
wire s0n736,s1n736,notn736;
or (n736,s0n736,s1n736);
not(notn736,n583);
and (s0n736,notn736,1'b0);
and (s1n736,n583,n737);
nand (n737,n738,n741);
or (n738,n739,n19);
not (n739,n740);
nand (n741,n569,n742);
or (n742,1'b0,n743,n745,n747,n749);
and (n743,n744,n560);
and (n745,n746,n575);
and (n747,n748,n579);
and (n749,n740,n581);
wire s0n750,s1n750,notn750;
or (n750,s0n750,s1n750);
not(notn750,n751);
and (s0n750,notn750,1'b0);
and (s1n750,n751,n15);
xor (n751,n752,n753);
not (n752,n686);
and (n753,n754,n755);
not (n754,n639);
not (n755,n584);
and (n756,n757,n759);
wire s0n757,s1n757,notn757;
or (n757,s0n757,s1n757);
not(notn757,n758);
and (s0n757,notn757,1'b0);
and (s1n757,n758,n15);
xor (n758,n754,n755);
or (n759,n760,n763,n874);
and (n760,n761,n762);
wire s0n761,s1n761,notn761;
or (n761,s0n761,s1n761);
not(notn761,n758);
and (s0n761,notn761,1'b0);
and (s1n761,n758,n737);
wire s0n762,s1n762,notn762;
or (n762,s0n762,s1n762);
not(notn762,n584);
and (s0n762,notn762,1'b0);
and (s1n762,n584,n15);
and (n763,n762,n764);
or (n764,n765,n781,n873);
and (n765,n766,n780);
wire s0n766,s1n766,notn766;
or (n766,s0n766,s1n766);
not(notn766,n758);
and (s0n766,notn766,1'b0);
and (s1n766,n758,n767);
nand (n767,n768,n771);
or (n768,n769,n19);
not (n769,n770);
nand (n771,n569,n772);
or (n772,1'b0,n773,n775,n777,n779);
and (n773,n774,n560);
and (n775,n776,n575);
and (n777,n778,n579);
and (n779,n770,n581);
wire s0n780,s1n780,notn780;
or (n780,s0n780,s1n780);
not(notn780,n584);
and (s0n780,notn780,1'b0);
and (s1n780,n584,n737);
and (n781,n780,n782);
or (n782,n783,n799,n872);
and (n783,n784,n798);
wire s0n784,s1n784,notn784;
or (n784,s0n784,s1n784);
not(notn784,n758);
and (s0n784,notn784,1'b0);
and (s1n784,n758,n785);
nand (n785,n786,n789);
or (n786,n787,n19);
not (n787,n788);
nand (n789,n569,n790);
or (n790,1'b0,n791,n793,n795,n797);
and (n791,n792,n560);
and (n793,n794,n575);
and (n795,n796,n579);
and (n797,n788,n581);
wire s0n798,s1n798,notn798;
or (n798,s0n798,s1n798);
not(notn798,n584);
and (s0n798,notn798,1'b0);
and (s1n798,n584,n767);
and (n799,n798,n800);
or (n800,n801,n817,n871);
and (n801,n802,n816);
wire s0n802,s1n802,notn802;
or (n802,s0n802,s1n802);
not(notn802,n758);
and (s0n802,notn802,1'b0);
and (s1n802,n758,n803);
nand (n803,n804,n807);
or (n804,n805,n19);
not (n805,n806);
nand (n807,n569,n808);
or (n808,1'b0,n809,n811,n813,n815);
and (n809,n810,n560);
and (n811,n812,n575);
and (n813,n814,n579);
and (n815,n806,n581);
wire s0n816,s1n816,notn816;
or (n816,s0n816,s1n816);
not(notn816,n584);
and (s0n816,notn816,1'b0);
and (s1n816,n584,n785);
and (n817,n816,n818);
or (n818,n819,n836,n838);
and (n819,n820,n835);
wire s0n820,s1n820,notn820;
or (n820,s0n820,s1n820);
not(notn820,n758);
and (s0n820,notn820,1'b0);
and (s1n820,n758,n821);
nand (n821,n822,n834);
or (n822,n823,n833);
not (n823,n824);
or (n824,1'b0,n825,n827,n829,n831);
and (n825,n826,n560);
and (n827,n828,n575);
and (n829,n830,n579);
and (n831,n832,n581);
not (n833,n569);
nand (n834,n20,n832);
wire s0n835,s1n835,notn835;
or (n835,s0n835,s1n835);
not(notn835,n584);
and (s0n835,notn835,1'b0);
and (s1n835,n584,n803);
and (n836,n835,n837);
or (n837,n838,n854,n855);
and (n838,n839,n853);
wire s0n839,s1n839,notn839;
or (n839,s0n839,s1n839);
not(notn839,n758);
and (s0n839,notn839,1'b0);
and (s1n839,n758,n840);
nand (n840,n841,n852);
or (n841,n842,n833);
not (n842,n843);
or (n843,1'b0,n844,n846,n848,n850);
and (n844,n845,n560);
and (n846,n847,n575);
and (n848,n849,n579);
and (n850,n851,n581);
nand (n852,n20,n851);
wire s0n853,s1n853,notn853;
or (n853,s0n853,s1n853);
not(notn853,n584);
and (s0n853,notn853,1'b0);
and (s1n853,n584,n821);
and (n854,n853,n855);
and (n855,n856,n870);
wire s0n856,s1n856,notn856;
or (n856,s0n856,s1n856);
not(notn856,n758);
and (s0n856,notn856,1'b0);
and (s1n856,n758,n857);
nand (n857,n858,n861);
or (n858,n859,n19);
not (n859,n860);
nand (n861,n569,n862);
or (n862,1'b0,n863,n865,n867,n869);
and (n863,n864,n560);
and (n865,n866,n575);
and (n867,n868,n579);
and (n869,n860,n581);
wire s0n870,s1n870,notn870;
or (n870,s0n870,s1n870);
not(notn870,n584);
and (s0n870,notn870,1'b0);
and (s1n870,n584,n840);
and (n871,n802,n818);
and (n872,n784,n800);
and (n873,n766,n782);
and (n874,n761,n764);
and (n875,n756,n876);
or (n876,n877,n882,n932);
and (n877,n878,n881);
xor (n878,n879,n880);
wire s0n879,s1n879,notn879;
or (n879,s0n879,s1n879);
not(notn879,n583);
and (s0n879,notn879,1'b0);
and (s1n879,n583,n767);
wire s0n880,s1n880,notn880;
or (n880,s0n880,s1n880);
not(notn880,n751);
and (s0n880,notn880,1'b0);
and (s1n880,n751,n737);
xor (n881,n757,n759);
and (n882,n881,n883);
or (n883,n884,n890,n931);
and (n884,n885,n888);
xor (n885,n886,n887);
wire s0n886,s1n886,notn886;
or (n886,s0n886,s1n886);
not(notn886,n583);
and (s0n886,notn886,1'b0);
and (s1n886,n583,n785);
wire s0n887,s1n887,notn887;
or (n887,s0n887,s1n887);
not(notn887,n751);
and (s0n887,notn887,1'b0);
and (s1n887,n751,n767);
xor (n888,n889,n764);
xor (n889,n761,n762);
and (n890,n888,n891);
or (n891,n892,n898,n930);
and (n892,n893,n896);
xor (n893,n894,n895);
wire s0n894,s1n894,notn894;
or (n894,s0n894,s1n894);
not(notn894,n583);
and (s0n894,notn894,1'b0);
and (s1n894,n583,n803);
wire s0n895,s1n895,notn895;
or (n895,s0n895,s1n895);
not(notn895,n751);
and (s0n895,notn895,1'b0);
and (s1n895,n751,n785);
xor (n896,n897,n782);
xor (n897,n766,n780);
and (n898,n896,n899);
or (n899,n900,n906,n929);
and (n900,n901,n904);
xor (n901,n902,n903);
wire s0n902,s1n902,notn902;
or (n902,s0n902,s1n902);
not(notn902,n583);
and (s0n902,notn902,1'b0);
and (s1n902,n583,n821);
wire s0n903,s1n903,notn903;
or (n903,s0n903,s1n903);
not(notn903,n751);
and (s0n903,notn903,1'b0);
and (s1n903,n751,n803);
xor (n904,n905,n800);
xor (n905,n784,n798);
and (n906,n904,n907);
or (n907,n908,n914,n928);
and (n908,n909,n912);
xor (n909,n910,n911);
wire s0n910,s1n910,notn910;
or (n910,s0n910,s1n910);
not(notn910,n583);
and (s0n910,notn910,1'b0);
and (s1n910,n583,n840);
wire s0n911,s1n911,notn911;
or (n911,s0n911,s1n911);
not(notn911,n751);
and (s0n911,notn911,1'b0);
and (s1n911,n751,n821);
xor (n912,n913,n818);
xor (n913,n802,n816);
and (n914,n912,n915);
or (n915,n916,n922,n927);
and (n916,n917,n920);
xor (n917,n918,n919);
wire s0n918,s1n918,notn918;
or (n918,s0n918,s1n918);
not(notn918,n583);
and (s0n918,notn918,1'b0);
and (s1n918,n583,n857);
wire s0n919,s1n919,notn919;
or (n919,s0n919,s1n919);
not(notn919,n751);
and (s0n919,notn919,1'b0);
and (s1n919,n751,n840);
xor (n920,n921,n837);
xor (n921,n820,n835);
and (n922,n920,n923);
and (n923,n924,n925);
wire s0n924,s1n924,notn924;
or (n924,s0n924,s1n924);
not(notn924,n751);
and (s0n924,notn924,1'b0);
and (s1n924,n751,n857);
xor (n925,n926,n855);
xor (n926,n839,n853);
and (n927,n917,n923);
and (n928,n909,n915);
and (n929,n901,n907);
and (n930,n893,n899);
and (n931,n885,n891);
and (n932,n878,n883);
and (n933,n735,n876);
wire s0n934,s1n934,notn934;
or (n934,s0n934,s1n934);
not(notn934,n566);
and (s0n934,notn934,1'b0);
and (s1n934,n566,n935);
wire s0n935,s1n935,notn935;
or (n935,s0n935,s1n935);
not(notn935,n638);
and (s0n935,notn935,n936);
and (s1n935,n638,n972);
or (n936,n937,n948,n959,n970);
and (n937,n938,n29);
wire s0n938,s1n938,notn938;
or (n938,s0n938,s1n938);
not(notn938,n23);
and (s0n938,notn938,n939);
and (s1n938,n23,n940);
or (n940,n941,n943,n945,n947);
and (n941,n942,n593);
and (n943,n944,n598);
and (n945,n946,n602);
and (n947,n939,n604);
and (n948,n949,n34);
wire s0n949,s1n949,notn949;
or (n949,s0n949,s1n949);
not(notn949,n23);
and (s0n949,notn949,n950);
and (s1n949,n23,n951);
or (n951,n952,n954,n956,n958);
and (n952,n953,n593);
and (n954,n955,n598);
and (n956,n957,n602);
and (n958,n950,n604);
and (n959,n960,n39);
wire s0n960,s1n960,notn960;
or (n960,s0n960,s1n960);
not(notn960,n23);
and (s0n960,notn960,n961);
and (s1n960,n23,n962);
or (n962,n963,n965,n967,n969);
and (n963,n964,n593);
and (n965,n966,n598);
and (n967,n968,n602);
and (n969,n961,n604);
and (n970,n971,n42);
wire s0n971,s1n971,notn971;
or (n971,s0n971,s1n971);
not(notn971,n23);
and (s0n971,notn971,n972);
and (s1n971,n23,n973);
or (n973,n974,n976,n978,n980);
and (n974,n975,n593);
and (n976,n977,n598);
and (n978,n979,n602);
and (n980,n972,n604);
wire s0n981,s1n981,notn981;
or (n981,s0n981,s1n981);
not(notn981,n934);
and (s0n981,notn981,1'b0);
and (s1n981,n934,n982);
or (n982,n983,n1129,n1181);
and (n983,n984,n999);
not (n984,n985);
nand (n985,n686,n986);
nand (n986,n987,n998);
or (n987,n988,n833);
not (n988,n989);
or (n989,1'b0,n990,n992,n994,n996);
and (n990,n991,n560);
and (n992,n993,n575);
and (n994,n995,n579);
and (n996,n997,n581);
nand (n998,n20,n997);
and (n999,n1000,n1001);
wire s0n1000,s1n1000,notn1000;
or (n1000,s0n1000,s1n1000);
not(notn1000,n639);
and (s0n1000,notn1000,1'b0);
and (s1n1000,n639,n986);
or (n1001,n1002,n1018,n1128);
and (n1002,n1003,n1017);
wire s0n1003,s1n1003,notn1003;
or (n1003,s0n1003,s1n1003);
not(notn1003,n639);
and (s0n1003,notn1003,1'b0);
and (s1n1003,n639,n1004);
nand (n1004,n1005,n1016);
or (n1005,n1006,n833);
not (n1006,n1007);
or (n1007,1'b0,n1008,n1010,n1012,n1014);
and (n1008,n1009,n560);
and (n1010,n1011,n575);
and (n1012,n1013,n579);
and (n1014,n1015,n581);
nand (n1016,n20,n1015);
wire s0n1017,s1n1017,notn1017;
or (n1017,s0n1017,s1n1017);
not(notn1017,n584);
and (s0n1017,notn1017,1'b0);
and (s1n1017,n584,n986);
and (n1018,n1017,n1019);
or (n1019,n1020,n1036,n1127);
and (n1020,n1021,n1035);
wire s0n1021,s1n1021,notn1021;
or (n1021,s0n1021,s1n1021);
not(notn1021,n639);
and (s0n1021,notn1021,1'b0);
and (s1n1021,n639,n1022);
nand (n1022,n1023,n1034);
or (n1023,n1024,n833);
not (n1024,n1025);
or (n1025,1'b0,n1026,n1028,n1030,n1032);
and (n1026,n1027,n560);
and (n1028,n1029,n575);
and (n1030,n1031,n579);
and (n1032,n1033,n581);
nand (n1034,n20,n1033);
wire s0n1035,s1n1035,notn1035;
or (n1035,s0n1035,s1n1035);
not(notn1035,n584);
and (s0n1035,notn1035,1'b0);
and (s1n1035,n584,n1004);
and (n1036,n1035,n1037);
or (n1037,n1038,n1054,n1126);
and (n1038,n1039,n1053);
wire s0n1039,s1n1039,notn1039;
or (n1039,s0n1039,s1n1039);
not(notn1039,n639);
and (s0n1039,notn1039,1'b0);
and (s1n1039,n639,n1040);
nand (n1040,n1041,n1052);
or (n1041,n1042,n833);
not (n1042,n1043);
or (n1043,1'b0,n1044,n1046,n1048,n1050);
and (n1044,n1045,n560);
and (n1046,n1047,n575);
and (n1048,n1049,n579);
and (n1050,n1051,n581);
nand (n1052,n20,n1051);
wire s0n1053,s1n1053,notn1053;
or (n1053,s0n1053,s1n1053);
not(notn1053,n584);
and (s0n1053,notn1053,1'b0);
and (s1n1053,n584,n1022);
and (n1054,n1053,n1055);
or (n1055,n1056,n1072,n1125);
and (n1056,n1057,n1071);
wire s0n1057,s1n1057,notn1057;
or (n1057,s0n1057,s1n1057);
not(notn1057,n639);
and (s0n1057,notn1057,1'b0);
and (s1n1057,n639,n1058);
nand (n1058,n1059,n1070);
or (n1059,n1060,n833);
not (n1060,n1061);
or (n1061,1'b0,n1062,n1064,n1066,n1068);
and (n1062,n1063,n560);
and (n1064,n1065,n575);
and (n1066,n1067,n579);
and (n1068,n1069,n581);
nand (n1070,n20,n1069);
wire s0n1071,s1n1071,notn1071;
or (n1071,s0n1071,s1n1071);
not(notn1071,n584);
and (s0n1071,notn1071,1'b0);
and (s1n1071,n584,n1040);
and (n1072,n1071,n1073);
or (n1073,n1074,n1090,n1092);
and (n1074,n1075,n1089);
wire s0n1075,s1n1075,notn1075;
or (n1075,s0n1075,s1n1075);
not(notn1075,n639);
and (s0n1075,notn1075,1'b0);
and (s1n1075,n639,n1076);
nand (n1076,n1077,n1080);
or (n1077,n1078,n19);
not (n1078,n1079);
nand (n1080,n569,n1081);
or (n1081,1'b0,n1082,n1084,n1086,n1088);
and (n1082,n1083,n560);
and (n1084,n1085,n575);
and (n1086,n1087,n579);
and (n1088,n1079,n581);
wire s0n1089,s1n1089,notn1089;
or (n1089,s0n1089,s1n1089);
not(notn1089,n584);
and (s0n1089,notn1089,1'b0);
and (s1n1089,n584,n1058);
and (n1090,n1089,n1091);
or (n1091,n1092,n1108,n1109);
and (n1092,n1093,n1107);
wire s0n1093,s1n1093,notn1093;
or (n1093,s0n1093,s1n1093);
not(notn1093,n639);
and (s0n1093,notn1093,1'b0);
and (s1n1093,n639,n1094);
nand (n1094,n1095,n1106);
or (n1095,n1096,n833);
not (n1096,n1097);
or (n1097,1'b0,n1098,n1100,n1102,n1104);
and (n1098,n1099,n560);
and (n1100,n1101,n575);
and (n1102,n1103,n579);
and (n1104,n1105,n581);
nand (n1106,n20,n1105);
wire s0n1107,s1n1107,notn1107;
or (n1107,s0n1107,s1n1107);
not(notn1107,n584);
and (s0n1107,notn1107,1'b0);
and (s1n1107,n584,n1076);
and (n1108,n1107,n1109);
and (n1109,n1110,n1124);
wire s0n1110,s1n1110,notn1110;
or (n1110,s0n1110,s1n1110);
not(notn1110,n639);
and (s0n1110,notn1110,1'b0);
and (s1n1110,n639,n1111);
nand (n1111,n1112,n1123);
or (n1112,n1113,n833);
not (n1113,n1114);
or (n1114,1'b0,n1115,n1117,n1119,n1121);
and (n1115,n1116,n560);
and (n1117,n1118,n575);
and (n1119,n1120,n579);
and (n1121,n1122,n581);
nand (n1123,n20,n1122);
wire s0n1124,s1n1124,notn1124;
or (n1124,s0n1124,s1n1124);
not(notn1124,n584);
and (s0n1124,notn1124,1'b0);
and (s1n1124,n584,n1094);
and (n1125,n1057,n1073);
and (n1126,n1039,n1055);
and (n1127,n1021,n1037);
and (n1128,n1003,n1019);
and (n1129,n999,n1130);
or (n1130,n1131,n1135,n1180);
and (n1131,n1132,n1134);
not (n1132,n1133);
nand (n1133,n686,n1004);
xor (n1134,n1000,n1001);
and (n1135,n1134,n1136);
or (n1136,n1137,n1142,n1179);
and (n1137,n1138,n1140);
not (n1138,n1139);
nand (n1139,n686,n1022);
xor (n1140,n1141,n1019);
xor (n1141,n1003,n1017);
and (n1142,n1140,n1143);
or (n1143,n1144,n1149,n1178);
and (n1144,n1145,n1147);
not (n1145,n1146);
nand (n1146,n686,n1040);
xor (n1147,n1148,n1037);
xor (n1148,n1021,n1035);
and (n1149,n1147,n1150);
or (n1150,n1151,n1155,n1177);
and (n1151,n1152,n1153);
and (n1152,n686,n1058);
xor (n1153,n1154,n1055);
xor (n1154,n1039,n1053);
and (n1155,n1153,n1156);
or (n1156,n1157,n1162,n1176);
and (n1157,n1158,n1160);
not (n1158,n1159);
nand (n1159,n686,n1076);
xor (n1160,n1161,n1073);
xor (n1161,n1057,n1071);
and (n1162,n1160,n1163);
or (n1163,n1164,n1169,n1175);
and (n1164,n1165,n1167);
not (n1165,n1166);
nand (n1166,n686,n1094);
xor (n1167,n1168,n1091);
xor (n1168,n1075,n1089);
and (n1169,n1167,n1170);
and (n1170,n1171,n1173);
not (n1171,n1172);
nand (n1172,n686,n1111);
xor (n1173,n1174,n1109);
xor (n1174,n1093,n1107);
and (n1175,n1165,n1170);
and (n1176,n1158,n1163);
and (n1177,n1152,n1156);
and (n1178,n1145,n1150);
and (n1179,n1138,n1143);
and (n1180,n1132,n1136);
and (n1181,n984,n1130);
wire s0n1182,s1n1182,notn1182;
or (n1182,s0n1182,s1n1182);
not(notn1182,n1392);
and (s0n1182,notn1182,1'b0);
and (s1n1182,n1392,n1183);
xor (n1183,n1184,n1198);
wire s0n1184,s1n1184,notn1184;
or (n1184,s0n1184,s1n1184);
not(notn1184,n583);
and (s0n1184,notn1184,1'b0);
and (s1n1184,n583,n1185);
nand (n1185,n1186,n1189);
or (n1186,n1187,n19);
not (n1187,n1188);
nand (n1189,n569,n1190);
or (n1190,1'b0,n1191,n1193,n1195,n1197);
and (n1191,n1192,n560);
and (n1193,n1194,n575);
and (n1195,n1196,n579);
and (n1197,n1188,n581);
or (n1198,n1199,n1333,n1391);
and (n1199,n1200,n1216);
xor (n1200,n1201,n1215);
wire s0n1201,s1n1201,notn1201;
or (n1201,s0n1201,s1n1201);
not(notn1201,n583);
and (s0n1201,notn1201,1'b0);
and (s1n1201,n583,n1202);
nand (n1202,n1203,n1206);
or (n1203,n1204,n19);
not (n1204,n1205);
nand (n1206,n569,n1207);
or (n1207,1'b0,n1208,n1210,n1212,n1214);
and (n1208,n1209,n560);
and (n1210,n1211,n575);
and (n1212,n1213,n579);
and (n1214,n1205,n581);
wire s0n1215,s1n1215,notn1215;
or (n1215,s0n1215,s1n1215);
not(notn1215,n751);
and (s0n1215,notn1215,1'b0);
and (s1n1215,n751,n1185);
and (n1216,n1217,n1218);
wire s0n1217,s1n1217,notn1217;
or (n1217,s0n1217,s1n1217);
not(notn1217,n758);
and (s0n1217,notn1217,1'b0);
and (s1n1217,n758,n1185);
or (n1218,n1219,n1222,n1332);
and (n1219,n1220,n1221);
wire s0n1220,s1n1220,notn1220;
or (n1220,s0n1220,s1n1220);
not(notn1220,n758);
and (s0n1220,notn1220,1'b0);
and (s1n1220,n758,n1202);
wire s0n1221,s1n1221,notn1221;
or (n1221,s0n1221,s1n1221);
not(notn1221,n584);
and (s0n1221,notn1221,1'b0);
and (s1n1221,n584,n1185);
and (n1222,n1221,n1223);
or (n1223,n1224,n1240,n1331);
and (n1224,n1225,n1239);
wire s0n1225,s1n1225,notn1225;
or (n1225,s0n1225,s1n1225);
not(notn1225,n758);
and (s0n1225,notn1225,1'b0);
and (s1n1225,n758,n1226);
nand (n1226,n1227,n1230);
or (n1227,n1228,n19);
not (n1228,n1229);
nand (n1230,n569,n1231);
or (n1231,1'b0,n1232,n1234,n1236,n1238);
and (n1232,n1233,n560);
and (n1234,n1235,n575);
and (n1236,n1237,n579);
and (n1238,n1229,n581);
wire s0n1239,s1n1239,notn1239;
or (n1239,s0n1239,s1n1239);
not(notn1239,n584);
and (s0n1239,notn1239,1'b0);
and (s1n1239,n584,n1202);
and (n1240,n1239,n1241);
or (n1241,n1242,n1258,n1330);
and (n1242,n1243,n1257);
wire s0n1243,s1n1243,notn1243;
or (n1243,s0n1243,s1n1243);
not(notn1243,n758);
and (s0n1243,notn1243,1'b0);
and (s1n1243,n758,n1244);
nand (n1244,n1245,n1248);
or (n1245,n1246,n19);
not (n1246,n1247);
nand (n1248,n569,n1249);
or (n1249,1'b0,n1250,n1252,n1254,n1256);
and (n1250,n1251,n560);
and (n1252,n1253,n575);
and (n1254,n1255,n579);
and (n1256,n1247,n581);
wire s0n1257,s1n1257,notn1257;
or (n1257,s0n1257,s1n1257);
not(notn1257,n584);
and (s0n1257,notn1257,1'b0);
and (s1n1257,n584,n1226);
and (n1258,n1257,n1259);
or (n1259,n1260,n1276,n1329);
and (n1260,n1261,n1275);
wire s0n1261,s1n1261,notn1261;
or (n1261,s0n1261,s1n1261);
not(notn1261,n758);
and (s0n1261,notn1261,1'b0);
and (s1n1261,n758,n1262);
nand (n1262,n1263,n1266);
or (n1263,n1264,n19);
not (n1264,n1265);
nand (n1266,n569,n1267);
or (n1267,1'b0,n1268,n1270,n1272,n1274);
and (n1268,n1269,n560);
and (n1270,n1271,n575);
and (n1272,n1273,n579);
and (n1274,n1265,n581);
wire s0n1275,s1n1275,notn1275;
or (n1275,s0n1275,s1n1275);
not(notn1275,n584);
and (s0n1275,notn1275,1'b0);
and (s1n1275,n584,n1244);
and (n1276,n1275,n1277);
or (n1277,n1278,n1294,n1296);
and (n1278,n1279,n1293);
wire s0n1279,s1n1279,notn1279;
or (n1279,s0n1279,s1n1279);
not(notn1279,n758);
and (s0n1279,notn1279,1'b0);
and (s1n1279,n758,n1280);
nand (n1280,n1281,n1284);
or (n1281,n1282,n19);
not (n1282,n1283);
nand (n1284,n569,n1285);
or (n1285,1'b0,n1286,n1288,n1290,n1292);
and (n1286,n1287,n560);
and (n1288,n1289,n575);
and (n1290,n1291,n579);
and (n1292,n1283,n581);
wire s0n1293,s1n1293,notn1293;
or (n1293,s0n1293,s1n1293);
not(notn1293,n584);
and (s0n1293,notn1293,1'b0);
and (s1n1293,n584,n1262);
and (n1294,n1293,n1295);
or (n1295,n1296,n1312,n1313);
and (n1296,n1297,n1311);
wire s0n1297,s1n1297,notn1297;
or (n1297,s0n1297,s1n1297);
not(notn1297,n758);
and (s0n1297,notn1297,1'b0);
and (s1n1297,n758,n1298);
nand (n1298,n1299,n1302);
or (n1299,n1300,n19);
not (n1300,n1301);
nand (n1302,n569,n1303);
or (n1303,1'b0,n1304,n1306,n1308,n1310);
and (n1304,n1305,n560);
and (n1306,n1307,n575);
and (n1308,n1309,n579);
and (n1310,n1301,n581);
wire s0n1311,s1n1311,notn1311;
or (n1311,s0n1311,s1n1311);
not(notn1311,n584);
and (s0n1311,notn1311,1'b0);
and (s1n1311,n584,n1280);
and (n1312,n1311,n1313);
and (n1313,n1314,n1328);
wire s0n1314,s1n1314,notn1314;
or (n1314,s0n1314,s1n1314);
not(notn1314,n758);
and (s0n1314,notn1314,1'b0);
and (s1n1314,n758,n1315);
nand (n1315,n1316,n1327);
or (n1316,n1317,n833);
not (n1317,n1318);
or (n1318,1'b0,n1319,n1321,n1323,n1325);
and (n1319,n1320,n560);
and (n1321,n1322,n575);
and (n1323,n1324,n579);
and (n1325,n1326,n581);
nand (n1327,n20,n1326);
wire s0n1328,s1n1328,notn1328;
or (n1328,s0n1328,s1n1328);
not(notn1328,n584);
and (s0n1328,notn1328,1'b0);
and (s1n1328,n584,n1298);
and (n1329,n1261,n1277);
and (n1330,n1243,n1259);
and (n1331,n1225,n1241);
and (n1332,n1220,n1223);
and (n1333,n1216,n1334);
or (n1334,n1335,n1340,n1390);
and (n1335,n1336,n1339);
xor (n1336,n1337,n1338);
wire s0n1337,s1n1337,notn1337;
or (n1337,s0n1337,s1n1337);
not(notn1337,n583);
and (s0n1337,notn1337,1'b0);
and (s1n1337,n583,n1226);
wire s0n1338,s1n1338,notn1338;
or (n1338,s0n1338,s1n1338);
not(notn1338,n751);
and (s0n1338,notn1338,1'b0);
and (s1n1338,n751,n1202);
xor (n1339,n1217,n1218);
and (n1340,n1339,n1341);
or (n1341,n1342,n1348,n1389);
and (n1342,n1343,n1346);
xor (n1343,n1344,n1345);
wire s0n1344,s1n1344,notn1344;
or (n1344,s0n1344,s1n1344);
not(notn1344,n583);
and (s0n1344,notn1344,1'b0);
and (s1n1344,n583,n1244);
wire s0n1345,s1n1345,notn1345;
or (n1345,s0n1345,s1n1345);
not(notn1345,n751);
and (s0n1345,notn1345,1'b0);
and (s1n1345,n751,n1226);
xor (n1346,n1347,n1223);
xor (n1347,n1220,n1221);
and (n1348,n1346,n1349);
or (n1349,n1350,n1356,n1388);
and (n1350,n1351,n1354);
xor (n1351,n1352,n1353);
wire s0n1352,s1n1352,notn1352;
or (n1352,s0n1352,s1n1352);
not(notn1352,n583);
and (s0n1352,notn1352,1'b0);
and (s1n1352,n583,n1262);
wire s0n1353,s1n1353,notn1353;
or (n1353,s0n1353,s1n1353);
not(notn1353,n751);
and (s0n1353,notn1353,1'b0);
and (s1n1353,n751,n1244);
xor (n1354,n1355,n1241);
xor (n1355,n1225,n1239);
and (n1356,n1354,n1357);
or (n1357,n1358,n1364,n1387);
and (n1358,n1359,n1362);
xor (n1359,n1360,n1361);
wire s0n1360,s1n1360,notn1360;
or (n1360,s0n1360,s1n1360);
not(notn1360,n583);
and (s0n1360,notn1360,1'b0);
and (s1n1360,n583,n1280);
wire s0n1361,s1n1361,notn1361;
or (n1361,s0n1361,s1n1361);
not(notn1361,n751);
and (s0n1361,notn1361,1'b0);
and (s1n1361,n751,n1262);
xor (n1362,n1363,n1259);
xor (n1363,n1243,n1257);
and (n1364,n1362,n1365);
or (n1365,n1366,n1372,n1386);
and (n1366,n1367,n1370);
xor (n1367,n1368,n1369);
wire s0n1368,s1n1368,notn1368;
or (n1368,s0n1368,s1n1368);
not(notn1368,n583);
and (s0n1368,notn1368,1'b0);
and (s1n1368,n583,n1298);
wire s0n1369,s1n1369,notn1369;
or (n1369,s0n1369,s1n1369);
not(notn1369,n751);
and (s0n1369,notn1369,1'b0);
and (s1n1369,n751,n1280);
xor (n1370,n1371,n1277);
xor (n1371,n1261,n1275);
and (n1372,n1370,n1373);
or (n1373,n1374,n1380,n1385);
and (n1374,n1375,n1378);
xor (n1375,n1376,n1377);
wire s0n1376,s1n1376,notn1376;
or (n1376,s0n1376,s1n1376);
not(notn1376,n583);
and (s0n1376,notn1376,1'b0);
and (s1n1376,n583,n1315);
wire s0n1377,s1n1377,notn1377;
or (n1377,s0n1377,s1n1377);
not(notn1377,n751);
and (s0n1377,notn1377,1'b0);
and (s1n1377,n751,n1298);
xor (n1378,n1379,n1295);
xor (n1379,n1279,n1293);
and (n1380,n1378,n1381);
and (n1381,n1382,n1383);
wire s0n1382,s1n1382,notn1382;
or (n1382,s0n1382,s1n1382);
not(notn1382,n751);
and (s0n1382,notn1382,1'b0);
and (s1n1382,n751,n1315);
xor (n1383,n1384,n1313);
xor (n1384,n1297,n1311);
and (n1385,n1375,n1381);
and (n1386,n1367,n1373);
and (n1387,n1359,n1365);
and (n1388,n1351,n1357);
and (n1389,n1343,n1349);
and (n1390,n1336,n1341);
and (n1391,n1200,n1334);
xor (n1392,n1393,n1394);
not (n1393,n934);
and (n1394,n1395,n1443);
not (n1395,n1396);
wire s0n1396,s1n1396,notn1396;
or (n1396,s0n1396,s1n1396);
not(notn1396,n566);
and (s0n1396,notn1396,1'b0);
and (s1n1396,n566,n1397);
wire s0n1397,s1n1397,notn1397;
or (n1397,s0n1397,s1n1397);
not(notn1397,n638);
and (s0n1397,notn1397,n1398);
and (s1n1397,n638,n1434);
or (n1398,n1399,n1410,n1421,n1432);
and (n1399,n1400,n29);
wire s0n1400,s1n1400,notn1400;
or (n1400,s0n1400,s1n1400);
not(notn1400,n23);
and (s0n1400,notn1400,n1401);
and (s1n1400,n23,n1402);
or (n1402,n1403,n1405,n1407,n1409);
and (n1403,n1404,n593);
and (n1405,n1406,n598);
and (n1407,n1408,n602);
and (n1409,n1401,n604);
and (n1410,n1411,n34);
wire s0n1411,s1n1411,notn1411;
or (n1411,s0n1411,s1n1411);
not(notn1411,n23);
and (s0n1411,notn1411,n1412);
and (s1n1411,n23,n1413);
or (n1413,n1414,n1416,n1418,n1420);
and (n1414,n1415,n593);
and (n1416,n1417,n598);
and (n1418,n1419,n602);
and (n1420,n1412,n604);
and (n1421,n1422,n39);
wire s0n1422,s1n1422,notn1422;
or (n1422,s0n1422,s1n1422);
not(notn1422,n23);
and (s0n1422,notn1422,n1423);
and (s1n1422,n23,n1424);
or (n1424,n1425,n1427,n1429,n1431);
and (n1425,n1426,n593);
and (n1427,n1428,n598);
and (n1429,n1430,n602);
and (n1431,n1423,n604);
and (n1432,n1433,n42);
wire s0n1433,s1n1433,notn1433;
or (n1433,s0n1433,s1n1433);
not(notn1433,n23);
and (s0n1433,notn1433,n1434);
and (s1n1433,n23,n1435);
or (n1435,n1436,n1438,n1440,n1442);
and (n1436,n1437,n593);
and (n1438,n1439,n598);
and (n1440,n1441,n602);
and (n1442,n1434,n604);
not (n1443,n1444);
wire s0n1444,s1n1444,notn1444;
or (n1444,s0n1444,s1n1444);
not(notn1444,n566);
and (s0n1444,notn1444,1'b0);
and (s1n1444,n566,n1445);
wire s0n1445,s1n1445,notn1445;
or (n1445,s0n1445,s1n1445);
not(notn1445,n638);
and (s0n1445,notn1445,n1446);
and (s1n1445,n638,n1482);
or (n1446,n1447,n1458,n1469,n1480);
and (n1447,n1448,n29);
wire s0n1448,s1n1448,notn1448;
or (n1448,s0n1448,s1n1448);
not(notn1448,n23);
and (s0n1448,notn1448,n1449);
and (s1n1448,n23,n1450);
or (n1450,n1451,n1453,n1455,n1457);
and (n1451,n1452,n593);
and (n1453,n1454,n598);
and (n1455,n1456,n602);
and (n1457,n1449,n604);
and (n1458,n1459,n34);
wire s0n1459,s1n1459,notn1459;
or (n1459,s0n1459,s1n1459);
not(notn1459,n23);
and (s0n1459,notn1459,n1460);
and (s1n1459,n23,n1461);
or (n1461,n1462,n1464,n1466,n1468);
and (n1462,n1463,n593);
and (n1464,n1465,n598);
and (n1466,n1467,n602);
and (n1468,n1460,n604);
and (n1469,n1470,n39);
wire s0n1470,s1n1470,notn1470;
or (n1470,s0n1470,s1n1470);
not(notn1470,n23);
and (s0n1470,notn1470,n1471);
and (s1n1470,n23,n1472);
or (n1472,n1473,n1475,n1477,n1479);
and (n1473,n1474,n593);
and (n1475,n1476,n598);
and (n1477,n1478,n602);
and (n1479,n1471,n604);
and (n1480,n1481,n42);
wire s0n1481,s1n1481,notn1481;
or (n1481,s0n1481,s1n1481);
not(notn1481,n23);
and (s0n1481,notn1481,n1482);
and (s1n1481,n23,n1483);
or (n1483,n1484,n1486,n1488,n1490);
and (n1484,n1485,n593);
and (n1486,n1487,n598);
and (n1488,n1489,n602);
and (n1490,n1482,n604);
not (n1491,n1492);
nor (n1492,n1493,n1702);
and (n1493,n1494,n1699);
xor (n1494,n1495,n1694);
wire s0n1495,s1n1495,notn1495;
or (n1495,s0n1495,s1n1495);
not(notn1495,n1693);
and (s0n1495,notn1495,1'b0);
and (s1n1495,n1693,n1496);
xor (n1496,n1497,n1642);
xor (n1497,n1498,n1512);
and (n1498,n686,n1499);
nand (n1499,n1500,n1503);
or (n1500,n1501,n19);
not (n1501,n1502);
nand (n1503,n569,n1504);
or (n1504,1'b0,n1505,n1507,n1509,n1511);
and (n1505,n1506,n560);
and (n1507,n1508,n575);
and (n1509,n1510,n579);
and (n1511,n1502,n581);
and (n1512,n1513,n1514);
wire s0n1513,s1n1513,notn1513;
or (n1513,s0n1513,s1n1513);
not(notn1513,n639);
and (s0n1513,notn1513,1'b0);
and (s1n1513,n639,n1499);
or (n1514,n1515,n1531,n1641);
and (n1515,n1516,n1530);
wire s0n1516,s1n1516,notn1516;
or (n1516,s0n1516,s1n1516);
not(notn1516,n639);
and (s0n1516,notn1516,1'b0);
and (s1n1516,n639,n1517);
nand (n1517,n1518,n1521);
or (n1518,n1519,n19);
not (n1519,n1520);
nand (n1521,n569,n1522);
or (n1522,1'b0,n1523,n1525,n1527,n1529);
and (n1523,n1524,n560);
and (n1525,n1526,n575);
and (n1527,n1528,n579);
and (n1529,n1520,n581);
wire s0n1530,s1n1530,notn1530;
or (n1530,s0n1530,s1n1530);
not(notn1530,n584);
and (s0n1530,notn1530,1'b0);
and (s1n1530,n584,n1499);
and (n1531,n1530,n1532);
or (n1532,n1533,n1549,n1640);
and (n1533,n1534,n1548);
wire s0n1534,s1n1534,notn1534;
or (n1534,s0n1534,s1n1534);
not(notn1534,n639);
and (s0n1534,notn1534,1'b0);
and (s1n1534,n639,n1535);
nand (n1535,n1536,n1547);
or (n1536,n1537,n833);
not (n1537,n1538);
or (n1538,1'b0,n1539,n1541,n1543,n1545);
and (n1539,n1540,n560);
and (n1541,n1542,n575);
and (n1543,n1544,n579);
and (n1545,n1546,n581);
nand (n1547,n20,n1546);
wire s0n1548,s1n1548,notn1548;
or (n1548,s0n1548,s1n1548);
not(notn1548,n584);
and (s0n1548,notn1548,1'b0);
and (s1n1548,n584,n1517);
and (n1549,n1548,n1550);
or (n1550,n1551,n1567,n1639);
and (n1551,n1552,n1566);
wire s0n1552,s1n1552,notn1552;
or (n1552,s0n1552,s1n1552);
not(notn1552,n639);
and (s0n1552,notn1552,1'b0);
and (s1n1552,n639,n1553);
nand (n1553,n1554,n1565);
or (n1554,n1555,n833);
not (n1555,n1556);
or (n1556,1'b0,n1557,n1559,n1561,n1563);
and (n1557,n1558,n560);
and (n1559,n1560,n575);
and (n1561,n1562,n579);
and (n1563,n1564,n581);
nand (n1565,n20,n1564);
wire s0n1566,s1n1566,notn1566;
or (n1566,s0n1566,s1n1566);
not(notn1566,n584);
and (s0n1566,notn1566,1'b0);
and (s1n1566,n584,n1535);
and (n1567,n1566,n1568);
or (n1568,n1569,n1585,n1638);
and (n1569,n1570,n1584);
wire s0n1570,s1n1570,notn1570;
or (n1570,s0n1570,s1n1570);
not(notn1570,n639);
and (s0n1570,notn1570,1'b0);
and (s1n1570,n639,n1571);
nand (n1571,n1572,n1575);
or (n1572,n1573,n19);
not (n1573,n1574);
nand (n1575,n569,n1576);
or (n1576,1'b0,n1577,n1579,n1581,n1583);
and (n1577,n1578,n560);
and (n1579,n1580,n575);
and (n1581,n1582,n579);
and (n1583,n1574,n581);
wire s0n1584,s1n1584,notn1584;
or (n1584,s0n1584,s1n1584);
not(notn1584,n584);
and (s0n1584,notn1584,1'b0);
and (s1n1584,n584,n1553);
and (n1585,n1584,n1586);
or (n1586,n1587,n1603,n1605);
and (n1587,n1588,n1602);
wire s0n1588,s1n1588,notn1588;
or (n1588,s0n1588,s1n1588);
not(notn1588,n639);
and (s0n1588,notn1588,1'b0);
and (s1n1588,n639,n1589);
nand (n1589,n1590,n1601);
or (n1590,n1591,n833);
not (n1591,n1592);
or (n1592,1'b0,n1593,n1595,n1597,n1599);
and (n1593,n1594,n560);
and (n1595,n1596,n575);
and (n1597,n1598,n579);
and (n1599,n1600,n581);
nand (n1601,n20,n1600);
wire s0n1602,s1n1602,notn1602;
or (n1602,s0n1602,s1n1602);
not(notn1602,n584);
and (s0n1602,notn1602,1'b0);
and (s1n1602,n584,n1571);
and (n1603,n1602,n1604);
or (n1604,n1605,n1621,n1622);
and (n1605,n1606,n1620);
wire s0n1606,s1n1606,notn1606;
or (n1606,s0n1606,s1n1606);
not(notn1606,n639);
and (s0n1606,notn1606,1'b0);
and (s1n1606,n639,n1607);
nand (n1607,n1608,n1611);
or (n1608,n1609,n19);
not (n1609,n1610);
nand (n1611,n569,n1612);
or (n1612,1'b0,n1613,n1615,n1617,n1619);
and (n1613,n1614,n560);
and (n1615,n1616,n575);
and (n1617,n1618,n579);
and (n1619,n1610,n581);
wire s0n1620,s1n1620,notn1620;
or (n1620,s0n1620,s1n1620);
not(notn1620,n584);
and (s0n1620,notn1620,1'b0);
and (s1n1620,n584,n1589);
and (n1621,n1620,n1622);
and (n1622,n1623,n1637);
wire s0n1623,s1n1623,notn1623;
or (n1623,s0n1623,s1n1623);
not(notn1623,n639);
and (s0n1623,notn1623,1'b0);
and (s1n1623,n639,n1624);
nand (n1624,n1625,n1628);
or (n1625,n1626,n19);
not (n1626,n1627);
nand (n1628,n569,n1629);
or (n1629,1'b0,n1630,n1632,n1634,n1636);
and (n1630,n1631,n560);
and (n1632,n1633,n575);
and (n1634,n1635,n579);
and (n1636,n1627,n581);
wire s0n1637,s1n1637,notn1637;
or (n1637,s0n1637,s1n1637);
not(notn1637,n584);
and (s0n1637,notn1637,1'b0);
and (s1n1637,n584,n1607);
and (n1638,n1570,n1586);
and (n1639,n1552,n1568);
and (n1640,n1534,n1550);
and (n1641,n1516,n1532);
or (n1642,n1643,n1647,n1692);
and (n1643,n1644,n1646);
not (n1644,n1645);
nand (n1645,n686,n1517);
xor (n1646,n1513,n1514);
and (n1647,n1646,n1648);
or (n1648,n1649,n1654,n1691);
and (n1649,n1650,n1652);
not (n1650,n1651);
nand (n1651,n686,n1535);
xor (n1652,n1653,n1532);
xor (n1653,n1516,n1530);
and (n1654,n1652,n1655);
or (n1655,n1656,n1661,n1690);
and (n1656,n1657,n1659);
not (n1657,n1658);
nand (n1658,n686,n1553);
xor (n1659,n1660,n1550);
xor (n1660,n1534,n1548);
and (n1661,n1659,n1662);
or (n1662,n1663,n1668,n1689);
and (n1663,n1664,n1666);
not (n1664,n1665);
nand (n1665,n686,n1571);
xor (n1666,n1667,n1568);
xor (n1667,n1552,n1566);
and (n1668,n1666,n1669);
or (n1669,n1670,n1675,n1688);
and (n1670,n1671,n1673);
not (n1671,n1672);
nand (n1672,n686,n1589);
xor (n1673,n1674,n1586);
xor (n1674,n1570,n1584);
and (n1675,n1673,n1676);
or (n1676,n1677,n1682,n1687);
and (n1677,n1678,n1680);
not (n1678,n1679);
nand (n1679,n686,n1607);
xor (n1680,n1681,n1604);
xor (n1681,n1588,n1602);
and (n1682,n1680,n1683);
and (n1683,n1684,n1685);
and (n1684,n686,n1624);
xor (n1685,n1686,n1622);
xor (n1686,n1606,n1620);
and (n1687,n1678,n1683);
and (n1688,n1671,n1676);
and (n1689,n1664,n1669);
and (n1690,n1657,n1662);
and (n1691,n1650,n1655);
and (n1692,n1644,n1648);
nor (n1693,n1444,n1396,n934);
wire s0n1694,s1n1694,notn1694;
or (n1694,s0n1694,s1n1694);
not(notn1694,n1392);
and (s0n1694,notn1694,1'b0);
and (s1n1694,n1392,n1695);
or (n1695,n1696,n1697,n1698);
and (n1696,n1498,n1512);
and (n1697,n1512,n1642);
and (n1698,n1498,n1642);
wire s0n1699,s1n1699,notn1699;
or (n1699,s0n1699,s1n1699);
not(notn1699,n1693);
and (s0n1699,notn1699,1'b0);
and (s1n1699,n1693,n1700);
xor (n1700,n1701,n1334);
xor (n1701,n1200,n1216);
not (n1702,n1703);
xnor (n1703,n1704,n1705);
wire s0n1704,s1n1704,notn1704;
or (n1704,s0n1704,s1n1704);
not(notn1704,n1693);
and (s0n1704,notn1704,1'b0);
and (s1n1704,n1693,n1183);
wire s0n1705,s1n1705,notn1705;
or (n1705,s0n1705,s1n1705);
not(notn1705,n1693);
and (s0n1705,notn1705,1'b0);
and (s1n1705,n1693,n1695);
or (n1706,n1707,n1768);
and (n1707,n1708,n1767);
xor (n1708,n1709,n1766);
or (n1709,n1710,n1765);
and (n1710,n1711,n1764);
xor (n1711,n1712,n1758);
or (n1712,n1713,n1757);
and (n1713,n1714,n1754);
xor (n1714,n1715,n1751);
and (n1715,n1716,n1748);
xor (n1716,n1717,n1720);
wire s0n1717,s1n1717,notn1717;
or (n1717,s0n1717,s1n1717);
not(notn1717,n1693);
and (s0n1717,notn1717,1'b0);
and (s1n1717,n1693,n1718);
xor (n1718,n1719,n1662);
xor (n1719,n1657,n1659);
xor (n1720,n1721,n1728);
xor (n1721,n1722,n1727);
xor (n1722,n1723,n1726);
xor (n1723,n1724,n1725);
nor (n1724,n985,n1443);
and (n1725,n1498,n1444);
and (n1726,n1725,n1516);
and (n1727,n1724,n1003);
or (n1728,n1729,n1747);
and (n1729,n1730,n1739);
xor (n1730,n1731,n1734);
nor (n1731,n1732,n1443);
xnor (n1732,n1133,n1733);
not (n1733,n1000);
and (n1734,n1735,n1444);
nand (n1735,n1736,n1738);
or (n1736,n1737,n1644);
not (n1737,n1513);
or (n1738,n1645,n1513);
and (n1739,n1740,n1444);
or (n1740,n1741,n1745);
nor (n1741,n1742,n1744);
and (n1742,n1139,n1743);
not (n1743,n1017);
not (n1744,n1003);
nor (n1745,n1746,n985);
not (n1746,n1053);
and (n1747,n1731,n1734);
wire s0n1748,s1n1748,notn1748;
or (n1748,s0n1748,s1n1748);
not(notn1748,n1392);
and (s0n1748,notn1748,1'b0);
and (s1n1748,n1392,n1749);
xor (n1749,n1750,n1655);
xor (n1750,n1650,n1652);
wire s0n1751,s1n1751,notn1751;
or (n1751,s0n1751,s1n1751);
not(notn1751,n1392);
and (s0n1751,notn1751,1'b0);
and (s1n1751,n1392,n1752);
xor (n1752,n1753,n1648);
xor (n1753,n1644,n1646);
wire s0n1754,s1n1754,notn1754;
or (n1754,s0n1754,s1n1754);
not(notn1754,n934);
and (s0n1754,notn1754,1'b0);
and (s1n1754,n934,n1755);
xor (n1755,n1756,n1136);
xor (n1756,n1132,n1134);
and (n1757,n1715,n1751);
xor (n1758,n1759,n1763);
xor (n1759,n1760,n1762);
wire s0n1760,s1n1760,notn1760;
or (n1760,s0n1760,s1n1760);
not(notn1760,n1761);
and (s0n1760,notn1760,1'b0);
and (s1n1760,n1761,n1695);
xor (n1761,n1395,n1443);
wire s0n1762,s1n1762,notn1762;
or (n1762,s0n1762,s1n1762);
not(notn1762,n1693);
and (s0n1762,notn1762,1'b0);
and (s1n1762,n1693,n1752);
wire s0n1763,s1n1763,notn1763;
or (n1763,s0n1763,s1n1763);
not(notn1763,n1392);
and (s0n1763,notn1763,1'b0);
and (s1n1763,n1392,n1496);
wire s0n1764,s1n1764,notn1764;
or (n1764,s0n1764,s1n1764);
not(notn1764,n1396);
and (s0n1764,notn1764,1'b0);
and (s1n1764,n1396,n982);
and (n1765,n1712,n1758);
xor (n1766,n1494,n1699);
xor (n1767,n10,n1182);
and (n1768,n1709,n1766);
or (n1769,n1770,n1945);
and (n1770,n1771,n1934);
xor (n1771,n1772,n1819);
or (n1772,n1773,n1818);
and (n1773,n1774,n1811);
xor (n1774,n1775,n1790);
xor (n1775,n1776,n1787);
xor (n1776,n1777,n1780);
wire s0n1777,s1n1777,notn1777;
or (n1777,s0n1777,s1n1777);
not(notn1777,n1693);
and (s0n1777,notn1777,1'b0);
and (s1n1777,n1693,n1778);
xor (n1778,n1779,n1341);
xor (n1779,n1336,n1339);
and (n1780,n1781,n1784);
or (n1781,n1782,n1783);
and (n1782,n1721,n1728);
and (n1783,n1722,n1727);
or (n1784,n1785,n1786);
and (n1785,n1723,n1726);
and (n1786,n1724,n1725);
wire s0n1787,s1n1787,notn1787;
or (n1787,s0n1787,s1n1787);
not(notn1787,n934);
and (s0n1787,notn1787,1'b0);
and (s1n1787,n934,n1788);
xor (n1788,n1789,n1130);
xor (n1789,n984,n999);
or (n1790,n1791,n1810);
and (n1791,n1792,n1809);
xor (n1792,n1793,n1806);
or (n1793,n1794,n1805);
and (n1794,n1795,n1804);
xor (n1795,n1796,n1797);
xor (n1796,n1716,n1748);
and (n1797,n1798,n1803);
xor (n1798,n1799,n1802);
wire s0n1799,s1n1799,notn1799;
or (n1799,s0n1799,s1n1799);
not(notn1799,n1693);
and (s0n1799,notn1799,1'b0);
and (s1n1799,n1693,n1800);
xor (n1800,n1801,n1669);
xor (n1801,n1664,n1666);
wire s0n1802,s1n1802,notn1802;
or (n1802,s0n1802,s1n1802);
not(notn1802,n1392);
and (s0n1802,notn1802,1'b0);
and (s1n1802,n1392,n1718);
wire s0n1803,s1n1803,notn1803;
or (n1803,s0n1803,s1n1803);
not(notn1803,n1761);
and (s0n1803,notn1803,1'b0);
and (s1n1803,n1761,n1749);
wire s0n1804,s1n1804,notn1804;
or (n1804,s0n1804,s1n1804);
not(notn1804,n1396);
and (s0n1804,notn1804,1'b0);
and (s1n1804,n1396,n1755);
and (n1805,n1796,n1797);
wire s0n1806,s1n1806,notn1806;
or (n1806,s0n1806,s1n1806);
not(notn1806,n934);
and (s0n1806,notn1806,1'b0);
and (s1n1806,n934,n1807);
xor (n1807,n1808,n883);
xor (n1808,n878,n881);
wire s0n1809,s1n1809,notn1809;
or (n1809,s0n1809,s1n1809);
not(notn1809,n1392);
and (s0n1809,notn1809,1'b0);
and (s1n1809,n1392,n1778);
and (n1810,n1793,n1806);
or (n1811,n1812,n1817);
and (n1812,n1813,n1816);
xor (n1813,n1814,n1815);
wire s0n1814,s1n1814,notn1814;
or (n1814,s0n1814,s1n1814);
not(notn1814,n1444);
and (s0n1814,notn1814,1'b0);
and (s1n1814,n1444,n1183);
wire s0n1815,s1n1815,notn1815;
or (n1815,s0n1815,s1n1815);
not(notn1815,n1444);
and (s0n1815,notn1815,1'b0);
and (s1n1815,n1444,n13);
wire s0n1816,s1n1816,notn1816;
or (n1816,s0n1816,s1n1816);
not(notn1816,n1761);
and (s0n1816,notn1816,1'b0);
and (s1n1816,n1761,n1700);
and (n1817,n1814,n1815);
and (n1818,n1775,n1790);
and (n1819,n1820,n1833);
xor (n1820,n1821,n1832);
or (n1821,n1822,n1831);
and (n1822,n1823,n1828);
xor (n1823,n1824,n1825);
wire s0n1824,s1n1824,notn1824;
or (n1824,s0n1824,s1n1824);
not(notn1824,n1761);
and (s0n1824,notn1824,1'b0);
and (s1n1824,n1761,n1496);
xor (n1825,n1826,n1827);
xor (n1826,n1781,n1784);
wire s0n1827,s1n1827,notn1827;
or (n1827,s0n1827,s1n1827);
not(notn1827,n1693);
and (s0n1827,notn1827,1'b0);
and (s1n1827,n1693,n1749);
wire s0n1828,s1n1828,notn1828;
or (n1828,s0n1828,s1n1828);
not(notn1828,n1396);
and (s0n1828,notn1828,1'b0);
and (s1n1828,n1396,n1829);
xor (n1829,n1830,n876);
xor (n1830,n735,n756);
and (n1831,n1824,n1825);
wire s0n1832,s1n1832,notn1832;
or (n1832,s0n1832,s1n1832);
not(notn1832,n1396);
and (s0n1832,notn1832,1'b0);
and (s1n1832,n1396,n13);
and (n1833,n1834,n1933);
xor (n1834,n1835,n1887);
and (n1835,n1836,n1693);
xor (n1836,n1837,n1849);
nor (n1837,n1838,n1848);
not (n1838,n1839);
or (n1839,n1840,n1843);
xor (n1840,n1841,n1224);
xor (n1841,n1345,n1842);
xor (n1842,n1347,n1344);
or (n1843,n1844,n1847);
and (n1844,n1845,n1242);
xor (n1845,n1353,n1846);
xor (n1846,n1355,n1352);
and (n1847,n1353,n1846);
and (n1848,n1840,n1843);
nand (n1849,n1850,n1886);
or (n1850,n1851,n1859);
not (n1851,n1852);
or (n1852,n1853,n1854);
xor (n1853,n1845,n1242);
or (n1854,n1855,n1858);
and (n1855,n1856,n1260);
xor (n1856,n1361,n1857);
xor (n1857,n1363,n1360);
and (n1858,n1361,n1857);
not (n1859,n1860);
nand (n1860,n1861,n1882,n1885);
nand (n1861,n1862,n1869,n1879);
or (n1862,n1863,n1864);
xor (n1863,n1856,n1260);
or (n1864,n1865,n1868);
and (n1865,n1866,n1867);
xor (n1866,n1369,n1278);
xor (n1867,n1371,n1368);
and (n1868,n1369,n1278);
or (n1869,n1870,n1878);
and (n1870,n1871,n1876);
xor (n1871,n1296,n1872);
or (n1872,n1873,n1875);
and (n1873,n1874,n1384);
xor (n1874,n1313,n1382);
and (n1875,n1313,n1382);
xor (n1876,n1877,n1377);
xor (n1877,n1376,n1379);
and (n1878,n1296,n1872);
or (n1879,n1880,n1881);
xor (n1880,n1866,n1867);
and (n1881,n1877,n1377);
nand (n1882,n1883,n1862);
not (n1883,n1884);
nand (n1884,n1880,n1881);
nand (n1885,n1863,n1864);
nand (n1886,n1853,n1854);
or (n1887,n1888,n1932);
and (n1888,n1889,n1929);
xor (n1889,n1890,n1891);
wire s0n1890,s1n1890,notn1890;
or (n1890,s0n1890,s1n1890);
not(notn1890,n1761);
and (s0n1890,notn1890,1'b0);
and (s1n1890,n1761,n1752);
or (n1891,n1892,n1928);
and (n1892,n1893,n1904);
xor (n1893,n1894,n1895);
xor (n1894,n1730,n1739);
and (n1895,n1896,n1444);
nand (n1896,n1897,n1901);
or (n1897,n1898,n1900);
and (n1898,n1899,n1651);
not (n1899,n1530);
not (n1900,n1516);
or (n1901,n1902,n1903);
not (n1902,n1566);
not (n1903,n1498);
or (n1904,n1905,n1927);
and (n1905,n1906,n1921);
xor (n1906,n1907,n1914);
and (n1907,n1908,n1444);
nand (n1908,n1909,n1911,n1912);
or (n1909,n1651,n1910);
not (n1910,n1552);
not (n1911,n1533);
or (n1912,n1658,n1913);
not (n1913,n1548);
and (n1914,n1915,n1444);
nand (n1915,n1916,n1920);
or (n1916,n1917,n1146);
and (n1917,n1918,n1919);
not (n1918,n1021);
not (n1919,n1035);
not (n1920,n1020);
and (n1921,n1922,n1444);
nor (n1922,n1923,n1925);
and (n1923,n1924,n1516);
xor (n1924,n1899,n1651);
and (n1925,n1926,n1900);
not (n1926,n1924);
and (n1927,n1907,n1914);
and (n1928,n1894,n1895);
wire s0n1929,s1n1929,notn1929;
or (n1929,s0n1929,s1n1929);
not(notn1929,n934);
and (s0n1929,notn1929,1'b0);
and (s1n1929,n934,n1930);
xor (n1930,n1931,n1143);
xor (n1931,n1138,n1140);
and (n1932,n1890,n1891);
wire s0n1933,s1n1933,notn1933;
or (n1933,s0n1933,s1n1933);
not(notn1933,n1396);
and (s0n1933,notn1933,1'b0);
and (s1n1933,n1396,n1788);
xor (n1934,n1935,n1938);
xor (n1935,n1936,n1937);
and (n1936,n1776,n1787);
and (n1937,n1759,n1763);
or (n1938,n1939,n1944);
and (n1939,n1940,n1943);
xor (n1940,n1941,n1942);
wire s0n1941,s1n1941,notn1941;
or (n1941,s0n1941,s1n1941);
not(notn1941,n1761);
and (s0n1941,notn1941,1'b0);
and (s1n1941,n1761,n1183);
wire s0n1942,s1n1942,notn1942;
or (n1942,s0n1942,s1n1942);
not(notn1942,n934);
and (s0n1942,notn1942,1'b0);
and (s1n1942,n934,n1829);
wire s0n1943,s1n1943,notn1943;
or (n1943,s0n1943,s1n1943);
not(notn1943,n1392);
and (s0n1943,notn1943,1'b0);
and (s1n1943,n1392,n1700);
and (n1944,n1941,n1942);
and (n1945,n1772,n1819);
or (n1946,n1947,n2095);
and (n1947,n1948,n2021);
xor (n1948,n1949,n2020);
or (n1949,n1950,n2019);
and (n1950,n1951,n1954);
xor (n1951,n1952,n1953);
xor (n1952,n1940,n1943);
xor (n1953,n1711,n1764);
or (n1954,n1955,n2018);
and (n1955,n1956,n1967);
xor (n1956,n1957,n1966);
or (n1957,n1958,n1965);
and (n1958,n1959,n1964);
xor (n1959,n1960,n1961);
wire s0n1960,s1n1960,notn1960;
or (n1960,s0n1960,s1n1960);
not(notn1960,n1396);
and (s0n1960,notn1960,1'b0);
and (s1n1960,n1396,n1807);
wire s0n1961,s1n1961,notn1961;
or (n1961,s0n1961,s1n1961);
not(notn1961,n934);
and (s0n1961,notn1961,1'b0);
and (s1n1961,n934,n1962);
xor (n1962,n1963,n891);
xor (n1963,n885,n888);
and (n1964,n1836,n1392);
and (n1965,n1960,n1961);
xor (n1966,n1714,n1754);
and (n1967,n1968,n2017);
xor (n1968,n1969,n1972);
and (n1969,n1970,n1693);
xnor (n1970,n1860,n1971);
nand (n1971,n1852,n1886);
or (n1972,n1973,n2016);
and (n1973,n1974,n2007);
xor (n1974,n1975,n1978);
wire s0n1975,s1n1975,notn1975;
or (n1975,s0n1975,s1n1975);
not(notn1975,n934);
and (s0n1975,notn1975,1'b0);
and (s1n1975,n934,n1976);
xor (n1976,n1977,n1150);
xor (n1977,n1145,n1147);
and (n1978,n1979,n2001);
or (n1979,n1980,n2000);
and (n1980,n1981,n1993);
xor (n1981,n1982,n1989);
and (n1982,n1983,n1444);
nand (n1983,n1984,n1986,n1988);
or (n1984,n1985,n1139);
not (n1985,n1089);
or (n1986,n1146,n1987);
not (n1987,n1057);
not (n1988,n1038);
nor (n1989,n1443,n1990);
nor (n1990,n1551,n1991);
nor (n1991,n1992,n1665);
and (n1992,n1902,n1910);
nor (n1993,n1994,n1443);
nor (n1994,n1995,n1998);
and (n1995,n1996,n1534);
not (n1996,n1997);
xor (n1997,n1658,n1913);
and (n1998,n1997,n1999);
not (n1999,n1534);
and (n2000,n1982,n1989);
and (n2001,n2002,n1444);
nor (n2002,n2003,n2005);
and (n2003,n2004,n1003);
xor (n2004,n1139,n1743);
and (n2005,n2006,n1744);
not (n2006,n2004);
or (n2007,n2008,n2015);
and (n2008,n2009,n2012);
xor (n2009,n2010,n2011);
wire s0n2010,s1n2010,notn2010;
or (n2010,s0n2010,s1n2010);
not(notn2010,n1392);
and (s0n2010,notn2010,1'b0);
and (s1n2010,n1392,n1800);
xor (n2011,n1906,n1921);
wire s0n2012,s1n2012,notn2012;
or (n2012,s0n2012,s1n2012);
not(notn2012,n934);
and (s0n2012,notn2012,1'b0);
and (s1n2012,n934,n2013);
xor (n2013,n2014,n1156);
xor (n2014,n1152,n1153);
and (n2015,n2010,n2011);
and (n2016,n1975,n1978);
wire s0n2017,s1n2017,notn2017;
or (n2017,s0n2017,s1n2017);
not(notn2017,n1761);
and (s0n2017,notn2017,1'b0);
and (s1n2017,n1761,n1778);
and (n2018,n1957,n1966);
and (n2019,n1952,n1953);
xor (n2020,n1708,n1767);
or (n2021,n2022,n2094);
and (n2022,n2023,n2038);
xor (n2023,n2024,n2037);
or (n2024,n2025,n2036);
and (n2025,n2026,n2029);
xor (n2026,n2027,n2028);
xor (n2027,n1792,n1809);
xor (n2028,n1823,n1828);
or (n2029,n2030,n2035);
and (n2030,n2031,n2034);
xor (n2031,n2032,n2033);
wire s0n2032,s1n2032,notn2032;
or (n2032,s0n2032,s1n2032);
not(notn2032,n1444);
and (s0n2032,notn2032,1'b0);
and (s1n2032,n1444,n1829);
xor (n2033,n1889,n1929);
wire s0n2034,s1n2034,notn2034;
or (n2034,s0n2034,s1n2034);
not(notn2034,n1444);
and (s0n2034,notn2034,1'b0);
and (s1n2034,n1444,n1700);
and (n2035,n2032,n2033);
and (n2036,n2027,n2028);
xor (n2037,n1820,n1833);
or (n2038,n2039,n2093);
and (n2039,n2040,n2092);
xor (n2040,n2041,n2042);
xor (n2041,n1834,n1933);
or (n2042,n2043,n2091);
and (n2043,n2044,n2080);
xor (n2044,n2045,n2046);
xor (n2045,n1795,n1804);
or (n2046,n2047,n2079);
and (n2047,n2048,n2078);
xor (n2048,n2049,n2077);
or (n2049,n2050,n2076);
and (n2050,n2051,n2075);
xor (n2051,n2052,n2053);
wire s0n2052,s1n2052,notn2052;
or (n2052,s0n2052,s1n2052);
not(notn2052,n1761);
and (s0n2052,notn2052,1'b0);
and (s1n2052,n1761,n1718);
or (n2053,n2054,n2074);
and (n2054,n2055,n2071);
xor (n2055,n2056,n2069);
or (n2056,n2057,n2064);
and (n2057,n2058,n1444);
nand (n2058,n2059,n2061,n2063);
or (n2059,n1658,n2060);
not (n2060,n1620);
or (n2061,n1665,n2062);
not (n2062,n1588);
not (n2063,n1569);
and (n2064,n2065,n1444);
or (n2065,n2066,n1056);
nor (n2066,n2067,n1159);
and (n2067,n2068,n1987);
not (n2068,n1071);
nor (n2069,n2070,n1443);
xor (n2070,n1148,n1146);
wire s0n2071,s1n2071,notn2071;
or (n2071,s0n2071,s1n2071);
not(notn2071,n1392);
and (s0n2071,notn2071,1'b0);
and (s1n2071,n1392,n2072);
xor (n2072,n2073,n1676);
xor (n2073,n1671,n1673);
and (n2074,n2056,n2069);
wire s0n2075,s1n2075,notn2075;
or (n2075,s0n2075,s1n2075);
not(notn2075,n1396);
and (s0n2075,notn2075,1'b0);
and (s1n2075,n1396,n1976);
and (n2076,n2052,n2053);
xor (n2077,n1893,n1904);
wire s0n2078,s1n2078,notn2078;
or (n2078,s0n2078,s1n2078);
not(notn2078,n1396);
and (s0n2078,notn2078,1'b0);
and (s1n2078,n1396,n1930);
and (n2079,n2049,n2077);
or (n2080,n2081,n2090);
and (n2081,n2082,n2087);
xor (n2082,n2083,n2086);
wire s0n2083,s1n2083,notn2083;
or (n2083,s0n2083,s1n2083);
not(notn2083,n1693);
and (s0n2083,notn2083,1'b0);
and (s1n2083,n1693,n2084);
xor (n2084,n2085,n1365);
xor (n2085,n1359,n1362);
xor (n2086,n1798,n1803);
wire s0n2087,s1n2087,notn2087;
or (n2087,s0n2087,s1n2087);
not(notn2087,n934);
and (s0n2087,notn2087,1'b0);
and (s1n2087,n934,n2088);
xor (n2088,n2089,n899);
xor (n2089,n893,n896);
and (n2090,n2083,n2086);
and (n2091,n2045,n2046);
xor (n2092,n1813,n1816);
and (n2093,n2041,n2042);
and (n2094,n2024,n2037);
and (n2095,n1949,n2020);
or (n2096,n2097,n2251);
and (n2097,n2098,n2250);
xor (n2098,n2099,n2249);
or (n2099,n2100,n2248);
and (n2100,n2101,n2104);
xor (n2101,n2102,n2103);
xor (n2102,n1951,n1954);
xor (n2103,n1774,n1811);
or (n2104,n2105,n2247);
and (n2105,n2106,n2145);
xor (n2106,n2107,n2108);
xor (n2107,n1956,n1967);
or (n2108,n2109,n2144);
and (n2109,n2110,n2119);
xor (n2110,n2111,n2112);
xor (n2111,n1968,n2017);
or (n2112,n2113,n2118);
and (n2113,n2114,n2117);
xor (n2114,n2115,n2116);
and (n2115,n1970,n1392);
xor (n2116,n1974,n2007);
wire s0n2117,s1n2117,notn2117;
or (n2117,s0n2117,s1n2117);
not(notn2117,n1444);
and (s0n2117,notn2117,1'b0);
and (s1n2117,n1444,n1807);
and (n2118,n2115,n2116);
or (n2119,n2120,n2143);
and (n2120,n2121,n2142);
xor (n2121,n2122,n2123);
wire s0n2122,s1n2122,notn2122;
or (n2122,s0n2122,s1n2122);
not(notn2122,n1396);
and (s0n2122,notn2122,1'b0);
and (s1n2122,n1396,n1962);
or (n2123,n2124,n2141);
and (n2124,n2125,n2138);
xor (n2125,n2126,n2129);
xor (n2126,n2127,n2128);
xor (n2127,n1979,n2001);
wire s0n2128,s1n2128,notn2128;
or (n2128,s0n2128,s1n2128);
not(notn2128,n1693);
and (s0n2128,notn2128,1'b0);
and (s1n2128,n1693,n2072);
and (n2129,n2130,n2135);
xor (n2130,n2131,n2132);
xor (n2131,n1981,n1993);
wire s0n2132,s1n2132,notn2132;
or (n2132,s0n2132,s1n2132);
not(notn2132,n1693);
and (s0n2132,notn2132,1'b0);
and (s1n2132,n1693,n2133);
xor (n2133,n2134,n1683);
xor (n2134,n1678,n1680);
wire s0n2135,s1n2135,notn2135;
or (n2135,s0n2135,s1n2135);
not(notn2135,n934);
and (s0n2135,notn2135,1'b0);
and (s1n2135,n934,n2136);
xor (n2136,n2137,n1163);
xor (n2137,n1158,n1160);
wire s0n2138,s1n2138,notn2138;
or (n2138,s0n2138,s1n2138);
not(notn2138,n1693);
and (s0n2138,notn2138,1'b0);
and (s1n2138,n1693,n2139);
xor (n2139,n2140,n1373);
xor (n2140,n1367,n1370);
and (n2141,n2126,n2129);
and (n2142,n1836,n1761);
and (n2143,n2122,n2123);
and (n2144,n2111,n2112);
or (n2145,n2146,n2246);
and (n2146,n2147,n2245);
xor (n2147,n2148,n2244);
or (n2148,n2149,n2243);
and (n2149,n2150,n2242);
xor (n2150,n2151,n2184);
or (n2151,n2152,n2183);
and (n2152,n2153,n2180);
xor (n2153,n2154,n2155);
xor (n2154,n2009,n2012);
or (n2155,n2156,n2179);
and (n2156,n2157,n2178);
xor (n2157,n2158,n2159);
wire s0n2158,s1n2158,notn2158;
or (n2158,s0n2158,s1n2158);
not(notn2158,n1761);
and (s0n2158,notn2158,1'b0);
and (s1n2158,n1761,n1800);
or (n2159,n2160,n2177);
and (n2160,n2161,n2176);
xor (n2161,n2162,n2172);
and (n2162,n2163,n1444);
nand (n2163,n2164,n2170);
or (n2164,n1039,n2165);
not (n2165,n2166);
nand (n2166,n2167,n2169);
or (n2167,n1053,n2168);
not (n2168,n1152);
or (n2169,n1152,n1746);
or (n2170,n2166,n2171);
not (n2171,n1039);
and (n2172,n2173,n1444);
nand (n2173,n2174,n2175);
or (n2174,n1665,n1667);
nand (n2175,n1667,n1665);
wire s0n2176,s1n2176,notn2176;
or (n2176,s0n2176,s1n2176);
not(notn2176,n1392);
and (s0n2176,notn2176,1'b0);
and (s1n2176,n1392,n2133);
and (n2177,n2162,n2172);
wire s0n2178,s1n2178,notn2178;
or (n2178,s0n2178,s1n2178);
not(notn2178,n1396);
and (s0n2178,notn2178,1'b0);
and (s1n2178,n1396,n2013);
and (n2179,n2158,n2159);
wire s0n2180,s1n2180,notn2180;
or (n2180,s0n2180,s1n2180);
not(notn2180,n934);
and (s0n2180,notn2180,1'b0);
and (s1n2180,n934,n2181);
xor (n2181,n2182,n907);
xor (n2182,n901,n904);
and (n2183,n2154,n2155);
or (n2184,n2185,n2241);
and (n2185,n2186,n2240);
xor (n2186,n2187,n2188);
xor (n2187,n2051,n2075);
and (n2188,n2189,n2239);
xor (n2189,n2190,n2233);
or (n2190,n2191,n2232);
and (n2191,n2192,n2229);
xor (n2192,n2193,n2207);
and (n2193,n2194,n2205);
xor (n2194,n2195,n2203);
and (n2195,n2196,n2200);
nor (n2196,n2197,n1159);
not (n2197,n2198);
wire s0n2198,s1n2198,notn2198;
or (n2198,s0n2198,s1n2198);
not(notn2198,n1444);
and (s0n2198,notn2198,1'b0);
and (s1n2198,n1444,n2199);
wire s0n2199,s1n2199,notn2199;
or (n2199,s0n2199,s1n2199);
not(notn2199,n584);
and (s0n2199,notn2199,1'b0);
and (s1n2199,n584,n1111);
and (n2200,n2201,n1444);
nor (n2201,n2202,n2060);
not (n2202,n1684);
wire s0n2203,s1n2203,notn2203;
or (n2203,s0n2203,s1n2203);
not(notn2203,n1693);
and (s0n2203,notn2203,1'b0);
and (s1n2203,n1693,n2204);
xor (n2204,n1623,n1637);
and (n2205,n2206,n1444);
xnor (n2206,n1159,n1161);
or (n2207,n2208,n2228);
and (n2208,n2209,n2223);
xor (n2209,n2210,n2216);
and (n2210,n2211,n1444);
nand (n2211,n2212,n2213,n2215);
or (n2212,n1679,n2062);
or (n2213,n1665,n2214);
not (n2214,n1637);
not (n2215,n1587);
and (n2216,n2217,n1444);
not (n2217,n2218);
nor (n2218,n2219,n2220);
and (n2219,n1158,n1093);
nor (n2220,n2221,n1985);
and (n2221,n1166,n2222);
not (n2222,n1075);
and (n2223,n2224,n1444);
xor (n2224,n2225,n2226);
not (n2225,n1570);
xnor (n2226,n1672,n2227);
not (n2227,n1584);
and (n2228,n2210,n2216);
wire s0n2229,s1n2229,notn2229;
or (n2229,s0n2229,s1n2229);
not(notn2229,n934);
and (s0n2229,notn2229,1'b0);
and (s1n2229,n934,n2230);
xor (n2230,n2231,n1170);
xor (n2231,n1165,n1167);
and (n2232,n2193,n2207);
and (n2233,n2234,n2238);
xor (n2234,n2235,n2236);
wire s0n2235,s1n2235,notn2235;
or (n2235,s0n2235,s1n2235);
not(notn2235,n1396);
and (s0n2235,notn2235,1'b0);
and (s1n2235,n1396,n2136);
wire s0n2236,s1n2236,notn2236;
or (n2236,s0n2236,s1n2236);
not(notn2236,n1693);
and (s0n2236,notn2236,1'b0);
and (s1n2236,n1693,n2237);
xor (n2237,n1684,n1685);
wire s0n2238,s1n2238,notn2238;
or (n2238,s0n2238,s1n2238);
not(notn2238,n1761);
and (s0n2238,notn2238,1'b0);
and (s1n2238,n1761,n2072);
xor (n2239,n2130,n2135);
wire s0n2240,s1n2240,notn2240;
or (n2240,s0n2240,s1n2240);
not(notn2240,n1392);
and (s0n2240,notn2240,1'b0);
and (s1n2240,n1392,n2084);
and (n2241,n2187,n2188);
wire s0n2242,s1n2242,notn2242;
or (n2242,s0n2242,s1n2242);
not(notn2242,n1444);
and (s0n2242,notn2242,1'b0);
and (s1n2242,n1444,n1778);
and (n2243,n2151,n2184);
xor (n2244,n1959,n1964);
xor (n2245,n2031,n2034);
and (n2246,n2148,n2244);
and (n2247,n2107,n2108);
and (n2248,n2102,n2103);
xor (n2249,n1771,n1934);
xor (n2250,n1948,n2021);
and (n2251,n2099,n2249);
or (n2252,n2253,n0);
or (n2253,n2254,n2805);
and (n2254,n2255,n2330);
xor (n2255,n2256,n2257);
xor (n2256,n2098,n2250);
or (n2257,n2258,n2329);
and (n2258,n2259,n2328);
xor (n2259,n2260,n2261);
xor (n2260,n2023,n2038);
or (n2261,n2262,n2327);
and (n2262,n2263,n2266);
xor (n2263,n2264,n2265);
xor (n2264,n2040,n2092);
xor (n2265,n2026,n2029);
or (n2266,n2267,n2326);
and (n2267,n2268,n2313);
xor (n2268,n2269,n2312);
or (n2269,n2270,n2311);
and (n2270,n2271,n2274);
xor (n2271,n2272,n2273);
xor (n2272,n2082,n2087);
xor (n2273,n2048,n2078);
or (n2274,n2275,n2310);
and (n2275,n2276,n2309);
xor (n2276,n2277,n2300);
or (n2277,n2278,n2299);
and (n2278,n2279,n2298);
xor (n2279,n2280,n2281);
xor (n2280,n2157,n2178);
or (n2281,n2282,n2297);
and (n2282,n2283,n2289);
xor (n2283,n2284,n2285);
xor (n2284,n2161,n2176);
nand (n2285,n2286,n2056);
or (n2286,n2287,n2288);
not (n2287,n2064);
not (n2288,n2057);
or (n2289,n2290,n2296);
and (n2290,n2291,n2295);
xor (n2291,n2292,n2293);
wire s0n2292,s1n2292,notn2292;
or (n2292,s0n2292,s1n2292);
not(notn2292,n1392);
and (s0n2292,notn2292,1'b0);
and (s1n2292,n1392,n2237);
wire s0n2293,s1n2293,notn2293;
or (n2293,s0n2293,s1n2293);
not(notn2293,n934);
and (s0n2293,notn2293,1'b0);
and (s1n2293,n934,n2294);
xor (n2294,n1171,n1173);
wire s0n2295,s1n2295,notn2295;
or (n2295,s0n2295,s1n2295);
not(notn2295,n1761);
and (s0n2295,notn2295,1'b0);
and (s1n2295,n1761,n2133);
and (n2296,n2292,n2293);
and (n2297,n2284,n2285);
wire s0n2298,s1n2298,notn2298;
or (n2298,s0n2298,s1n2298);
not(notn2298,n1392);
and (s0n2298,notn2298,1'b0);
and (s1n2298,n1392,n2139);
and (n2299,n2280,n2281);
and (n2300,n2301,n2306);
xor (n2301,n2302,n2305);
wire s0n2302,s1n2302,notn2302;
or (n2302,s0n2302,s1n2302);
not(notn2302,n1693);
and (s0n2302,notn2302,1'b0);
and (s1n2302,n1693,n2303);
xor (n2303,n2304,n1381);
xor (n2304,n1375,n1378);
xor (n2305,n2055,n2071);
wire s0n2306,s1n2306,notn2306;
or (n2306,s0n2306,s1n2306);
not(notn2306,n934);
and (s0n2306,notn2306,1'b0);
and (s1n2306,n934,n2307);
xor (n2307,n2308,n915);
xor (n2308,n909,n912);
wire s0n2309,s1n2309,notn2309;
or (n2309,s0n2309,s1n2309);
not(notn2309,n1444);
and (s0n2309,notn2309,1'b0);
and (s1n2309,n1444,n1962);
and (n2310,n2277,n2300);
and (n2311,n2272,n2273);
xor (n2312,n2044,n2080);
or (n2313,n2314,n2325);
and (n2314,n2315,n2324);
xor (n2315,n2316,n2317);
xor (n2316,n2114,n2117);
or (n2317,n2318,n2323);
and (n2318,n2319,n2322);
xor (n2319,n2320,n2321);
and (n2320,n1970,n1761);
wire s0n2321,s1n2321,notn2321;
or (n2321,s0n2321,s1n2321);
not(notn2321,n1396);
and (s0n2321,notn2321,1'b0);
and (s1n2321,n1396,n2088);
and (n2322,n1836,n1444);
and (n2323,n2320,n2321);
xor (n2324,n2121,n2142);
and (n2325,n2316,n2317);
and (n2326,n2269,n2312);
and (n2327,n2264,n2265);
xor (n2328,n2101,n2104);
and (n2329,n2260,n2261);
or (n2330,n2331,n2804);
and (n2331,n2332,n2409);
xor (n2332,n2333,n2334);
xor (n2333,n2259,n2328);
or (n2334,n2335,n2408);
and (n2335,n2336,n2407);
xor (n2336,n2337,n2338);
xor (n2337,n2106,n2145);
or (n2338,n2339,n2406);
and (n2339,n2340,n2343);
xor (n2340,n2341,n2342);
xor (n2341,n2110,n2119);
xor (n2342,n2147,n2245);
or (n2343,n2344,n2405);
and (n2344,n2345,n2384);
xor (n2345,n2346,n2347);
xor (n2346,n2150,n2242);
or (n2347,n2348,n2383);
and (n2348,n2349,n2352);
xor (n2349,n2350,n2351);
xor (n2350,n2153,n2180);
xor (n2351,n2125,n2138);
or (n2352,n2353,n2382);
and (n2353,n2354,n2381);
xor (n2354,n2355,n2380);
and (n2355,n2356,n2357);
xor (n2356,n2192,n2229);
or (n2357,n2358,n2379);
and (n2358,n2359,n2378);
xor (n2359,n2360,n2377);
or (n2360,n2361,n2376);
and (n2361,n2362,n2369);
xor (n2362,n2363,n2365);
wire s0n2363,s1n2363,notn2363;
or (n2363,s0n2363,s1n2363);
not(notn2363,n934);
and (s0n2363,notn2363,1'b0);
and (s1n2363,n934,n2364);
xor (n2364,n1110,n1124);
and (n2365,n2366,n2367);
wire s0n2366,s1n2366,notn2366;
or (n2366,s0n2366,s1n2366);
not(notn2366,n934);
and (s0n2366,notn2366,1'b0);
and (s1n2366,n934,n2199);
wire s0n2367,s1n2367,notn2367;
or (n2367,s0n2367,s1n2367);
not(notn2367,n934);
and (s0n2367,notn2367,1'b0);
and (s1n2367,n934,n2368);
wire s0n2368,s1n2368,notn2368;
or (n2368,s0n2368,s1n2368);
not(notn2368,n584);
and (s0n2368,notn2368,1'b0);
and (s1n2368,n584,n857);
and (n2369,n2370,n1444);
nand (n2370,n2371,n2375);
or (n2371,n2222,n2372);
nand (n2372,n2373,n2374);
or (n2373,n1089,n1166);
nand (n2374,n1089,n1166);
nand (n2375,n2372,n2222);
and (n2376,n2363,n2365);
xor (n2377,n2209,n2223);
wire s0n2378,s1n2378,notn2378;
or (n2378,s0n2378,s1n2378);
not(notn2378,n1396);
and (s0n2378,notn2378,1'b0);
and (s1n2378,n1396,n2230);
and (n2379,n2360,n2377);
wire s0n2380,s1n2380,notn2380;
or (n2380,s0n2380,s1n2380);
not(notn2380,n1761);
and (s0n2380,notn2380,1'b0);
and (s1n2380,n1761,n2084);
wire s0n2381,s1n2381,notn2381;
or (n2381,s0n2381,s1n2381);
not(notn2381,n1396);
and (s0n2381,notn2381,1'b0);
and (s1n2381,n1396,n2181);
and (n2382,n2355,n2380);
and (n2383,n2350,n2351);
or (n2384,n2385,n2404);
and (n2385,n2386,n2403);
xor (n2386,n2387,n2388);
xor (n2387,n2186,n2240);
or (n2388,n2389,n2402);
and (n2389,n2390,n2401);
xor (n2390,n2391,n2400);
or (n2391,n2392,n2399);
and (n2392,n2393,n2398);
xor (n2393,n2394,n2395);
xor (n2394,n2234,n2238);
wire s0n2395,s1n2395,notn2395;
or (n2395,s0n2395,s1n2395);
not(notn2395,n934);
and (s0n2395,notn2395,1'b0);
and (s1n2395,n934,n2396);
xor (n2396,n2397,n923);
xor (n2397,n917,n920);
wire s0n2398,s1n2398,notn2398;
or (n2398,s0n2398,s1n2398);
not(notn2398,n1392);
and (s0n2398,notn2398,1'b0);
and (s1n2398,n1392,n2303);
and (n2399,n2394,n2395);
xor (n2400,n2189,n2239);
and (n2401,n1970,n1444);
and (n2402,n2391,n2400);
xor (n2403,n2319,n2322);
and (n2404,n2387,n2388);
and (n2405,n2346,n2347);
and (n2406,n2341,n2342);
xor (n2407,n2263,n2266);
and (n2408,n2337,n2338);
or (n2409,n2410,n2803);
and (n2410,n2411,n2541);
xor (n2411,n2412,n2413);
xor (n2412,n2336,n2407);
or (n2413,n2414,n2540);
and (n2414,n2415,n2539);
xor (n2415,n2416,n2417);
xor (n2416,n2268,n2313);
or (n2417,n2418,n2538);
and (n2418,n2419,n2537);
xor (n2419,n2420,n2421);
xor (n2420,n2271,n2274);
or (n2421,n2422,n2536);
and (n2422,n2423,n2468);
xor (n2423,n2424,n2467);
or (n2424,n2425,n2466);
and (n2425,n2426,n2429);
xor (n2426,n2427,n2428);
xor (n2427,n2301,n2306);
wire s0n2428,s1n2428,notn2428;
or (n2428,s0n2428,s1n2428);
not(notn2428,n1444);
and (s0n2428,notn2428,1'b0);
and (s1n2428,n1444,n2088);
or (n2429,n2430,n2465);
and (n2430,n2431,n2464);
xor (n2431,n2432,n2446);
or (n2432,n2433,n2445);
and (n2433,n2434,n2443);
xor (n2434,n2435,n2437);
wire s0n2435,s1n2435,notn2435;
or (n2435,s0n2435,s1n2435);
not(notn2435,n934);
and (s0n2435,notn2435,1'b0);
and (s1n2435,n934,n2436);
xor (n2436,n924,n925);
and (n2437,n2438,n2442);
xor (n2438,n2439,n2440);
xor (n2439,n2196,n2200);
wire s0n2440,s1n2440,notn2440;
or (n2440,s0n2440,s1n2440);
not(notn2440,n1693);
and (s0n2440,notn2440,1'b0);
and (s1n2440,n1693,n2441);
wire s0n2441,s1n2441,notn2441;
or (n2441,s0n2441,s1n2441);
not(notn2441,n584);
and (s0n2441,notn2441,1'b0);
and (s1n2441,n584,n1624);
wire s0n2442,s1n2442,notn2442;
or (n2442,s0n2442,s1n2442);
not(notn2442,n1396);
and (s0n2442,notn2442,1'b0);
and (s1n2442,n1396,n2294);
wire s0n2443,s1n2443,notn2443;
or (n2443,s0n2443,s1n2443);
not(notn2443,n1392);
and (s0n2443,notn2443,1'b0);
and (s1n2443,n1392,n2444);
xor (n2444,n1382,n1383);
and (n2445,n2435,n2437);
or (n2446,n2447,n2463);
and (n2447,n2448,n2461);
xor (n2448,n2449,n2450);
xor (n2449,n2194,n2205);
and (n2450,n2451,n2460);
xor (n2451,n2452,n2458);
and (n2452,n2453,n1444);
xnor (n2453,n2454,n2062);
nand (n2454,n2455,n2457);
or (n2455,n1678,n2456);
not (n2456,n1602);
nand (n2457,n1678,n2456);
wire s0n2458,s1n2458,notn2458;
or (n2458,s0n2458,s1n2458);
not(notn2458,n1693);
and (s0n2458,notn2458,1'b0);
and (s1n2458,n1693,n2459);
wire s0n2459,s1n2459,notn2459;
or (n2459,s0n2459,s1n2459);
not(notn2459,n584);
and (s0n2459,notn2459,1'b0);
and (s1n2459,n584,n1315);
wire s0n2460,s1n2460,notn2460;
or (n2460,s0n2460,s1n2460);
not(notn2460,n1392);
and (s0n2460,notn2460,1'b0);
and (s1n2460,n1392,n2204);
wire s0n2461,s1n2461,notn2461;
or (n2461,s0n2461,s1n2461);
not(notn2461,n1693);
and (s0n2461,notn2461,1'b0);
and (s1n2461,n1693,n2462);
xor (n2462,n1314,n1328);
and (n2463,n2449,n2450);
wire s0n2464,s1n2464,notn2464;
or (n2464,s0n2464,s1n2464);
not(notn2464,n1761);
and (s0n2464,notn2464,1'b0);
and (s1n2464,n1761,n2139);
and (n2465,n2432,n2446);
and (n2466,n2427,n2428);
xor (n2467,n2276,n2309);
or (n2468,n2469,n2535);
and (n2469,n2470,n2534);
xor (n2470,n2471,n2533);
or (n2471,n2472,n2532);
and (n2472,n2473,n2531);
xor (n2473,n2474,n2475);
xor (n2474,n2283,n2289);
or (n2475,n2476,n2530);
and (n2476,n2477,n2505);
xor (n2477,n2478,n2479);
xor (n2478,n2291,n2295);
or (n2479,n2480,n2504);
and (n2480,n2481,n2503);
xor (n2481,n2482,n2492);
or (n2482,n2483,n2491);
and (n2483,n2484,n2487);
xor (n2484,n2485,n2486);
wire s0n2485,s1n2485,notn2485;
or (n2485,s0n2485,s1n2485);
not(notn2485,n1396);
and (s0n2485,notn2485,1'b0);
and (s1n2485,n1396,n2364);
xor (n2486,n2366,n2367);
and (n2487,n2488,n1444);
nand (n2488,n2489,n2490);
or (n2489,n1620,n2202);
or (n2490,n1684,n2060);
and (n2491,n2485,n2486);
or (n2492,n2493,n2502);
and (n2493,n2494,n2497);
xor (n2494,n2495,n2496);
and (n2495,n1606,n1444);
and (n2496,n1093,n1444);
and (n2497,n2498,n1444);
nand (n2498,n2499,n2501);
or (n2499,n1171,n2500);
not (n2500,n1107);
nand (n2501,n1171,n2500);
and (n2502,n2495,n2496);
wire s0n2503,s1n2503,notn2503;
or (n2503,s0n2503,s1n2503);
not(notn2503,n1761);
and (s0n2503,notn2503,1'b0);
and (s1n2503,n1761,n2237);
and (n2504,n2482,n2492);
or (n2505,n2506,n2529);
and (n2506,n2507,n2527);
xor (n2507,n2508,n2509);
xor (n2508,n2362,n2369);
or (n2509,n2510,n2526);
and (n2510,n2511,n2525);
xor (n2511,n2512,n2520);
or (n2512,n2513,n2519);
and (n2513,n2514,n2517);
xor (n2514,n2515,n2516);
nor (n2515,n2214,n1443);
wire s0n2516,s1n2516,notn2516;
or (n2516,s0n2516,s1n2516);
not(notn2516,n1396);
and (s0n2516,notn2516,1'b0);
and (s1n2516,n1396,n2199);
nor (n2517,n2518,n1443);
not (n2518,n1124);
and (n2519,n2515,n2516);
and (n2520,n2521,n2523);
nor (n2521,n2522,n1443);
not (n2522,n1623);
nor (n2523,n2524,n1443);
not (n2524,n1110);
wire s0n2525,s1n2525,notn2525;
or (n2525,s0n2525,s1n2525);
not(notn2525,n1392);
and (s0n2525,notn2525,1'b0);
and (s1n2525,n1392,n2459);
and (n2526,n2512,n2520);
wire s0n2527,s1n2527,notn2527;
or (n2527,s0n2527,s1n2527);
not(notn2527,n934);
and (s0n2527,notn2527,1'b0);
and (s1n2527,n934,n2528);
xor (n2528,n856,n870);
and (n2529,n2508,n2509);
and (n2530,n2478,n2479);
wire s0n2531,s1n2531,notn2531;
or (n2531,s0n2531,s1n2531);
not(notn2531,n1396);
and (s0n2531,notn2531,1'b0);
and (s1n2531,n1396,n2307);
and (n2532,n2474,n2475);
xor (n2533,n2279,n2298);
xor (n2534,n2354,n2381);
and (n2535,n2471,n2533);
and (n2536,n2424,n2467);
xor (n2537,n2315,n2324);
and (n2538,n2420,n2421);
xor (n2539,n2340,n2343);
and (n2540,n2416,n2417);
or (n2541,n2542,n2802);
and (n2542,n2543,n2602);
xor (n2543,n2544,n2545);
xor (n2544,n2415,n2539);
or (n2545,n2546,n2601);
and (n2546,n2547,n2600);
xor (n2547,n2548,n2549);
xor (n2548,n2345,n2384);
or (n2549,n2550,n2599);
and (n2550,n2551,n2598);
xor (n2551,n2552,n2553);
xor (n2552,n2349,n2352);
or (n2553,n2554,n2597);
and (n2554,n2555,n2596);
xor (n2555,n2556,n2565);
or (n2556,n2557,n2564);
and (n2557,n2558,n2563);
xor (n2558,n2559,n2562);
xor (n2559,n2560,n2561);
xor (n2560,n2356,n2357);
wire s0n2561,s1n2561,notn2561;
or (n2561,s0n2561,s1n2561);
not(notn2561,n1693);
and (s0n2561,notn2561,1'b0);
and (s1n2561,n1693,n2444);
wire s0n2562,s1n2562,notn2562;
or (n2562,s0n2562,s1n2562);
not(notn2562,n1444);
and (s0n2562,notn2562,1'b0);
and (s1n2562,n1444,n2084);
wire s0n2563,s1n2563,notn2563;
or (n2563,s0n2563,s1n2563);
not(notn2563,n1444);
and (s0n2563,notn2563,1'b0);
and (s1n2563,n1444,n2181);
and (n2564,n2559,n2562);
or (n2565,n2566,n2595);
and (n2566,n2567,n2588);
xor (n2567,n2568,n2587);
or (n2568,n2569,n2586);
and (n2569,n2570,n2585);
xor (n2570,n2571,n2572);
xor (n2571,n2448,n2461);
or (n2572,n2573,n2584);
and (n2573,n2574,n2583);
xor (n2574,n2575,n2576);
wire s0n2575,s1n2575,notn2575;
or (n2575,s0n2575,s1n2575);
not(notn2575,n1392);
and (s0n2575,notn2575,1'b0);
and (s1n2575,n1392,n2462);
or (n2576,n2577,n2582);
and (n2577,n2578,n2581);
xor (n2578,n2579,n2580);
xor (n2579,n2494,n2497);
wire s0n2580,s1n2580,notn2580;
or (n2580,s0n2580,s1n2580);
not(notn2580,n1761);
and (s0n2580,notn2580,1'b0);
and (s1n2580,n1761,n2204);
wire s0n2581,s1n2581,notn2581;
or (n2581,s0n2581,s1n2581);
not(notn2581,n1392);
and (s0n2581,notn2581,1'b0);
and (s1n2581,n1392,n2441);
and (n2582,n2579,n2580);
xor (n2583,n2438,n2442);
and (n2584,n2575,n2576);
wire s0n2585,s1n2585,notn2585;
or (n2585,s0n2585,s1n2585);
not(notn2585,n1761);
and (s0n2585,notn2585,1'b0);
and (s1n2585,n1761,n2303);
and (n2586,n2571,n2572);
xor (n2587,n2393,n2398);
or (n2588,n2589,n2594);
and (n2589,n2590,n2593);
xor (n2590,n2591,n2592);
wire s0n2591,s1n2591,notn2591;
or (n2591,s0n2591,s1n2591);
not(notn2591,n1396);
and (s0n2591,notn2591,1'b0);
and (s1n2591,n1396,n2396);
xor (n2592,n2359,n2378);
wire s0n2593,s1n2593,notn2593;
or (n2593,s0n2593,s1n2593);
not(notn2593,n1444);
and (s0n2593,notn2593,1'b0);
and (s1n2593,n1444,n2139);
and (n2594,n2591,n2592);
and (n2595,n2568,n2587);
xor (n2596,n2390,n2401);
and (n2597,n2556,n2565);
xor (n2598,n2386,n2403);
and (n2599,n2552,n2553);
xor (n2600,n2419,n2537);
and (n2601,n2548,n2549);
or (n2602,n2603,n2801);
and (n2603,n2604,n2637);
xor (n2604,n2605,n2636);
or (n2605,n2606,n2635);
and (n2606,n2607,n2634);
xor (n2607,n2608,n2633);
or (n2608,n2609,n2632);
and (n2609,n2610,n2631);
xor (n2610,n2611,n2630);
or (n2611,n2612,n2629);
and (n2612,n2613,n2616);
xor (n2613,n2614,n2615);
xor (n2614,n2431,n2464);
xor (n2615,n2473,n2531);
or (n2616,n2617,n2628);
and (n2617,n2618,n2627);
xor (n2618,n2619,n2620);
xor (n2619,n2434,n2443);
or (n2620,n2621,n2626);
and (n2621,n2622,n2625);
xor (n2622,n2623,n2624);
xor (n2623,n2451,n2460);
wire s0n2624,s1n2624,notn2624;
or (n2624,s0n2624,s1n2624);
not(notn2624,n1396);
and (s0n2624,notn2624,1'b0);
and (s1n2624,n1396,n2436);
wire s0n2625,s1n2625,notn2625;
or (n2625,s0n2625,s1n2625);
not(notn2625,n1761);
and (s0n2625,notn2625,1'b0);
and (s1n2625,n1761,n2444);
and (n2626,n2623,n2624);
wire s0n2627,s1n2627,notn2627;
or (n2627,s0n2627,s1n2627);
not(notn2627,n1444);
and (s0n2627,notn2627,1'b0);
and (s1n2627,n1444,n2307);
and (n2628,n2619,n2620);
and (n2629,n2614,n2615);
xor (n2630,n2426,n2429);
xor (n2631,n2470,n2534);
and (n2632,n2611,n2630);
xor (n2633,n2423,n2468);
xor (n2634,n2551,n2598);
and (n2635,n2608,n2633);
xor (n2636,n2547,n2600);
or (n2637,n2638,n2800);
and (n2638,n2639,n2704);
xor (n2639,n2640,n2703);
or (n2640,n2641,n2702);
and (n2641,n2642,n2701);
xor (n2642,n2643,n2700);
or (n2643,n2644,n2699);
and (n2644,n2645,n2692);
xor (n2645,n2646,n2691);
or (n2646,n2647,n2690);
and (n2647,n2648,n2671);
xor (n2648,n2649,n2670);
or (n2649,n2650,n2669);
and (n2650,n2651,n2668);
xor (n2651,n2652,n2667);
or (n2652,n2653,n2666);
and (n2653,n2654,n2665);
xor (n2654,n2655,n2656);
xor (n2655,n2484,n2487);
or (n2656,n2657,n2664);
and (n2657,n2658,n2663);
xor (n2658,n2659,n2662);
and (n2659,n2660,n2661);
wire s0n2660,s1n2660,notn2660;
or (n2660,s0n2660,s1n2660);
not(notn2660,n1444);
and (s0n2660,notn2660,1'b0);
and (s1n2660,n1444,n2441);
wire s0n2661,s1n2661,notn2661;
or (n2661,s0n2661,s1n2661);
not(notn2661,n1444);
and (s0n2661,notn2661,1'b0);
and (s1n2661,n1444,n2368);
wire s0n2662,s1n2662,notn2662;
or (n2662,s0n2662,s1n2662);
not(notn2662,n1396);
and (s0n2662,notn2662,1'b0);
and (s1n2662,n1396,n2368);
xor (n2663,n2521,n2523);
and (n2664,n2659,n2662);
wire s0n2665,s1n2665,notn2665;
or (n2665,s0n2665,s1n2665);
not(notn2665,n1761);
and (s0n2665,notn2665,1'b0);
and (s1n2665,n1761,n2462);
and (n2666,n2655,n2656);
xor (n2667,n2481,n2503);
xor (n2668,n2507,n2527);
and (n2669,n2652,n2667);
xor (n2670,n2477,n2505);
or (n2671,n2672,n2689);
and (n2672,n2673,n2688);
xor (n2673,n2674,n2687);
or (n2674,n2675,n2686);
and (n2675,n2676,n2685);
xor (n2676,n2677,n2678);
wire s0n2677,s1n2677,notn2677;
or (n2677,s0n2677,s1n2677);
not(notn2677,n1396);
and (s0n2677,notn2677,1'b0);
and (s1n2677,n1396,n2528);
or (n2678,n2679,n2684);
and (n2679,n2680,n2683);
xor (n2680,n2681,n2682);
wire s0n2681,s1n2681,notn2681;
or (n2681,s0n2681,s1n2681);
not(notn2681,n1761);
and (s0n2681,notn2681,1'b0);
and (s1n2681,n1761,n2459);
xor (n2682,n2514,n2517);
wire s0n2683,s1n2683,notn2683;
or (n2683,s0n2683,s1n2683);
not(notn2683,n1761);
and (s0n2683,notn2683,1'b0);
and (s1n2683,n1761,n2441);
and (n2684,n2681,n2682);
xor (n2685,n2578,n2581);
and (n2686,n2677,n2678);
wire s0n2687,s1n2687,notn2687;
or (n2687,s0n2687,s1n2687);
not(notn2687,n1444);
and (s0n2687,notn2687,1'b0);
and (s1n2687,n1444,n2396);
wire s0n2688,s1n2688,notn2688;
or (n2688,s0n2688,s1n2688);
not(notn2688,n1444);
and (s0n2688,notn2688,1'b0);
and (s1n2688,n1444,n2303);
and (n2689,n2674,n2687);
and (n2690,n2649,n2670);
xor (n2691,n2558,n2563);
or (n2692,n2693,n2698);
and (n2693,n2694,n2697);
xor (n2694,n2695,n2696);
xor (n2695,n2570,n2585);
xor (n2696,n2590,n2593);
xor (n2697,n2618,n2627);
and (n2698,n2695,n2696);
and (n2699,n2646,n2691);
xor (n2700,n2555,n2596);
xor (n2701,n2610,n2631);
and (n2702,n2643,n2700);
xor (n2703,n2607,n2634);
or (n2704,n2705,n2799);
and (n2705,n2706,n2798);
xor (n2706,n2707,n2750);
or (n2707,n2708,n2749);
and (n2708,n2709,n2748);
xor (n2709,n2710,n2747);
or (n2710,n2711,n2746);
and (n2711,n2712,n2727);
xor (n2712,n2713,n2726);
or (n2713,n2714,n2725);
and (n2714,n2715,n2724);
xor (n2715,n2716,n2723);
or (n2716,n2717,n2722);
and (n2717,n2718,n2721);
xor (n2718,n2719,n2720);
wire s0n2719,s1n2719,notn2719;
or (n2719,s0n2719,s1n2719);
not(notn2719,n1444);
and (s0n2719,notn2719,1'b0);
and (s1n2719,n1444,n2436);
xor (n2720,n2511,n2525);
wire s0n2721,s1n2721,notn2721;
or (n2721,s0n2721,s1n2721);
not(notn2721,n1444);
and (s0n2721,notn2721,1'b0);
and (s1n2721,n1444,n2444);
and (n2722,n2719,n2720);
xor (n2723,n2574,n2583);
xor (n2724,n2622,n2625);
and (n2725,n2716,n2723);
xor (n2726,n2648,n2671);
or (n2727,n2728,n2745);
and (n2728,n2729,n2744);
xor (n2729,n2730,n2731);
xor (n2730,n2651,n2668);
or (n2731,n2732,n2743);
and (n2732,n2733,n2742);
xor (n2733,n2734,n2741);
or (n2734,n2735,n2740);
and (n2735,n2736,n2739);
xor (n2736,n2737,n2738);
wire s0n2737,s1n2737,notn2737;
or (n2737,s0n2737,s1n2737);
not(notn2737,n1444);
and (s0n2737,notn2737,1'b0);
and (s1n2737,n1444,n2462);
xor (n2738,n2658,n2663);
wire s0n2739,s1n2739,notn2739;
or (n2739,s0n2739,s1n2739);
not(notn2739,n1444);
and (s0n2739,notn2739,1'b0);
and (s1n2739,n1444,n2528);
and (n2740,n2737,n2738);
xor (n2741,n2654,n2665);
xor (n2742,n2676,n2685);
and (n2743,n2734,n2741);
xor (n2744,n2673,n2688);
and (n2745,n2730,n2731);
and (n2746,n2713,n2726);
xor (n2747,n2567,n2588);
xor (n2748,n2613,n2616);
and (n2749,n2710,n2747);
nand (n2750,n2751,n2794);
or (n2751,n2752,n2792);
not (n2752,n2753);
nand (n2753,n2754,n2756,n2791);
not (n2754,n2755);
xor (n2755,n2645,n2692);
nand (n2756,n2757,n2790);
or (n2757,n2758,n2759);
xor (n2758,n2712,n2727);
nand (n2759,n2760,n2787);
or (n2760,n2761,n2785);
not (n2761,n2762);
nand (n2762,n2763,n2782);
or (n2763,n2764,n2780);
not (n2764,n2765);
nand (n2765,n2766,n2777);
or (n2766,n2767,n2775);
not (n2767,n2768);
nand (n2768,n2769,n2772);
or (n2769,n2197,n2770);
not (n2770,n2771);
wire s0n2771,s1n2771,notn2771;
or (n2771,s0n2771,s1n2771);
not(notn2771,n1444);
and (s0n2771,notn2771,1'b0);
and (s1n2771,n1444,n2459);
nand (n2772,n2773,n2774);
or (n2773,n2771,n2198);
xor (n2774,n2660,n2661);
not (n2775,n2776);
xor (n2776,n2680,n2683);
nand (n2777,n2778,n2779);
or (n2778,n2776,n2768);
xor (n2779,n2736,n2739);
not (n2780,n2781);
xor (n2781,n2718,n2721);
nand (n2782,n2783,n2784);
or (n2783,n2781,n2765);
xor (n2784,n2733,n2742);
not (n2785,n2786);
xor (n2786,n2715,n2724);
nand (n2787,n2788,n2789);
or (n2788,n2786,n2762);
xor (n2789,n2729,n2744);
xor (n2790,n2694,n2697);
nand (n2791,n2758,n2759);
not (n2792,n2793);
xor (n2793,n2709,n2748);
nand (n2794,n2795,n2755);
or (n2795,n2796,n2797);
not (n2796,n2791);
not (n2797,n2756);
xor (n2798,n2642,n2701);
and (n2799,n2707,n2750);
and (n2800,n2640,n2703);
and (n2801,n2605,n2636);
and (n2802,n2544,n2545);
and (n2803,n2412,n2413);
and (n2804,n2333,n2334);
and (n2805,n2256,n2257);
endmodule
