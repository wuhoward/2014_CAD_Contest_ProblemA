module top (out,n18,n19,n25,n27,n34,n48,n49,n55,n59
        ,n65,n74,n75,n83,n89,n100,n106,n110,n128,n134
        ,n138,n152,n160,n168,n174,n182,n203,n210,n212,n217
        ,n221,n241,n275);
output out;
input n18;
input n19;
input n25;
input n27;
input n34;
input n48;
input n49;
input n55;
input n59;
input n65;
input n74;
input n75;
input n83;
input n89;
input n100;
input n106;
input n110;
input n128;
input n134;
input n138;
input n152;
input n160;
input n168;
input n174;
input n182;
input n203;
input n210;
input n212;
input n217;
input n221;
input n241;
input n275;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n20;
wire n21;
wire n22;
wire n23;
wire n24;
wire n26;
wire n28;
wire n29;
wire n30;
wire n31;
wire n32;
wire n33;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n56;
wire n57;
wire n58;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n107;
wire n108;
wire n109;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n135;
wire n136;
wire n137;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n211;
wire n213;
wire n214;
wire n215;
wire n216;
wire n218;
wire n219;
wire n220;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
xor (out,n0,n1058);
nand (n0,n1,n1057);
or (n1,n2,n484);
not (n2,n3);
nand (n3,n4,n483);
not (n4,n5);
nor (n5,n6,n391);
xor (n6,n7,n343);
xor (n7,n8,n185);
xor (n8,n9,n145);
xor (n9,n10,n93);
or (n10,n11,n92);
and (n11,n12,n68);
xor (n12,n13,n42);
nand (n13,n14,n30);
or (n14,n15,n22);
nor (n15,n16,n20);
and (n16,n17,n19);
not (n17,n18);
and (n20,n18,n21);
not (n21,n19);
not (n22,n23);
nand (n23,n24,n28);
or (n24,n25,n26);
not (n26,n27);
or (n28,n29,n27);
not (n29,n25);
nand (n30,n31,n37);
not (n31,n32);
nor (n32,n33,n35);
and (n33,n34,n29);
and (n35,n36,n25);
not (n36,n34);
not (n37,n38);
nand (n38,n15,n39);
nand (n39,n40,n41);
or (n40,n18,n29);
nand (n41,n29,n18);
nand (n42,n43,n62);
or (n43,n44,n57);
nand (n44,n45,n52);
nor (n45,n46,n50);
and (n46,n47,n49);
not (n47,n48);
and (n50,n48,n51);
not (n51,n49);
nand (n52,n53,n56);
nand (n53,n54,n49);
not (n54,n55);
nand (n56,n55,n51);
nor (n57,n58,n60);
and (n58,n59,n54);
and (n60,n55,n61);
not (n61,n59);
or (n62,n63,n45);
nor (n63,n64,n66);
and (n64,n65,n54);
and (n66,n55,n67);
not (n67,n65);
nand (n68,n69,n86);
or (n69,n70,n81);
nand (n70,n71,n78);
or (n71,n72,n76);
and (n72,n73,n75);
not (n73,n74);
and (n76,n74,n77);
not (n77,n75);
nor (n78,n79,n80);
and (n79,n55,n73);
and (n80,n54,n74);
nor (n81,n82,n84);
and (n82,n83,n77);
and (n84,n75,n85);
not (n85,n83);
or (n86,n87,n78);
nor (n87,n88,n90);
and (n88,n89,n77);
and (n90,n75,n91);
not (n91,n89);
and (n92,n13,n42);
xor (n93,n94,n123);
xor (n94,n95,n117);
nand (n95,n96,n113);
or (n96,n97,n108);
nand (n97,n98,n103);
nor (n98,n99,n101);
and (n99,n29,n100);
and (n101,n25,n102);
not (n102,n100);
nand (n103,n104,n107);
or (n104,n100,n105);
not (n105,n106);
nand (n107,n105,n100);
nor (n108,n109,n111);
and (n109,n105,n110);
and (n111,n106,n112);
not (n112,n110);
or (n113,n98,n114);
nor (n114,n115,n116);
and (n115,n105,n34);
and (n116,n106,n36);
nand (n117,n118,n119);
or (n118,n70,n87);
or (n119,n120,n78);
nor (n120,n121,n122);
and (n121,n59,n77);
and (n122,n75,n61);
nand (n123,n124,n141);
or (n124,n125,n136);
nand (n125,n126,n131);
nor (n126,n127,n129);
and (n127,n77,n128);
and (n129,n75,n130);
not (n130,n128);
nand (n131,n132,n135);
or (n132,n133,n128);
not (n133,n134);
nand (n135,n133,n128);
nor (n136,n137,n139);
and (n137,n138,n133);
and (n139,n134,n140);
not (n140,n138);
or (n141,n142,n126);
nor (n142,n143,n144);
and (n143,n83,n133);
and (n144,n134,n85);
xor (n145,n146,n177);
xor (n146,n147,n155);
nand (n147,n148,n149);
or (n148,n22,n38);
or (n149,n15,n150);
nor (n150,n151,n153);
and (n151,n29,n152);
and (n153,n25,n154);
not (n154,n152);
nand (n155,n156,n171);
or (n156,n157,n166);
nand (n157,n158,n163);
nor (n158,n159,n161);
and (n159,n105,n160);
and (n161,n106,n162);
not (n162,n160);
nand (n163,n164,n165);
or (n164,n47,n160);
nand (n165,n47,n160);
nor (n166,n167,n169);
and (n167,n47,n168);
and (n169,n48,n170);
not (n170,n168);
or (n171,n158,n172);
nor (n172,n173,n175);
and (n173,n47,n174);
and (n175,n48,n176);
not (n176,n174);
nand (n177,n178,n179);
or (n178,n44,n63);
or (n179,n45,n180);
nor (n180,n181,n183);
and (n181,n182,n54);
and (n183,n55,n184);
not (n184,n182);
or (n185,n186,n342);
and (n186,n187,n314);
xor (n187,n188,n255);
or (n188,n189,n254);
and (n189,n190,n224);
xor (n190,n191,n198);
nand (n191,n192,n197);
or (n192,n70,n193);
not (n193,n194);
nand (n194,n195,n196);
or (n195,n140,n75);
or (n196,n77,n138);
or (n197,n81,n78);
xor (n198,n199,n206);
nor (n199,n200,n133);
nor (n200,n201,n204);
and (n201,n202,n77);
nand (n202,n203,n128);
and (n204,n205,n130);
not (n205,n203);
nand (n206,n207,n218);
or (n207,n208,n215);
nor (n208,n209,n213);
and (n209,n210,n211);
not (n211,n212);
and (n213,n214,n212);
not (n214,n210);
nand (n215,n216,n212);
not (n216,n217);
or (n218,n219,n216);
nor (n219,n220,n222);
and (n220,n211,n221);
and (n222,n212,n223);
not (n223,n221);
or (n224,n225,n253);
and (n225,n226,n234);
xor (n226,n227,n228);
nor (n227,n126,n205);
nand (n228,n229,n233);
or (n229,n230,n215);
nor (n230,n231,n232);
and (n231,n212,n154);
nor (n232,n212,n154);
or (n233,n208,n216);
nand (n234,n235,n249);
or (n235,n236,n246);
nand (n236,n237,n243);
not (n237,n238);
nand (n238,n239,n242);
or (n239,n240,n212);
not (n240,n241);
nand (n242,n240,n212);
nand (n243,n244,n245);
or (n244,n240,n19);
nand (n245,n19,n240);
nor (n246,n247,n248);
and (n247,n21,n34);
and (n248,n19,n36);
or (n249,n237,n250);
nor (n250,n251,n252);
and (n251,n21,n27);
and (n252,n19,n26);
and (n253,n227,n228);
and (n254,n191,n198);
xor (n255,n256,n288);
xor (n256,n257,n258);
and (n257,n199,n206);
or (n258,n259,n287);
and (n259,n260,n278);
xor (n260,n261,n267);
nand (n261,n262,n263);
or (n262,n236,n250);
or (n263,n237,n264);
nor (n264,n265,n266);
and (n265,n21,n152);
and (n266,n19,n154);
nand (n267,n268,n272);
or (n268,n125,n269);
nor (n269,n270,n271);
and (n270,n205,n134);
and (n271,n203,n133);
or (n272,n273,n126);
nor (n273,n274,n276);
and (n274,n275,n133);
and (n276,n277,n134);
not (n277,n275);
nand (n278,n279,n283);
or (n279,n97,n280);
nor (n280,n281,n282);
and (n281,n105,n168);
and (n282,n106,n170);
or (n283,n98,n284);
nor (n284,n285,n286);
and (n285,n105,n174);
and (n286,n106,n176);
and (n287,n261,n267);
or (n288,n289,n313);
and (n289,n290,n307);
xor (n290,n291,n301);
nand (n291,n292,n297);
or (n292,n158,n293);
not (n293,n294);
nor (n294,n295,n296);
and (n295,n184,n47);
and (n296,n182,n48);
or (n297,n157,n298);
nor (n298,n299,n300);
and (n299,n47,n65);
and (n300,n48,n67);
nand (n301,n302,n306);
or (n302,n38,n303);
nor (n303,n304,n305);
and (n304,n29,n110);
and (n305,n25,n112);
or (n306,n15,n32);
nand (n307,n308,n312);
or (n308,n44,n309);
nor (n309,n310,n311);
and (n310,n54,n89);
and (n311,n55,n91);
or (n312,n45,n57);
and (n313,n291,n301);
or (n314,n315,n341);
and (n315,n316,n340);
xor (n316,n317,n339);
or (n317,n318,n338);
and (n318,n319,n332);
xor (n319,n320,n326);
nand (n320,n321,n325);
or (n321,n97,n322);
nor (n322,n323,n324);
and (n323,n182,n105);
and (n324,n106,n184);
or (n325,n280,n98);
nand (n326,n327,n331);
or (n327,n157,n328);
nor (n328,n329,n330);
and (n329,n47,n59);
and (n330,n48,n61);
or (n331,n298,n158);
nand (n332,n333,n337);
or (n333,n38,n334);
nor (n334,n335,n336);
and (n335,n29,n174);
and (n336,n25,n176);
or (n337,n15,n303);
and (n338,n320,n326);
xor (n339,n290,n307);
xor (n340,n260,n278);
and (n341,n317,n339);
and (n342,n188,n255);
xor (n343,n344,n383);
xor (n344,n345,n348);
or (n345,n346,n347);
and (n346,n256,n288);
and (n347,n257,n258);
xor (n348,n349,n370);
xor (n349,n350,n360);
not (n350,n351);
nand (n351,n352,n356);
or (n352,n236,n353);
nor (n353,n354,n355);
and (n354,n21,n210);
and (n355,n19,n214);
or (n356,n237,n357);
nor (n357,n358,n359);
and (n358,n21,n221);
and (n359,n19,n223);
nand (n360,n361,n366);
not (n361,n362);
nand (n362,n363,n365);
or (n363,n364,n217);
not (n364,n215);
not (n365,n219);
not (n366,n367);
nand (n367,n368,n369);
or (n368,n236,n264);
or (n369,n237,n353);
or (n370,n371,n382);
and (n371,n372,n379);
xor (n372,n373,n376);
nand (n373,n374,n375);
or (n374,n125,n273);
or (n375,n136,n126);
nand (n376,n377,n378);
or (n377,n97,n284);
or (n378,n98,n108);
nand (n379,n380,n381);
or (n380,n157,n293);
or (n381,n166,n158);
and (n382,n373,n376);
or (n383,n384,n390);
and (n384,n385,n389);
xor (n385,n386,n387);
xor (n386,n12,n68);
nand (n387,n388,n360);
or (n388,n361,n366);
xor (n389,n372,n379);
and (n390,n386,n387);
or (n391,n392,n482);
and (n392,n393,n481);
xor (n393,n394,n395);
xor (n394,n385,n389);
or (n395,n396,n480);
and (n396,n397,n429);
xor (n397,n398,n428);
or (n398,n399,n427);
and (n399,n400,n415);
xor (n400,n401,n407);
nand (n401,n402,n406);
or (n402,n44,n403);
nor (n403,n404,n405);
and (n404,n83,n54);
and (n405,n55,n85);
or (n406,n45,n309);
nand (n407,n408,n409);
or (n408,n78,n193);
nand (n409,n410,n414);
not (n410,n411);
nor (n411,n412,n413);
and (n412,n77,n275);
and (n413,n277,n75);
not (n414,n70);
and (n415,n416,n421);
nor (n416,n417,n77);
nor (n417,n418,n420);
and (n418,n419,n54);
nand (n419,n74,n203);
and (n420,n205,n73);
nand (n421,n422,n426);
or (n422,n423,n215);
nor (n423,n424,n425);
and (n424,n211,n27);
and (n425,n212,n26);
or (n426,n230,n216);
and (n427,n401,n407);
xor (n428,n190,n224);
or (n429,n430,n479);
and (n430,n431,n478);
xor (n431,n432,n456);
or (n432,n433,n455);
and (n433,n434,n448);
xor (n434,n435,n441);
nand (n435,n436,n440);
or (n436,n236,n437);
nor (n437,n438,n439);
and (n438,n110,n21);
and (n439,n112,n19);
or (n440,n237,n246);
nand (n441,n442,n447);
or (n442,n443,n97);
not (n443,n444);
nand (n444,n445,n446);
or (n445,n106,n67);
or (n446,n105,n65);
or (n447,n322,n98);
nand (n448,n449,n454);
or (n449,n157,n450);
not (n450,n451);
nor (n451,n452,n453);
and (n452,n91,n47);
and (n453,n89,n48);
or (n454,n328,n158);
and (n455,n435,n441);
or (n456,n457,n477);
and (n457,n458,n471);
xor (n458,n459,n465);
nand (n459,n460,n464);
or (n460,n38,n461);
nor (n461,n462,n463);
and (n462,n29,n168);
and (n463,n25,n170);
or (n464,n15,n334);
nand (n465,n466,n470);
or (n466,n44,n467);
nor (n467,n468,n469);
and (n468,n138,n54);
and (n469,n55,n140);
or (n470,n403,n45);
nand (n471,n472,n476);
or (n472,n70,n473);
nor (n473,n474,n475);
and (n474,n205,n75);
and (n475,n203,n77);
or (n476,n411,n78);
and (n477,n459,n465);
xor (n478,n226,n234);
and (n479,n432,n456);
and (n480,n398,n428);
xor (n481,n187,n314);
and (n482,n394,n395);
nand (n483,n6,n391);
not (n484,n485);
nand (n485,n486,n1056);
or (n486,n487,n1051);
not (n487,n488);
or (n488,n489,n1050);
and (n489,n490,n613);
xor (n490,n491,n606);
or (n491,n492,n605);
and (n492,n493,n549);
xor (n493,n494,n495);
xor (n494,n431,n478);
xor (n495,n496,n499);
xor (n496,n497,n498);
xor (n497,n319,n332);
xor (n498,n400,n415);
or (n499,n500,n548);
and (n500,n501,n524);
xor (n501,n502,n503);
xor (n502,n416,n421);
or (n503,n504,n523);
and (n504,n505,n516);
xor (n505,n506,n508);
and (n506,n507,n203);
not (n507,n78);
nand (n508,n509,n514);
or (n509,n510,n236);
not (n510,n511);
nand (n511,n512,n513);
or (n512,n19,n176);
or (n513,n21,n174);
nand (n514,n515,n238);
not (n515,n437);
nand (n516,n517,n522);
or (n517,n97,n518);
not (n518,n519);
nand (n519,n520,n521);
or (n520,n106,n61);
or (n521,n105,n59);
or (n522,n98,n443);
and (n523,n506,n508);
or (n524,n525,n547);
and (n525,n526,n541);
xor (n526,n527,n535);
nand (n527,n528,n533);
or (n528,n529,n157);
not (n529,n530);
nand (n530,n531,n532);
or (n531,n48,n85);
or (n532,n47,n83);
nand (n533,n451,n534);
not (n534,n158);
nand (n535,n536,n537);
or (n536,n216,n423);
or (n537,n538,n215);
nor (n538,n539,n540);
and (n539,n211,n34);
and (n540,n212,n36);
nand (n541,n542,n546);
or (n542,n543,n44);
nor (n543,n544,n545);
and (n544,n275,n54);
and (n545,n55,n277);
or (n546,n467,n45);
and (n547,n527,n535);
and (n548,n502,n503);
or (n549,n550,n604);
and (n550,n551,n554);
xor (n551,n552,n553);
xor (n552,n458,n471);
xor (n553,n434,n448);
or (n554,n555,n603);
and (n555,n556,n577);
xor (n556,n557,n563);
nand (n557,n558,n562);
or (n558,n38,n559);
nor (n559,n560,n561);
and (n560,n29,n182);
and (n561,n25,n184);
or (n562,n15,n461);
nor (n563,n564,n571);
not (n564,n565);
nand (n565,n566,n570);
or (n566,n567,n236);
nor (n567,n568,n569);
and (n568,n168,n21);
and (n569,n170,n19);
nand (n570,n238,n511);
nand (n571,n572,n55);
nand (n572,n573,n574);
or (n573,n203,n49);
nand (n574,n575,n47);
not (n575,n576);
and (n576,n203,n49);
or (n577,n578,n602);
and (n578,n579,n595);
xor (n579,n580,n588);
nand (n580,n581,n582);
or (n581,n98,n518);
nand (n582,n583,n587);
not (n583,n584);
nor (n584,n585,n586);
and (n585,n91,n106);
and (n586,n89,n105);
not (n587,n97);
nand (n588,n589,n594);
or (n589,n590,n157);
not (n590,n591);
nor (n591,n592,n593);
and (n592,n47,n140);
and (n593,n48,n138);
nand (n594,n534,n530);
nand (n595,n596,n601);
or (n596,n597,n215);
not (n597,n598);
or (n598,n599,n600);
and (n599,n112,n212);
and (n600,n110,n211);
or (n601,n538,n216);
and (n602,n580,n588);
and (n603,n557,n563);
and (n604,n552,n553);
and (n605,n494,n495);
xor (n606,n607,n612);
xor (n607,n608,n609);
xor (n608,n316,n340);
or (n609,n610,n611);
and (n610,n496,n499);
and (n611,n497,n498);
xor (n612,n397,n429);
or (n613,n614,n1049);
and (n614,n615,n649);
xor (n615,n616,n648);
or (n616,n617,n647);
and (n617,n618,n646);
xor (n618,n619,n620);
xor (n619,n501,n524);
or (n620,n621,n645);
and (n621,n622,n625);
xor (n622,n623,n624);
xor (n623,n526,n541);
xor (n624,n505,n516);
or (n625,n626,n644);
and (n626,n627,n640);
xor (n627,n628,n634);
nand (n628,n629,n633);
or (n629,n44,n630);
nor (n630,n631,n632);
and (n631,n205,n55);
and (n632,n203,n54);
or (n633,n543,n45);
nand (n634,n635,n639);
or (n635,n38,n636);
nor (n636,n637,n638);
and (n637,n29,n65);
and (n638,n25,n67);
or (n639,n15,n559);
nand (n640,n641,n643);
or (n641,n642,n564);
not (n642,n571);
or (n643,n565,n571);
and (n644,n628,n634);
and (n645,n623,n624);
xor (n646,n551,n554);
and (n647,n619,n620);
xor (n648,n493,n549);
nand (n649,n650,n1045);
or (n650,n651,n1023);
nor (n651,n652,n1022);
and (n652,n653,n1003);
or (n653,n654,n1002);
and (n654,n655,n798);
xor (n655,n656,n767);
or (n656,n657,n766);
and (n657,n658,n728);
xor (n658,n659,n689);
xor (n659,n660,n679);
xor (n660,n661,n670);
nand (n661,n662,n666);
or (n662,n97,n663);
nor (n663,n664,n665);
and (n664,n138,n105);
and (n665,n140,n106);
or (n666,n667,n98);
nor (n667,n668,n669);
and (n668,n105,n83);
and (n669,n106,n85);
nand (n670,n671,n675);
or (n671,n157,n672);
nor (n672,n673,n674);
and (n673,n205,n48);
and (n674,n203,n47);
or (n675,n676,n158);
nor (n676,n677,n678);
and (n677,n275,n47);
and (n678,n277,n48);
nand (n679,n680,n685);
or (n680,n215,n681);
not (n681,n682);
nor (n682,n683,n684);
and (n683,n168,n212);
and (n684,n170,n211);
or (n685,n686,n216);
nor (n686,n687,n688);
and (n687,n174,n211);
and (n688,n176,n212);
or (n689,n690,n727);
and (n690,n691,n710);
xor (n691,n692,n701);
nand (n692,n693,n697);
or (n693,n236,n694);
nor (n694,n695,n696);
and (n695,n21,n59);
and (n696,n19,n61);
or (n697,n237,n698);
nor (n698,n699,n700);
and (n699,n67,n19);
and (n700,n65,n21);
nand (n701,n702,n706);
or (n702,n38,n703);
nor (n703,n704,n705);
and (n704,n83,n29);
and (n705,n25,n85);
or (n706,n15,n707);
nor (n707,n708,n709);
and (n708,n29,n89);
and (n709,n25,n91);
and (n710,n711,n717);
nor (n711,n712,n105);
nor (n712,n713,n716);
and (n713,n714,n29);
not (n714,n715);
and (n715,n203,n100);
and (n716,n205,n102);
nand (n717,n718,n723);
or (n718,n719,n215);
not (n719,n720);
nor (n720,n721,n722);
and (n721,n67,n211);
and (n722,n65,n212);
or (n723,n724,n216);
nor (n724,n725,n726);
and (n725,n182,n211);
and (n726,n184,n212);
and (n727,n692,n701);
xor (n728,n729,n751);
xor (n729,n730,n736);
nand (n730,n731,n732);
or (n731,n38,n707);
or (n732,n15,n733);
nor (n733,n734,n735);
and (n734,n29,n59);
and (n735,n25,n61);
xor (n736,n737,n742);
nor (n737,n738,n47);
nor (n738,n739,n741);
and (n739,n740,n105);
nand (n740,n203,n160);
and (n741,n205,n162);
nand (n742,n743,n748);
or (n743,n237,n744);
not (n744,n745);
nand (n745,n746,n747);
or (n746,n19,n184);
or (n747,n21,n182);
nand (n748,n749,n750);
not (n749,n698);
not (n750,n236);
or (n751,n752,n765);
and (n752,n753,n758);
xor (n753,n754,n755);
nor (n754,n158,n205);
nand (n755,n756,n757);
or (n756,n216,n681);
or (n757,n724,n215);
nand (n758,n759,n760);
or (n759,n98,n663);
nand (n760,n761,n587);
not (n761,n762);
or (n762,n763,n764);
and (n763,n277,n105);
and (n764,n275,n106);
and (n765,n754,n755);
and (n766,n659,n689);
xor (n767,n768,n783);
xor (n768,n769,n780);
xor (n769,n770,n777);
xor (n770,n771,n774);
nand (n771,n772,n773);
or (n772,n158,n590);
or (n773,n157,n676);
nand (n774,n775,n776);
or (n775,n686,n215);
nand (n776,n598,n217);
nand (n777,n778,n779);
or (n778,n38,n733);
or (n779,n15,n636);
or (n780,n781,n782);
and (n781,n729,n751);
and (n782,n730,n736);
xor (n783,n784,n789);
xor (n784,n785,n786);
and (n785,n737,n742);
or (n786,n787,n788);
and (n787,n660,n679);
and (n788,n661,n670);
xor (n789,n790,n795);
xor (n790,n791,n792);
nor (n791,n45,n205);
nand (n792,n793,n794);
or (n793,n744,n236);
or (n794,n237,n567);
nand (n795,n796,n797);
or (n796,n97,n667);
or (n797,n98,n584);
nand (n798,n799,n998,n1001);
nand (n799,n800,n855,n991);
not (n800,n801);
nor (n801,n802,n829);
xor (n802,n803,n828);
xor (n803,n804,n827);
or (n804,n805,n826);
and (n805,n806,n820);
xor (n806,n807,n813);
nand (n807,n808,n812);
or (n808,n97,n809);
nor (n809,n810,n811);
and (n810,n205,n106);
and (n811,n203,n105);
or (n812,n762,n98);
nand (n813,n814,n819);
or (n814,n815,n236);
not (n815,n816);
nor (n816,n817,n818);
and (n817,n89,n19);
and (n818,n91,n21);
or (n819,n237,n694);
nand (n820,n821,n825);
or (n821,n38,n822);
nor (n822,n823,n824);
and (n823,n138,n29);
and (n824,n25,n140);
or (n825,n15,n703);
and (n826,n807,n813);
xor (n827,n753,n758);
xor (n828,n691,n710);
or (n829,n830,n854);
and (n830,n831,n853);
xor (n831,n832,n833);
xor (n832,n711,n717);
or (n833,n834,n852);
and (n834,n835,n845);
xor (n835,n836,n838);
and (n836,n837,n203);
not (n837,n98);
nand (n838,n839,n844);
or (n839,n215,n840);
not (n840,n841);
nor (n841,n842,n843);
and (n842,n61,n211);
and (n843,n59,n212);
nand (n844,n720,n217);
nand (n845,n846,n851);
or (n846,n847,n236);
not (n847,n848);
nor (n848,n849,n850);
and (n849,n85,n21);
and (n850,n83,n19);
nand (n851,n816,n238);
and (n852,n836,n838);
xor (n853,n806,n820);
and (n854,n832,n833);
or (n855,n856,n990);
and (n856,n857,n883);
xor (n857,n858,n882);
or (n858,n859,n881);
and (n859,n860,n880);
xor (n860,n861,n867);
nand (n861,n862,n866);
or (n862,n38,n863);
nor (n863,n864,n865);
and (n864,n29,n275);
and (n865,n25,n277);
or (n866,n822,n15);
and (n867,n868,n874);
and (n868,n869,n25);
nand (n869,n870,n871);
or (n870,n203,n18);
nand (n871,n872,n21);
not (n872,n873);
and (n873,n203,n18);
nand (n874,n875,n876);
or (n875,n216,n840);
or (n876,n877,n215);
nor (n877,n878,n879);
and (n878,n211,n89);
and (n879,n212,n91);
xor (n880,n835,n845);
and (n881,n861,n867);
xor (n882,n831,n853);
nand (n883,n884,n989);
or (n884,n885,n984);
nor (n885,n886,n983);
and (n886,n887,n962);
nand (n887,n888,n960);
or (n888,n889,n943);
not (n889,n890);
or (n890,n891,n942);
and (n891,n892,n921);
xor (n892,n893,n902);
nand (n893,n894,n898);
or (n894,n236,n895);
nor (n895,n896,n897);
and (n896,n19,n205);
and (n897,n203,n21);
or (n898,n237,n899);
nor (n899,n900,n901);
and (n900,n277,n19);
and (n901,n275,n21);
nand (n902,n903,n920);
or (n903,n904,n910);
not (n904,n905);
nand (n905,n906,n19);
nand (n906,n907,n909);
or (n907,n908,n212);
and (n908,n203,n241);
nand (n909,n205,n240);
not (n910,n911);
nand (n911,n912,n916);
or (n912,n913,n215);
or (n913,n914,n915);
and (n914,n138,n212);
and (n915,n140,n211);
or (n916,n917,n216);
nor (n917,n918,n919);
and (n918,n85,n212);
and (n919,n83,n211);
or (n920,n911,n905);
or (n921,n922,n941);
and (n922,n923,n931);
xor (n923,n924,n925);
nor (n924,n237,n205);
nand (n925,n926,n930);
or (n926,n927,n215);
nor (n927,n928,n929);
and (n928,n277,n212);
and (n929,n275,n211);
or (n930,n913,n216);
nor (n931,n932,n939);
nor (n932,n933,n935);
and (n933,n934,n217);
not (n934,n927);
and (n935,n936,n364);
nand (n936,n937,n938);
or (n937,n205,n212);
nand (n938,n212,n205);
or (n939,n940,n211);
and (n940,n203,n217);
and (n941,n924,n925);
and (n942,n893,n902);
not (n943,n944);
nand (n944,n945,n959);
not (n945,n946);
xor (n946,n947,n956);
xor (n947,n948,n950);
and (n948,n949,n203);
not (n949,n15);
nand (n950,n951,n952);
or (n951,n899,n236);
nand (n952,n953,n238);
nor (n953,n954,n955);
and (n954,n140,n21);
and (n955,n138,n19);
nand (n956,n957,n958);
or (n957,n917,n215);
or (n958,n877,n216);
nand (n959,n904,n911);
nand (n960,n961,n946);
not (n961,n959);
nand (n962,n963,n979);
not (n963,n964);
xor (n964,n965,n978);
xor (n965,n966,n970);
nand (n966,n967,n969);
or (n967,n968,n236);
not (n968,n953);
nand (n969,n848,n238);
nand (n970,n971,n976);
or (n971,n972,n38);
not (n972,n973);
nand (n973,n974,n975);
or (n974,n203,n29);
or (n975,n205,n25);
nand (n976,n977,n949);
not (n977,n863);
xor (n978,n868,n874);
not (n979,n980);
or (n980,n981,n982);
and (n981,n947,n956);
and (n982,n948,n950);
nor (n983,n963,n979);
nor (n984,n985,n986);
xor (n985,n860,n880);
or (n986,n987,n988);
and (n987,n965,n978);
and (n988,n966,n970);
nand (n989,n985,n986);
and (n990,n858,n882);
nand (n991,n992,n996);
not (n992,n993);
or (n993,n994,n995);
and (n994,n803,n828);
and (n995,n804,n827);
not (n996,n997);
xor (n997,n658,n728);
nand (n998,n999,n991);
not (n999,n1000);
nand (n1000,n802,n829);
nand (n1001,n997,n993);
and (n1002,n656,n767);
or (n1003,n1004,n1019);
xor (n1004,n1005,n1016);
xor (n1005,n1006,n1007);
xor (n1006,n627,n640);
xor (n1007,n1008,n1015);
xor (n1008,n1009,n1012);
or (n1009,n1010,n1011);
and (n1010,n790,n795);
and (n1011,n791,n792);
or (n1012,n1013,n1014);
and (n1013,n770,n777);
and (n1014,n771,n774);
xor (n1015,n579,n595);
or (n1016,n1017,n1018);
and (n1017,n784,n789);
and (n1018,n785,n786);
or (n1019,n1020,n1021);
and (n1020,n768,n783);
and (n1021,n769,n780);
and (n1022,n1004,n1019);
nand (n1023,n1024,n1038);
not (n1024,n1025);
and (n1025,n1026,n1034);
not (n1026,n1027);
xor (n1027,n1028,n1033);
xor (n1028,n1029,n1030);
xor (n1029,n556,n577);
or (n1030,n1031,n1032);
and (n1031,n1008,n1015);
and (n1032,n1009,n1012);
xor (n1033,n622,n625);
not (n1034,n1035);
or (n1035,n1036,n1037);
and (n1036,n1005,n1016);
and (n1037,n1006,n1007);
nand (n1038,n1039,n1041);
not (n1039,n1040);
xor (n1040,n618,n646);
not (n1041,n1042);
or (n1042,n1043,n1044);
and (n1043,n1028,n1033);
and (n1044,n1029,n1030);
nor (n1045,n1046,n1048);
and (n1046,n1038,n1047);
nor (n1047,n1026,n1034);
nor (n1048,n1039,n1041);
and (n1049,n616,n648);
and (n1050,n491,n606);
nor (n1051,n1052,n1055);
or (n1052,n1053,n1054);
and (n1053,n607,n612);
and (n1054,n608,n609);
xor (n1055,n393,n481);
nand (n1056,n1055,n1052);
or (n1057,n485,n3);
xor (n1058,n1059,n1850);
xor (n1059,n1060,n1851);
xor (n1060,n1061,n1845);
xor (n1061,n1062,n1842);
xor (n1062,n1063,n1841);
xor (n1063,n1064,n1826);
xor (n1064,n1065,n1825);
xor (n1065,n1066,n1804);
xor (n1066,n1067,n1803);
xor (n1067,n1068,n1776);
xor (n1068,n1069,n1775);
xor (n1069,n1070,n1742);
xor (n1070,n1071,n1741);
xor (n1071,n1072,n1703);
xor (n1072,n1073,n1702);
xor (n1073,n1074,n1660);
xor (n1074,n1075,n1659);
xor (n1075,n1076,n1608);
xor (n1076,n1077,n1607);
xor (n1077,n1078,n1551);
xor (n1078,n1079,n1550);
xor (n1079,n1080,n1488);
xor (n1080,n1081,n1487);
xor (n1081,n1082,n1418);
xor (n1082,n1083,n1417);
xor (n1083,n1084,n1343);
xor (n1084,n1085,n1342);
xor (n1085,n1086,n1264);
xor (n1086,n1087,n1263);
xor (n1087,n1088,n1095);
xor (n1088,n1089,n1094);
xor (n1089,n1090,n1093);
xor (n1090,n1091,n1092);
and (n1091,n221,n217);
and (n1092,n221,n212);
and (n1093,n1091,n1092);
and (n1094,n221,n241);
or (n1095,n1096,n1181);
and (n1096,n1097,n1180);
xor (n1097,n1090,n1098);
or (n1098,n1099,n1101);
and (n1099,n1091,n1100);
and (n1100,n210,n212);
and (n1101,n1102,n1103);
xor (n1102,n1091,n1100);
or (n1103,n1104,n1107);
and (n1104,n1105,n1106);
and (n1105,n210,n217);
and (n1106,n152,n212);
and (n1107,n1108,n1109);
xor (n1108,n1105,n1106);
or (n1109,n1110,n1113);
and (n1110,n1111,n1112);
and (n1111,n152,n217);
and (n1112,n27,n212);
and (n1113,n1114,n1115);
xor (n1114,n1111,n1112);
or (n1115,n1116,n1119);
and (n1116,n1117,n1118);
and (n1117,n27,n217);
and (n1118,n34,n212);
and (n1119,n1120,n1121);
xor (n1120,n1117,n1118);
or (n1121,n1122,n1125);
and (n1122,n1123,n1124);
and (n1123,n34,n217);
and (n1124,n110,n212);
and (n1125,n1126,n1127);
xor (n1126,n1123,n1124);
or (n1127,n1128,n1131);
and (n1128,n1129,n1130);
and (n1129,n110,n217);
and (n1130,n174,n212);
and (n1131,n1132,n1133);
xor (n1132,n1129,n1130);
or (n1133,n1134,n1136);
and (n1134,n1135,n683);
and (n1135,n174,n217);
and (n1136,n1137,n1138);
xor (n1137,n1135,n683);
or (n1138,n1139,n1142);
and (n1139,n1140,n1141);
and (n1140,n168,n217);
and (n1141,n182,n212);
and (n1142,n1143,n1144);
xor (n1143,n1140,n1141);
or (n1144,n1145,n1147);
and (n1145,n1146,n722);
and (n1146,n182,n217);
and (n1147,n1148,n1149);
xor (n1148,n1146,n722);
or (n1149,n1150,n1152);
and (n1150,n1151,n843);
and (n1151,n65,n217);
and (n1152,n1153,n1154);
xor (n1153,n1151,n843);
or (n1154,n1155,n1158);
and (n1155,n1156,n1157);
and (n1156,n59,n217);
and (n1157,n89,n212);
and (n1158,n1159,n1160);
xor (n1159,n1156,n1157);
or (n1160,n1161,n1164);
and (n1161,n1162,n1163);
and (n1162,n89,n217);
and (n1163,n83,n212);
and (n1164,n1165,n1166);
xor (n1165,n1162,n1163);
or (n1166,n1167,n1169);
and (n1167,n1168,n914);
and (n1168,n83,n217);
and (n1169,n1170,n1171);
xor (n1170,n1168,n914);
or (n1171,n1172,n1175);
and (n1172,n1173,n1174);
and (n1173,n138,n217);
and (n1174,n275,n212);
and (n1175,n1176,n1177);
xor (n1176,n1173,n1174);
and (n1177,n1178,n1179);
and (n1178,n275,n217);
and (n1179,n203,n212);
and (n1180,n210,n241);
and (n1181,n1182,n1183);
xor (n1182,n1097,n1180);
or (n1183,n1184,n1187);
and (n1184,n1185,n1186);
xor (n1185,n1102,n1103);
and (n1186,n152,n241);
and (n1187,n1188,n1189);
xor (n1188,n1185,n1186);
or (n1189,n1190,n1193);
and (n1190,n1191,n1192);
xor (n1191,n1108,n1109);
and (n1192,n27,n241);
and (n1193,n1194,n1195);
xor (n1194,n1191,n1192);
or (n1195,n1196,n1199);
and (n1196,n1197,n1198);
xor (n1197,n1114,n1115);
and (n1198,n34,n241);
and (n1199,n1200,n1201);
xor (n1200,n1197,n1198);
or (n1201,n1202,n1205);
and (n1202,n1203,n1204);
xor (n1203,n1120,n1121);
and (n1204,n110,n241);
and (n1205,n1206,n1207);
xor (n1206,n1203,n1204);
or (n1207,n1208,n1211);
and (n1208,n1209,n1210);
xor (n1209,n1126,n1127);
and (n1210,n174,n241);
and (n1211,n1212,n1213);
xor (n1212,n1209,n1210);
or (n1213,n1214,n1217);
and (n1214,n1215,n1216);
xor (n1215,n1132,n1133);
and (n1216,n168,n241);
and (n1217,n1218,n1219);
xor (n1218,n1215,n1216);
or (n1219,n1220,n1223);
and (n1220,n1221,n1222);
xor (n1221,n1137,n1138);
and (n1222,n182,n241);
and (n1223,n1224,n1225);
xor (n1224,n1221,n1222);
or (n1225,n1226,n1229);
and (n1226,n1227,n1228);
xor (n1227,n1143,n1144);
and (n1228,n65,n241);
and (n1229,n1230,n1231);
xor (n1230,n1227,n1228);
or (n1231,n1232,n1235);
and (n1232,n1233,n1234);
xor (n1233,n1148,n1149);
and (n1234,n59,n241);
and (n1235,n1236,n1237);
xor (n1236,n1233,n1234);
or (n1237,n1238,n1241);
and (n1238,n1239,n1240);
xor (n1239,n1153,n1154);
and (n1240,n89,n241);
and (n1241,n1242,n1243);
xor (n1242,n1239,n1240);
or (n1243,n1244,n1247);
and (n1244,n1245,n1246);
xor (n1245,n1159,n1160);
and (n1246,n83,n241);
and (n1247,n1248,n1249);
xor (n1248,n1245,n1246);
or (n1249,n1250,n1253);
and (n1250,n1251,n1252);
xor (n1251,n1165,n1166);
and (n1252,n138,n241);
and (n1253,n1254,n1255);
xor (n1254,n1251,n1252);
or (n1255,n1256,n1259);
and (n1256,n1257,n1258);
xor (n1257,n1170,n1171);
and (n1258,n275,n241);
and (n1259,n1260,n1261);
xor (n1260,n1257,n1258);
and (n1261,n1262,n908);
xor (n1262,n1176,n1177);
and (n1263,n210,n19);
or (n1264,n1265,n1268);
and (n1265,n1266,n1267);
xor (n1266,n1182,n1183);
and (n1267,n152,n19);
and (n1268,n1269,n1270);
xor (n1269,n1266,n1267);
or (n1270,n1271,n1274);
and (n1271,n1272,n1273);
xor (n1272,n1188,n1189);
and (n1273,n27,n19);
and (n1274,n1275,n1276);
xor (n1275,n1272,n1273);
or (n1276,n1277,n1280);
and (n1277,n1278,n1279);
xor (n1278,n1194,n1195);
and (n1279,n34,n19);
and (n1280,n1281,n1282);
xor (n1281,n1278,n1279);
or (n1282,n1283,n1286);
and (n1283,n1284,n1285);
xor (n1284,n1200,n1201);
and (n1285,n110,n19);
and (n1286,n1287,n1288);
xor (n1287,n1284,n1285);
or (n1288,n1289,n1292);
and (n1289,n1290,n1291);
xor (n1290,n1206,n1207);
and (n1291,n174,n19);
and (n1292,n1293,n1294);
xor (n1293,n1290,n1291);
or (n1294,n1295,n1298);
and (n1295,n1296,n1297);
xor (n1296,n1212,n1213);
and (n1297,n168,n19);
and (n1298,n1299,n1300);
xor (n1299,n1296,n1297);
or (n1300,n1301,n1304);
and (n1301,n1302,n1303);
xor (n1302,n1218,n1219);
and (n1303,n182,n19);
and (n1304,n1305,n1306);
xor (n1305,n1302,n1303);
or (n1306,n1307,n1310);
and (n1307,n1308,n1309);
xor (n1308,n1224,n1225);
and (n1309,n65,n19);
and (n1310,n1311,n1312);
xor (n1311,n1308,n1309);
or (n1312,n1313,n1316);
and (n1313,n1314,n1315);
xor (n1314,n1230,n1231);
and (n1315,n59,n19);
and (n1316,n1317,n1318);
xor (n1317,n1314,n1315);
or (n1318,n1319,n1321);
and (n1319,n1320,n817);
xor (n1320,n1236,n1237);
and (n1321,n1322,n1323);
xor (n1322,n1320,n817);
or (n1323,n1324,n1326);
and (n1324,n1325,n850);
xor (n1325,n1242,n1243);
and (n1326,n1327,n1328);
xor (n1327,n1325,n850);
or (n1328,n1329,n1331);
and (n1329,n1330,n955);
xor (n1330,n1248,n1249);
and (n1331,n1332,n1333);
xor (n1332,n1330,n955);
or (n1333,n1334,n1337);
and (n1334,n1335,n1336);
xor (n1335,n1254,n1255);
and (n1336,n275,n19);
and (n1337,n1338,n1339);
xor (n1338,n1335,n1336);
and (n1339,n1340,n1341);
xor (n1340,n1260,n1261);
and (n1341,n203,n19);
and (n1342,n152,n18);
or (n1343,n1344,n1347);
and (n1344,n1345,n1346);
xor (n1345,n1269,n1270);
and (n1346,n27,n18);
and (n1347,n1348,n1349);
xor (n1348,n1345,n1346);
or (n1349,n1350,n1353);
and (n1350,n1351,n1352);
xor (n1351,n1275,n1276);
and (n1352,n34,n18);
and (n1353,n1354,n1355);
xor (n1354,n1351,n1352);
or (n1355,n1356,n1359);
and (n1356,n1357,n1358);
xor (n1357,n1281,n1282);
and (n1358,n110,n18);
and (n1359,n1360,n1361);
xor (n1360,n1357,n1358);
or (n1361,n1362,n1365);
and (n1362,n1363,n1364);
xor (n1363,n1287,n1288);
and (n1364,n174,n18);
and (n1365,n1366,n1367);
xor (n1366,n1363,n1364);
or (n1367,n1368,n1371);
and (n1368,n1369,n1370);
xor (n1369,n1293,n1294);
and (n1370,n168,n18);
and (n1371,n1372,n1373);
xor (n1372,n1369,n1370);
or (n1373,n1374,n1377);
and (n1374,n1375,n1376);
xor (n1375,n1299,n1300);
and (n1376,n182,n18);
and (n1377,n1378,n1379);
xor (n1378,n1375,n1376);
or (n1379,n1380,n1383);
and (n1380,n1381,n1382);
xor (n1381,n1305,n1306);
and (n1382,n65,n18);
and (n1383,n1384,n1385);
xor (n1384,n1381,n1382);
or (n1385,n1386,n1389);
and (n1386,n1387,n1388);
xor (n1387,n1311,n1312);
and (n1388,n59,n18);
and (n1389,n1390,n1391);
xor (n1390,n1387,n1388);
or (n1391,n1392,n1395);
and (n1392,n1393,n1394);
xor (n1393,n1317,n1318);
and (n1394,n89,n18);
and (n1395,n1396,n1397);
xor (n1396,n1393,n1394);
or (n1397,n1398,n1401);
and (n1398,n1399,n1400);
xor (n1399,n1322,n1323);
and (n1400,n83,n18);
and (n1401,n1402,n1403);
xor (n1402,n1399,n1400);
or (n1403,n1404,n1407);
and (n1404,n1405,n1406);
xor (n1405,n1327,n1328);
and (n1406,n138,n18);
and (n1407,n1408,n1409);
xor (n1408,n1405,n1406);
or (n1409,n1410,n1413);
and (n1410,n1411,n1412);
xor (n1411,n1332,n1333);
and (n1412,n275,n18);
and (n1413,n1414,n1415);
xor (n1414,n1411,n1412);
and (n1415,n1416,n873);
xor (n1416,n1338,n1339);
and (n1417,n27,n25);
or (n1418,n1419,n1422);
and (n1419,n1420,n1421);
xor (n1420,n1348,n1349);
and (n1421,n34,n25);
and (n1422,n1423,n1424);
xor (n1423,n1420,n1421);
or (n1424,n1425,n1428);
and (n1425,n1426,n1427);
xor (n1426,n1354,n1355);
and (n1427,n110,n25);
and (n1428,n1429,n1430);
xor (n1429,n1426,n1427);
or (n1430,n1431,n1434);
and (n1431,n1432,n1433);
xor (n1432,n1360,n1361);
and (n1433,n174,n25);
and (n1434,n1435,n1436);
xor (n1435,n1432,n1433);
or (n1436,n1437,n1440);
and (n1437,n1438,n1439);
xor (n1438,n1366,n1367);
and (n1439,n168,n25);
and (n1440,n1441,n1442);
xor (n1441,n1438,n1439);
or (n1442,n1443,n1446);
and (n1443,n1444,n1445);
xor (n1444,n1372,n1373);
and (n1445,n182,n25);
and (n1446,n1447,n1448);
xor (n1447,n1444,n1445);
or (n1448,n1449,n1452);
and (n1449,n1450,n1451);
xor (n1450,n1378,n1379);
and (n1451,n65,n25);
and (n1452,n1453,n1454);
xor (n1453,n1450,n1451);
or (n1454,n1455,n1458);
and (n1455,n1456,n1457);
xor (n1456,n1384,n1385);
and (n1457,n59,n25);
and (n1458,n1459,n1460);
xor (n1459,n1456,n1457);
or (n1460,n1461,n1464);
and (n1461,n1462,n1463);
xor (n1462,n1390,n1391);
and (n1463,n89,n25);
and (n1464,n1465,n1466);
xor (n1465,n1462,n1463);
or (n1466,n1467,n1470);
and (n1467,n1468,n1469);
xor (n1468,n1396,n1397);
and (n1469,n83,n25);
and (n1470,n1471,n1472);
xor (n1471,n1468,n1469);
or (n1472,n1473,n1476);
and (n1473,n1474,n1475);
xor (n1474,n1402,n1403);
and (n1475,n138,n25);
and (n1476,n1477,n1478);
xor (n1477,n1474,n1475);
or (n1478,n1479,n1482);
and (n1479,n1480,n1481);
xor (n1480,n1408,n1409);
and (n1481,n275,n25);
and (n1482,n1483,n1484);
xor (n1483,n1480,n1481);
and (n1484,n1485,n1486);
xor (n1485,n1414,n1415);
and (n1486,n203,n25);
and (n1487,n34,n100);
or (n1488,n1489,n1492);
and (n1489,n1490,n1491);
xor (n1490,n1423,n1424);
and (n1491,n110,n100);
and (n1492,n1493,n1494);
xor (n1493,n1490,n1491);
or (n1494,n1495,n1498);
and (n1495,n1496,n1497);
xor (n1496,n1429,n1430);
and (n1497,n174,n100);
and (n1498,n1499,n1500);
xor (n1499,n1496,n1497);
or (n1500,n1501,n1504);
and (n1501,n1502,n1503);
xor (n1502,n1435,n1436);
and (n1503,n168,n100);
and (n1504,n1505,n1506);
xor (n1505,n1502,n1503);
or (n1506,n1507,n1510);
and (n1507,n1508,n1509);
xor (n1508,n1441,n1442);
and (n1509,n182,n100);
and (n1510,n1511,n1512);
xor (n1511,n1508,n1509);
or (n1512,n1513,n1516);
and (n1513,n1514,n1515);
xor (n1514,n1447,n1448);
and (n1515,n65,n100);
and (n1516,n1517,n1518);
xor (n1517,n1514,n1515);
or (n1518,n1519,n1522);
and (n1519,n1520,n1521);
xor (n1520,n1453,n1454);
and (n1521,n59,n100);
and (n1522,n1523,n1524);
xor (n1523,n1520,n1521);
or (n1524,n1525,n1528);
and (n1525,n1526,n1527);
xor (n1526,n1459,n1460);
and (n1527,n89,n100);
and (n1528,n1529,n1530);
xor (n1529,n1526,n1527);
or (n1530,n1531,n1534);
and (n1531,n1532,n1533);
xor (n1532,n1465,n1466);
and (n1533,n83,n100);
and (n1534,n1535,n1536);
xor (n1535,n1532,n1533);
or (n1536,n1537,n1540);
and (n1537,n1538,n1539);
xor (n1538,n1471,n1472);
and (n1539,n138,n100);
and (n1540,n1541,n1542);
xor (n1541,n1538,n1539);
or (n1542,n1543,n1546);
and (n1543,n1544,n1545);
xor (n1544,n1477,n1478);
and (n1545,n275,n100);
and (n1546,n1547,n1548);
xor (n1547,n1544,n1545);
and (n1548,n1549,n715);
xor (n1549,n1483,n1484);
and (n1550,n110,n106);
or (n1551,n1552,n1555);
and (n1552,n1553,n1554);
xor (n1553,n1493,n1494);
and (n1554,n174,n106);
and (n1555,n1556,n1557);
xor (n1556,n1553,n1554);
or (n1557,n1558,n1561);
and (n1558,n1559,n1560);
xor (n1559,n1499,n1500);
and (n1560,n168,n106);
and (n1561,n1562,n1563);
xor (n1562,n1559,n1560);
or (n1563,n1564,n1567);
and (n1564,n1565,n1566);
xor (n1565,n1505,n1506);
and (n1566,n182,n106);
and (n1567,n1568,n1569);
xor (n1568,n1565,n1566);
or (n1569,n1570,n1573);
and (n1570,n1571,n1572);
xor (n1571,n1511,n1512);
and (n1572,n65,n106);
and (n1573,n1574,n1575);
xor (n1574,n1571,n1572);
or (n1575,n1576,n1579);
and (n1576,n1577,n1578);
xor (n1577,n1517,n1518);
and (n1578,n59,n106);
and (n1579,n1580,n1581);
xor (n1580,n1577,n1578);
or (n1581,n1582,n1585);
and (n1582,n1583,n1584);
xor (n1583,n1523,n1524);
and (n1584,n89,n106);
and (n1585,n1586,n1587);
xor (n1586,n1583,n1584);
or (n1587,n1588,n1591);
and (n1588,n1589,n1590);
xor (n1589,n1529,n1530);
and (n1590,n83,n106);
and (n1591,n1592,n1593);
xor (n1592,n1589,n1590);
or (n1593,n1594,n1597);
and (n1594,n1595,n1596);
xor (n1595,n1535,n1536);
and (n1596,n138,n106);
and (n1597,n1598,n1599);
xor (n1598,n1595,n1596);
or (n1599,n1600,n1602);
and (n1600,n1601,n764);
xor (n1601,n1541,n1542);
and (n1602,n1603,n1604);
xor (n1603,n1601,n764);
and (n1604,n1605,n1606);
xor (n1605,n1547,n1548);
and (n1606,n203,n106);
and (n1607,n174,n160);
or (n1608,n1609,n1612);
and (n1609,n1610,n1611);
xor (n1610,n1556,n1557);
and (n1611,n168,n160);
and (n1612,n1613,n1614);
xor (n1613,n1610,n1611);
or (n1614,n1615,n1618);
and (n1615,n1616,n1617);
xor (n1616,n1562,n1563);
and (n1617,n182,n160);
and (n1618,n1619,n1620);
xor (n1619,n1616,n1617);
or (n1620,n1621,n1624);
and (n1621,n1622,n1623);
xor (n1622,n1568,n1569);
and (n1623,n65,n160);
and (n1624,n1625,n1626);
xor (n1625,n1622,n1623);
or (n1626,n1627,n1630);
and (n1627,n1628,n1629);
xor (n1628,n1574,n1575);
and (n1629,n59,n160);
and (n1630,n1631,n1632);
xor (n1631,n1628,n1629);
or (n1632,n1633,n1636);
and (n1633,n1634,n1635);
xor (n1634,n1580,n1581);
and (n1635,n89,n160);
and (n1636,n1637,n1638);
xor (n1637,n1634,n1635);
or (n1638,n1639,n1642);
and (n1639,n1640,n1641);
xor (n1640,n1586,n1587);
and (n1641,n83,n160);
and (n1642,n1643,n1644);
xor (n1643,n1640,n1641);
or (n1644,n1645,n1648);
and (n1645,n1646,n1647);
xor (n1646,n1592,n1593);
and (n1647,n138,n160);
and (n1648,n1649,n1650);
xor (n1649,n1646,n1647);
or (n1650,n1651,n1654);
and (n1651,n1652,n1653);
xor (n1652,n1598,n1599);
and (n1653,n275,n160);
and (n1654,n1655,n1656);
xor (n1655,n1652,n1653);
and (n1656,n1657,n1658);
xor (n1657,n1603,n1604);
not (n1658,n740);
and (n1659,n168,n48);
or (n1660,n1661,n1663);
and (n1661,n1662,n296);
xor (n1662,n1613,n1614);
and (n1663,n1664,n1665);
xor (n1664,n1662,n296);
or (n1665,n1666,n1669);
and (n1666,n1667,n1668);
xor (n1667,n1619,n1620);
and (n1668,n65,n48);
and (n1669,n1670,n1671);
xor (n1670,n1667,n1668);
or (n1671,n1672,n1675);
and (n1672,n1673,n1674);
xor (n1673,n1625,n1626);
and (n1674,n59,n48);
and (n1675,n1676,n1677);
xor (n1676,n1673,n1674);
or (n1677,n1678,n1680);
and (n1678,n1679,n453);
xor (n1679,n1631,n1632);
and (n1680,n1681,n1682);
xor (n1681,n1679,n453);
or (n1682,n1683,n1686);
and (n1683,n1684,n1685);
xor (n1684,n1637,n1638);
and (n1685,n83,n48);
and (n1686,n1687,n1688);
xor (n1687,n1684,n1685);
or (n1688,n1689,n1691);
and (n1689,n1690,n593);
xor (n1690,n1643,n1644);
and (n1691,n1692,n1693);
xor (n1692,n1690,n593);
or (n1693,n1694,n1697);
and (n1694,n1695,n1696);
xor (n1695,n1649,n1650);
and (n1696,n275,n48);
and (n1697,n1698,n1699);
xor (n1698,n1695,n1696);
and (n1699,n1700,n1701);
xor (n1700,n1655,n1656);
and (n1701,n203,n48);
and (n1702,n182,n49);
or (n1703,n1704,n1707);
and (n1704,n1705,n1706);
xor (n1705,n1664,n1665);
and (n1706,n65,n49);
and (n1707,n1708,n1709);
xor (n1708,n1705,n1706);
or (n1709,n1710,n1713);
and (n1710,n1711,n1712);
xor (n1711,n1670,n1671);
and (n1712,n59,n49);
and (n1713,n1714,n1715);
xor (n1714,n1711,n1712);
or (n1715,n1716,n1719);
and (n1716,n1717,n1718);
xor (n1717,n1676,n1677);
and (n1718,n89,n49);
and (n1719,n1720,n1721);
xor (n1720,n1717,n1718);
or (n1721,n1722,n1725);
and (n1722,n1723,n1724);
xor (n1723,n1681,n1682);
and (n1724,n83,n49);
and (n1725,n1726,n1727);
xor (n1726,n1723,n1724);
or (n1727,n1728,n1731);
and (n1728,n1729,n1730);
xor (n1729,n1687,n1688);
and (n1730,n138,n49);
and (n1731,n1732,n1733);
xor (n1732,n1729,n1730);
or (n1733,n1734,n1737);
and (n1734,n1735,n1736);
xor (n1735,n1692,n1693);
and (n1736,n275,n49);
and (n1737,n1738,n1739);
xor (n1738,n1735,n1736);
and (n1739,n1740,n576);
xor (n1740,n1698,n1699);
and (n1741,n65,n55);
or (n1742,n1743,n1746);
and (n1743,n1744,n1745);
xor (n1744,n1708,n1709);
and (n1745,n59,n55);
and (n1746,n1747,n1748);
xor (n1747,n1744,n1745);
or (n1748,n1749,n1752);
and (n1749,n1750,n1751);
xor (n1750,n1714,n1715);
and (n1751,n89,n55);
and (n1752,n1753,n1754);
xor (n1753,n1750,n1751);
or (n1754,n1755,n1758);
and (n1755,n1756,n1757);
xor (n1756,n1720,n1721);
and (n1757,n83,n55);
and (n1758,n1759,n1760);
xor (n1759,n1756,n1757);
or (n1760,n1761,n1764);
and (n1761,n1762,n1763);
xor (n1762,n1726,n1727);
and (n1763,n138,n55);
and (n1764,n1765,n1766);
xor (n1765,n1762,n1763);
or (n1766,n1767,n1770);
and (n1767,n1768,n1769);
xor (n1768,n1732,n1733);
and (n1769,n275,n55);
and (n1770,n1771,n1772);
xor (n1771,n1768,n1769);
and (n1772,n1773,n1774);
xor (n1773,n1738,n1739);
and (n1774,n203,n55);
and (n1775,n59,n74);
or (n1776,n1777,n1780);
and (n1777,n1778,n1779);
xor (n1778,n1747,n1748);
and (n1779,n89,n74);
and (n1780,n1781,n1782);
xor (n1781,n1778,n1779);
or (n1782,n1783,n1786);
and (n1783,n1784,n1785);
xor (n1784,n1753,n1754);
and (n1785,n83,n74);
and (n1786,n1787,n1788);
xor (n1787,n1784,n1785);
or (n1788,n1789,n1792);
and (n1789,n1790,n1791);
xor (n1790,n1759,n1760);
and (n1791,n138,n74);
and (n1792,n1793,n1794);
xor (n1793,n1790,n1791);
or (n1794,n1795,n1798);
and (n1795,n1796,n1797);
xor (n1796,n1765,n1766);
and (n1797,n275,n74);
and (n1798,n1799,n1800);
xor (n1799,n1796,n1797);
and (n1800,n1801,n1802);
xor (n1801,n1771,n1772);
not (n1802,n419);
and (n1803,n89,n75);
or (n1804,n1805,n1808);
and (n1805,n1806,n1807);
xor (n1806,n1781,n1782);
and (n1807,n83,n75);
and (n1808,n1809,n1810);
xor (n1809,n1806,n1807);
or (n1810,n1811,n1814);
and (n1811,n1812,n1813);
xor (n1812,n1787,n1788);
and (n1813,n138,n75);
and (n1814,n1815,n1816);
xor (n1815,n1812,n1813);
or (n1816,n1817,n1820);
and (n1817,n1818,n1819);
xor (n1818,n1793,n1794);
and (n1819,n275,n75);
and (n1820,n1821,n1822);
xor (n1821,n1818,n1819);
and (n1822,n1823,n1824);
xor (n1823,n1799,n1800);
and (n1824,n203,n75);
and (n1825,n83,n128);
or (n1826,n1827,n1830);
and (n1827,n1828,n1829);
xor (n1828,n1809,n1810);
and (n1829,n138,n128);
and (n1830,n1831,n1832);
xor (n1831,n1828,n1829);
or (n1832,n1833,n1836);
and (n1833,n1834,n1835);
xor (n1834,n1815,n1816);
and (n1835,n275,n128);
and (n1836,n1837,n1838);
xor (n1837,n1834,n1835);
and (n1838,n1839,n1840);
xor (n1839,n1821,n1822);
not (n1840,n202);
and (n1841,n138,n134);
or (n1842,n1843,n1846);
and (n1843,n1844,n1845);
xor (n1844,n1831,n1832);
and (n1845,n275,n134);
and (n1846,n1847,n1848);
xor (n1847,n1844,n1845);
and (n1848,n1849,n1850);
xor (n1849,n1837,n1838);
and (n1850,n203,n134);
and (n1851,n1852,n1850);
xor (n1852,n1847,n1848);
endmodule
