module top (out,n3,n4,n5,n22,n24,n31,n32,n42,n49
        ,n50,n55,n59,n68,n70,n75,n80,n86,n97,n105
        ,n115,n121,n143,n154,n182,n202);
output out;
input n3;
input n4;
input n5;
input n22;
input n24;
input n31;
input n32;
input n42;
input n49;
input n50;
input n55;
input n59;
input n68;
input n70;
input n75;
input n80;
input n86;
input n97;
input n105;
input n115;
input n121;
input n143;
input n154;
input n182;
input n202;
wire n0;
wire n1;
wire n2;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n23;
wire n25;
wire n26;
wire n27;
wire n28;
wire n29;
wire n30;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n51;
wire n52;
wire n53;
wire n54;
wire n56;
wire n57;
wire n58;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n69;
wire n71;
wire n72;
wire n73;
wire n74;
wire n76;
wire n77;
wire n78;
wire n79;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
xnor (out,n0,n464);
nor (n0,n1,n6);
and (n1,n2,n5);
nor (n2,n3,n4);
and (n6,n7,n461);
nand (n7,n8,n460);
or (n8,n9,n256);
not (n9,n10);
and (n10,n11,n255);
or (n11,n12,n218);
xor (n12,n13,n170);
xor (n13,n14,n90);
xor (n14,n15,n62);
xor (n15,n16,n44);
nand (n16,n17,n38);
or (n17,n18,n26);
not (n18,n19);
nor (n19,n20,n25);
and (n20,n21,n23);
not (n21,n22);
not (n23,n24);
and (n25,n22,n24);
not (n26,n27);
nor (n27,n28,n34);
nand (n28,n29,n33);
or (n29,n30,n32);
not (n30,n31);
nand (n33,n30,n32);
nor (n34,n35,n36);
and (n35,n23,n32);
and (n36,n24,n37);
not (n37,n32);
nand (n38,n28,n39);
nand (n39,n40,n43);
or (n40,n24,n41);
not (n41,n42);
or (n43,n23,n42);
nand (n44,n45,n56);
or (n45,n46,n53);
nor (n46,n47,n51);
and (n47,n48,n50);
not (n48,n49);
and (n51,n49,n52);
not (n52,n50);
nand (n53,n54,n49);
not (n54,n55);
or (n56,n57,n54);
nor (n57,n58,n60);
and (n58,n48,n59);
and (n60,n49,n61);
not (n61,n59);
nand (n62,n63,n83);
or (n63,n64,n78);
not (n64,n65);
nor (n65,n66,n72);
nand (n66,n67,n71);
or (n67,n68,n69);
not (n69,n70);
nand (n71,n68,n69);
nor (n72,n73,n76);
and (n73,n74,n75);
not (n74,n68);
and (n76,n68,n77);
not (n77,n75);
nor (n78,n79,n81);
and (n79,n77,n80);
and (n81,n75,n82);
not (n82,n80);
or (n83,n84,n89);
nor (n84,n85,n87);
and (n85,n77,n86);
and (n87,n75,n88);
not (n88,n86);
not (n89,n66);
or (n90,n91,n169);
and (n91,n92,n133);
xor (n92,n93,n101);
nand (n93,n94,n100);
or (n94,n64,n95);
nor (n95,n96,n98);
and (n96,n77,n97);
and (n98,n75,n99);
not (n99,n97);
or (n100,n89,n78);
xor (n101,n102,n109);
and (n102,n103,n24);
nand (n103,n104,n106);
or (n104,n105,n32);
nand (n106,n107,n30);
not (n107,n108);
and (n108,n105,n32);
nand (n109,n110,n123);
or (n110,n111,n117);
not (n111,n112);
nand (n112,n113,n116);
or (n113,n70,n114);
not (n114,n115);
or (n116,n69,n115);
not (n117,n118);
nand (n118,n119,n122);
or (n119,n120,n49);
not (n120,n121);
nand (n122,n49,n120);
nand (n123,n124,n128);
not (n124,n125);
nor (n125,n126,n127);
and (n126,n69,n86);
and (n127,n70,n88);
not (n128,n129);
nand (n129,n117,n130);
nand (n130,n131,n132);
or (n131,n120,n70);
nand (n132,n120,n70);
or (n133,n134,n168);
and (n134,n135,n149);
xor (n135,n136,n137);
and (n136,n28,n105);
nand (n137,n138,n145);
or (n138,n54,n139);
not (n139,n140);
nor (n140,n141,n144);
and (n141,n142,n48);
not (n142,n143);
and (n144,n143,n49);
or (n145,n146,n53);
nor (n146,n147,n148);
and (n147,n48,n115);
and (n148,n49,n114);
nand (n149,n150,n163);
or (n150,n151,n160);
nand (n151,n152,n156);
nand (n152,n153,n155);
or (n153,n154,n30);
nand (n155,n30,n154);
not (n156,n157);
nand (n157,n158,n159);
or (n158,n77,n154);
nand (n159,n154,n77);
nor (n160,n161,n162);
and (n161,n30,n22);
and (n162,n31,n21);
or (n163,n156,n164);
not (n164,n165);
nor (n165,n166,n167);
and (n166,n42,n31);
and (n167,n41,n30);
and (n168,n136,n137);
and (n169,n93,n101);
xor (n170,n171,n196);
xor (n171,n172,n173);
and (n172,n102,n109);
or (n173,n174,n195);
and (n174,n175,n192);
xor (n175,n176,n184);
nand (n176,n177,n178);
or (n177,n164,n151);
nand (n178,n157,n179);
nor (n179,n180,n183);
and (n180,n181,n30);
not (n181,n182);
and (n183,n182,n31);
nand (n184,n185,n191);
or (n185,n186,n26);
not (n186,n187);
nand (n187,n188,n189);
or (n188,n23,n105);
or (n189,n190,n24);
not (n190,n105);
nand (n191,n28,n19);
nand (n192,n193,n194);
or (n193,n53,n139);
or (n194,n46,n54);
and (n195,n176,n184);
xor (n196,n197,n210);
xor (n197,n198,n204);
and (n198,n199,n105);
nand (n199,n200,n203);
or (n200,n201,n24);
not (n201,n202);
nand (n203,n24,n201);
nand (n204,n205,n206);
or (n205,n111,n129);
nand (n206,n118,n207);
nand (n207,n208,n209);
or (n208,n70,n142);
or (n209,n69,n143);
nand (n210,n211,n213);
or (n211,n212,n151);
not (n212,n179);
nand (n213,n214,n157);
not (n214,n215);
nor (n215,n216,n217);
and (n216,n30,n97);
and (n217,n31,n99);
or (n218,n219,n254);
and (n219,n220,n253);
xor (n220,n221,n222);
xor (n221,n175,n192);
or (n222,n223,n252);
and (n223,n224,n237);
xor (n224,n225,n231);
nand (n225,n226,n230);
or (n226,n129,n227);
nor (n227,n228,n229);
and (n228,n69,n80);
and (n229,n70,n82);
or (n230,n117,n125);
nand (n231,n232,n236);
or (n232,n64,n233);
nor (n233,n234,n235);
and (n234,n77,n182);
and (n235,n75,n181);
or (n236,n95,n89);
and (n237,n238,n245);
nor (n238,n239,n30);
nor (n239,n240,n243);
and (n240,n241,n77);
not (n241,n242);
and (n242,n105,n154);
and (n243,n190,n244);
not (n244,n154);
nand (n245,n246,n251);
or (n246,n247,n53);
not (n247,n248);
nor (n248,n249,n250);
and (n249,n88,n48);
and (n250,n86,n49);
or (n251,n146,n54);
and (n252,n225,n231);
xor (n253,n92,n133);
and (n254,n221,n222);
nand (n255,n12,n218);
not (n256,n257);
nor (n257,n258,n456);
and (n258,n259,n322);
not (n259,n260);
nand (n260,n261,n316);
not (n261,n262);
nor (n262,n263,n291);
xor (n263,n264,n290);
xor (n264,n265,n289);
or (n265,n266,n288);
and (n266,n267,n282);
xor (n267,n268,n276);
nand (n268,n269,n274);
or (n269,n270,n151);
not (n270,n271);
nand (n271,n272,n273);
or (n272,n30,n105);
or (n273,n31,n190);
nand (n274,n275,n157);
not (n275,n160);
nand (n276,n277,n281);
or (n277,n129,n278);
nor (n278,n279,n280);
and (n279,n69,n97);
and (n280,n70,n99);
or (n281,n227,n117);
nand (n282,n283,n287);
or (n283,n64,n284);
nor (n284,n285,n286);
and (n285,n77,n42);
and (n286,n75,n41);
or (n287,n233,n89);
and (n288,n268,n276);
xor (n289,n135,n149);
xor (n290,n224,n237);
or (n291,n292,n315);
and (n292,n293,n314);
xor (n293,n294,n295);
xor (n294,n238,n245);
or (n295,n296,n313);
and (n296,n297,n306);
xor (n297,n298,n299);
and (n298,n157,n105);
nand (n299,n300,n305);
or (n300,n53,n301);
not (n301,n302);
nor (n302,n303,n304);
and (n303,n80,n49);
and (n304,n82,n48);
nand (n305,n248,n55);
nand (n306,n307,n312);
or (n307,n129,n308);
not (n308,n309);
nor (n309,n310,n311);
and (n310,n181,n69);
and (n311,n182,n70);
or (n312,n117,n278);
and (n313,n298,n299);
xor (n314,n267,n282);
and (n315,n294,n295);
not (n316,n317);
nor (n317,n318,n319);
xor (n318,n220,n253);
or (n319,n320,n321);
and (n320,n264,n290);
and (n321,n265,n289);
or (n322,n323,n455);
and (n323,n324,n352);
xor (n324,n325,n351);
or (n325,n326,n350);
and (n326,n327,n349);
xor (n327,n328,n335);
nand (n328,n329,n334);
or (n329,n64,n330);
not (n330,n331);
nor (n331,n332,n333);
and (n332,n22,n75);
and (n333,n21,n77);
or (n334,n284,n89);
and (n335,n336,n342);
nor (n336,n337,n77);
nor (n337,n338,n341);
and (n338,n339,n69);
not (n339,n340);
and (n340,n105,n68);
and (n341,n190,n74);
nand (n342,n343,n344);
or (n343,n54,n301);
nand (n344,n345,n348);
nand (n345,n346,n347);
or (n346,n97,n48);
nand (n347,n48,n97);
not (n348,n53);
xor (n349,n297,n306);
and (n350,n328,n335);
xor (n351,n293,n314);
or (n352,n353,n454);
and (n353,n354,n373);
xor (n354,n355,n372);
or (n355,n356,n371);
and (n356,n357,n370);
xor (n357,n358,n363);
nand (n358,n359,n362);
or (n359,n360,n129);
not (n360,n361);
xor (n361,n41,n69);
nand (n362,n118,n309);
nand (n363,n364,n369);
or (n364,n365,n64);
not (n365,n366);
nand (n366,n367,n368);
or (n367,n77,n105);
or (n368,n190,n75);
nand (n369,n331,n66);
xor (n370,n336,n342);
and (n371,n358,n363);
xor (n372,n327,n349);
or (n373,n374,n453);
and (n374,n375,n397);
xor (n375,n376,n396);
or (n376,n377,n395);
and (n377,n378,n387);
xor (n378,n379,n380);
and (n379,n66,n105);
nand (n380,n381,n386);
or (n381,n382,n129);
not (n382,n383);
nor (n383,n384,n385);
and (n384,n21,n69);
and (n385,n22,n70);
nand (n386,n118,n361);
nand (n387,n388,n393);
or (n388,n53,n389);
not (n389,n390);
nand (n390,n391,n392);
or (n391,n182,n48);
nand (n392,n48,n182);
or (n393,n394,n54);
not (n394,n345);
and (n395,n379,n380);
xor (n396,n357,n370);
nand (n397,n398,n452);
or (n398,n399,n414);
nor (n399,n400,n401);
xor (n400,n378,n387);
nor (n401,n402,n409);
not (n402,n403);
nand (n403,n404,n408);
or (n404,n53,n405);
nor (n405,n406,n407);
and (n406,n41,n49);
and (n407,n42,n48);
nand (n408,n390,n55);
nand (n409,n410,n70);
nand (n410,n411,n413);
or (n411,n412,n49);
and (n412,n105,n121);
or (n413,n105,n121);
nor (n414,n415,n451);
and (n415,n416,n427);
nand (n416,n417,n421);
nor (n417,n418,n419);
and (n418,n409,n403);
and (n419,n420,n402);
not (n420,n409);
nor (n421,n422,n426);
and (n422,n128,n423);
nand (n423,n424,n425);
or (n424,n69,n105);
or (n425,n190,n70);
and (n426,n118,n383);
nand (n427,n428,n450);
or (n428,n429,n444);
not (n429,n430);
nor (n430,n431,n442);
not (n431,n432);
nand (n432,n433,n438);
or (n433,n54,n434);
not (n434,n435);
nor (n435,n436,n437);
and (n436,n21,n48);
and (n437,n22,n49);
nand (n438,n439,n348);
nor (n439,n440,n441);
and (n440,n190,n48);
and (n441,n105,n49);
nand (n442,n443,n49);
nand (n443,n105,n55);
not (n444,n445);
nand (n445,n446,n449);
nor (n446,n447,n448);
nor (n447,n434,n53);
nor (n448,n405,n54);
nand (n449,n105,n118);
or (n450,n446,n449);
nor (n451,n421,n417);
nand (n452,n400,n401);
and (n453,n376,n396);
and (n454,n355,n372);
and (n455,n325,n351);
nand (n456,n457,n459);
or (n457,n317,n458);
nand (n458,n263,n291);
nand (n459,n318,n319);
or (n460,n257,n10);
not (n461,n462);
nand (n462,n463,n3);
not (n463,n4);
wire s0n464,s1n464,notn464;
or (n464,s0n464,s1n464);
not(notn464,n4);
and (s0n464,notn464,n465);
and (s1n464,n4,1'b0);
wire s0n465,s1n465,notn465;
or (n465,s0n465,s1n465);
not(notn465,n3);
and (s0n465,notn465,n5);
and (s1n465,n3,n466);
xor (n466,n467,n723);
xor (n467,n468,n720);
xor (n468,n469,n25);
xor (n469,n470,n712);
xor (n470,n471,n711);
xor (n471,n472,n697);
xor (n472,n473,n183);
xor (n473,n474,n677);
xor (n474,n475,n676);
xor (n475,n476,n650);
xor (n476,n477,n649);
xor (n477,n478,n617);
xor (n478,n479,n616);
xor (n479,n480,n579);
xor (n480,n481,n578);
xor (n481,n482,n534);
xor (n482,n483,n533);
xor (n483,n484,n487);
xor (n484,n485,n486);
and (n485,n59,n55);
and (n486,n50,n49);
or (n487,n488,n490);
and (n488,n489,n144);
and (n489,n50,n55);
and (n490,n491,n492);
xor (n491,n489,n144);
or (n492,n493,n496);
and (n493,n494,n495);
and (n494,n143,n55);
and (n495,n115,n49);
and (n496,n497,n498);
xor (n497,n494,n495);
or (n498,n499,n501);
and (n499,n500,n250);
and (n500,n115,n55);
and (n501,n502,n503);
xor (n502,n500,n250);
or (n503,n504,n506);
and (n504,n505,n303);
and (n505,n86,n55);
and (n506,n507,n508);
xor (n507,n505,n303);
or (n508,n509,n512);
and (n509,n510,n511);
and (n510,n80,n55);
and (n511,n97,n49);
and (n512,n513,n514);
xor (n513,n510,n511);
or (n514,n515,n518);
and (n515,n516,n517);
and (n516,n97,n55);
and (n517,n182,n49);
and (n518,n519,n520);
xor (n519,n516,n517);
or (n520,n521,n524);
and (n521,n522,n523);
and (n522,n182,n55);
and (n523,n42,n49);
and (n524,n525,n526);
xor (n525,n522,n523);
or (n526,n527,n529);
and (n527,n528,n437);
and (n528,n42,n55);
and (n529,n530,n531);
xor (n530,n528,n437);
and (n531,n532,n441);
and (n532,n22,n55);
and (n533,n143,n121);
or (n534,n535,n538);
and (n535,n536,n537);
xor (n536,n491,n492);
and (n537,n115,n121);
and (n538,n539,n540);
xor (n539,n536,n537);
or (n540,n541,n544);
and (n541,n542,n543);
xor (n542,n497,n498);
and (n543,n86,n121);
and (n544,n545,n546);
xor (n545,n542,n543);
or (n546,n547,n550);
and (n547,n548,n549);
xor (n548,n502,n503);
and (n549,n80,n121);
and (n550,n551,n552);
xor (n551,n548,n549);
or (n552,n553,n556);
and (n553,n554,n555);
xor (n554,n507,n508);
and (n555,n97,n121);
and (n556,n557,n558);
xor (n557,n554,n555);
or (n558,n559,n562);
and (n559,n560,n561);
xor (n560,n513,n514);
and (n561,n182,n121);
and (n562,n563,n564);
xor (n563,n560,n561);
or (n564,n565,n568);
and (n565,n566,n567);
xor (n566,n519,n520);
and (n567,n42,n121);
and (n568,n569,n570);
xor (n569,n566,n567);
or (n570,n571,n574);
and (n571,n572,n573);
xor (n572,n525,n526);
and (n573,n22,n121);
and (n574,n575,n576);
xor (n575,n572,n573);
and (n576,n577,n412);
xor (n577,n530,n531);
and (n578,n115,n70);
or (n579,n580,n583);
and (n580,n581,n582);
xor (n581,n539,n540);
and (n582,n86,n70);
and (n583,n584,n585);
xor (n584,n581,n582);
or (n585,n586,n589);
and (n586,n587,n588);
xor (n587,n545,n546);
and (n588,n80,n70);
and (n589,n590,n591);
xor (n590,n587,n588);
or (n591,n592,n595);
and (n592,n593,n594);
xor (n593,n551,n552);
and (n594,n97,n70);
and (n595,n596,n597);
xor (n596,n593,n594);
or (n597,n598,n600);
and (n598,n599,n311);
xor (n599,n557,n558);
and (n600,n601,n602);
xor (n601,n599,n311);
or (n602,n603,n606);
and (n603,n604,n605);
xor (n604,n563,n564);
and (n605,n42,n70);
and (n606,n607,n608);
xor (n607,n604,n605);
or (n608,n609,n611);
and (n609,n610,n385);
xor (n610,n569,n570);
and (n611,n612,n613);
xor (n612,n610,n385);
and (n613,n614,n615);
xor (n614,n575,n576);
and (n615,n105,n70);
and (n616,n86,n68);
or (n617,n618,n621);
and (n618,n619,n620);
xor (n619,n584,n585);
and (n620,n80,n68);
and (n621,n622,n623);
xor (n622,n619,n620);
or (n623,n624,n627);
and (n624,n625,n626);
xor (n625,n590,n591);
and (n626,n97,n68);
and (n627,n628,n629);
xor (n628,n625,n626);
or (n629,n630,n633);
and (n630,n631,n632);
xor (n631,n596,n597);
and (n632,n182,n68);
and (n633,n634,n635);
xor (n634,n631,n632);
or (n635,n636,n639);
and (n636,n637,n638);
xor (n637,n601,n602);
and (n638,n42,n68);
and (n639,n640,n641);
xor (n640,n637,n638);
or (n641,n642,n645);
and (n642,n643,n644);
xor (n643,n607,n608);
and (n644,n22,n68);
and (n645,n646,n647);
xor (n646,n643,n644);
and (n647,n648,n340);
xor (n648,n612,n613);
and (n649,n80,n75);
or (n650,n651,n654);
and (n651,n652,n653);
xor (n652,n622,n623);
and (n653,n97,n75);
and (n654,n655,n656);
xor (n655,n652,n653);
or (n656,n657,n660);
and (n657,n658,n659);
xor (n658,n628,n629);
and (n659,n182,n75);
and (n660,n661,n662);
xor (n661,n658,n659);
or (n662,n663,n666);
and (n663,n664,n665);
xor (n664,n634,n635);
and (n665,n42,n75);
and (n666,n667,n668);
xor (n667,n664,n665);
or (n668,n669,n671);
and (n669,n670,n332);
xor (n670,n640,n641);
and (n671,n672,n673);
xor (n672,n670,n332);
and (n673,n674,n675);
xor (n674,n646,n647);
and (n675,n105,n75);
and (n676,n97,n154);
or (n677,n678,n681);
and (n678,n679,n680);
xor (n679,n655,n656);
and (n680,n182,n154);
and (n681,n682,n683);
xor (n682,n679,n680);
or (n683,n684,n687);
and (n684,n685,n686);
xor (n685,n661,n662);
and (n686,n42,n154);
and (n687,n688,n689);
xor (n688,n685,n686);
or (n689,n690,n693);
and (n690,n691,n692);
xor (n691,n667,n668);
and (n692,n22,n154);
and (n693,n694,n695);
xor (n694,n691,n692);
and (n695,n696,n242);
xor (n696,n672,n673);
or (n697,n698,n700);
and (n698,n699,n166);
xor (n699,n682,n683);
and (n700,n701,n702);
xor (n701,n699,n166);
or (n702,n703,n706);
and (n703,n704,n705);
xor (n704,n688,n689);
and (n705,n22,n31);
and (n706,n707,n708);
xor (n707,n704,n705);
and (n708,n709,n710);
xor (n709,n694,n695);
and (n710,n105,n31);
and (n711,n42,n32);
or (n712,n713,n716);
and (n713,n714,n715);
xor (n714,n701,n702);
and (n715,n22,n32);
and (n716,n717,n718);
xor (n717,n714,n715);
and (n718,n719,n108);
xor (n719,n707,n708);
and (n720,n721,n722);
xor (n721,n717,n718);
and (n722,n105,n24);
and (n723,n105,n202);
endmodule
