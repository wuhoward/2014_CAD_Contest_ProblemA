module top (out,n23,n24,n28,n30,n37,n44,n51,n58,n65
        ,n72,n79,n86,n93,n99,n101,n168,n235,n302,n369
        ,n436,n503,n568,n627,n680,n748,n749,n753,n755,n762
        ,n769,n776,n783,n790,n797,n804,n811,n818,n824,n826
        ,n893,n960,n1027,n1094,n1161,n1228,n1293,n1352,n1405,n1451);
output out;
input n23;
input n24;
input n28;
input n30;
input n37;
input n44;
input n51;
input n58;
input n65;
input n72;
input n79;
input n86;
input n93;
input n99;
input n101;
input n168;
input n235;
input n302;
input n369;
input n436;
input n503;
input n568;
input n627;
input n680;
input n748;
input n749;
input n753;
input n755;
input n762;
input n769;
input n776;
input n783;
input n790;
input n797;
input n804;
input n811;
input n818;
input n824;
input n826;
input n893;
input n960;
input n1027;
input n1094;
input n1161;
input n1228;
input n1293;
input n1352;
input n1405;
input n1451;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n25;
wire n26;
wire n27;
wire n29;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n100;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n750;
wire n751;
wire n752;
wire n754;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n825;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
xor (out,n0,n1452);
wire s0n0,s1n0,notn0;
or (n0,s0n0,s1n0);
not(notn0,n1451);
and (s0n0,notn0,n1);
and (s1n0,n1451,n726);
xor (n1,n2,n681);
xor (n2,n3,n679);
xor (n3,n4,n628);
xor (n4,n5,n626);
xor (n5,n6,n569);
xor (n6,n7,n567);
xor (n7,n8,n504);
xor (n8,n9,n502);
or (n9,n10,n437);
and (n10,n11,n435);
or (n11,n12,n370);
and (n12,n13,n368);
or (n13,n14,n303);
and (n14,n15,n301);
or (n15,n16,n236);
and (n16,n17,n234);
or (n17,n18,n169);
and (n18,n19,n167);
or (n19,n20,n102);
and (n20,n21,n100);
and (n21,n22,n25);
and (n22,n23,n24);
or (n25,n26,n31);
and (n26,n27,n29);
and (n27,n23,n28);
and (n29,n30,n24);
and (n31,n32,n33);
xor (n32,n27,n29);
or (n33,n34,n38);
and (n34,n35,n36);
and (n35,n30,n28);
and (n36,n37,n24);
and (n38,n39,n40);
xor (n39,n35,n36);
or (n40,n41,n45);
and (n41,n42,n43);
and (n42,n37,n28);
and (n43,n44,n24);
and (n45,n46,n47);
xor (n46,n42,n43);
or (n47,n48,n52);
and (n48,n49,n50);
and (n49,n44,n28);
and (n50,n51,n24);
and (n52,n53,n54);
xor (n53,n49,n50);
or (n54,n55,n59);
and (n55,n56,n57);
and (n56,n51,n28);
and (n57,n58,n24);
and (n59,n60,n61);
xor (n60,n56,n57);
or (n61,n62,n66);
and (n62,n63,n64);
and (n63,n58,n28);
and (n64,n65,n24);
and (n66,n67,n68);
xor (n67,n63,n64);
or (n68,n69,n73);
and (n69,n70,n71);
and (n70,n65,n28);
and (n71,n72,n24);
and (n73,n74,n75);
xor (n74,n70,n71);
or (n75,n76,n80);
and (n76,n77,n78);
and (n77,n72,n28);
and (n78,n79,n24);
and (n80,n81,n82);
xor (n81,n77,n78);
or (n82,n83,n87);
and (n83,n84,n85);
and (n84,n79,n28);
and (n85,n86,n24);
and (n87,n88,n89);
xor (n88,n84,n85);
or (n89,n90,n94);
and (n90,n91,n92);
and (n91,n86,n28);
and (n92,n93,n24);
and (n94,n95,n96);
xor (n95,n91,n92);
and (n96,n97,n98);
and (n97,n93,n28);
and (n98,n99,n24);
and (n100,n23,n101);
and (n102,n103,n104);
xor (n103,n21,n100);
or (n104,n105,n108);
and (n105,n106,n107);
xor (n106,n22,n25);
and (n107,n30,n101);
and (n108,n109,n110);
xor (n109,n106,n107);
or (n110,n111,n114);
and (n111,n112,n113);
xor (n112,n32,n33);
and (n113,n37,n101);
and (n114,n115,n116);
xor (n115,n112,n113);
or (n116,n117,n120);
and (n117,n118,n119);
xor (n118,n39,n40);
and (n119,n44,n101);
and (n120,n121,n122);
xor (n121,n118,n119);
or (n122,n123,n126);
and (n123,n124,n125);
xor (n124,n46,n47);
and (n125,n51,n101);
and (n126,n127,n128);
xor (n127,n124,n125);
or (n128,n129,n132);
and (n129,n130,n131);
xor (n130,n53,n54);
and (n131,n58,n101);
and (n132,n133,n134);
xor (n133,n130,n131);
or (n134,n135,n138);
and (n135,n136,n137);
xor (n136,n60,n61);
and (n137,n65,n101);
and (n138,n139,n140);
xor (n139,n136,n137);
or (n140,n141,n144);
and (n141,n142,n143);
xor (n142,n67,n68);
and (n143,n72,n101);
and (n144,n145,n146);
xor (n145,n142,n143);
or (n146,n147,n150);
and (n147,n148,n149);
xor (n148,n74,n75);
and (n149,n79,n101);
and (n150,n151,n152);
xor (n151,n148,n149);
or (n152,n153,n156);
and (n153,n154,n155);
xor (n154,n81,n82);
and (n155,n86,n101);
and (n156,n157,n158);
xor (n157,n154,n155);
or (n158,n159,n162);
and (n159,n160,n161);
xor (n160,n88,n89);
and (n161,n93,n101);
and (n162,n163,n164);
xor (n163,n160,n161);
and (n164,n165,n166);
xor (n165,n95,n96);
and (n166,n99,n101);
and (n167,n23,n168);
and (n169,n170,n171);
xor (n170,n19,n167);
or (n171,n172,n175);
and (n172,n173,n174);
xor (n173,n103,n104);
and (n174,n30,n168);
and (n175,n176,n177);
xor (n176,n173,n174);
or (n177,n178,n181);
and (n178,n179,n180);
xor (n179,n109,n110);
and (n180,n37,n168);
and (n181,n182,n183);
xor (n182,n179,n180);
or (n183,n184,n187);
and (n184,n185,n186);
xor (n185,n115,n116);
and (n186,n44,n168);
and (n187,n188,n189);
xor (n188,n185,n186);
or (n189,n190,n193);
and (n190,n191,n192);
xor (n191,n121,n122);
and (n192,n51,n168);
and (n193,n194,n195);
xor (n194,n191,n192);
or (n195,n196,n199);
and (n196,n197,n198);
xor (n197,n127,n128);
and (n198,n58,n168);
and (n199,n200,n201);
xor (n200,n197,n198);
or (n201,n202,n205);
and (n202,n203,n204);
xor (n203,n133,n134);
and (n204,n65,n168);
and (n205,n206,n207);
xor (n206,n203,n204);
or (n207,n208,n211);
and (n208,n209,n210);
xor (n209,n139,n140);
and (n210,n72,n168);
and (n211,n212,n213);
xor (n212,n209,n210);
or (n213,n214,n217);
and (n214,n215,n216);
xor (n215,n145,n146);
and (n216,n79,n168);
and (n217,n218,n219);
xor (n218,n215,n216);
or (n219,n220,n223);
and (n220,n221,n222);
xor (n221,n151,n152);
and (n222,n86,n168);
and (n223,n224,n225);
xor (n224,n221,n222);
or (n225,n226,n229);
and (n226,n227,n228);
xor (n227,n157,n158);
and (n228,n93,n168);
and (n229,n230,n231);
xor (n230,n227,n228);
and (n231,n232,n233);
xor (n232,n163,n164);
and (n233,n99,n168);
and (n234,n23,n235);
and (n236,n237,n238);
xor (n237,n17,n234);
or (n238,n239,n242);
and (n239,n240,n241);
xor (n240,n170,n171);
and (n241,n30,n235);
and (n242,n243,n244);
xor (n243,n240,n241);
or (n244,n245,n248);
and (n245,n246,n247);
xor (n246,n176,n177);
and (n247,n37,n235);
and (n248,n249,n250);
xor (n249,n246,n247);
or (n250,n251,n254);
and (n251,n252,n253);
xor (n252,n182,n183);
and (n253,n44,n235);
and (n254,n255,n256);
xor (n255,n252,n253);
or (n256,n257,n260);
and (n257,n258,n259);
xor (n258,n188,n189);
and (n259,n51,n235);
and (n260,n261,n262);
xor (n261,n258,n259);
or (n262,n263,n266);
and (n263,n264,n265);
xor (n264,n194,n195);
and (n265,n58,n235);
and (n266,n267,n268);
xor (n267,n264,n265);
or (n268,n269,n272);
and (n269,n270,n271);
xor (n270,n200,n201);
and (n271,n65,n235);
and (n272,n273,n274);
xor (n273,n270,n271);
or (n274,n275,n278);
and (n275,n276,n277);
xor (n276,n206,n207);
and (n277,n72,n235);
and (n278,n279,n280);
xor (n279,n276,n277);
or (n280,n281,n284);
and (n281,n282,n283);
xor (n282,n212,n213);
and (n283,n79,n235);
and (n284,n285,n286);
xor (n285,n282,n283);
or (n286,n287,n290);
and (n287,n288,n289);
xor (n288,n218,n219);
and (n289,n86,n235);
and (n290,n291,n292);
xor (n291,n288,n289);
or (n292,n293,n296);
and (n293,n294,n295);
xor (n294,n224,n225);
and (n295,n93,n235);
and (n296,n297,n298);
xor (n297,n294,n295);
and (n298,n299,n300);
xor (n299,n230,n231);
and (n300,n99,n235);
and (n301,n23,n302);
and (n303,n304,n305);
xor (n304,n15,n301);
or (n305,n306,n309);
and (n306,n307,n308);
xor (n307,n237,n238);
and (n308,n30,n302);
and (n309,n310,n311);
xor (n310,n307,n308);
or (n311,n312,n315);
and (n312,n313,n314);
xor (n313,n243,n244);
and (n314,n37,n302);
and (n315,n316,n317);
xor (n316,n313,n314);
or (n317,n318,n321);
and (n318,n319,n320);
xor (n319,n249,n250);
and (n320,n44,n302);
and (n321,n322,n323);
xor (n322,n319,n320);
or (n323,n324,n327);
and (n324,n325,n326);
xor (n325,n255,n256);
and (n326,n51,n302);
and (n327,n328,n329);
xor (n328,n325,n326);
or (n329,n330,n333);
and (n330,n331,n332);
xor (n331,n261,n262);
and (n332,n58,n302);
and (n333,n334,n335);
xor (n334,n331,n332);
or (n335,n336,n339);
and (n336,n337,n338);
xor (n337,n267,n268);
and (n338,n65,n302);
and (n339,n340,n341);
xor (n340,n337,n338);
or (n341,n342,n345);
and (n342,n343,n344);
xor (n343,n273,n274);
and (n344,n72,n302);
and (n345,n346,n347);
xor (n346,n343,n344);
or (n347,n348,n351);
and (n348,n349,n350);
xor (n349,n279,n280);
and (n350,n79,n302);
and (n351,n352,n353);
xor (n352,n349,n350);
or (n353,n354,n357);
and (n354,n355,n356);
xor (n355,n285,n286);
and (n356,n86,n302);
and (n357,n358,n359);
xor (n358,n355,n356);
or (n359,n360,n363);
and (n360,n361,n362);
xor (n361,n291,n292);
and (n362,n93,n302);
and (n363,n364,n365);
xor (n364,n361,n362);
and (n365,n366,n367);
xor (n366,n297,n298);
and (n367,n99,n302);
and (n368,n23,n369);
and (n370,n371,n372);
xor (n371,n13,n368);
or (n372,n373,n376);
and (n373,n374,n375);
xor (n374,n304,n305);
and (n375,n30,n369);
and (n376,n377,n378);
xor (n377,n374,n375);
or (n378,n379,n382);
and (n379,n380,n381);
xor (n380,n310,n311);
and (n381,n37,n369);
and (n382,n383,n384);
xor (n383,n380,n381);
or (n384,n385,n388);
and (n385,n386,n387);
xor (n386,n316,n317);
and (n387,n44,n369);
and (n388,n389,n390);
xor (n389,n386,n387);
or (n390,n391,n394);
and (n391,n392,n393);
xor (n392,n322,n323);
and (n393,n51,n369);
and (n394,n395,n396);
xor (n395,n392,n393);
or (n396,n397,n400);
and (n397,n398,n399);
xor (n398,n328,n329);
and (n399,n58,n369);
and (n400,n401,n402);
xor (n401,n398,n399);
or (n402,n403,n406);
and (n403,n404,n405);
xor (n404,n334,n335);
and (n405,n65,n369);
and (n406,n407,n408);
xor (n407,n404,n405);
or (n408,n409,n412);
and (n409,n410,n411);
xor (n410,n340,n341);
and (n411,n72,n369);
and (n412,n413,n414);
xor (n413,n410,n411);
or (n414,n415,n418);
and (n415,n416,n417);
xor (n416,n346,n347);
and (n417,n79,n369);
and (n418,n419,n420);
xor (n419,n416,n417);
or (n420,n421,n424);
and (n421,n422,n423);
xor (n422,n352,n353);
and (n423,n86,n369);
and (n424,n425,n426);
xor (n425,n422,n423);
or (n426,n427,n430);
and (n427,n428,n429);
xor (n428,n358,n359);
and (n429,n93,n369);
and (n430,n431,n432);
xor (n431,n428,n429);
and (n432,n433,n434);
xor (n433,n364,n365);
and (n434,n99,n369);
and (n435,n23,n436);
and (n437,n438,n439);
xor (n438,n11,n435);
or (n439,n440,n443);
and (n440,n441,n442);
xor (n441,n371,n372);
and (n442,n30,n436);
and (n443,n444,n445);
xor (n444,n441,n442);
or (n445,n446,n449);
and (n446,n447,n448);
xor (n447,n377,n378);
and (n448,n37,n436);
and (n449,n450,n451);
xor (n450,n447,n448);
or (n451,n452,n455);
and (n452,n453,n454);
xor (n453,n383,n384);
and (n454,n44,n436);
and (n455,n456,n457);
xor (n456,n453,n454);
or (n457,n458,n461);
and (n458,n459,n460);
xor (n459,n389,n390);
and (n460,n51,n436);
and (n461,n462,n463);
xor (n462,n459,n460);
or (n463,n464,n467);
and (n464,n465,n466);
xor (n465,n395,n396);
and (n466,n58,n436);
and (n467,n468,n469);
xor (n468,n465,n466);
or (n469,n470,n473);
and (n470,n471,n472);
xor (n471,n401,n402);
and (n472,n65,n436);
and (n473,n474,n475);
xor (n474,n471,n472);
or (n475,n476,n479);
and (n476,n477,n478);
xor (n477,n407,n408);
and (n478,n72,n436);
and (n479,n480,n481);
xor (n480,n477,n478);
or (n481,n482,n485);
and (n482,n483,n484);
xor (n483,n413,n414);
and (n484,n79,n436);
and (n485,n486,n487);
xor (n486,n483,n484);
or (n487,n488,n491);
and (n488,n489,n490);
xor (n489,n419,n420);
and (n490,n86,n436);
and (n491,n492,n493);
xor (n492,n489,n490);
or (n493,n494,n497);
and (n494,n495,n496);
xor (n495,n425,n426);
and (n496,n93,n436);
and (n497,n498,n499);
xor (n498,n495,n496);
and (n499,n500,n501);
xor (n500,n431,n432);
and (n501,n99,n436);
and (n502,n23,n503);
or (n504,n505,n508);
and (n505,n506,n507);
xor (n506,n438,n439);
and (n507,n30,n503);
and (n508,n509,n510);
xor (n509,n506,n507);
or (n510,n511,n514);
and (n511,n512,n513);
xor (n512,n444,n445);
and (n513,n37,n503);
and (n514,n515,n516);
xor (n515,n512,n513);
or (n516,n517,n520);
and (n517,n518,n519);
xor (n518,n450,n451);
and (n519,n44,n503);
and (n520,n521,n522);
xor (n521,n518,n519);
or (n522,n523,n526);
and (n523,n524,n525);
xor (n524,n456,n457);
and (n525,n51,n503);
and (n526,n527,n528);
xor (n527,n524,n525);
or (n528,n529,n532);
and (n529,n530,n531);
xor (n530,n462,n463);
and (n531,n58,n503);
and (n532,n533,n534);
xor (n533,n530,n531);
or (n534,n535,n538);
and (n535,n536,n537);
xor (n536,n468,n469);
and (n537,n65,n503);
and (n538,n539,n540);
xor (n539,n536,n537);
or (n540,n541,n544);
and (n541,n542,n543);
xor (n542,n474,n475);
and (n543,n72,n503);
and (n544,n545,n546);
xor (n545,n542,n543);
or (n546,n547,n550);
and (n547,n548,n549);
xor (n548,n480,n481);
and (n549,n79,n503);
and (n550,n551,n552);
xor (n551,n548,n549);
or (n552,n553,n556);
and (n553,n554,n555);
xor (n554,n486,n487);
and (n555,n86,n503);
and (n556,n557,n558);
xor (n557,n554,n555);
or (n558,n559,n562);
and (n559,n560,n561);
xor (n560,n492,n493);
and (n561,n93,n503);
and (n562,n563,n564);
xor (n563,n560,n561);
and (n564,n565,n566);
xor (n565,n498,n499);
and (n566,n99,n503);
and (n567,n30,n568);
or (n569,n570,n573);
and (n570,n571,n572);
xor (n571,n509,n510);
and (n572,n37,n568);
and (n573,n574,n575);
xor (n574,n571,n572);
or (n575,n576,n579);
and (n576,n577,n578);
xor (n577,n515,n516);
and (n578,n44,n568);
and (n579,n580,n581);
xor (n580,n577,n578);
or (n581,n582,n585);
and (n582,n583,n584);
xor (n583,n521,n522);
and (n584,n51,n568);
and (n585,n586,n587);
xor (n586,n583,n584);
or (n587,n588,n591);
and (n588,n589,n590);
xor (n589,n527,n528);
and (n590,n58,n568);
and (n591,n592,n593);
xor (n592,n589,n590);
or (n593,n594,n597);
and (n594,n595,n596);
xor (n595,n533,n534);
and (n596,n65,n568);
and (n597,n598,n599);
xor (n598,n595,n596);
or (n599,n600,n603);
and (n600,n601,n602);
xor (n601,n539,n540);
and (n602,n72,n568);
and (n603,n604,n605);
xor (n604,n601,n602);
or (n605,n606,n609);
and (n606,n607,n608);
xor (n607,n545,n546);
and (n608,n79,n568);
and (n609,n610,n611);
xor (n610,n607,n608);
or (n611,n612,n615);
and (n612,n613,n614);
xor (n613,n551,n552);
and (n614,n86,n568);
and (n615,n616,n617);
xor (n616,n613,n614);
or (n617,n618,n621);
and (n618,n619,n620);
xor (n619,n557,n558);
and (n620,n93,n568);
and (n621,n622,n623);
xor (n622,n619,n620);
and (n623,n624,n625);
xor (n624,n563,n564);
and (n625,n99,n568);
and (n626,n37,n627);
or (n628,n629,n632);
and (n629,n630,n631);
xor (n630,n574,n575);
and (n631,n44,n627);
and (n632,n633,n634);
xor (n633,n630,n631);
or (n634,n635,n638);
and (n635,n636,n637);
xor (n636,n580,n581);
and (n637,n51,n627);
and (n638,n639,n640);
xor (n639,n636,n637);
or (n640,n641,n644);
and (n641,n642,n643);
xor (n642,n586,n587);
and (n643,n58,n627);
and (n644,n645,n646);
xor (n645,n642,n643);
or (n646,n647,n650);
and (n647,n648,n649);
xor (n648,n592,n593);
and (n649,n65,n627);
and (n650,n651,n652);
xor (n651,n648,n649);
or (n652,n653,n656);
and (n653,n654,n655);
xor (n654,n598,n599);
and (n655,n72,n627);
and (n656,n657,n658);
xor (n657,n654,n655);
or (n658,n659,n662);
and (n659,n660,n661);
xor (n660,n604,n605);
and (n661,n79,n627);
and (n662,n663,n664);
xor (n663,n660,n661);
or (n664,n665,n668);
and (n665,n666,n667);
xor (n666,n610,n611);
and (n667,n86,n627);
and (n668,n669,n670);
xor (n669,n666,n667);
or (n670,n671,n674);
and (n671,n672,n673);
xor (n672,n616,n617);
and (n673,n93,n627);
and (n674,n675,n676);
xor (n675,n672,n673);
and (n676,n677,n678);
xor (n677,n622,n623);
and (n678,n99,n627);
and (n679,n44,n680);
or (n681,n682,n685);
and (n682,n683,n684);
xor (n683,n633,n634);
and (n684,n51,n680);
and (n685,n686,n687);
xor (n686,n683,n684);
or (n687,n688,n691);
and (n688,n689,n690);
xor (n689,n639,n640);
and (n690,n58,n680);
and (n691,n692,n693);
xor (n692,n689,n690);
or (n693,n694,n697);
and (n694,n695,n696);
xor (n695,n645,n646);
and (n696,n65,n680);
and (n697,n698,n699);
xor (n698,n695,n696);
or (n699,n700,n703);
and (n700,n701,n702);
xor (n701,n651,n652);
and (n702,n72,n680);
and (n703,n704,n705);
xor (n704,n701,n702);
or (n705,n706,n709);
and (n706,n707,n708);
xor (n707,n657,n658);
and (n708,n79,n680);
and (n709,n710,n711);
xor (n710,n707,n708);
or (n711,n712,n715);
and (n712,n713,n714);
xor (n713,n663,n664);
and (n714,n86,n680);
and (n715,n716,n717);
xor (n716,n713,n714);
or (n717,n718,n721);
and (n718,n719,n720);
xor (n719,n669,n670);
and (n720,n93,n680);
and (n721,n722,n723);
xor (n722,n719,n720);
and (n723,n724,n725);
xor (n724,n675,n676);
and (n725,n99,n680);
xor (n726,n727,n1406);
xor (n727,n728,n1404);
xor (n728,n729,n1353);
xor (n729,n730,n1351);
xor (n730,n731,n1294);
xor (n731,n732,n1292);
xor (n732,n733,n1229);
xor (n733,n734,n1227);
or (n734,n735,n1162);
and (n735,n736,n1160);
or (n736,n737,n1095);
and (n737,n738,n1093);
or (n738,n739,n1028);
and (n739,n740,n1026);
or (n740,n741,n961);
and (n741,n742,n959);
or (n742,n743,n894);
and (n743,n744,n892);
or (n744,n745,n827);
and (n745,n746,n825);
and (n746,n747,n750);
and (n747,n748,n749);
or (n750,n751,n756);
and (n751,n752,n754);
and (n752,n748,n753);
and (n754,n755,n749);
and (n756,n757,n758);
xor (n757,n752,n754);
or (n758,n759,n763);
and (n759,n760,n761);
and (n760,n755,n753);
and (n761,n762,n749);
and (n763,n764,n765);
xor (n764,n760,n761);
or (n765,n766,n770);
and (n766,n767,n768);
and (n767,n762,n753);
and (n768,n769,n749);
and (n770,n771,n772);
xor (n771,n767,n768);
or (n772,n773,n777);
and (n773,n774,n775);
and (n774,n769,n753);
and (n775,n776,n749);
and (n777,n778,n779);
xor (n778,n774,n775);
or (n779,n780,n784);
and (n780,n781,n782);
and (n781,n776,n753);
and (n782,n783,n749);
and (n784,n785,n786);
xor (n785,n781,n782);
or (n786,n787,n791);
and (n787,n788,n789);
and (n788,n783,n753);
and (n789,n790,n749);
and (n791,n792,n793);
xor (n792,n788,n789);
or (n793,n794,n798);
and (n794,n795,n796);
and (n795,n790,n753);
and (n796,n797,n749);
and (n798,n799,n800);
xor (n799,n795,n796);
or (n800,n801,n805);
and (n801,n802,n803);
and (n802,n797,n753);
and (n803,n804,n749);
and (n805,n806,n807);
xor (n806,n802,n803);
or (n807,n808,n812);
and (n808,n809,n810);
and (n809,n804,n753);
and (n810,n811,n749);
and (n812,n813,n814);
xor (n813,n809,n810);
or (n814,n815,n819);
and (n815,n816,n817);
and (n816,n811,n753);
and (n817,n818,n749);
and (n819,n820,n821);
xor (n820,n816,n817);
and (n821,n822,n823);
and (n822,n818,n753);
and (n823,n824,n749);
and (n825,n748,n826);
and (n827,n828,n829);
xor (n828,n746,n825);
or (n829,n830,n833);
and (n830,n831,n832);
xor (n831,n747,n750);
and (n832,n755,n826);
and (n833,n834,n835);
xor (n834,n831,n832);
or (n835,n836,n839);
and (n836,n837,n838);
xor (n837,n757,n758);
and (n838,n762,n826);
and (n839,n840,n841);
xor (n840,n837,n838);
or (n841,n842,n845);
and (n842,n843,n844);
xor (n843,n764,n765);
and (n844,n769,n826);
and (n845,n846,n847);
xor (n846,n843,n844);
or (n847,n848,n851);
and (n848,n849,n850);
xor (n849,n771,n772);
and (n850,n776,n826);
and (n851,n852,n853);
xor (n852,n849,n850);
or (n853,n854,n857);
and (n854,n855,n856);
xor (n855,n778,n779);
and (n856,n783,n826);
and (n857,n858,n859);
xor (n858,n855,n856);
or (n859,n860,n863);
and (n860,n861,n862);
xor (n861,n785,n786);
and (n862,n790,n826);
and (n863,n864,n865);
xor (n864,n861,n862);
or (n865,n866,n869);
and (n866,n867,n868);
xor (n867,n792,n793);
and (n868,n797,n826);
and (n869,n870,n871);
xor (n870,n867,n868);
or (n871,n872,n875);
and (n872,n873,n874);
xor (n873,n799,n800);
and (n874,n804,n826);
and (n875,n876,n877);
xor (n876,n873,n874);
or (n877,n878,n881);
and (n878,n879,n880);
xor (n879,n806,n807);
and (n880,n811,n826);
and (n881,n882,n883);
xor (n882,n879,n880);
or (n883,n884,n887);
and (n884,n885,n886);
xor (n885,n813,n814);
and (n886,n818,n826);
and (n887,n888,n889);
xor (n888,n885,n886);
and (n889,n890,n891);
xor (n890,n820,n821);
and (n891,n824,n826);
and (n892,n748,n893);
and (n894,n895,n896);
xor (n895,n744,n892);
or (n896,n897,n900);
and (n897,n898,n899);
xor (n898,n828,n829);
and (n899,n755,n893);
and (n900,n901,n902);
xor (n901,n898,n899);
or (n902,n903,n906);
and (n903,n904,n905);
xor (n904,n834,n835);
and (n905,n762,n893);
and (n906,n907,n908);
xor (n907,n904,n905);
or (n908,n909,n912);
and (n909,n910,n911);
xor (n910,n840,n841);
and (n911,n769,n893);
and (n912,n913,n914);
xor (n913,n910,n911);
or (n914,n915,n918);
and (n915,n916,n917);
xor (n916,n846,n847);
and (n917,n776,n893);
and (n918,n919,n920);
xor (n919,n916,n917);
or (n920,n921,n924);
and (n921,n922,n923);
xor (n922,n852,n853);
and (n923,n783,n893);
and (n924,n925,n926);
xor (n925,n922,n923);
or (n926,n927,n930);
and (n927,n928,n929);
xor (n928,n858,n859);
and (n929,n790,n893);
and (n930,n931,n932);
xor (n931,n928,n929);
or (n932,n933,n936);
and (n933,n934,n935);
xor (n934,n864,n865);
and (n935,n797,n893);
and (n936,n937,n938);
xor (n937,n934,n935);
or (n938,n939,n942);
and (n939,n940,n941);
xor (n940,n870,n871);
and (n941,n804,n893);
and (n942,n943,n944);
xor (n943,n940,n941);
or (n944,n945,n948);
and (n945,n946,n947);
xor (n946,n876,n877);
and (n947,n811,n893);
and (n948,n949,n950);
xor (n949,n946,n947);
or (n950,n951,n954);
and (n951,n952,n953);
xor (n952,n882,n883);
and (n953,n818,n893);
and (n954,n955,n956);
xor (n955,n952,n953);
and (n956,n957,n958);
xor (n957,n888,n889);
and (n958,n824,n893);
and (n959,n748,n960);
and (n961,n962,n963);
xor (n962,n742,n959);
or (n963,n964,n967);
and (n964,n965,n966);
xor (n965,n895,n896);
and (n966,n755,n960);
and (n967,n968,n969);
xor (n968,n965,n966);
or (n969,n970,n973);
and (n970,n971,n972);
xor (n971,n901,n902);
and (n972,n762,n960);
and (n973,n974,n975);
xor (n974,n971,n972);
or (n975,n976,n979);
and (n976,n977,n978);
xor (n977,n907,n908);
and (n978,n769,n960);
and (n979,n980,n981);
xor (n980,n977,n978);
or (n981,n982,n985);
and (n982,n983,n984);
xor (n983,n913,n914);
and (n984,n776,n960);
and (n985,n986,n987);
xor (n986,n983,n984);
or (n987,n988,n991);
and (n988,n989,n990);
xor (n989,n919,n920);
and (n990,n783,n960);
and (n991,n992,n993);
xor (n992,n989,n990);
or (n993,n994,n997);
and (n994,n995,n996);
xor (n995,n925,n926);
and (n996,n790,n960);
and (n997,n998,n999);
xor (n998,n995,n996);
or (n999,n1000,n1003);
and (n1000,n1001,n1002);
xor (n1001,n931,n932);
and (n1002,n797,n960);
and (n1003,n1004,n1005);
xor (n1004,n1001,n1002);
or (n1005,n1006,n1009);
and (n1006,n1007,n1008);
xor (n1007,n937,n938);
and (n1008,n804,n960);
and (n1009,n1010,n1011);
xor (n1010,n1007,n1008);
or (n1011,n1012,n1015);
and (n1012,n1013,n1014);
xor (n1013,n943,n944);
and (n1014,n811,n960);
and (n1015,n1016,n1017);
xor (n1016,n1013,n1014);
or (n1017,n1018,n1021);
and (n1018,n1019,n1020);
xor (n1019,n949,n950);
and (n1020,n818,n960);
and (n1021,n1022,n1023);
xor (n1022,n1019,n1020);
and (n1023,n1024,n1025);
xor (n1024,n955,n956);
and (n1025,n824,n960);
and (n1026,n748,n1027);
and (n1028,n1029,n1030);
xor (n1029,n740,n1026);
or (n1030,n1031,n1034);
and (n1031,n1032,n1033);
xor (n1032,n962,n963);
and (n1033,n755,n1027);
and (n1034,n1035,n1036);
xor (n1035,n1032,n1033);
or (n1036,n1037,n1040);
and (n1037,n1038,n1039);
xor (n1038,n968,n969);
and (n1039,n762,n1027);
and (n1040,n1041,n1042);
xor (n1041,n1038,n1039);
or (n1042,n1043,n1046);
and (n1043,n1044,n1045);
xor (n1044,n974,n975);
and (n1045,n769,n1027);
and (n1046,n1047,n1048);
xor (n1047,n1044,n1045);
or (n1048,n1049,n1052);
and (n1049,n1050,n1051);
xor (n1050,n980,n981);
and (n1051,n776,n1027);
and (n1052,n1053,n1054);
xor (n1053,n1050,n1051);
or (n1054,n1055,n1058);
and (n1055,n1056,n1057);
xor (n1056,n986,n987);
and (n1057,n783,n1027);
and (n1058,n1059,n1060);
xor (n1059,n1056,n1057);
or (n1060,n1061,n1064);
and (n1061,n1062,n1063);
xor (n1062,n992,n993);
and (n1063,n790,n1027);
and (n1064,n1065,n1066);
xor (n1065,n1062,n1063);
or (n1066,n1067,n1070);
and (n1067,n1068,n1069);
xor (n1068,n998,n999);
and (n1069,n797,n1027);
and (n1070,n1071,n1072);
xor (n1071,n1068,n1069);
or (n1072,n1073,n1076);
and (n1073,n1074,n1075);
xor (n1074,n1004,n1005);
and (n1075,n804,n1027);
and (n1076,n1077,n1078);
xor (n1077,n1074,n1075);
or (n1078,n1079,n1082);
and (n1079,n1080,n1081);
xor (n1080,n1010,n1011);
and (n1081,n811,n1027);
and (n1082,n1083,n1084);
xor (n1083,n1080,n1081);
or (n1084,n1085,n1088);
and (n1085,n1086,n1087);
xor (n1086,n1016,n1017);
and (n1087,n818,n1027);
and (n1088,n1089,n1090);
xor (n1089,n1086,n1087);
and (n1090,n1091,n1092);
xor (n1091,n1022,n1023);
and (n1092,n824,n1027);
and (n1093,n748,n1094);
and (n1095,n1096,n1097);
xor (n1096,n738,n1093);
or (n1097,n1098,n1101);
and (n1098,n1099,n1100);
xor (n1099,n1029,n1030);
and (n1100,n755,n1094);
and (n1101,n1102,n1103);
xor (n1102,n1099,n1100);
or (n1103,n1104,n1107);
and (n1104,n1105,n1106);
xor (n1105,n1035,n1036);
and (n1106,n762,n1094);
and (n1107,n1108,n1109);
xor (n1108,n1105,n1106);
or (n1109,n1110,n1113);
and (n1110,n1111,n1112);
xor (n1111,n1041,n1042);
and (n1112,n769,n1094);
and (n1113,n1114,n1115);
xor (n1114,n1111,n1112);
or (n1115,n1116,n1119);
and (n1116,n1117,n1118);
xor (n1117,n1047,n1048);
and (n1118,n776,n1094);
and (n1119,n1120,n1121);
xor (n1120,n1117,n1118);
or (n1121,n1122,n1125);
and (n1122,n1123,n1124);
xor (n1123,n1053,n1054);
and (n1124,n783,n1094);
and (n1125,n1126,n1127);
xor (n1126,n1123,n1124);
or (n1127,n1128,n1131);
and (n1128,n1129,n1130);
xor (n1129,n1059,n1060);
and (n1130,n790,n1094);
and (n1131,n1132,n1133);
xor (n1132,n1129,n1130);
or (n1133,n1134,n1137);
and (n1134,n1135,n1136);
xor (n1135,n1065,n1066);
and (n1136,n797,n1094);
and (n1137,n1138,n1139);
xor (n1138,n1135,n1136);
or (n1139,n1140,n1143);
and (n1140,n1141,n1142);
xor (n1141,n1071,n1072);
and (n1142,n804,n1094);
and (n1143,n1144,n1145);
xor (n1144,n1141,n1142);
or (n1145,n1146,n1149);
and (n1146,n1147,n1148);
xor (n1147,n1077,n1078);
and (n1148,n811,n1094);
and (n1149,n1150,n1151);
xor (n1150,n1147,n1148);
or (n1151,n1152,n1155);
and (n1152,n1153,n1154);
xor (n1153,n1083,n1084);
and (n1154,n818,n1094);
and (n1155,n1156,n1157);
xor (n1156,n1153,n1154);
and (n1157,n1158,n1159);
xor (n1158,n1089,n1090);
and (n1159,n824,n1094);
and (n1160,n748,n1161);
and (n1162,n1163,n1164);
xor (n1163,n736,n1160);
or (n1164,n1165,n1168);
and (n1165,n1166,n1167);
xor (n1166,n1096,n1097);
and (n1167,n755,n1161);
and (n1168,n1169,n1170);
xor (n1169,n1166,n1167);
or (n1170,n1171,n1174);
and (n1171,n1172,n1173);
xor (n1172,n1102,n1103);
and (n1173,n762,n1161);
and (n1174,n1175,n1176);
xor (n1175,n1172,n1173);
or (n1176,n1177,n1180);
and (n1177,n1178,n1179);
xor (n1178,n1108,n1109);
and (n1179,n769,n1161);
and (n1180,n1181,n1182);
xor (n1181,n1178,n1179);
or (n1182,n1183,n1186);
and (n1183,n1184,n1185);
xor (n1184,n1114,n1115);
and (n1185,n776,n1161);
and (n1186,n1187,n1188);
xor (n1187,n1184,n1185);
or (n1188,n1189,n1192);
and (n1189,n1190,n1191);
xor (n1190,n1120,n1121);
and (n1191,n783,n1161);
and (n1192,n1193,n1194);
xor (n1193,n1190,n1191);
or (n1194,n1195,n1198);
and (n1195,n1196,n1197);
xor (n1196,n1126,n1127);
and (n1197,n790,n1161);
and (n1198,n1199,n1200);
xor (n1199,n1196,n1197);
or (n1200,n1201,n1204);
and (n1201,n1202,n1203);
xor (n1202,n1132,n1133);
and (n1203,n797,n1161);
and (n1204,n1205,n1206);
xor (n1205,n1202,n1203);
or (n1206,n1207,n1210);
and (n1207,n1208,n1209);
xor (n1208,n1138,n1139);
and (n1209,n804,n1161);
and (n1210,n1211,n1212);
xor (n1211,n1208,n1209);
or (n1212,n1213,n1216);
and (n1213,n1214,n1215);
xor (n1214,n1144,n1145);
and (n1215,n811,n1161);
and (n1216,n1217,n1218);
xor (n1217,n1214,n1215);
or (n1218,n1219,n1222);
and (n1219,n1220,n1221);
xor (n1220,n1150,n1151);
and (n1221,n818,n1161);
and (n1222,n1223,n1224);
xor (n1223,n1220,n1221);
and (n1224,n1225,n1226);
xor (n1225,n1156,n1157);
and (n1226,n824,n1161);
and (n1227,n748,n1228);
or (n1229,n1230,n1233);
and (n1230,n1231,n1232);
xor (n1231,n1163,n1164);
and (n1232,n755,n1228);
and (n1233,n1234,n1235);
xor (n1234,n1231,n1232);
or (n1235,n1236,n1239);
and (n1236,n1237,n1238);
xor (n1237,n1169,n1170);
and (n1238,n762,n1228);
and (n1239,n1240,n1241);
xor (n1240,n1237,n1238);
or (n1241,n1242,n1245);
and (n1242,n1243,n1244);
xor (n1243,n1175,n1176);
and (n1244,n769,n1228);
and (n1245,n1246,n1247);
xor (n1246,n1243,n1244);
or (n1247,n1248,n1251);
and (n1248,n1249,n1250);
xor (n1249,n1181,n1182);
and (n1250,n776,n1228);
and (n1251,n1252,n1253);
xor (n1252,n1249,n1250);
or (n1253,n1254,n1257);
and (n1254,n1255,n1256);
xor (n1255,n1187,n1188);
and (n1256,n783,n1228);
and (n1257,n1258,n1259);
xor (n1258,n1255,n1256);
or (n1259,n1260,n1263);
and (n1260,n1261,n1262);
xor (n1261,n1193,n1194);
and (n1262,n790,n1228);
and (n1263,n1264,n1265);
xor (n1264,n1261,n1262);
or (n1265,n1266,n1269);
and (n1266,n1267,n1268);
xor (n1267,n1199,n1200);
and (n1268,n797,n1228);
and (n1269,n1270,n1271);
xor (n1270,n1267,n1268);
or (n1271,n1272,n1275);
and (n1272,n1273,n1274);
xor (n1273,n1205,n1206);
and (n1274,n804,n1228);
and (n1275,n1276,n1277);
xor (n1276,n1273,n1274);
or (n1277,n1278,n1281);
and (n1278,n1279,n1280);
xor (n1279,n1211,n1212);
and (n1280,n811,n1228);
and (n1281,n1282,n1283);
xor (n1282,n1279,n1280);
or (n1283,n1284,n1287);
and (n1284,n1285,n1286);
xor (n1285,n1217,n1218);
and (n1286,n818,n1228);
and (n1287,n1288,n1289);
xor (n1288,n1285,n1286);
and (n1289,n1290,n1291);
xor (n1290,n1223,n1224);
and (n1291,n824,n1228);
and (n1292,n755,n1293);
or (n1294,n1295,n1298);
and (n1295,n1296,n1297);
xor (n1296,n1234,n1235);
and (n1297,n762,n1293);
and (n1298,n1299,n1300);
xor (n1299,n1296,n1297);
or (n1300,n1301,n1304);
and (n1301,n1302,n1303);
xor (n1302,n1240,n1241);
and (n1303,n769,n1293);
and (n1304,n1305,n1306);
xor (n1305,n1302,n1303);
or (n1306,n1307,n1310);
and (n1307,n1308,n1309);
xor (n1308,n1246,n1247);
and (n1309,n776,n1293);
and (n1310,n1311,n1312);
xor (n1311,n1308,n1309);
or (n1312,n1313,n1316);
and (n1313,n1314,n1315);
xor (n1314,n1252,n1253);
and (n1315,n783,n1293);
and (n1316,n1317,n1318);
xor (n1317,n1314,n1315);
or (n1318,n1319,n1322);
and (n1319,n1320,n1321);
xor (n1320,n1258,n1259);
and (n1321,n790,n1293);
and (n1322,n1323,n1324);
xor (n1323,n1320,n1321);
or (n1324,n1325,n1328);
and (n1325,n1326,n1327);
xor (n1326,n1264,n1265);
and (n1327,n797,n1293);
and (n1328,n1329,n1330);
xor (n1329,n1326,n1327);
or (n1330,n1331,n1334);
and (n1331,n1332,n1333);
xor (n1332,n1270,n1271);
and (n1333,n804,n1293);
and (n1334,n1335,n1336);
xor (n1335,n1332,n1333);
or (n1336,n1337,n1340);
and (n1337,n1338,n1339);
xor (n1338,n1276,n1277);
and (n1339,n811,n1293);
and (n1340,n1341,n1342);
xor (n1341,n1338,n1339);
or (n1342,n1343,n1346);
and (n1343,n1344,n1345);
xor (n1344,n1282,n1283);
and (n1345,n818,n1293);
and (n1346,n1347,n1348);
xor (n1347,n1344,n1345);
and (n1348,n1349,n1350);
xor (n1349,n1288,n1289);
and (n1350,n824,n1293);
and (n1351,n762,n1352);
or (n1353,n1354,n1357);
and (n1354,n1355,n1356);
xor (n1355,n1299,n1300);
and (n1356,n769,n1352);
and (n1357,n1358,n1359);
xor (n1358,n1355,n1356);
or (n1359,n1360,n1363);
and (n1360,n1361,n1362);
xor (n1361,n1305,n1306);
and (n1362,n776,n1352);
and (n1363,n1364,n1365);
xor (n1364,n1361,n1362);
or (n1365,n1366,n1369);
and (n1366,n1367,n1368);
xor (n1367,n1311,n1312);
and (n1368,n783,n1352);
and (n1369,n1370,n1371);
xor (n1370,n1367,n1368);
or (n1371,n1372,n1375);
and (n1372,n1373,n1374);
xor (n1373,n1317,n1318);
and (n1374,n790,n1352);
and (n1375,n1376,n1377);
xor (n1376,n1373,n1374);
or (n1377,n1378,n1381);
and (n1378,n1379,n1380);
xor (n1379,n1323,n1324);
and (n1380,n797,n1352);
and (n1381,n1382,n1383);
xor (n1382,n1379,n1380);
or (n1383,n1384,n1387);
and (n1384,n1385,n1386);
xor (n1385,n1329,n1330);
and (n1386,n804,n1352);
and (n1387,n1388,n1389);
xor (n1388,n1385,n1386);
or (n1389,n1390,n1393);
and (n1390,n1391,n1392);
xor (n1391,n1335,n1336);
and (n1392,n811,n1352);
and (n1393,n1394,n1395);
xor (n1394,n1391,n1392);
or (n1395,n1396,n1399);
and (n1396,n1397,n1398);
xor (n1397,n1341,n1342);
and (n1398,n818,n1352);
and (n1399,n1400,n1401);
xor (n1400,n1397,n1398);
and (n1401,n1402,n1403);
xor (n1402,n1347,n1348);
and (n1403,n824,n1352);
and (n1404,n769,n1405);
or (n1406,n1407,n1410);
and (n1407,n1408,n1409);
xor (n1408,n1358,n1359);
and (n1409,n776,n1405);
and (n1410,n1411,n1412);
xor (n1411,n1408,n1409);
or (n1412,n1413,n1416);
and (n1413,n1414,n1415);
xor (n1414,n1364,n1365);
and (n1415,n783,n1405);
and (n1416,n1417,n1418);
xor (n1417,n1414,n1415);
or (n1418,n1419,n1422);
and (n1419,n1420,n1421);
xor (n1420,n1370,n1371);
and (n1421,n790,n1405);
and (n1422,n1423,n1424);
xor (n1423,n1420,n1421);
or (n1424,n1425,n1428);
and (n1425,n1426,n1427);
xor (n1426,n1376,n1377);
and (n1427,n797,n1405);
and (n1428,n1429,n1430);
xor (n1429,n1426,n1427);
or (n1430,n1431,n1434);
and (n1431,n1432,n1433);
xor (n1432,n1382,n1383);
and (n1433,n804,n1405);
and (n1434,n1435,n1436);
xor (n1435,n1432,n1433);
or (n1436,n1437,n1440);
and (n1437,n1438,n1439);
xor (n1438,n1388,n1389);
and (n1439,n811,n1405);
and (n1440,n1441,n1442);
xor (n1441,n1438,n1439);
or (n1442,n1443,n1446);
and (n1443,n1444,n1445);
xor (n1444,n1394,n1395);
and (n1445,n818,n1405);
and (n1446,n1447,n1448);
xor (n1447,n1444,n1445);
and (n1448,n1449,n1450);
xor (n1449,n1400,n1401);
and (n1450,n824,n1405);
xor (n1452,n1453,n2132);
xor (n1453,n1454,n2130);
xor (n1454,n1455,n2079);
xor (n1455,n1456,n2077);
xor (n1456,n1457,n2020);
xor (n1457,n1458,n2018);
xor (n1458,n1459,n1955);
xor (n1459,n1460,n1953);
or (n1460,n1461,n1888);
and (n1461,n1462,n1886);
or (n1462,n1463,n1821);
and (n1463,n1464,n1819);
or (n1464,n1465,n1754);
and (n1465,n1466,n1752);
or (n1466,n1467,n1687);
and (n1467,n1468,n1685);
or (n1468,n1469,n1620);
and (n1469,n1470,n1618);
or (n1470,n1471,n1553);
and (n1471,n1472,n1551);
and (n1472,n1473,n1476);
and (n1473,n1474,n1475);
wire s0n1474,s1n1474,notn1474;
or (n1474,s0n1474,s1n1474);
not(notn1474,n1451);
and (s0n1474,notn1474,n23);
and (s1n1474,n1451,n748);
wire s0n1475,s1n1475,notn1475;
or (n1475,s0n1475,s1n1475);
not(notn1475,n1451);
and (s0n1475,notn1475,n24);
and (s1n1475,n1451,n749);
or (n1476,n1477,n1482);
and (n1477,n1478,n1480);
and (n1478,n1474,n1479);
wire s0n1479,s1n1479,notn1479;
or (n1479,s0n1479,s1n1479);
not(notn1479,n1451);
and (s0n1479,notn1479,n28);
and (s1n1479,n1451,n753);
and (n1480,n1481,n1475);
wire s0n1481,s1n1481,notn1481;
or (n1481,s0n1481,s1n1481);
not(notn1481,n1451);
and (s0n1481,notn1481,n30);
and (s1n1481,n1451,n755);
and (n1482,n1483,n1484);
xor (n1483,n1478,n1480);
or (n1484,n1485,n1489);
and (n1485,n1486,n1487);
and (n1486,n1481,n1479);
and (n1487,n1488,n1475);
wire s0n1488,s1n1488,notn1488;
or (n1488,s0n1488,s1n1488);
not(notn1488,n1451);
and (s0n1488,notn1488,n37);
and (s1n1488,n1451,n762);
and (n1489,n1490,n1491);
xor (n1490,n1486,n1487);
or (n1491,n1492,n1496);
and (n1492,n1493,n1494);
and (n1493,n1488,n1479);
and (n1494,n1495,n1475);
wire s0n1495,s1n1495,notn1495;
or (n1495,s0n1495,s1n1495);
not(notn1495,n1451);
and (s0n1495,notn1495,n44);
and (s1n1495,n1451,n769);
and (n1496,n1497,n1498);
xor (n1497,n1493,n1494);
or (n1498,n1499,n1503);
and (n1499,n1500,n1501);
and (n1500,n1495,n1479);
and (n1501,n1502,n1475);
wire s0n1502,s1n1502,notn1502;
or (n1502,s0n1502,s1n1502);
not(notn1502,n1451);
and (s0n1502,notn1502,n51);
and (s1n1502,n1451,n776);
and (n1503,n1504,n1505);
xor (n1504,n1500,n1501);
or (n1505,n1506,n1510);
and (n1506,n1507,n1508);
and (n1507,n1502,n1479);
and (n1508,n1509,n1475);
wire s0n1509,s1n1509,notn1509;
or (n1509,s0n1509,s1n1509);
not(notn1509,n1451);
and (s0n1509,notn1509,n58);
and (s1n1509,n1451,n783);
and (n1510,n1511,n1512);
xor (n1511,n1507,n1508);
or (n1512,n1513,n1517);
and (n1513,n1514,n1515);
and (n1514,n1509,n1479);
and (n1515,n1516,n1475);
wire s0n1516,s1n1516,notn1516;
or (n1516,s0n1516,s1n1516);
not(notn1516,n1451);
and (s0n1516,notn1516,n65);
and (s1n1516,n1451,n790);
and (n1517,n1518,n1519);
xor (n1518,n1514,n1515);
or (n1519,n1520,n1524);
and (n1520,n1521,n1522);
and (n1521,n1516,n1479);
and (n1522,n1523,n1475);
wire s0n1523,s1n1523,notn1523;
or (n1523,s0n1523,s1n1523);
not(notn1523,n1451);
and (s0n1523,notn1523,n72);
and (s1n1523,n1451,n797);
and (n1524,n1525,n1526);
xor (n1525,n1521,n1522);
or (n1526,n1527,n1531);
and (n1527,n1528,n1529);
and (n1528,n1523,n1479);
and (n1529,n1530,n1475);
wire s0n1530,s1n1530,notn1530;
or (n1530,s0n1530,s1n1530);
not(notn1530,n1451);
and (s0n1530,notn1530,n79);
and (s1n1530,n1451,n804);
and (n1531,n1532,n1533);
xor (n1532,n1528,n1529);
or (n1533,n1534,n1538);
and (n1534,n1535,n1536);
and (n1535,n1530,n1479);
and (n1536,n1537,n1475);
wire s0n1537,s1n1537,notn1537;
or (n1537,s0n1537,s1n1537);
not(notn1537,n1451);
and (s0n1537,notn1537,n86);
and (s1n1537,n1451,n811);
and (n1538,n1539,n1540);
xor (n1539,n1535,n1536);
or (n1540,n1541,n1545);
and (n1541,n1542,n1543);
and (n1542,n1537,n1479);
and (n1543,n1544,n1475);
wire s0n1544,s1n1544,notn1544;
or (n1544,s0n1544,s1n1544);
not(notn1544,n1451);
and (s0n1544,notn1544,n93);
and (s1n1544,n1451,n818);
and (n1545,n1546,n1547);
xor (n1546,n1542,n1543);
and (n1547,n1548,n1549);
and (n1548,n1544,n1479);
and (n1549,n1550,n1475);
wire s0n1550,s1n1550,notn1550;
or (n1550,s0n1550,s1n1550);
not(notn1550,n1451);
and (s0n1550,notn1550,n99);
and (s1n1550,n1451,n824);
and (n1551,n1474,n1552);
wire s0n1552,s1n1552,notn1552;
or (n1552,s0n1552,s1n1552);
not(notn1552,n1451);
and (s0n1552,notn1552,n101);
and (s1n1552,n1451,n826);
and (n1553,n1554,n1555);
xor (n1554,n1472,n1551);
or (n1555,n1556,n1559);
and (n1556,n1557,n1558);
xor (n1557,n1473,n1476);
and (n1558,n1481,n1552);
and (n1559,n1560,n1561);
xor (n1560,n1557,n1558);
or (n1561,n1562,n1565);
and (n1562,n1563,n1564);
xor (n1563,n1483,n1484);
and (n1564,n1488,n1552);
and (n1565,n1566,n1567);
xor (n1566,n1563,n1564);
or (n1567,n1568,n1571);
and (n1568,n1569,n1570);
xor (n1569,n1490,n1491);
and (n1570,n1495,n1552);
and (n1571,n1572,n1573);
xor (n1572,n1569,n1570);
or (n1573,n1574,n1577);
and (n1574,n1575,n1576);
xor (n1575,n1497,n1498);
and (n1576,n1502,n1552);
and (n1577,n1578,n1579);
xor (n1578,n1575,n1576);
or (n1579,n1580,n1583);
and (n1580,n1581,n1582);
xor (n1581,n1504,n1505);
and (n1582,n1509,n1552);
and (n1583,n1584,n1585);
xor (n1584,n1581,n1582);
or (n1585,n1586,n1589);
and (n1586,n1587,n1588);
xor (n1587,n1511,n1512);
and (n1588,n1516,n1552);
and (n1589,n1590,n1591);
xor (n1590,n1587,n1588);
or (n1591,n1592,n1595);
and (n1592,n1593,n1594);
xor (n1593,n1518,n1519);
and (n1594,n1523,n1552);
and (n1595,n1596,n1597);
xor (n1596,n1593,n1594);
or (n1597,n1598,n1601);
and (n1598,n1599,n1600);
xor (n1599,n1525,n1526);
and (n1600,n1530,n1552);
and (n1601,n1602,n1603);
xor (n1602,n1599,n1600);
or (n1603,n1604,n1607);
and (n1604,n1605,n1606);
xor (n1605,n1532,n1533);
and (n1606,n1537,n1552);
and (n1607,n1608,n1609);
xor (n1608,n1605,n1606);
or (n1609,n1610,n1613);
and (n1610,n1611,n1612);
xor (n1611,n1539,n1540);
and (n1612,n1544,n1552);
and (n1613,n1614,n1615);
xor (n1614,n1611,n1612);
and (n1615,n1616,n1617);
xor (n1616,n1546,n1547);
and (n1617,n1550,n1552);
and (n1618,n1474,n1619);
wire s0n1619,s1n1619,notn1619;
or (n1619,s0n1619,s1n1619);
not(notn1619,n1451);
and (s0n1619,notn1619,n168);
and (s1n1619,n1451,n893);
and (n1620,n1621,n1622);
xor (n1621,n1470,n1618);
or (n1622,n1623,n1626);
and (n1623,n1624,n1625);
xor (n1624,n1554,n1555);
and (n1625,n1481,n1619);
and (n1626,n1627,n1628);
xor (n1627,n1624,n1625);
or (n1628,n1629,n1632);
and (n1629,n1630,n1631);
xor (n1630,n1560,n1561);
and (n1631,n1488,n1619);
and (n1632,n1633,n1634);
xor (n1633,n1630,n1631);
or (n1634,n1635,n1638);
and (n1635,n1636,n1637);
xor (n1636,n1566,n1567);
and (n1637,n1495,n1619);
and (n1638,n1639,n1640);
xor (n1639,n1636,n1637);
or (n1640,n1641,n1644);
and (n1641,n1642,n1643);
xor (n1642,n1572,n1573);
and (n1643,n1502,n1619);
and (n1644,n1645,n1646);
xor (n1645,n1642,n1643);
or (n1646,n1647,n1650);
and (n1647,n1648,n1649);
xor (n1648,n1578,n1579);
and (n1649,n1509,n1619);
and (n1650,n1651,n1652);
xor (n1651,n1648,n1649);
or (n1652,n1653,n1656);
and (n1653,n1654,n1655);
xor (n1654,n1584,n1585);
and (n1655,n1516,n1619);
and (n1656,n1657,n1658);
xor (n1657,n1654,n1655);
or (n1658,n1659,n1662);
and (n1659,n1660,n1661);
xor (n1660,n1590,n1591);
and (n1661,n1523,n1619);
and (n1662,n1663,n1664);
xor (n1663,n1660,n1661);
or (n1664,n1665,n1668);
and (n1665,n1666,n1667);
xor (n1666,n1596,n1597);
and (n1667,n1530,n1619);
and (n1668,n1669,n1670);
xor (n1669,n1666,n1667);
or (n1670,n1671,n1674);
and (n1671,n1672,n1673);
xor (n1672,n1602,n1603);
and (n1673,n1537,n1619);
and (n1674,n1675,n1676);
xor (n1675,n1672,n1673);
or (n1676,n1677,n1680);
and (n1677,n1678,n1679);
xor (n1678,n1608,n1609);
and (n1679,n1544,n1619);
and (n1680,n1681,n1682);
xor (n1681,n1678,n1679);
and (n1682,n1683,n1684);
xor (n1683,n1614,n1615);
and (n1684,n1550,n1619);
and (n1685,n1474,n1686);
wire s0n1686,s1n1686,notn1686;
or (n1686,s0n1686,s1n1686);
not(notn1686,n1451);
and (s0n1686,notn1686,n235);
and (s1n1686,n1451,n960);
and (n1687,n1688,n1689);
xor (n1688,n1468,n1685);
or (n1689,n1690,n1693);
and (n1690,n1691,n1692);
xor (n1691,n1621,n1622);
and (n1692,n1481,n1686);
and (n1693,n1694,n1695);
xor (n1694,n1691,n1692);
or (n1695,n1696,n1699);
and (n1696,n1697,n1698);
xor (n1697,n1627,n1628);
and (n1698,n1488,n1686);
and (n1699,n1700,n1701);
xor (n1700,n1697,n1698);
or (n1701,n1702,n1705);
and (n1702,n1703,n1704);
xor (n1703,n1633,n1634);
and (n1704,n1495,n1686);
and (n1705,n1706,n1707);
xor (n1706,n1703,n1704);
or (n1707,n1708,n1711);
and (n1708,n1709,n1710);
xor (n1709,n1639,n1640);
and (n1710,n1502,n1686);
and (n1711,n1712,n1713);
xor (n1712,n1709,n1710);
or (n1713,n1714,n1717);
and (n1714,n1715,n1716);
xor (n1715,n1645,n1646);
and (n1716,n1509,n1686);
and (n1717,n1718,n1719);
xor (n1718,n1715,n1716);
or (n1719,n1720,n1723);
and (n1720,n1721,n1722);
xor (n1721,n1651,n1652);
and (n1722,n1516,n1686);
and (n1723,n1724,n1725);
xor (n1724,n1721,n1722);
or (n1725,n1726,n1729);
and (n1726,n1727,n1728);
xor (n1727,n1657,n1658);
and (n1728,n1523,n1686);
and (n1729,n1730,n1731);
xor (n1730,n1727,n1728);
or (n1731,n1732,n1735);
and (n1732,n1733,n1734);
xor (n1733,n1663,n1664);
and (n1734,n1530,n1686);
and (n1735,n1736,n1737);
xor (n1736,n1733,n1734);
or (n1737,n1738,n1741);
and (n1738,n1739,n1740);
xor (n1739,n1669,n1670);
and (n1740,n1537,n1686);
and (n1741,n1742,n1743);
xor (n1742,n1739,n1740);
or (n1743,n1744,n1747);
and (n1744,n1745,n1746);
xor (n1745,n1675,n1676);
and (n1746,n1544,n1686);
and (n1747,n1748,n1749);
xor (n1748,n1745,n1746);
and (n1749,n1750,n1751);
xor (n1750,n1681,n1682);
and (n1751,n1550,n1686);
and (n1752,n1474,n1753);
wire s0n1753,s1n1753,notn1753;
or (n1753,s0n1753,s1n1753);
not(notn1753,n1451);
and (s0n1753,notn1753,n302);
and (s1n1753,n1451,n1027);
and (n1754,n1755,n1756);
xor (n1755,n1466,n1752);
or (n1756,n1757,n1760);
and (n1757,n1758,n1759);
xor (n1758,n1688,n1689);
and (n1759,n1481,n1753);
and (n1760,n1761,n1762);
xor (n1761,n1758,n1759);
or (n1762,n1763,n1766);
and (n1763,n1764,n1765);
xor (n1764,n1694,n1695);
and (n1765,n1488,n1753);
and (n1766,n1767,n1768);
xor (n1767,n1764,n1765);
or (n1768,n1769,n1772);
and (n1769,n1770,n1771);
xor (n1770,n1700,n1701);
and (n1771,n1495,n1753);
and (n1772,n1773,n1774);
xor (n1773,n1770,n1771);
or (n1774,n1775,n1778);
and (n1775,n1776,n1777);
xor (n1776,n1706,n1707);
and (n1777,n1502,n1753);
and (n1778,n1779,n1780);
xor (n1779,n1776,n1777);
or (n1780,n1781,n1784);
and (n1781,n1782,n1783);
xor (n1782,n1712,n1713);
and (n1783,n1509,n1753);
and (n1784,n1785,n1786);
xor (n1785,n1782,n1783);
or (n1786,n1787,n1790);
and (n1787,n1788,n1789);
xor (n1788,n1718,n1719);
and (n1789,n1516,n1753);
and (n1790,n1791,n1792);
xor (n1791,n1788,n1789);
or (n1792,n1793,n1796);
and (n1793,n1794,n1795);
xor (n1794,n1724,n1725);
and (n1795,n1523,n1753);
and (n1796,n1797,n1798);
xor (n1797,n1794,n1795);
or (n1798,n1799,n1802);
and (n1799,n1800,n1801);
xor (n1800,n1730,n1731);
and (n1801,n1530,n1753);
and (n1802,n1803,n1804);
xor (n1803,n1800,n1801);
or (n1804,n1805,n1808);
and (n1805,n1806,n1807);
xor (n1806,n1736,n1737);
and (n1807,n1537,n1753);
and (n1808,n1809,n1810);
xor (n1809,n1806,n1807);
or (n1810,n1811,n1814);
and (n1811,n1812,n1813);
xor (n1812,n1742,n1743);
and (n1813,n1544,n1753);
and (n1814,n1815,n1816);
xor (n1815,n1812,n1813);
and (n1816,n1817,n1818);
xor (n1817,n1748,n1749);
and (n1818,n1550,n1753);
and (n1819,n1474,n1820);
wire s0n1820,s1n1820,notn1820;
or (n1820,s0n1820,s1n1820);
not(notn1820,n1451);
and (s0n1820,notn1820,n369);
and (s1n1820,n1451,n1094);
and (n1821,n1822,n1823);
xor (n1822,n1464,n1819);
or (n1823,n1824,n1827);
and (n1824,n1825,n1826);
xor (n1825,n1755,n1756);
and (n1826,n1481,n1820);
and (n1827,n1828,n1829);
xor (n1828,n1825,n1826);
or (n1829,n1830,n1833);
and (n1830,n1831,n1832);
xor (n1831,n1761,n1762);
and (n1832,n1488,n1820);
and (n1833,n1834,n1835);
xor (n1834,n1831,n1832);
or (n1835,n1836,n1839);
and (n1836,n1837,n1838);
xor (n1837,n1767,n1768);
and (n1838,n1495,n1820);
and (n1839,n1840,n1841);
xor (n1840,n1837,n1838);
or (n1841,n1842,n1845);
and (n1842,n1843,n1844);
xor (n1843,n1773,n1774);
and (n1844,n1502,n1820);
and (n1845,n1846,n1847);
xor (n1846,n1843,n1844);
or (n1847,n1848,n1851);
and (n1848,n1849,n1850);
xor (n1849,n1779,n1780);
and (n1850,n1509,n1820);
and (n1851,n1852,n1853);
xor (n1852,n1849,n1850);
or (n1853,n1854,n1857);
and (n1854,n1855,n1856);
xor (n1855,n1785,n1786);
and (n1856,n1516,n1820);
and (n1857,n1858,n1859);
xor (n1858,n1855,n1856);
or (n1859,n1860,n1863);
and (n1860,n1861,n1862);
xor (n1861,n1791,n1792);
and (n1862,n1523,n1820);
and (n1863,n1864,n1865);
xor (n1864,n1861,n1862);
or (n1865,n1866,n1869);
and (n1866,n1867,n1868);
xor (n1867,n1797,n1798);
and (n1868,n1530,n1820);
and (n1869,n1870,n1871);
xor (n1870,n1867,n1868);
or (n1871,n1872,n1875);
and (n1872,n1873,n1874);
xor (n1873,n1803,n1804);
and (n1874,n1537,n1820);
and (n1875,n1876,n1877);
xor (n1876,n1873,n1874);
or (n1877,n1878,n1881);
and (n1878,n1879,n1880);
xor (n1879,n1809,n1810);
and (n1880,n1544,n1820);
and (n1881,n1882,n1883);
xor (n1882,n1879,n1880);
and (n1883,n1884,n1885);
xor (n1884,n1815,n1816);
and (n1885,n1550,n1820);
and (n1886,n1474,n1887);
wire s0n1887,s1n1887,notn1887;
or (n1887,s0n1887,s1n1887);
not(notn1887,n1451);
and (s0n1887,notn1887,n436);
and (s1n1887,n1451,n1161);
and (n1888,n1889,n1890);
xor (n1889,n1462,n1886);
or (n1890,n1891,n1894);
and (n1891,n1892,n1893);
xor (n1892,n1822,n1823);
and (n1893,n1481,n1887);
and (n1894,n1895,n1896);
xor (n1895,n1892,n1893);
or (n1896,n1897,n1900);
and (n1897,n1898,n1899);
xor (n1898,n1828,n1829);
and (n1899,n1488,n1887);
and (n1900,n1901,n1902);
xor (n1901,n1898,n1899);
or (n1902,n1903,n1906);
and (n1903,n1904,n1905);
xor (n1904,n1834,n1835);
and (n1905,n1495,n1887);
and (n1906,n1907,n1908);
xor (n1907,n1904,n1905);
or (n1908,n1909,n1912);
and (n1909,n1910,n1911);
xor (n1910,n1840,n1841);
and (n1911,n1502,n1887);
and (n1912,n1913,n1914);
xor (n1913,n1910,n1911);
or (n1914,n1915,n1918);
and (n1915,n1916,n1917);
xor (n1916,n1846,n1847);
and (n1917,n1509,n1887);
and (n1918,n1919,n1920);
xor (n1919,n1916,n1917);
or (n1920,n1921,n1924);
and (n1921,n1922,n1923);
xor (n1922,n1852,n1853);
and (n1923,n1516,n1887);
and (n1924,n1925,n1926);
xor (n1925,n1922,n1923);
or (n1926,n1927,n1930);
and (n1927,n1928,n1929);
xor (n1928,n1858,n1859);
and (n1929,n1523,n1887);
and (n1930,n1931,n1932);
xor (n1931,n1928,n1929);
or (n1932,n1933,n1936);
and (n1933,n1934,n1935);
xor (n1934,n1864,n1865);
and (n1935,n1530,n1887);
and (n1936,n1937,n1938);
xor (n1937,n1934,n1935);
or (n1938,n1939,n1942);
and (n1939,n1940,n1941);
xor (n1940,n1870,n1871);
and (n1941,n1537,n1887);
and (n1942,n1943,n1944);
xor (n1943,n1940,n1941);
or (n1944,n1945,n1948);
and (n1945,n1946,n1947);
xor (n1946,n1876,n1877);
and (n1947,n1544,n1887);
and (n1948,n1949,n1950);
xor (n1949,n1946,n1947);
and (n1950,n1951,n1952);
xor (n1951,n1882,n1883);
and (n1952,n1550,n1887);
and (n1953,n1474,n1954);
wire s0n1954,s1n1954,notn1954;
or (n1954,s0n1954,s1n1954);
not(notn1954,n1451);
and (s0n1954,notn1954,n503);
and (s1n1954,n1451,n1228);
or (n1955,n1956,n1959);
and (n1956,n1957,n1958);
xor (n1957,n1889,n1890);
and (n1958,n1481,n1954);
and (n1959,n1960,n1961);
xor (n1960,n1957,n1958);
or (n1961,n1962,n1965);
and (n1962,n1963,n1964);
xor (n1963,n1895,n1896);
and (n1964,n1488,n1954);
and (n1965,n1966,n1967);
xor (n1966,n1963,n1964);
or (n1967,n1968,n1971);
and (n1968,n1969,n1970);
xor (n1969,n1901,n1902);
and (n1970,n1495,n1954);
and (n1971,n1972,n1973);
xor (n1972,n1969,n1970);
or (n1973,n1974,n1977);
and (n1974,n1975,n1976);
xor (n1975,n1907,n1908);
and (n1976,n1502,n1954);
and (n1977,n1978,n1979);
xor (n1978,n1975,n1976);
or (n1979,n1980,n1983);
and (n1980,n1981,n1982);
xor (n1981,n1913,n1914);
and (n1982,n1509,n1954);
and (n1983,n1984,n1985);
xor (n1984,n1981,n1982);
or (n1985,n1986,n1989);
and (n1986,n1987,n1988);
xor (n1987,n1919,n1920);
and (n1988,n1516,n1954);
and (n1989,n1990,n1991);
xor (n1990,n1987,n1988);
or (n1991,n1992,n1995);
and (n1992,n1993,n1994);
xor (n1993,n1925,n1926);
and (n1994,n1523,n1954);
and (n1995,n1996,n1997);
xor (n1996,n1993,n1994);
or (n1997,n1998,n2001);
and (n1998,n1999,n2000);
xor (n1999,n1931,n1932);
and (n2000,n1530,n1954);
and (n2001,n2002,n2003);
xor (n2002,n1999,n2000);
or (n2003,n2004,n2007);
and (n2004,n2005,n2006);
xor (n2005,n1937,n1938);
and (n2006,n1537,n1954);
and (n2007,n2008,n2009);
xor (n2008,n2005,n2006);
or (n2009,n2010,n2013);
and (n2010,n2011,n2012);
xor (n2011,n1943,n1944);
and (n2012,n1544,n1954);
and (n2013,n2014,n2015);
xor (n2014,n2011,n2012);
and (n2015,n2016,n2017);
xor (n2016,n1949,n1950);
and (n2017,n1550,n1954);
and (n2018,n1481,n2019);
wire s0n2019,s1n2019,notn2019;
or (n2019,s0n2019,s1n2019);
not(notn2019,n1451);
and (s0n2019,notn2019,n568);
and (s1n2019,n1451,n1293);
or (n2020,n2021,n2024);
and (n2021,n2022,n2023);
xor (n2022,n1960,n1961);
and (n2023,n1488,n2019);
and (n2024,n2025,n2026);
xor (n2025,n2022,n2023);
or (n2026,n2027,n2030);
and (n2027,n2028,n2029);
xor (n2028,n1966,n1967);
and (n2029,n1495,n2019);
and (n2030,n2031,n2032);
xor (n2031,n2028,n2029);
or (n2032,n2033,n2036);
and (n2033,n2034,n2035);
xor (n2034,n1972,n1973);
and (n2035,n1502,n2019);
and (n2036,n2037,n2038);
xor (n2037,n2034,n2035);
or (n2038,n2039,n2042);
and (n2039,n2040,n2041);
xor (n2040,n1978,n1979);
and (n2041,n1509,n2019);
and (n2042,n2043,n2044);
xor (n2043,n2040,n2041);
or (n2044,n2045,n2048);
and (n2045,n2046,n2047);
xor (n2046,n1984,n1985);
and (n2047,n1516,n2019);
and (n2048,n2049,n2050);
xor (n2049,n2046,n2047);
or (n2050,n2051,n2054);
and (n2051,n2052,n2053);
xor (n2052,n1990,n1991);
and (n2053,n1523,n2019);
and (n2054,n2055,n2056);
xor (n2055,n2052,n2053);
or (n2056,n2057,n2060);
and (n2057,n2058,n2059);
xor (n2058,n1996,n1997);
and (n2059,n1530,n2019);
and (n2060,n2061,n2062);
xor (n2061,n2058,n2059);
or (n2062,n2063,n2066);
and (n2063,n2064,n2065);
xor (n2064,n2002,n2003);
and (n2065,n1537,n2019);
and (n2066,n2067,n2068);
xor (n2067,n2064,n2065);
or (n2068,n2069,n2072);
and (n2069,n2070,n2071);
xor (n2070,n2008,n2009);
and (n2071,n1544,n2019);
and (n2072,n2073,n2074);
xor (n2073,n2070,n2071);
and (n2074,n2075,n2076);
xor (n2075,n2014,n2015);
and (n2076,n1550,n2019);
and (n2077,n1488,n2078);
wire s0n2078,s1n2078,notn2078;
or (n2078,s0n2078,s1n2078);
not(notn2078,n1451);
and (s0n2078,notn2078,n627);
and (s1n2078,n1451,n1352);
or (n2079,n2080,n2083);
and (n2080,n2081,n2082);
xor (n2081,n2025,n2026);
and (n2082,n1495,n2078);
and (n2083,n2084,n2085);
xor (n2084,n2081,n2082);
or (n2085,n2086,n2089);
and (n2086,n2087,n2088);
xor (n2087,n2031,n2032);
and (n2088,n1502,n2078);
and (n2089,n2090,n2091);
xor (n2090,n2087,n2088);
or (n2091,n2092,n2095);
and (n2092,n2093,n2094);
xor (n2093,n2037,n2038);
and (n2094,n1509,n2078);
and (n2095,n2096,n2097);
xor (n2096,n2093,n2094);
or (n2097,n2098,n2101);
and (n2098,n2099,n2100);
xor (n2099,n2043,n2044);
and (n2100,n1516,n2078);
and (n2101,n2102,n2103);
xor (n2102,n2099,n2100);
or (n2103,n2104,n2107);
and (n2104,n2105,n2106);
xor (n2105,n2049,n2050);
and (n2106,n1523,n2078);
and (n2107,n2108,n2109);
xor (n2108,n2105,n2106);
or (n2109,n2110,n2113);
and (n2110,n2111,n2112);
xor (n2111,n2055,n2056);
and (n2112,n1530,n2078);
and (n2113,n2114,n2115);
xor (n2114,n2111,n2112);
or (n2115,n2116,n2119);
and (n2116,n2117,n2118);
xor (n2117,n2061,n2062);
and (n2118,n1537,n2078);
and (n2119,n2120,n2121);
xor (n2120,n2117,n2118);
or (n2121,n2122,n2125);
and (n2122,n2123,n2124);
xor (n2123,n2067,n2068);
and (n2124,n1544,n2078);
and (n2125,n2126,n2127);
xor (n2126,n2123,n2124);
and (n2127,n2128,n2129);
xor (n2128,n2073,n2074);
and (n2129,n1550,n2078);
and (n2130,n1495,n2131);
wire s0n2131,s1n2131,notn2131;
or (n2131,s0n2131,s1n2131);
not(notn2131,n1451);
and (s0n2131,notn2131,n680);
and (s1n2131,n1451,n1405);
or (n2132,n2133,n2136);
and (n2133,n2134,n2135);
xor (n2134,n2084,n2085);
and (n2135,n1502,n2131);
and (n2136,n2137,n2138);
xor (n2137,n2134,n2135);
or (n2138,n2139,n2142);
and (n2139,n2140,n2141);
xor (n2140,n2090,n2091);
and (n2141,n1509,n2131);
and (n2142,n2143,n2144);
xor (n2143,n2140,n2141);
or (n2144,n2145,n2148);
and (n2145,n2146,n2147);
xor (n2146,n2096,n2097);
and (n2147,n1516,n2131);
and (n2148,n2149,n2150);
xor (n2149,n2146,n2147);
or (n2150,n2151,n2154);
and (n2151,n2152,n2153);
xor (n2152,n2102,n2103);
and (n2153,n1523,n2131);
and (n2154,n2155,n2156);
xor (n2155,n2152,n2153);
or (n2156,n2157,n2160);
and (n2157,n2158,n2159);
xor (n2158,n2108,n2109);
and (n2159,n1530,n2131);
and (n2160,n2161,n2162);
xor (n2161,n2158,n2159);
or (n2162,n2163,n2166);
and (n2163,n2164,n2165);
xor (n2164,n2114,n2115);
and (n2165,n1537,n2131);
and (n2166,n2167,n2168);
xor (n2167,n2164,n2165);
or (n2168,n2169,n2172);
and (n2169,n2170,n2171);
xor (n2170,n2120,n2121);
and (n2171,n1544,n2131);
and (n2172,n2173,n2174);
xor (n2173,n2170,n2171);
and (n2174,n2175,n2176);
xor (n2175,n2126,n2127);
and (n2176,n1550,n2131);
endmodule
