module top (out,n23,n24,n28,n30,n37,n44,n51,n58,n65
        ,n72,n79,n86,n93,n99,n101,n168,n233,n292,n345
        ,n392,n433,n468,n497,n520,n558,n559,n563,n565,n572
        ,n579,n586,n593,n600,n607,n614,n621,n628,n634,n636
        ,n703,n768,n827,n880,n927,n968,n1003,n1032,n1055,n1071);
output out;
input n23;
input n24;
input n28;
input n30;
input n37;
input n44;
input n51;
input n58;
input n65;
input n72;
input n79;
input n86;
input n93;
input n99;
input n101;
input n168;
input n233;
input n292;
input n345;
input n392;
input n433;
input n468;
input n497;
input n520;
input n558;
input n559;
input n563;
input n565;
input n572;
input n579;
input n586;
input n593;
input n600;
input n607;
input n614;
input n621;
input n628;
input n634;
input n636;
input n703;
input n768;
input n827;
input n880;
input n927;
input n968;
input n1003;
input n1032;
input n1055;
input n1071;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n25;
wire n26;
wire n27;
wire n29;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n100;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n560;
wire n561;
wire n562;
wire n564;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n635;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
xor (out,n0,n1072);
wire s0n0,s1n0,notn0;
or (n0,s0n0,s1n0);
not(notn0,n1071);
and (s0n0,notn0,n1);
and (s1n0,n1071,n536);
xor (n1,n2,n521);
xor (n2,n3,n519);
xor (n3,n4,n498);
xor (n4,n5,n496);
xor (n5,n6,n469);
xor (n6,n7,n467);
xor (n7,n8,n434);
xor (n8,n9,n432);
xor (n9,n10,n393);
xor (n10,n11,n391);
xor (n11,n12,n346);
xor (n12,n13,n344);
xor (n13,n14,n293);
xor (n14,n15,n291);
xor (n15,n16,n234);
xor (n16,n17,n232);
xor (n17,n18,n169);
xor (n18,n19,n167);
or (n19,n20,n102);
and (n20,n21,n100);
and (n21,n22,n25);
and (n22,n23,n24);
or (n25,n26,n31);
and (n26,n27,n29);
and (n27,n23,n28);
and (n29,n30,n24);
and (n31,n32,n33);
xor (n32,n27,n29);
or (n33,n34,n38);
and (n34,n35,n36);
and (n35,n30,n28);
and (n36,n37,n24);
and (n38,n39,n40);
xor (n39,n35,n36);
or (n40,n41,n45);
and (n41,n42,n43);
and (n42,n37,n28);
and (n43,n44,n24);
and (n45,n46,n47);
xor (n46,n42,n43);
or (n47,n48,n52);
and (n48,n49,n50);
and (n49,n44,n28);
and (n50,n51,n24);
and (n52,n53,n54);
xor (n53,n49,n50);
or (n54,n55,n59);
and (n55,n56,n57);
and (n56,n51,n28);
and (n57,n58,n24);
and (n59,n60,n61);
xor (n60,n56,n57);
or (n61,n62,n66);
and (n62,n63,n64);
and (n63,n58,n28);
and (n64,n65,n24);
and (n66,n67,n68);
xor (n67,n63,n64);
or (n68,n69,n73);
and (n69,n70,n71);
and (n70,n65,n28);
and (n71,n72,n24);
and (n73,n74,n75);
xor (n74,n70,n71);
or (n75,n76,n80);
and (n76,n77,n78);
and (n77,n72,n28);
and (n78,n79,n24);
and (n80,n81,n82);
xor (n81,n77,n78);
or (n82,n83,n87);
and (n83,n84,n85);
and (n84,n79,n28);
and (n85,n86,n24);
and (n87,n88,n89);
xor (n88,n84,n85);
or (n89,n90,n94);
and (n90,n91,n92);
and (n91,n86,n28);
and (n92,n93,n24);
and (n94,n95,n96);
xor (n95,n91,n92);
and (n96,n97,n98);
and (n97,n93,n28);
and (n98,n99,n24);
and (n100,n23,n101);
and (n102,n103,n104);
xor (n103,n21,n100);
or (n104,n105,n108);
and (n105,n106,n107);
xor (n106,n22,n25);
and (n107,n30,n101);
and (n108,n109,n110);
xor (n109,n106,n107);
or (n110,n111,n114);
and (n111,n112,n113);
xor (n112,n32,n33);
and (n113,n37,n101);
and (n114,n115,n116);
xor (n115,n112,n113);
or (n116,n117,n120);
and (n117,n118,n119);
xor (n118,n39,n40);
and (n119,n44,n101);
and (n120,n121,n122);
xor (n121,n118,n119);
or (n122,n123,n126);
and (n123,n124,n125);
xor (n124,n46,n47);
and (n125,n51,n101);
and (n126,n127,n128);
xor (n127,n124,n125);
or (n128,n129,n132);
and (n129,n130,n131);
xor (n130,n53,n54);
and (n131,n58,n101);
and (n132,n133,n134);
xor (n133,n130,n131);
or (n134,n135,n138);
and (n135,n136,n137);
xor (n136,n60,n61);
and (n137,n65,n101);
and (n138,n139,n140);
xor (n139,n136,n137);
or (n140,n141,n144);
and (n141,n142,n143);
xor (n142,n67,n68);
and (n143,n72,n101);
and (n144,n145,n146);
xor (n145,n142,n143);
or (n146,n147,n150);
and (n147,n148,n149);
xor (n148,n74,n75);
and (n149,n79,n101);
and (n150,n151,n152);
xor (n151,n148,n149);
or (n152,n153,n156);
and (n153,n154,n155);
xor (n154,n81,n82);
and (n155,n86,n101);
and (n156,n157,n158);
xor (n157,n154,n155);
or (n158,n159,n162);
and (n159,n160,n161);
xor (n160,n88,n89);
and (n161,n93,n101);
and (n162,n163,n164);
xor (n163,n160,n161);
and (n164,n165,n166);
xor (n165,n95,n96);
and (n166,n99,n101);
and (n167,n23,n168);
or (n169,n170,n173);
and (n170,n171,n172);
xor (n171,n103,n104);
and (n172,n30,n168);
and (n173,n174,n175);
xor (n174,n171,n172);
or (n175,n176,n179);
and (n176,n177,n178);
xor (n177,n109,n110);
and (n178,n37,n168);
and (n179,n180,n181);
xor (n180,n177,n178);
or (n181,n182,n185);
and (n182,n183,n184);
xor (n183,n115,n116);
and (n184,n44,n168);
and (n185,n186,n187);
xor (n186,n183,n184);
or (n187,n188,n191);
and (n188,n189,n190);
xor (n189,n121,n122);
and (n190,n51,n168);
and (n191,n192,n193);
xor (n192,n189,n190);
or (n193,n194,n197);
and (n194,n195,n196);
xor (n195,n127,n128);
and (n196,n58,n168);
and (n197,n198,n199);
xor (n198,n195,n196);
or (n199,n200,n203);
and (n200,n201,n202);
xor (n201,n133,n134);
and (n202,n65,n168);
and (n203,n204,n205);
xor (n204,n201,n202);
or (n205,n206,n209);
and (n206,n207,n208);
xor (n207,n139,n140);
and (n208,n72,n168);
and (n209,n210,n211);
xor (n210,n207,n208);
or (n211,n212,n215);
and (n212,n213,n214);
xor (n213,n145,n146);
and (n214,n79,n168);
and (n215,n216,n217);
xor (n216,n213,n214);
or (n217,n218,n221);
and (n218,n219,n220);
xor (n219,n151,n152);
and (n220,n86,n168);
and (n221,n222,n223);
xor (n222,n219,n220);
or (n223,n224,n227);
and (n224,n225,n226);
xor (n225,n157,n158);
and (n226,n93,n168);
and (n227,n228,n229);
xor (n228,n225,n226);
and (n229,n230,n231);
xor (n230,n163,n164);
and (n231,n99,n168);
and (n232,n30,n233);
or (n234,n235,n238);
and (n235,n236,n237);
xor (n236,n174,n175);
and (n237,n37,n233);
and (n238,n239,n240);
xor (n239,n236,n237);
or (n240,n241,n244);
and (n241,n242,n243);
xor (n242,n180,n181);
and (n243,n44,n233);
and (n244,n245,n246);
xor (n245,n242,n243);
or (n246,n247,n250);
and (n247,n248,n249);
xor (n248,n186,n187);
and (n249,n51,n233);
and (n250,n251,n252);
xor (n251,n248,n249);
or (n252,n253,n256);
and (n253,n254,n255);
xor (n254,n192,n193);
and (n255,n58,n233);
and (n256,n257,n258);
xor (n257,n254,n255);
or (n258,n259,n262);
and (n259,n260,n261);
xor (n260,n198,n199);
and (n261,n65,n233);
and (n262,n263,n264);
xor (n263,n260,n261);
or (n264,n265,n268);
and (n265,n266,n267);
xor (n266,n204,n205);
and (n267,n72,n233);
and (n268,n269,n270);
xor (n269,n266,n267);
or (n270,n271,n274);
and (n271,n272,n273);
xor (n272,n210,n211);
and (n273,n79,n233);
and (n274,n275,n276);
xor (n275,n272,n273);
or (n276,n277,n280);
and (n277,n278,n279);
xor (n278,n216,n217);
and (n279,n86,n233);
and (n280,n281,n282);
xor (n281,n278,n279);
or (n282,n283,n286);
and (n283,n284,n285);
xor (n284,n222,n223);
and (n285,n93,n233);
and (n286,n287,n288);
xor (n287,n284,n285);
and (n288,n289,n290);
xor (n289,n228,n229);
and (n290,n99,n233);
and (n291,n37,n292);
or (n293,n294,n297);
and (n294,n295,n296);
xor (n295,n239,n240);
and (n296,n44,n292);
and (n297,n298,n299);
xor (n298,n295,n296);
or (n299,n300,n303);
and (n300,n301,n302);
xor (n301,n245,n246);
and (n302,n51,n292);
and (n303,n304,n305);
xor (n304,n301,n302);
or (n305,n306,n309);
and (n306,n307,n308);
xor (n307,n251,n252);
and (n308,n58,n292);
and (n309,n310,n311);
xor (n310,n307,n308);
or (n311,n312,n315);
and (n312,n313,n314);
xor (n313,n257,n258);
and (n314,n65,n292);
and (n315,n316,n317);
xor (n316,n313,n314);
or (n317,n318,n321);
and (n318,n319,n320);
xor (n319,n263,n264);
and (n320,n72,n292);
and (n321,n322,n323);
xor (n322,n319,n320);
or (n323,n324,n327);
and (n324,n325,n326);
xor (n325,n269,n270);
and (n326,n79,n292);
and (n327,n328,n329);
xor (n328,n325,n326);
or (n329,n330,n333);
and (n330,n331,n332);
xor (n331,n275,n276);
and (n332,n86,n292);
and (n333,n334,n335);
xor (n334,n331,n332);
or (n335,n336,n339);
and (n336,n337,n338);
xor (n337,n281,n282);
and (n338,n93,n292);
and (n339,n340,n341);
xor (n340,n337,n338);
and (n341,n342,n343);
xor (n342,n287,n288);
and (n343,n99,n292);
and (n344,n44,n345);
or (n346,n347,n350);
and (n347,n348,n349);
xor (n348,n298,n299);
and (n349,n51,n345);
and (n350,n351,n352);
xor (n351,n348,n349);
or (n352,n353,n356);
and (n353,n354,n355);
xor (n354,n304,n305);
and (n355,n58,n345);
and (n356,n357,n358);
xor (n357,n354,n355);
or (n358,n359,n362);
and (n359,n360,n361);
xor (n360,n310,n311);
and (n361,n65,n345);
and (n362,n363,n364);
xor (n363,n360,n361);
or (n364,n365,n368);
and (n365,n366,n367);
xor (n366,n316,n317);
and (n367,n72,n345);
and (n368,n369,n370);
xor (n369,n366,n367);
or (n370,n371,n374);
and (n371,n372,n373);
xor (n372,n322,n323);
and (n373,n79,n345);
and (n374,n375,n376);
xor (n375,n372,n373);
or (n376,n377,n380);
and (n377,n378,n379);
xor (n378,n328,n329);
and (n379,n86,n345);
and (n380,n381,n382);
xor (n381,n378,n379);
or (n382,n383,n386);
and (n383,n384,n385);
xor (n384,n334,n335);
and (n385,n93,n345);
and (n386,n387,n388);
xor (n387,n384,n385);
and (n388,n389,n390);
xor (n389,n340,n341);
and (n390,n99,n345);
and (n391,n51,n392);
or (n393,n394,n397);
and (n394,n395,n396);
xor (n395,n351,n352);
and (n396,n58,n392);
and (n397,n398,n399);
xor (n398,n395,n396);
or (n399,n400,n403);
and (n400,n401,n402);
xor (n401,n357,n358);
and (n402,n65,n392);
and (n403,n404,n405);
xor (n404,n401,n402);
or (n405,n406,n409);
and (n406,n407,n408);
xor (n407,n363,n364);
and (n408,n72,n392);
and (n409,n410,n411);
xor (n410,n407,n408);
or (n411,n412,n415);
and (n412,n413,n414);
xor (n413,n369,n370);
and (n414,n79,n392);
and (n415,n416,n417);
xor (n416,n413,n414);
or (n417,n418,n421);
and (n418,n419,n420);
xor (n419,n375,n376);
and (n420,n86,n392);
and (n421,n422,n423);
xor (n422,n419,n420);
or (n423,n424,n427);
and (n424,n425,n426);
xor (n425,n381,n382);
and (n426,n93,n392);
and (n427,n428,n429);
xor (n428,n425,n426);
and (n429,n430,n431);
xor (n430,n387,n388);
and (n431,n99,n392);
and (n432,n58,n433);
or (n434,n435,n438);
and (n435,n436,n437);
xor (n436,n398,n399);
and (n437,n65,n433);
and (n438,n439,n440);
xor (n439,n436,n437);
or (n440,n441,n444);
and (n441,n442,n443);
xor (n442,n404,n405);
and (n443,n72,n433);
and (n444,n445,n446);
xor (n445,n442,n443);
or (n446,n447,n450);
and (n447,n448,n449);
xor (n448,n410,n411);
and (n449,n79,n433);
and (n450,n451,n452);
xor (n451,n448,n449);
or (n452,n453,n456);
and (n453,n454,n455);
xor (n454,n416,n417);
and (n455,n86,n433);
and (n456,n457,n458);
xor (n457,n454,n455);
or (n458,n459,n462);
and (n459,n460,n461);
xor (n460,n422,n423);
and (n461,n93,n433);
and (n462,n463,n464);
xor (n463,n460,n461);
and (n464,n465,n466);
xor (n465,n428,n429);
and (n466,n99,n433);
and (n467,n65,n468);
or (n469,n470,n473);
and (n470,n471,n472);
xor (n471,n439,n440);
and (n472,n72,n468);
and (n473,n474,n475);
xor (n474,n471,n472);
or (n475,n476,n479);
and (n476,n477,n478);
xor (n477,n445,n446);
and (n478,n79,n468);
and (n479,n480,n481);
xor (n480,n477,n478);
or (n481,n482,n485);
and (n482,n483,n484);
xor (n483,n451,n452);
and (n484,n86,n468);
and (n485,n486,n487);
xor (n486,n483,n484);
or (n487,n488,n491);
and (n488,n489,n490);
xor (n489,n457,n458);
and (n490,n93,n468);
and (n491,n492,n493);
xor (n492,n489,n490);
and (n493,n494,n495);
xor (n494,n463,n464);
and (n495,n99,n468);
and (n496,n72,n497);
or (n498,n499,n502);
and (n499,n500,n501);
xor (n500,n474,n475);
and (n501,n79,n497);
and (n502,n503,n504);
xor (n503,n500,n501);
or (n504,n505,n508);
and (n505,n506,n507);
xor (n506,n480,n481);
and (n507,n86,n497);
and (n508,n509,n510);
xor (n509,n506,n507);
or (n510,n511,n514);
and (n511,n512,n513);
xor (n512,n486,n487);
and (n513,n93,n497);
and (n514,n515,n516);
xor (n515,n512,n513);
and (n516,n517,n518);
xor (n517,n492,n493);
and (n518,n99,n497);
and (n519,n79,n520);
or (n521,n522,n525);
and (n522,n523,n524);
xor (n523,n503,n504);
and (n524,n86,n520);
and (n525,n526,n527);
xor (n526,n523,n524);
or (n527,n528,n531);
and (n528,n529,n530);
xor (n529,n509,n510);
and (n530,n93,n520);
and (n531,n532,n533);
xor (n532,n529,n530);
and (n533,n534,n535);
xor (n534,n515,n516);
and (n535,n99,n520);
xor (n536,n537,n1056);
xor (n537,n538,n1054);
xor (n538,n539,n1033);
xor (n539,n540,n1031);
xor (n540,n541,n1004);
xor (n541,n542,n1002);
xor (n542,n543,n969);
xor (n543,n544,n967);
xor (n544,n545,n928);
xor (n545,n546,n926);
xor (n546,n547,n881);
xor (n547,n548,n879);
xor (n548,n549,n828);
xor (n549,n550,n826);
xor (n550,n551,n769);
xor (n551,n552,n767);
xor (n552,n553,n704);
xor (n553,n554,n702);
or (n554,n555,n637);
and (n555,n556,n635);
and (n556,n557,n560);
and (n557,n558,n559);
or (n560,n561,n566);
and (n561,n562,n564);
and (n562,n558,n563);
and (n564,n565,n559);
and (n566,n567,n568);
xor (n567,n562,n564);
or (n568,n569,n573);
and (n569,n570,n571);
and (n570,n565,n563);
and (n571,n572,n559);
and (n573,n574,n575);
xor (n574,n570,n571);
or (n575,n576,n580);
and (n576,n577,n578);
and (n577,n572,n563);
and (n578,n579,n559);
and (n580,n581,n582);
xor (n581,n577,n578);
or (n582,n583,n587);
and (n583,n584,n585);
and (n584,n579,n563);
and (n585,n586,n559);
and (n587,n588,n589);
xor (n588,n584,n585);
or (n589,n590,n594);
and (n590,n591,n592);
and (n591,n586,n563);
and (n592,n593,n559);
and (n594,n595,n596);
xor (n595,n591,n592);
or (n596,n597,n601);
and (n597,n598,n599);
and (n598,n593,n563);
and (n599,n600,n559);
and (n601,n602,n603);
xor (n602,n598,n599);
or (n603,n604,n608);
and (n604,n605,n606);
and (n605,n600,n563);
and (n606,n607,n559);
and (n608,n609,n610);
xor (n609,n605,n606);
or (n610,n611,n615);
and (n611,n612,n613);
and (n612,n607,n563);
and (n613,n614,n559);
and (n615,n616,n617);
xor (n616,n612,n613);
or (n617,n618,n622);
and (n618,n619,n620);
and (n619,n614,n563);
and (n620,n621,n559);
and (n622,n623,n624);
xor (n623,n619,n620);
or (n624,n625,n629);
and (n625,n626,n627);
and (n626,n621,n563);
and (n627,n628,n559);
and (n629,n630,n631);
xor (n630,n626,n627);
and (n631,n632,n633);
and (n632,n628,n563);
and (n633,n634,n559);
and (n635,n558,n636);
and (n637,n638,n639);
xor (n638,n556,n635);
or (n639,n640,n643);
and (n640,n641,n642);
xor (n641,n557,n560);
and (n642,n565,n636);
and (n643,n644,n645);
xor (n644,n641,n642);
or (n645,n646,n649);
and (n646,n647,n648);
xor (n647,n567,n568);
and (n648,n572,n636);
and (n649,n650,n651);
xor (n650,n647,n648);
or (n651,n652,n655);
and (n652,n653,n654);
xor (n653,n574,n575);
and (n654,n579,n636);
and (n655,n656,n657);
xor (n656,n653,n654);
or (n657,n658,n661);
and (n658,n659,n660);
xor (n659,n581,n582);
and (n660,n586,n636);
and (n661,n662,n663);
xor (n662,n659,n660);
or (n663,n664,n667);
and (n664,n665,n666);
xor (n665,n588,n589);
and (n666,n593,n636);
and (n667,n668,n669);
xor (n668,n665,n666);
or (n669,n670,n673);
and (n670,n671,n672);
xor (n671,n595,n596);
and (n672,n600,n636);
and (n673,n674,n675);
xor (n674,n671,n672);
or (n675,n676,n679);
and (n676,n677,n678);
xor (n677,n602,n603);
and (n678,n607,n636);
and (n679,n680,n681);
xor (n680,n677,n678);
or (n681,n682,n685);
and (n682,n683,n684);
xor (n683,n609,n610);
and (n684,n614,n636);
and (n685,n686,n687);
xor (n686,n683,n684);
or (n687,n688,n691);
and (n688,n689,n690);
xor (n689,n616,n617);
and (n690,n621,n636);
and (n691,n692,n693);
xor (n692,n689,n690);
or (n693,n694,n697);
and (n694,n695,n696);
xor (n695,n623,n624);
and (n696,n628,n636);
and (n697,n698,n699);
xor (n698,n695,n696);
and (n699,n700,n701);
xor (n700,n630,n631);
and (n701,n634,n636);
and (n702,n558,n703);
or (n704,n705,n708);
and (n705,n706,n707);
xor (n706,n638,n639);
and (n707,n565,n703);
and (n708,n709,n710);
xor (n709,n706,n707);
or (n710,n711,n714);
and (n711,n712,n713);
xor (n712,n644,n645);
and (n713,n572,n703);
and (n714,n715,n716);
xor (n715,n712,n713);
or (n716,n717,n720);
and (n717,n718,n719);
xor (n718,n650,n651);
and (n719,n579,n703);
and (n720,n721,n722);
xor (n721,n718,n719);
or (n722,n723,n726);
and (n723,n724,n725);
xor (n724,n656,n657);
and (n725,n586,n703);
and (n726,n727,n728);
xor (n727,n724,n725);
or (n728,n729,n732);
and (n729,n730,n731);
xor (n730,n662,n663);
and (n731,n593,n703);
and (n732,n733,n734);
xor (n733,n730,n731);
or (n734,n735,n738);
and (n735,n736,n737);
xor (n736,n668,n669);
and (n737,n600,n703);
and (n738,n739,n740);
xor (n739,n736,n737);
or (n740,n741,n744);
and (n741,n742,n743);
xor (n742,n674,n675);
and (n743,n607,n703);
and (n744,n745,n746);
xor (n745,n742,n743);
or (n746,n747,n750);
and (n747,n748,n749);
xor (n748,n680,n681);
and (n749,n614,n703);
and (n750,n751,n752);
xor (n751,n748,n749);
or (n752,n753,n756);
and (n753,n754,n755);
xor (n754,n686,n687);
and (n755,n621,n703);
and (n756,n757,n758);
xor (n757,n754,n755);
or (n758,n759,n762);
and (n759,n760,n761);
xor (n760,n692,n693);
and (n761,n628,n703);
and (n762,n763,n764);
xor (n763,n760,n761);
and (n764,n765,n766);
xor (n765,n698,n699);
and (n766,n634,n703);
and (n767,n565,n768);
or (n769,n770,n773);
and (n770,n771,n772);
xor (n771,n709,n710);
and (n772,n572,n768);
and (n773,n774,n775);
xor (n774,n771,n772);
or (n775,n776,n779);
and (n776,n777,n778);
xor (n777,n715,n716);
and (n778,n579,n768);
and (n779,n780,n781);
xor (n780,n777,n778);
or (n781,n782,n785);
and (n782,n783,n784);
xor (n783,n721,n722);
and (n784,n586,n768);
and (n785,n786,n787);
xor (n786,n783,n784);
or (n787,n788,n791);
and (n788,n789,n790);
xor (n789,n727,n728);
and (n790,n593,n768);
and (n791,n792,n793);
xor (n792,n789,n790);
or (n793,n794,n797);
and (n794,n795,n796);
xor (n795,n733,n734);
and (n796,n600,n768);
and (n797,n798,n799);
xor (n798,n795,n796);
or (n799,n800,n803);
and (n800,n801,n802);
xor (n801,n739,n740);
and (n802,n607,n768);
and (n803,n804,n805);
xor (n804,n801,n802);
or (n805,n806,n809);
and (n806,n807,n808);
xor (n807,n745,n746);
and (n808,n614,n768);
and (n809,n810,n811);
xor (n810,n807,n808);
or (n811,n812,n815);
and (n812,n813,n814);
xor (n813,n751,n752);
and (n814,n621,n768);
and (n815,n816,n817);
xor (n816,n813,n814);
or (n817,n818,n821);
and (n818,n819,n820);
xor (n819,n757,n758);
and (n820,n628,n768);
and (n821,n822,n823);
xor (n822,n819,n820);
and (n823,n824,n825);
xor (n824,n763,n764);
and (n825,n634,n768);
and (n826,n572,n827);
or (n828,n829,n832);
and (n829,n830,n831);
xor (n830,n774,n775);
and (n831,n579,n827);
and (n832,n833,n834);
xor (n833,n830,n831);
or (n834,n835,n838);
and (n835,n836,n837);
xor (n836,n780,n781);
and (n837,n586,n827);
and (n838,n839,n840);
xor (n839,n836,n837);
or (n840,n841,n844);
and (n841,n842,n843);
xor (n842,n786,n787);
and (n843,n593,n827);
and (n844,n845,n846);
xor (n845,n842,n843);
or (n846,n847,n850);
and (n847,n848,n849);
xor (n848,n792,n793);
and (n849,n600,n827);
and (n850,n851,n852);
xor (n851,n848,n849);
or (n852,n853,n856);
and (n853,n854,n855);
xor (n854,n798,n799);
and (n855,n607,n827);
and (n856,n857,n858);
xor (n857,n854,n855);
or (n858,n859,n862);
and (n859,n860,n861);
xor (n860,n804,n805);
and (n861,n614,n827);
and (n862,n863,n864);
xor (n863,n860,n861);
or (n864,n865,n868);
and (n865,n866,n867);
xor (n866,n810,n811);
and (n867,n621,n827);
and (n868,n869,n870);
xor (n869,n866,n867);
or (n870,n871,n874);
and (n871,n872,n873);
xor (n872,n816,n817);
and (n873,n628,n827);
and (n874,n875,n876);
xor (n875,n872,n873);
and (n876,n877,n878);
xor (n877,n822,n823);
and (n878,n634,n827);
and (n879,n579,n880);
or (n881,n882,n885);
and (n882,n883,n884);
xor (n883,n833,n834);
and (n884,n586,n880);
and (n885,n886,n887);
xor (n886,n883,n884);
or (n887,n888,n891);
and (n888,n889,n890);
xor (n889,n839,n840);
and (n890,n593,n880);
and (n891,n892,n893);
xor (n892,n889,n890);
or (n893,n894,n897);
and (n894,n895,n896);
xor (n895,n845,n846);
and (n896,n600,n880);
and (n897,n898,n899);
xor (n898,n895,n896);
or (n899,n900,n903);
and (n900,n901,n902);
xor (n901,n851,n852);
and (n902,n607,n880);
and (n903,n904,n905);
xor (n904,n901,n902);
or (n905,n906,n909);
and (n906,n907,n908);
xor (n907,n857,n858);
and (n908,n614,n880);
and (n909,n910,n911);
xor (n910,n907,n908);
or (n911,n912,n915);
and (n912,n913,n914);
xor (n913,n863,n864);
and (n914,n621,n880);
and (n915,n916,n917);
xor (n916,n913,n914);
or (n917,n918,n921);
and (n918,n919,n920);
xor (n919,n869,n870);
and (n920,n628,n880);
and (n921,n922,n923);
xor (n922,n919,n920);
and (n923,n924,n925);
xor (n924,n875,n876);
and (n925,n634,n880);
and (n926,n586,n927);
or (n928,n929,n932);
and (n929,n930,n931);
xor (n930,n886,n887);
and (n931,n593,n927);
and (n932,n933,n934);
xor (n933,n930,n931);
or (n934,n935,n938);
and (n935,n936,n937);
xor (n936,n892,n893);
and (n937,n600,n927);
and (n938,n939,n940);
xor (n939,n936,n937);
or (n940,n941,n944);
and (n941,n942,n943);
xor (n942,n898,n899);
and (n943,n607,n927);
and (n944,n945,n946);
xor (n945,n942,n943);
or (n946,n947,n950);
and (n947,n948,n949);
xor (n948,n904,n905);
and (n949,n614,n927);
and (n950,n951,n952);
xor (n951,n948,n949);
or (n952,n953,n956);
and (n953,n954,n955);
xor (n954,n910,n911);
and (n955,n621,n927);
and (n956,n957,n958);
xor (n957,n954,n955);
or (n958,n959,n962);
and (n959,n960,n961);
xor (n960,n916,n917);
and (n961,n628,n927);
and (n962,n963,n964);
xor (n963,n960,n961);
and (n964,n965,n966);
xor (n965,n922,n923);
and (n966,n634,n927);
and (n967,n593,n968);
or (n969,n970,n973);
and (n970,n971,n972);
xor (n971,n933,n934);
and (n972,n600,n968);
and (n973,n974,n975);
xor (n974,n971,n972);
or (n975,n976,n979);
and (n976,n977,n978);
xor (n977,n939,n940);
and (n978,n607,n968);
and (n979,n980,n981);
xor (n980,n977,n978);
or (n981,n982,n985);
and (n982,n983,n984);
xor (n983,n945,n946);
and (n984,n614,n968);
and (n985,n986,n987);
xor (n986,n983,n984);
or (n987,n988,n991);
and (n988,n989,n990);
xor (n989,n951,n952);
and (n990,n621,n968);
and (n991,n992,n993);
xor (n992,n989,n990);
or (n993,n994,n997);
and (n994,n995,n996);
xor (n995,n957,n958);
and (n996,n628,n968);
and (n997,n998,n999);
xor (n998,n995,n996);
and (n999,n1000,n1001);
xor (n1000,n963,n964);
and (n1001,n634,n968);
and (n1002,n600,n1003);
or (n1004,n1005,n1008);
and (n1005,n1006,n1007);
xor (n1006,n974,n975);
and (n1007,n607,n1003);
and (n1008,n1009,n1010);
xor (n1009,n1006,n1007);
or (n1010,n1011,n1014);
and (n1011,n1012,n1013);
xor (n1012,n980,n981);
and (n1013,n614,n1003);
and (n1014,n1015,n1016);
xor (n1015,n1012,n1013);
or (n1016,n1017,n1020);
and (n1017,n1018,n1019);
xor (n1018,n986,n987);
and (n1019,n621,n1003);
and (n1020,n1021,n1022);
xor (n1021,n1018,n1019);
or (n1022,n1023,n1026);
and (n1023,n1024,n1025);
xor (n1024,n992,n993);
and (n1025,n628,n1003);
and (n1026,n1027,n1028);
xor (n1027,n1024,n1025);
and (n1028,n1029,n1030);
xor (n1029,n998,n999);
and (n1030,n634,n1003);
and (n1031,n607,n1032);
or (n1033,n1034,n1037);
and (n1034,n1035,n1036);
xor (n1035,n1009,n1010);
and (n1036,n614,n1032);
and (n1037,n1038,n1039);
xor (n1038,n1035,n1036);
or (n1039,n1040,n1043);
and (n1040,n1041,n1042);
xor (n1041,n1015,n1016);
and (n1042,n621,n1032);
and (n1043,n1044,n1045);
xor (n1044,n1041,n1042);
or (n1045,n1046,n1049);
and (n1046,n1047,n1048);
xor (n1047,n1021,n1022);
and (n1048,n628,n1032);
and (n1049,n1050,n1051);
xor (n1050,n1047,n1048);
and (n1051,n1052,n1053);
xor (n1052,n1027,n1028);
and (n1053,n634,n1032);
and (n1054,n614,n1055);
or (n1056,n1057,n1060);
and (n1057,n1058,n1059);
xor (n1058,n1038,n1039);
and (n1059,n621,n1055);
and (n1060,n1061,n1062);
xor (n1061,n1058,n1059);
or (n1062,n1063,n1066);
and (n1063,n1064,n1065);
xor (n1064,n1044,n1045);
and (n1065,n628,n1055);
and (n1066,n1067,n1068);
xor (n1067,n1064,n1065);
and (n1068,n1069,n1070);
xor (n1069,n1050,n1051);
and (n1070,n634,n1055);
xor (n1072,n1073,n1592);
xor (n1073,n1074,n1590);
xor (n1074,n1075,n1569);
xor (n1075,n1076,n1567);
xor (n1076,n1077,n1540);
xor (n1077,n1078,n1538);
xor (n1078,n1079,n1505);
xor (n1079,n1080,n1503);
xor (n1080,n1081,n1464);
xor (n1081,n1082,n1462);
xor (n1082,n1083,n1417);
xor (n1083,n1084,n1415);
xor (n1084,n1085,n1364);
xor (n1085,n1086,n1362);
xor (n1086,n1087,n1305);
xor (n1087,n1088,n1303);
xor (n1088,n1089,n1240);
xor (n1089,n1090,n1238);
or (n1090,n1091,n1173);
and (n1091,n1092,n1171);
and (n1092,n1093,n1096);
and (n1093,n1094,n1095);
wire s0n1094,s1n1094,notn1094;
or (n1094,s0n1094,s1n1094);
not(notn1094,n1071);
and (s0n1094,notn1094,n23);
and (s1n1094,n1071,n558);
wire s0n1095,s1n1095,notn1095;
or (n1095,s0n1095,s1n1095);
not(notn1095,n1071);
and (s0n1095,notn1095,n24);
and (s1n1095,n1071,n559);
or (n1096,n1097,n1102);
and (n1097,n1098,n1100);
and (n1098,n1094,n1099);
wire s0n1099,s1n1099,notn1099;
or (n1099,s0n1099,s1n1099);
not(notn1099,n1071);
and (s0n1099,notn1099,n28);
and (s1n1099,n1071,n563);
and (n1100,n1101,n1095);
wire s0n1101,s1n1101,notn1101;
or (n1101,s0n1101,s1n1101);
not(notn1101,n1071);
and (s0n1101,notn1101,n30);
and (s1n1101,n1071,n565);
and (n1102,n1103,n1104);
xor (n1103,n1098,n1100);
or (n1104,n1105,n1109);
and (n1105,n1106,n1107);
and (n1106,n1101,n1099);
and (n1107,n1108,n1095);
wire s0n1108,s1n1108,notn1108;
or (n1108,s0n1108,s1n1108);
not(notn1108,n1071);
and (s0n1108,notn1108,n37);
and (s1n1108,n1071,n572);
and (n1109,n1110,n1111);
xor (n1110,n1106,n1107);
or (n1111,n1112,n1116);
and (n1112,n1113,n1114);
and (n1113,n1108,n1099);
and (n1114,n1115,n1095);
wire s0n1115,s1n1115,notn1115;
or (n1115,s0n1115,s1n1115);
not(notn1115,n1071);
and (s0n1115,notn1115,n44);
and (s1n1115,n1071,n579);
and (n1116,n1117,n1118);
xor (n1117,n1113,n1114);
or (n1118,n1119,n1123);
and (n1119,n1120,n1121);
and (n1120,n1115,n1099);
and (n1121,n1122,n1095);
wire s0n1122,s1n1122,notn1122;
or (n1122,s0n1122,s1n1122);
not(notn1122,n1071);
and (s0n1122,notn1122,n51);
and (s1n1122,n1071,n586);
and (n1123,n1124,n1125);
xor (n1124,n1120,n1121);
or (n1125,n1126,n1130);
and (n1126,n1127,n1128);
and (n1127,n1122,n1099);
and (n1128,n1129,n1095);
wire s0n1129,s1n1129,notn1129;
or (n1129,s0n1129,s1n1129);
not(notn1129,n1071);
and (s0n1129,notn1129,n58);
and (s1n1129,n1071,n593);
and (n1130,n1131,n1132);
xor (n1131,n1127,n1128);
or (n1132,n1133,n1137);
and (n1133,n1134,n1135);
and (n1134,n1129,n1099);
and (n1135,n1136,n1095);
wire s0n1136,s1n1136,notn1136;
or (n1136,s0n1136,s1n1136);
not(notn1136,n1071);
and (s0n1136,notn1136,n65);
and (s1n1136,n1071,n600);
and (n1137,n1138,n1139);
xor (n1138,n1134,n1135);
or (n1139,n1140,n1144);
and (n1140,n1141,n1142);
and (n1141,n1136,n1099);
and (n1142,n1143,n1095);
wire s0n1143,s1n1143,notn1143;
or (n1143,s0n1143,s1n1143);
not(notn1143,n1071);
and (s0n1143,notn1143,n72);
and (s1n1143,n1071,n607);
and (n1144,n1145,n1146);
xor (n1145,n1141,n1142);
or (n1146,n1147,n1151);
and (n1147,n1148,n1149);
and (n1148,n1143,n1099);
and (n1149,n1150,n1095);
wire s0n1150,s1n1150,notn1150;
or (n1150,s0n1150,s1n1150);
not(notn1150,n1071);
and (s0n1150,notn1150,n79);
and (s1n1150,n1071,n614);
and (n1151,n1152,n1153);
xor (n1152,n1148,n1149);
or (n1153,n1154,n1158);
and (n1154,n1155,n1156);
and (n1155,n1150,n1099);
and (n1156,n1157,n1095);
wire s0n1157,s1n1157,notn1157;
or (n1157,s0n1157,s1n1157);
not(notn1157,n1071);
and (s0n1157,notn1157,n86);
and (s1n1157,n1071,n621);
and (n1158,n1159,n1160);
xor (n1159,n1155,n1156);
or (n1160,n1161,n1165);
and (n1161,n1162,n1163);
and (n1162,n1157,n1099);
and (n1163,n1164,n1095);
wire s0n1164,s1n1164,notn1164;
or (n1164,s0n1164,s1n1164);
not(notn1164,n1071);
and (s0n1164,notn1164,n93);
and (s1n1164,n1071,n628);
and (n1165,n1166,n1167);
xor (n1166,n1162,n1163);
and (n1167,n1168,n1169);
and (n1168,n1164,n1099);
and (n1169,n1170,n1095);
wire s0n1170,s1n1170,notn1170;
or (n1170,s0n1170,s1n1170);
not(notn1170,n1071);
and (s0n1170,notn1170,n99);
and (s1n1170,n1071,n634);
and (n1171,n1094,n1172);
wire s0n1172,s1n1172,notn1172;
or (n1172,s0n1172,s1n1172);
not(notn1172,n1071);
and (s0n1172,notn1172,n101);
and (s1n1172,n1071,n636);
and (n1173,n1174,n1175);
xor (n1174,n1092,n1171);
or (n1175,n1176,n1179);
and (n1176,n1177,n1178);
xor (n1177,n1093,n1096);
and (n1178,n1101,n1172);
and (n1179,n1180,n1181);
xor (n1180,n1177,n1178);
or (n1181,n1182,n1185);
and (n1182,n1183,n1184);
xor (n1183,n1103,n1104);
and (n1184,n1108,n1172);
and (n1185,n1186,n1187);
xor (n1186,n1183,n1184);
or (n1187,n1188,n1191);
and (n1188,n1189,n1190);
xor (n1189,n1110,n1111);
and (n1190,n1115,n1172);
and (n1191,n1192,n1193);
xor (n1192,n1189,n1190);
or (n1193,n1194,n1197);
and (n1194,n1195,n1196);
xor (n1195,n1117,n1118);
and (n1196,n1122,n1172);
and (n1197,n1198,n1199);
xor (n1198,n1195,n1196);
or (n1199,n1200,n1203);
and (n1200,n1201,n1202);
xor (n1201,n1124,n1125);
and (n1202,n1129,n1172);
and (n1203,n1204,n1205);
xor (n1204,n1201,n1202);
or (n1205,n1206,n1209);
and (n1206,n1207,n1208);
xor (n1207,n1131,n1132);
and (n1208,n1136,n1172);
and (n1209,n1210,n1211);
xor (n1210,n1207,n1208);
or (n1211,n1212,n1215);
and (n1212,n1213,n1214);
xor (n1213,n1138,n1139);
and (n1214,n1143,n1172);
and (n1215,n1216,n1217);
xor (n1216,n1213,n1214);
or (n1217,n1218,n1221);
and (n1218,n1219,n1220);
xor (n1219,n1145,n1146);
and (n1220,n1150,n1172);
and (n1221,n1222,n1223);
xor (n1222,n1219,n1220);
or (n1223,n1224,n1227);
and (n1224,n1225,n1226);
xor (n1225,n1152,n1153);
and (n1226,n1157,n1172);
and (n1227,n1228,n1229);
xor (n1228,n1225,n1226);
or (n1229,n1230,n1233);
and (n1230,n1231,n1232);
xor (n1231,n1159,n1160);
and (n1232,n1164,n1172);
and (n1233,n1234,n1235);
xor (n1234,n1231,n1232);
and (n1235,n1236,n1237);
xor (n1236,n1166,n1167);
and (n1237,n1170,n1172);
and (n1238,n1094,n1239);
wire s0n1239,s1n1239,notn1239;
or (n1239,s0n1239,s1n1239);
not(notn1239,n1071);
and (s0n1239,notn1239,n168);
and (s1n1239,n1071,n703);
or (n1240,n1241,n1244);
and (n1241,n1242,n1243);
xor (n1242,n1174,n1175);
and (n1243,n1101,n1239);
and (n1244,n1245,n1246);
xor (n1245,n1242,n1243);
or (n1246,n1247,n1250);
and (n1247,n1248,n1249);
xor (n1248,n1180,n1181);
and (n1249,n1108,n1239);
and (n1250,n1251,n1252);
xor (n1251,n1248,n1249);
or (n1252,n1253,n1256);
and (n1253,n1254,n1255);
xor (n1254,n1186,n1187);
and (n1255,n1115,n1239);
and (n1256,n1257,n1258);
xor (n1257,n1254,n1255);
or (n1258,n1259,n1262);
and (n1259,n1260,n1261);
xor (n1260,n1192,n1193);
and (n1261,n1122,n1239);
and (n1262,n1263,n1264);
xor (n1263,n1260,n1261);
or (n1264,n1265,n1268);
and (n1265,n1266,n1267);
xor (n1266,n1198,n1199);
and (n1267,n1129,n1239);
and (n1268,n1269,n1270);
xor (n1269,n1266,n1267);
or (n1270,n1271,n1274);
and (n1271,n1272,n1273);
xor (n1272,n1204,n1205);
and (n1273,n1136,n1239);
and (n1274,n1275,n1276);
xor (n1275,n1272,n1273);
or (n1276,n1277,n1280);
and (n1277,n1278,n1279);
xor (n1278,n1210,n1211);
and (n1279,n1143,n1239);
and (n1280,n1281,n1282);
xor (n1281,n1278,n1279);
or (n1282,n1283,n1286);
and (n1283,n1284,n1285);
xor (n1284,n1216,n1217);
and (n1285,n1150,n1239);
and (n1286,n1287,n1288);
xor (n1287,n1284,n1285);
or (n1288,n1289,n1292);
and (n1289,n1290,n1291);
xor (n1290,n1222,n1223);
and (n1291,n1157,n1239);
and (n1292,n1293,n1294);
xor (n1293,n1290,n1291);
or (n1294,n1295,n1298);
and (n1295,n1296,n1297);
xor (n1296,n1228,n1229);
and (n1297,n1164,n1239);
and (n1298,n1299,n1300);
xor (n1299,n1296,n1297);
and (n1300,n1301,n1302);
xor (n1301,n1234,n1235);
and (n1302,n1170,n1239);
and (n1303,n1101,n1304);
wire s0n1304,s1n1304,notn1304;
or (n1304,s0n1304,s1n1304);
not(notn1304,n1071);
and (s0n1304,notn1304,n233);
and (s1n1304,n1071,n768);
or (n1305,n1306,n1309);
and (n1306,n1307,n1308);
xor (n1307,n1245,n1246);
and (n1308,n1108,n1304);
and (n1309,n1310,n1311);
xor (n1310,n1307,n1308);
or (n1311,n1312,n1315);
and (n1312,n1313,n1314);
xor (n1313,n1251,n1252);
and (n1314,n1115,n1304);
and (n1315,n1316,n1317);
xor (n1316,n1313,n1314);
or (n1317,n1318,n1321);
and (n1318,n1319,n1320);
xor (n1319,n1257,n1258);
and (n1320,n1122,n1304);
and (n1321,n1322,n1323);
xor (n1322,n1319,n1320);
or (n1323,n1324,n1327);
and (n1324,n1325,n1326);
xor (n1325,n1263,n1264);
and (n1326,n1129,n1304);
and (n1327,n1328,n1329);
xor (n1328,n1325,n1326);
or (n1329,n1330,n1333);
and (n1330,n1331,n1332);
xor (n1331,n1269,n1270);
and (n1332,n1136,n1304);
and (n1333,n1334,n1335);
xor (n1334,n1331,n1332);
or (n1335,n1336,n1339);
and (n1336,n1337,n1338);
xor (n1337,n1275,n1276);
and (n1338,n1143,n1304);
and (n1339,n1340,n1341);
xor (n1340,n1337,n1338);
or (n1341,n1342,n1345);
and (n1342,n1343,n1344);
xor (n1343,n1281,n1282);
and (n1344,n1150,n1304);
and (n1345,n1346,n1347);
xor (n1346,n1343,n1344);
or (n1347,n1348,n1351);
and (n1348,n1349,n1350);
xor (n1349,n1287,n1288);
and (n1350,n1157,n1304);
and (n1351,n1352,n1353);
xor (n1352,n1349,n1350);
or (n1353,n1354,n1357);
and (n1354,n1355,n1356);
xor (n1355,n1293,n1294);
and (n1356,n1164,n1304);
and (n1357,n1358,n1359);
xor (n1358,n1355,n1356);
and (n1359,n1360,n1361);
xor (n1360,n1299,n1300);
and (n1361,n1170,n1304);
and (n1362,n1108,n1363);
wire s0n1363,s1n1363,notn1363;
or (n1363,s0n1363,s1n1363);
not(notn1363,n1071);
and (s0n1363,notn1363,n292);
and (s1n1363,n1071,n827);
or (n1364,n1365,n1368);
and (n1365,n1366,n1367);
xor (n1366,n1310,n1311);
and (n1367,n1115,n1363);
and (n1368,n1369,n1370);
xor (n1369,n1366,n1367);
or (n1370,n1371,n1374);
and (n1371,n1372,n1373);
xor (n1372,n1316,n1317);
and (n1373,n1122,n1363);
and (n1374,n1375,n1376);
xor (n1375,n1372,n1373);
or (n1376,n1377,n1380);
and (n1377,n1378,n1379);
xor (n1378,n1322,n1323);
and (n1379,n1129,n1363);
and (n1380,n1381,n1382);
xor (n1381,n1378,n1379);
or (n1382,n1383,n1386);
and (n1383,n1384,n1385);
xor (n1384,n1328,n1329);
and (n1385,n1136,n1363);
and (n1386,n1387,n1388);
xor (n1387,n1384,n1385);
or (n1388,n1389,n1392);
and (n1389,n1390,n1391);
xor (n1390,n1334,n1335);
and (n1391,n1143,n1363);
and (n1392,n1393,n1394);
xor (n1393,n1390,n1391);
or (n1394,n1395,n1398);
and (n1395,n1396,n1397);
xor (n1396,n1340,n1341);
and (n1397,n1150,n1363);
and (n1398,n1399,n1400);
xor (n1399,n1396,n1397);
or (n1400,n1401,n1404);
and (n1401,n1402,n1403);
xor (n1402,n1346,n1347);
and (n1403,n1157,n1363);
and (n1404,n1405,n1406);
xor (n1405,n1402,n1403);
or (n1406,n1407,n1410);
and (n1407,n1408,n1409);
xor (n1408,n1352,n1353);
and (n1409,n1164,n1363);
and (n1410,n1411,n1412);
xor (n1411,n1408,n1409);
and (n1412,n1413,n1414);
xor (n1413,n1358,n1359);
and (n1414,n1170,n1363);
and (n1415,n1115,n1416);
wire s0n1416,s1n1416,notn1416;
or (n1416,s0n1416,s1n1416);
not(notn1416,n1071);
and (s0n1416,notn1416,n345);
and (s1n1416,n1071,n880);
or (n1417,n1418,n1421);
and (n1418,n1419,n1420);
xor (n1419,n1369,n1370);
and (n1420,n1122,n1416);
and (n1421,n1422,n1423);
xor (n1422,n1419,n1420);
or (n1423,n1424,n1427);
and (n1424,n1425,n1426);
xor (n1425,n1375,n1376);
and (n1426,n1129,n1416);
and (n1427,n1428,n1429);
xor (n1428,n1425,n1426);
or (n1429,n1430,n1433);
and (n1430,n1431,n1432);
xor (n1431,n1381,n1382);
and (n1432,n1136,n1416);
and (n1433,n1434,n1435);
xor (n1434,n1431,n1432);
or (n1435,n1436,n1439);
and (n1436,n1437,n1438);
xor (n1437,n1387,n1388);
and (n1438,n1143,n1416);
and (n1439,n1440,n1441);
xor (n1440,n1437,n1438);
or (n1441,n1442,n1445);
and (n1442,n1443,n1444);
xor (n1443,n1393,n1394);
and (n1444,n1150,n1416);
and (n1445,n1446,n1447);
xor (n1446,n1443,n1444);
or (n1447,n1448,n1451);
and (n1448,n1449,n1450);
xor (n1449,n1399,n1400);
and (n1450,n1157,n1416);
and (n1451,n1452,n1453);
xor (n1452,n1449,n1450);
or (n1453,n1454,n1457);
and (n1454,n1455,n1456);
xor (n1455,n1405,n1406);
and (n1456,n1164,n1416);
and (n1457,n1458,n1459);
xor (n1458,n1455,n1456);
and (n1459,n1460,n1461);
xor (n1460,n1411,n1412);
and (n1461,n1170,n1416);
and (n1462,n1122,n1463);
wire s0n1463,s1n1463,notn1463;
or (n1463,s0n1463,s1n1463);
not(notn1463,n1071);
and (s0n1463,notn1463,n392);
and (s1n1463,n1071,n927);
or (n1464,n1465,n1468);
and (n1465,n1466,n1467);
xor (n1466,n1422,n1423);
and (n1467,n1129,n1463);
and (n1468,n1469,n1470);
xor (n1469,n1466,n1467);
or (n1470,n1471,n1474);
and (n1471,n1472,n1473);
xor (n1472,n1428,n1429);
and (n1473,n1136,n1463);
and (n1474,n1475,n1476);
xor (n1475,n1472,n1473);
or (n1476,n1477,n1480);
and (n1477,n1478,n1479);
xor (n1478,n1434,n1435);
and (n1479,n1143,n1463);
and (n1480,n1481,n1482);
xor (n1481,n1478,n1479);
or (n1482,n1483,n1486);
and (n1483,n1484,n1485);
xor (n1484,n1440,n1441);
and (n1485,n1150,n1463);
and (n1486,n1487,n1488);
xor (n1487,n1484,n1485);
or (n1488,n1489,n1492);
and (n1489,n1490,n1491);
xor (n1490,n1446,n1447);
and (n1491,n1157,n1463);
and (n1492,n1493,n1494);
xor (n1493,n1490,n1491);
or (n1494,n1495,n1498);
and (n1495,n1496,n1497);
xor (n1496,n1452,n1453);
and (n1497,n1164,n1463);
and (n1498,n1499,n1500);
xor (n1499,n1496,n1497);
and (n1500,n1501,n1502);
xor (n1501,n1458,n1459);
and (n1502,n1170,n1463);
and (n1503,n1129,n1504);
wire s0n1504,s1n1504,notn1504;
or (n1504,s0n1504,s1n1504);
not(notn1504,n1071);
and (s0n1504,notn1504,n433);
and (s1n1504,n1071,n968);
or (n1505,n1506,n1509);
and (n1506,n1507,n1508);
xor (n1507,n1469,n1470);
and (n1508,n1136,n1504);
and (n1509,n1510,n1511);
xor (n1510,n1507,n1508);
or (n1511,n1512,n1515);
and (n1512,n1513,n1514);
xor (n1513,n1475,n1476);
and (n1514,n1143,n1504);
and (n1515,n1516,n1517);
xor (n1516,n1513,n1514);
or (n1517,n1518,n1521);
and (n1518,n1519,n1520);
xor (n1519,n1481,n1482);
and (n1520,n1150,n1504);
and (n1521,n1522,n1523);
xor (n1522,n1519,n1520);
or (n1523,n1524,n1527);
and (n1524,n1525,n1526);
xor (n1525,n1487,n1488);
and (n1526,n1157,n1504);
and (n1527,n1528,n1529);
xor (n1528,n1525,n1526);
or (n1529,n1530,n1533);
and (n1530,n1531,n1532);
xor (n1531,n1493,n1494);
and (n1532,n1164,n1504);
and (n1533,n1534,n1535);
xor (n1534,n1531,n1532);
and (n1535,n1536,n1537);
xor (n1536,n1499,n1500);
and (n1537,n1170,n1504);
and (n1538,n1136,n1539);
wire s0n1539,s1n1539,notn1539;
or (n1539,s0n1539,s1n1539);
not(notn1539,n1071);
and (s0n1539,notn1539,n468);
and (s1n1539,n1071,n1003);
or (n1540,n1541,n1544);
and (n1541,n1542,n1543);
xor (n1542,n1510,n1511);
and (n1543,n1143,n1539);
and (n1544,n1545,n1546);
xor (n1545,n1542,n1543);
or (n1546,n1547,n1550);
and (n1547,n1548,n1549);
xor (n1548,n1516,n1517);
and (n1549,n1150,n1539);
and (n1550,n1551,n1552);
xor (n1551,n1548,n1549);
or (n1552,n1553,n1556);
and (n1553,n1554,n1555);
xor (n1554,n1522,n1523);
and (n1555,n1157,n1539);
and (n1556,n1557,n1558);
xor (n1557,n1554,n1555);
or (n1558,n1559,n1562);
and (n1559,n1560,n1561);
xor (n1560,n1528,n1529);
and (n1561,n1164,n1539);
and (n1562,n1563,n1564);
xor (n1563,n1560,n1561);
and (n1564,n1565,n1566);
xor (n1565,n1534,n1535);
and (n1566,n1170,n1539);
and (n1567,n1143,n1568);
wire s0n1568,s1n1568,notn1568;
or (n1568,s0n1568,s1n1568);
not(notn1568,n1071);
and (s0n1568,notn1568,n497);
and (s1n1568,n1071,n1032);
or (n1569,n1570,n1573);
and (n1570,n1571,n1572);
xor (n1571,n1545,n1546);
and (n1572,n1150,n1568);
and (n1573,n1574,n1575);
xor (n1574,n1571,n1572);
or (n1575,n1576,n1579);
and (n1576,n1577,n1578);
xor (n1577,n1551,n1552);
and (n1578,n1157,n1568);
and (n1579,n1580,n1581);
xor (n1580,n1577,n1578);
or (n1581,n1582,n1585);
and (n1582,n1583,n1584);
xor (n1583,n1557,n1558);
and (n1584,n1164,n1568);
and (n1585,n1586,n1587);
xor (n1586,n1583,n1584);
and (n1587,n1588,n1589);
xor (n1588,n1563,n1564);
and (n1589,n1170,n1568);
and (n1590,n1150,n1591);
wire s0n1591,s1n1591,notn1591;
or (n1591,s0n1591,s1n1591);
not(notn1591,n1071);
and (s0n1591,notn1591,n520);
and (s1n1591,n1071,n1055);
or (n1592,n1593,n1596);
and (n1593,n1594,n1595);
xor (n1594,n1574,n1575);
and (n1595,n1157,n1591);
and (n1596,n1597,n1598);
xor (n1597,n1594,n1595);
or (n1598,n1599,n1602);
and (n1599,n1600,n1601);
xor (n1600,n1580,n1581);
and (n1601,n1164,n1591);
and (n1602,n1603,n1604);
xor (n1603,n1600,n1601);
and (n1604,n1605,n1606);
xor (n1605,n1586,n1587);
and (n1606,n1170,n1591);
endmodule
