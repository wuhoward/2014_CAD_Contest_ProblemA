module top (out,n4,n6,n7,n8,n28,n29,n33,n40,n47
        ,n48,n56,n58,n68,n76,n78,n84,n89,n94,n106
        ,n107,n113,n119,n134,n135,n142,n146,n152,n161,n166
        ,n170,n176,n189,n197,n207,n208,n215,n219,n225,n246
        ,n255,n276,n286,n287,n298,n311,n323,n348,n358,n369
        ,n374,n395,n422,n432,n444);
output out;
input n4;
input n6;
input n7;
input n8;
input n28;
input n29;
input n33;
input n40;
input n47;
input n48;
input n56;
input n58;
input n68;
input n76;
input n78;
input n84;
input n89;
input n94;
input n106;
input n107;
input n113;
input n119;
input n134;
input n135;
input n142;
input n146;
input n152;
input n161;
input n166;
input n170;
input n176;
input n189;
input n197;
input n207;
input n208;
input n215;
input n219;
input n225;
input n246;
input n255;
input n276;
input n286;
input n287;
input n298;
input n311;
input n323;
input n348;
input n358;
input n369;
input n374;
input n395;
input n422;
input n432;
input n444;
wire n0;
wire n1;
wire n2;
wire n3;
wire n5;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n24;
wire n25;
wire n26;
wire n27;
wire n30;
wire n31;
wire n32;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n57;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n77;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n85;
wire n86;
wire n87;
wire n88;
wire n90;
wire n91;
wire n92;
wire n93;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n143;
wire n144;
wire n145;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n162;
wire n163;
wire n164;
wire n165;
wire n167;
wire n168;
wire n169;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n216;
wire n217;
wire n218;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n370;
wire n371;
wire n372;
wire n373;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2988;
wire n2989;
wire n2990;
wire n2991;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2996;
wire n2997;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3003;
wire n3004;
wire n3005;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3010;
wire n3011;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3038;
wire n3039;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
wire n3056;
wire n3057;
wire n3058;
wire n3059;
wire n3060;
wire n3061;
wire n3062;
wire n3063;
wire n3064;
wire n3065;
wire n3066;
wire n3067;
wire n3068;
wire n3069;
wire n3070;
wire n3071;
wire n3072;
wire n3073;
wire n3074;
wire n3075;
wire n3076;
wire n3077;
wire n3078;
wire n3079;
wire n3080;
wire n3081;
wire n3082;
wire n3083;
wire n3084;
wire n3085;
wire n3086;
wire n3087;
wire n3088;
wire n3089;
wire n3090;
wire n3091;
wire n3092;
wire n3093;
wire n3094;
wire n3095;
wire n3096;
wire n3097;
wire n3098;
wire n3099;
wire n3100;
wire n3101;
wire n3102;
wire n3103;
wire n3104;
wire n3105;
wire n3106;
wire n3107;
wire n3108;
wire n3109;
wire n3110;
wire n3111;
wire n3112;
wire n3113;
wire n3114;
wire n3115;
wire n3116;
wire n3117;
wire n3118;
wire n3119;
wire n3120;
wire n3121;
wire n3122;
wire n3123;
wire n3124;
wire n3125;
wire n3126;
wire n3127;
wire n3128;
wire n3129;
wire n3130;
wire n3131;
wire n3132;
wire n3133;
wire n3134;
wire n3135;
wire n3136;
wire n3137;
wire n3138;
wire n3139;
wire n3140;
wire n3141;
wire n3142;
wire n3143;
wire n3144;
wire n3145;
wire n3146;
wire n3147;
wire n3148;
wire n3149;
wire n3150;
wire n3151;
wire n3152;
wire n3153;
wire n3154;
wire n3155;
wire n3156;
wire n3157;
wire n3158;
wire n3159;
wire n3160;
wire n3161;
wire n3162;
wire n3163;
wire n3164;
wire n3165;
wire n3166;
wire n3167;
wire n3168;
wire n3169;
wire n3170;
wire n3171;
wire n3172;
wire n3173;
wire n3174;
wire n3175;
wire n3176;
wire n3177;
wire n3178;
wire n3179;
wire n3180;
wire n3181;
wire n3182;
wire n3183;
wire n3184;
wire n3185;
wire n3186;
wire n3187;
wire n3188;
wire n3189;
wire n3190;
wire n3191;
wire n3192;
wire n3193;
wire n3194;
wire n3195;
wire n3196;
wire n3197;
wire n3198;
wire n3199;
wire n3200;
wire n3201;
wire n3202;
wire n3203;
wire n3204;
wire n3205;
wire n3206;
wire n3207;
wire n3208;
wire n3209;
wire n3210;
wire n3211;
wire n3212;
wire n3213;
wire n3214;
wire n3215;
wire n3216;
wire n3217;
wire n3218;
wire n3219;
wire n3220;
wire n3221;
wire n3222;
wire n3223;
wire n3224;
wire n3225;
wire n3226;
wire n3227;
wire n3228;
wire n3229;
wire n3230;
wire n3231;
wire n3232;
wire n3233;
wire n3234;
wire n3235;
wire n3236;
wire n3237;
wire n3238;
wire n3239;
wire n3240;
wire n3241;
wire n3242;
wire n3243;
wire n3244;
wire n3245;
wire n3246;
wire n3247;
wire n3248;
wire n3249;
wire n3250;
wire n3251;
wire n3252;
wire n3253;
wire n3254;
wire n3255;
wire n3256;
wire n3257;
wire n3258;
wire n3259;
wire n3260;
wire n3261;
wire n3262;
wire n3263;
wire n3264;
wire n3265;
wire n3266;
wire n3267;
wire n3268;
wire n3269;
wire n3270;
wire n3271;
wire n3272;
wire n3273;
wire n3274;
wire n3275;
wire n3276;
wire n3277;
wire n3278;
wire n3279;
wire n3280;
wire n3281;
wire n3282;
wire n3283;
wire n3284;
wire n3285;
wire n3286;
wire n3287;
wire n3288;
wire n3289;
wire n3290;
wire n3291;
wire n3292;
wire n3293;
wire n3294;
wire n3295;
wire n3296;
wire n3297;
wire n3298;
wire n3299;
wire n3300;
wire n3301;
wire n3302;
wire n3303;
wire n3304;
wire n3305;
wire n3306;
wire n3307;
wire n3308;
wire n3309;
wire n3310;
wire n3311;
wire n3312;
wire n3313;
wire n3314;
wire n3315;
wire n3316;
wire n3317;
wire n3318;
wire n3319;
wire n3320;
wire n3321;
wire n3322;
wire n3323;
wire n3324;
wire n3325;
wire n3326;
wire n3327;
wire n3328;
wire n3329;
wire n3330;
wire n3331;
wire n3332;
wire n3333;
wire n3334;
wire n3335;
wire n3336;
wire n3337;
wire n3338;
wire n3339;
wire n3340;
wire n3341;
wire n3342;
wire n3343;
wire n3344;
wire n3345;
wire n3346;
wire n3347;
wire n3348;
wire n3349;
wire n3350;
wire n3351;
wire n3352;
wire n3353;
wire n3354;
wire n3355;
wire n3356;
wire n3357;
wire n3358;
wire n3359;
wire n3360;
wire n3361;
wire n3362;
wire n3363;
wire n3364;
wire n3365;
wire n3366;
wire n3367;
wire n3368;
wire n3369;
wire n3370;
wire n3371;
wire n3372;
wire n3373;
wire n3374;
wire n3375;
wire n3376;
wire n3377;
wire n3378;
wire n3379;
wire n3380;
wire n3381;
wire n3382;
wire n3383;
wire n3384;
wire n3385;
wire n3386;
wire n3387;
wire n3388;
wire n3389;
wire n3390;
wire n3391;
wire n3392;
wire n3393;
wire n3394;
wire n3395;
wire n3396;
wire n3397;
wire n3398;
wire n3399;
wire n3400;
wire n3401;
wire n3402;
wire n3403;
wire n3404;
wire n3405;
wire n3406;
wire n3407;
wire n3408;
wire n3409;
wire n3410;
wire n3411;
wire n3412;
wire n3413;
wire n3414;
wire n3415;
wire n3416;
wire n3417;
wire n3418;
wire n3419;
wire n3420;
wire n3421;
wire n3422;
wire n3423;
wire n3424;
wire n3425;
wire n3426;
wire n3427;
wire n3428;
wire n3429;
wire n3430;
wire n3431;
wire n3432;
wire n3433;
wire n3434;
wire n3435;
wire n3436;
wire n3437;
wire n3438;
wire n3439;
wire n3440;
wire n3441;
wire n3442;
wire n3443;
wire n3444;
wire n3445;
wire n3446;
wire n3447;
wire n3448;
wire n3449;
wire n3450;
wire n3451;
wire n3452;
wire n3453;
wire n3454;
wire n3455;
wire n3456;
wire n3457;
wire n3458;
wire n3459;
wire n3460;
wire n3461;
wire n3462;
wire n3463;
wire n3464;
wire n3465;
wire n3466;
wire n3467;
wire n3468;
wire n3469;
wire n3470;
wire n3471;
wire n3472;
wire n3473;
wire n3474;
wire n3475;
wire n3476;
wire n3477;
wire n3478;
wire n3479;
wire n3480;
wire n3481;
wire n3482;
wire n3483;
wire n3484;
wire n3485;
wire n3486;
wire n3487;
wire n3488;
wire n3489;
wire n3490;
wire n3491;
wire n3492;
wire n3493;
wire n3494;
wire n3495;
wire n3496;
wire n3497;
wire n3498;
wire n3499;
wire n3500;
wire n3501;
wire n3502;
wire n3503;
wire n3504;
wire n3505;
wire n3506;
wire n3507;
wire n3508;
wire n3509;
wire n3510;
wire n3511;
wire n3512;
wire n3513;
wire n3514;
wire n3515;
wire n3516;
wire n3517;
wire n3518;
wire n3519;
wire n3520;
wire n3521;
wire n3522;
wire n3523;
wire n3524;
wire n3525;
wire n3526;
wire n3527;
wire n3528;
wire n3529;
wire n3530;
wire n3531;
wire n3532;
wire n3533;
wire n3534;
wire n3535;
wire n3536;
wire n3537;
wire n3538;
wire n3539;
wire n3540;
wire n3541;
wire n3542;
wire n3543;
wire n3544;
wire n3545;
wire n3546;
wire n3547;
wire n3548;
wire n3549;
wire n3550;
wire n3551;
wire n3552;
wire n3553;
wire n3554;
wire n3555;
wire n3556;
wire n3557;
wire n3558;
wire n3559;
wire n3560;
wire n3561;
wire n3562;
wire n3563;
wire n3564;
wire n3565;
wire n3566;
wire n3567;
wire n3568;
wire n3569;
wire n3570;
wire n3571;
wire n3572;
wire n3573;
wire n3574;
wire n3575;
wire n3576;
wire n3577;
wire n3578;
wire n3579;
wire n3580;
wire n3581;
wire n3582;
wire n3583;
wire n3584;
wire n3585;
wire n3586;
wire n3587;
wire n3588;
wire n3589;
wire n3590;
wire n3591;
wire n3592;
wire n3593;
wire n3594;
wire n3595;
wire n3596;
wire n3597;
wire n3598;
wire n3599;
wire n3600;
wire n3601;
wire n3602;
wire n3603;
wire n3604;
wire n3605;
wire n3606;
wire n3607;
wire n3608;
wire n3609;
wire n3610;
wire n3611;
wire n3612;
wire n3613;
wire n3614;
wire n3615;
wire n3616;
wire n3617;
wire n3618;
wire n3619;
wire n3620;
wire n3621;
wire n3622;
wire n3623;
wire n3624;
wire n3625;
wire n3626;
wire n3627;
wire n3628;
wire n3629;
wire n3630;
wire n3631;
wire n3632;
wire n3633;
wire n3634;
wire n3635;
wire n3636;
wire n3637;
wire n3638;
wire n3639;
wire n3640;
wire n3641;
wire n3642;
wire n3643;
wire n3644;
wire n3645;
wire n3646;
wire n3647;
wire n3648;
wire n3649;
wire n3650;
wire n3651;
wire n3652;
wire n3653;
wire n3654;
wire n3655;
wire n3656;
wire n3657;
wire n3658;
wire n3659;
wire n3660;
wire n3661;
wire n3662;
wire n3663;
wire n3664;
wire n3665;
wire n3666;
wire n3667;
wire n3668;
wire n3669;
wire n3670;
wire n3671;
wire n3672;
wire n3673;
wire n3674;
wire n3675;
xor (out,n0,n2038);
or (n0,n1,n9);
and (n1,n2,n8);
nand (n2,n3,n5,n7);
not (n3,n4);
not (n5,n6);
and (n9,n10,n11);
not (n10,n2);
xnor (n11,n12,n871);
nand (n12,n13,n870);
not (n13,n14);
nor (n14,n15,n696);
xor (n15,n16,n648);
xor (n16,n17,n410);
xor (n17,n18,n327);
xor (n18,n19,n228);
xor (n19,n20,n180);
xor (n20,n21,n98);
or (n21,n22,n97);
and (n22,n23,n70);
xor (n23,n24,n42);
nand (n24,n25,n36);
or (n25,n26,n30);
nand (n26,n27,n29);
not (n27,n28);
nor (n30,n31,n34);
and (n31,n32,n29);
not (n32,n33);
and (n34,n33,n35);
not (n35,n29);
or (n36,n37,n27);
nor (n37,n38,n41);
and (n38,n39,n29);
not (n39,n40);
and (n41,n40,n35);
nand (n42,n43,n64);
or (n43,n44,n52);
not (n44,n45);
nor (n45,n46,n49);
and (n46,n47,n48);
and (n49,n50,n51);
not (n50,n47);
not (n51,n48);
not (n52,n53);
nor (n53,n54,n61);
nand (n54,n55,n59);
or (n55,n56,n57);
not (n57,n58);
or (n59,n58,n60);
not (n60,n56);
nor (n61,n62,n63);
and (n62,n51,n56);
and (n63,n48,n60);
nand (n64,n54,n65);
nand (n65,n66,n69);
or (n66,n48,n67);
not (n67,n68);
or (n69,n51,n68);
nand (n70,n71,n91);
or (n71,n72,n86);
not (n72,n73);
and (n73,n74,n81);
and (n74,n75,n79);
nand (n75,n76,n77);
not (n77,n78);
nand (n79,n78,n80);
not (n80,n76);
nor (n81,n82,n85);
and (n82,n77,n83);
not (n83,n84);
and (n85,n78,n84);
nor (n86,n87,n90);
and (n87,n88,n84);
not (n88,n89);
and (n90,n89,n83);
or (n91,n74,n92);
nor (n92,n93,n95);
and (n93,n83,n94);
and (n95,n84,n96);
not (n96,n94);
and (n97,n24,n42);
or (n98,n99,n179);
and (n99,n100,n155);
xor (n100,n101,n127);
nand (n101,n102,n115);
or (n102,n103,n110);
nor (n103,n104,n108);
and (n104,n105,n107);
not (n105,n106);
and (n108,n106,n109);
not (n109,n107);
not (n110,n111);
nand (n111,n112,n114);
or (n112,n113,n51);
nand (n114,n113,n51);
nand (n115,n116,n122);
not (n116,n117);
nor (n117,n118,n120);
and (n118,n119,n105);
and (n120,n121,n106);
not (n121,n119);
nor (n122,n111,n123);
nor (n123,n124,n125);
and (n124,n105,n113);
and (n125,n106,n126);
not (n126,n113);
nand (n127,n128,n149);
or (n128,n129,n144);
nand (n129,n130,n138);
not (n130,n131);
nor (n131,n132,n136);
and (n132,n133,n135);
not (n133,n134);
and (n136,n134,n137);
not (n137,n135);
not (n138,n139);
nand (n139,n140,n143);
or (n140,n141,n134);
not (n141,n142);
nand (n143,n134,n141);
nor (n144,n145,n147);
and (n145,n137,n146);
and (n147,n135,n148);
not (n148,n146);
or (n149,n138,n150);
nor (n150,n151,n153);
and (n151,n137,n152);
and (n153,n135,n154);
not (n154,n152);
nand (n155,n156,n173);
or (n156,n157,n168);
nand (n157,n158,n163);
and (n158,n159,n162);
nand (n159,n135,n160);
not (n160,n161);
nand (n162,n161,n137);
nand (n163,n164,n167);
or (n164,n161,n165);
not (n165,n166);
nand (n167,n161,n165);
nor (n168,n169,n171);
and (n169,n165,n170);
and (n171,n166,n172);
not (n172,n170);
or (n173,n158,n174);
nor (n174,n175,n177);
and (n175,n165,n176);
and (n177,n166,n178);
not (n178,n176);
and (n179,n101,n127);
xor (n180,n181,n200);
xor (n181,n182,n192);
nand (n182,n183,n185);
or (n183,n184,n52);
not (n184,n65);
nand (n185,n186,n54);
not (n186,n187);
nor (n187,n188,n190);
and (n188,n51,n189);
and (n190,n48,n191);
not (n191,n189);
nand (n192,n193,n194);
or (n193,n72,n92);
or (n194,n74,n195);
nor (n195,n196,n198);
and (n196,n197,n83);
and (n198,n84,n199);
not (n199,n197);
nand (n200,n201,n222);
or (n201,n202,n217);
not (n202,n203);
nor (n203,n204,n211);
nor (n204,n205,n209);
and (n205,n206,n208);
not (n206,n207);
and (n209,n207,n210);
not (n210,n208);
not (n211,n212);
nor (n212,n213,n216);
and (n213,n214,n208);
not (n214,n215);
and (n216,n215,n210);
nor (n217,n218,n220);
and (n218,n206,n219);
and (n220,n207,n221);
not (n221,n219);
or (n222,n212,n223);
nor (n223,n224,n226);
and (n224,n206,n225);
and (n226,n207,n227);
not (n227,n225);
or (n228,n229,n326);
and (n229,n230,n269);
xor (n230,n231,n268);
or (n231,n232,n267);
and (n232,n233,n249);
xor (n233,n234,n240);
nand (n234,n235,n239);
or (n235,n129,n236);
nor (n236,n237,n238);
and (n237,n178,n135);
and (n238,n176,n137);
or (n239,n144,n138);
nand (n240,n241,n248);
or (n241,n242,n157);
not (n242,n243);
nand (n243,n244,n247);
or (n244,n166,n245);
not (n245,n246);
or (n247,n165,n246);
or (n248,n158,n168);
nand (n249,n250,n263);
or (n250,n251,n260);
nand (n251,n252,n257);
and (n252,n253,n256);
nand (n253,n106,n254);
not (n254,n255);
nand (n256,n255,n105);
nand (n257,n258,n259);
or (n258,n255,n214);
nand (n259,n214,n255);
nor (n260,n261,n262);
and (n261,n214,n219);
and (n262,n215,n221);
or (n263,n252,n264);
nor (n264,n265,n266);
and (n265,n214,n225);
and (n266,n215,n227);
and (n267,n234,n240);
xor (n268,n23,n70);
xor (n269,n270,n304);
xor (n270,n271,n279);
nand (n271,n272,n273);
or (n272,n251,n264);
or (n273,n252,n274);
nor (n274,n275,n277);
and (n275,n214,n276);
and (n277,n215,n278);
not (n278,n276);
nand (n279,n280,n300);
or (n280,n281,n294);
nand (n281,n282,n290);
not (n282,n283);
nor (n283,n284,n288);
and (n284,n285,n287);
not (n285,n286);
and (n288,n286,n289);
not (n289,n287);
not (n290,n291);
nand (n291,n292,n293);
or (n292,n287,n165);
nand (n293,n165,n287);
not (n294,n295);
nor (n295,n296,n299);
and (n296,n297,n285);
not (n297,n298);
and (n299,n298,n286);
or (n300,n290,n301);
nor (n301,n302,n303);
and (n302,n285,n246);
and (n303,n286,n245);
nand (n304,n305,n319);
or (n305,n306,n316);
not (n306,n307);
nor (n307,n308,n313);
nand (n308,n309,n312);
or (n309,n286,n310);
not (n310,n311);
nand (n312,n286,n310);
nor (n313,n314,n315);
and (n314,n311,n80);
and (n315,n76,n310);
nor (n316,n317,n318);
and (n317,n80,n197);
and (n318,n76,n199);
or (n319,n320,n321);
not (n320,n308);
nor (n321,n322,n324);
and (n322,n80,n323);
and (n324,n76,n325);
not (n325,n323);
and (n326,n231,n268);
xor (n327,n328,n388);
xor (n328,n329,n351);
xor (n329,n330,n343);
xor (n330,n331,n337);
nand (n331,n332,n333);
or (n332,n281,n301);
or (n333,n290,n334);
nor (n334,n335,n336);
and (n335,n285,n170);
and (n336,n286,n172);
nand (n337,n338,n339);
or (n338,n306,n321);
or (n339,n320,n340);
nor (n340,n341,n342);
and (n341,n80,n298);
and (n342,n76,n297);
nand (n343,n344,n345);
or (n344,n26,n37);
or (n345,n346,n27);
nor (n346,n347,n349);
and (n347,n35,n348);
and (n349,n29,n350);
not (n350,n348);
xor (n351,n352,n381);
xor (n352,n353,n360);
nor (n353,n354,n88);
not (n354,n355);
nand (n355,n356,n359);
or (n356,n357,n84);
not (n357,n358);
nand (n359,n84,n357);
nand (n360,n361,n371);
or (n361,n362,n366);
not (n362,n363);
nand (n363,n364,n365);
or (n364,n58,n32);
or (n365,n57,n33);
nor (n366,n367,n370);
and (n367,n29,n368);
not (n368,n369);
and (n370,n35,n369);
or (n371,n372,n377);
nor (n372,n373,n375);
and (n373,n57,n374);
and (n375,n58,n376);
not (n376,n374);
nand (n377,n366,n378);
nand (n378,n379,n380);
or (n379,n369,n57);
nand (n380,n57,n369);
nand (n381,n382,n384);
or (n382,n383,n103);
not (n383,n122);
or (n384,n110,n385);
nor (n385,n386,n387);
and (n386,n105,n47);
and (n387,n106,n50);
xor (n388,n389,n404);
xor (n389,n390,n398);
nand (n390,n391,n392);
or (n391,n129,n150);
or (n392,n138,n393);
nor (n393,n394,n396);
and (n394,n137,n395);
and (n396,n135,n397);
not (n397,n395);
nand (n398,n399,n400);
or (n399,n157,n174);
or (n400,n158,n401);
nor (n401,n402,n403);
and (n402,n165,n146);
and (n403,n166,n148);
nand (n404,n405,n406);
or (n405,n251,n274);
or (n406,n252,n407);
nor (n407,n408,n409);
and (n408,n214,n119);
and (n409,n215,n121);
xor (n410,n411,n612);
xor (n411,n412,n544);
or (n412,n413,n543);
and (n413,n414,n460);
xor (n414,n415,n416);
xor (n415,n100,n155);
xor (n416,n417,n447);
xor (n417,n418,n426);
nand (n418,n419,n425);
or (n419,n202,n420);
nor (n420,n421,n423);
and (n421,n206,n422);
and (n423,n207,n424);
not (n424,n422);
or (n425,n212,n217);
nand (n426,n427,n441);
or (n427,n428,n438);
nand (n428,n429,n434);
not (n429,n430);
nand (n430,n431,n433);
or (n431,n432,n206);
nand (n433,n206,n432);
nand (n434,n435,n437);
or (n435,n142,n436);
not (n436,n432);
nand (n437,n142,n436);
nor (n438,n439,n440);
and (n439,n141,n395);
and (n440,n142,n397);
or (n441,n429,n442);
nor (n442,n443,n445);
and (n443,n141,n444);
and (n445,n142,n446);
not (n446,n444);
xor (n447,n448,n454);
and (n448,n449,n84);
nand (n449,n450,n451);
or (n450,n89,n78);
nand (n451,n452,n80);
not (n452,n453);
and (n453,n89,n78);
nand (n454,n455,n459);
or (n455,n377,n456);
nor (n456,n457,n458);
and (n457,n57,n189);
and (n458,n58,n191);
or (n459,n366,n372);
or (n460,n461,n542);
and (n461,n462,n513);
xor (n462,n463,n481);
nor (n463,n464,n475);
not (n464,n465);
nand (n465,n466,n470);
or (n466,n467,n377);
nor (n467,n468,n469);
and (n468,n57,n47);
and (n469,n58,n50);
nand (n470,n471,n472);
not (n471,n366);
nand (n472,n473,n474);
or (n473,n58,n67);
or (n474,n57,n68);
nand (n475,n476,n76);
nand (n476,n477,n478);
or (n477,n89,n311);
nand (n478,n479,n285);
not (n479,n480);
and (n480,n89,n311);
or (n481,n482,n512);
and (n482,n483,n503);
xor (n483,n484,n494);
nand (n484,n485,n490);
or (n485,n26,n486);
not (n486,n487);
nor (n487,n488,n489);
and (n488,n191,n35);
and (n489,n189,n29);
or (n490,n491,n27);
nor (n491,n492,n493);
and (n492,n35,n374);
and (n493,n29,n376);
nand (n494,n495,n499);
or (n495,n52,n496);
nor (n496,n497,n498);
and (n497,n51,n119);
and (n498,n48,n121);
nand (n499,n54,n500);
nand (n500,n501,n502);
or (n501,n48,n109);
or (n502,n51,n107);
nand (n503,n504,n508);
or (n504,n202,n505);
nor (n505,n506,n507);
and (n506,n206,n395);
and (n507,n207,n397);
or (n508,n212,n509);
nor (n509,n510,n511);
and (n510,n206,n444);
and (n511,n207,n446);
and (n512,n484,n494);
or (n513,n514,n541);
and (n514,n515,n532);
xor (n515,n516,n522);
nand (n516,n517,n521);
or (n517,n251,n518);
nor (n518,n519,n520);
and (n519,n424,n215);
and (n520,n422,n214);
or (n521,n252,n260);
nand (n522,n523,n527);
or (n523,n281,n524);
nor (n524,n525,n526);
and (n525,n285,n197);
and (n526,n286,n199);
or (n527,n290,n528);
not (n528,n529);
nand (n529,n530,n531);
or (n530,n286,n325);
or (n531,n285,n323);
nand (n532,n533,n537);
or (n533,n306,n534);
nor (n534,n535,n536);
and (n535,n88,n76);
and (n536,n89,n80);
or (n537,n320,n538);
nor (n538,n539,n540);
and (n539,n96,n76);
and (n540,n94,n80);
and (n541,n516,n522);
and (n542,n463,n481);
and (n543,n415,n416);
xor (n544,n545,n600);
xor (n545,n546,n549);
or (n546,n547,n548);
and (n547,n417,n447);
and (n548,n418,n426);
or (n549,n550,n599);
and (n550,n551,n583);
xor (n551,n552,n566);
or (n552,n553,n565);
and (n553,n554,n562);
xor (n554,n555,n558);
nand (n555,n556,n557);
or (n556,n528,n281);
nand (n557,n295,n291);
nand (n558,n559,n560);
or (n559,n320,n316);
nand (n560,n561,n307);
not (n561,n538);
nand (n562,n563,n564);
or (n563,n26,n491);
or (n564,n30,n27);
and (n565,n555,n558);
or (n566,n567,n582);
and (n567,n568,n576);
xor (n568,n569,n573);
nand (n569,n570,n572);
or (n570,n571,n52);
not (n571,n500);
nand (n572,n54,n45);
nand (n573,n574,n575);
or (n574,n509,n202);
or (n575,n212,n420);
nand (n576,n577,n581);
or (n577,n428,n578);
nor (n578,n579,n580);
and (n579,n141,n152);
and (n580,n142,n154);
or (n581,n429,n438);
and (n582,n569,n573);
or (n583,n584,n598);
and (n584,n585,n592);
xor (n585,n586,n587);
nor (n586,n74,n88);
nand (n587,n588,n590);
or (n588,n589,n377);
not (n589,n472);
nand (n590,n591,n471);
not (n591,n456);
nand (n592,n593,n597);
or (n593,n383,n594);
nor (n594,n595,n596);
and (n595,n105,n276);
and (n596,n106,n278);
or (n597,n110,n117);
and (n598,n586,n587);
and (n599,n552,n566);
xor (n600,n601,n609);
xor (n601,n602,n608);
nand (n602,n603,n604);
or (n603,n428,n442);
or (n604,n429,n605);
nor (n605,n606,n607);
and (n606,n141,n422);
and (n607,n142,n424);
and (n608,n448,n454);
or (n609,n610,n611);
and (n610,n270,n304);
and (n611,n271,n279);
or (n612,n613,n647);
and (n613,n614,n646);
xor (n614,n615,n616);
xor (n615,n551,n583);
or (n616,n617,n645);
and (n617,n618,n644);
xor (n618,n619,n643);
or (n619,n620,n642);
and (n620,n621,n636);
xor (n621,n622,n630);
nand (n622,n623,n628);
or (n623,n624,n383);
not (n624,n625);
nand (n625,n626,n627);
or (n626,n106,n227);
or (n627,n105,n225);
nand (n628,n629,n111);
not (n629,n594);
nand (n630,n631,n635);
or (n631,n129,n632);
nor (n632,n633,n634);
and (n633,n137,n170);
and (n634,n135,n172);
or (n635,n138,n236);
nand (n636,n637,n641);
or (n637,n157,n638);
nor (n638,n639,n640);
and (n639,n165,n298);
and (n640,n166,n297);
or (n641,n158,n242);
and (n642,n622,n630);
xor (n643,n568,n576);
xor (n644,n233,n249);
and (n645,n619,n643);
xor (n646,n230,n269);
and (n647,n615,n616);
or (n648,n649,n695);
and (n649,n650,n694);
xor (n650,n651,n652);
xor (n651,n414,n460);
or (n652,n653,n693);
and (n653,n654,n657);
xor (n654,n655,n656);
xor (n655,n554,n562);
xor (n656,n585,n592);
or (n657,n658,n692);
and (n658,n659,n670);
xor (n659,n660,n666);
nand (n660,n661,n665);
or (n661,n428,n662);
nor (n662,n663,n664);
and (n663,n141,n146);
and (n664,n148,n142);
or (n665,n429,n578);
nand (n666,n667,n669);
or (n667,n668,n464);
not (n668,n475);
or (n669,n465,n475);
or (n670,n671,n691);
and (n671,n672,n685);
xor (n672,n673,n679);
nand (n673,n674,n678);
or (n674,n129,n675);
nor (n675,n676,n677);
and (n676,n137,n246);
and (n677,n135,n245);
or (n678,n138,n632);
nand (n679,n680,n684);
or (n680,n157,n681);
nor (n681,n682,n683);
and (n682,n165,n323);
and (n683,n166,n325);
or (n684,n158,n638);
nand (n685,n686,n690);
or (n686,n377,n687);
nor (n687,n688,n689);
and (n688,n57,n107);
and (n689,n58,n109);
or (n690,n366,n467);
and (n691,n673,n679);
and (n692,n660,n666);
and (n693,n655,n656);
xor (n694,n614,n646);
and (n695,n651,n652);
or (n696,n697,n869);
and (n697,n698,n868);
xor (n698,n699,n784);
or (n699,n700,n783);
and (n700,n701,n747);
xor (n701,n702,n746);
or (n702,n703,n745);
and (n703,n704,n744);
xor (n704,n705,n721);
or (n705,n706,n720);
and (n706,n707,n715);
xor (n707,n708,n709);
nor (n708,n320,n88);
nand (n709,n710,n711);
or (n710,n27,n486);
or (n711,n26,n712);
nor (n712,n713,n714);
and (n713,n35,n68);
and (n714,n29,n67);
nand (n715,n716,n719);
or (n716,n383,n717);
not (n717,n718);
xor (n718,n219,n106);
or (n719,n110,n624);
and (n720,n708,n709);
or (n721,n722,n743);
and (n722,n723,n736);
xor (n723,n724,n730);
nand (n724,n725,n729);
or (n725,n281,n726);
nor (n726,n727,n728);
and (n727,n285,n94);
and (n728,n286,n96);
or (n729,n290,n524);
nand (n730,n731,n735);
or (n731,n251,n732);
nor (n732,n733,n734);
and (n733,n214,n444);
and (n734,n215,n446);
or (n735,n252,n518);
nand (n736,n737,n741);
or (n737,n52,n738);
nor (n738,n739,n740);
and (n739,n51,n276);
and (n740,n48,n278);
or (n741,n742,n496);
not (n742,n54);
and (n743,n724,n730);
xor (n744,n483,n503);
and (n745,n705,n721);
xor (n746,n462,n513);
or (n747,n748,n782);
and (n748,n749,n752);
xor (n749,n750,n751);
xor (n750,n621,n636);
xor (n751,n515,n532);
or (n752,n753,n781);
and (n753,n754,n767);
xor (n754,n755,n761);
nand (n755,n756,n760);
or (n756,n202,n757);
nor (n757,n758,n759);
and (n758,n206,n152);
and (n759,n207,n154);
or (n760,n212,n505);
nand (n761,n762,n766);
or (n762,n428,n763);
nor (n763,n764,n765);
and (n764,n141,n176);
and (n765,n142,n178);
or (n766,n429,n662);
and (n767,n768,n774);
nor (n768,n769,n285);
nor (n769,n770,n773);
and (n770,n771,n165);
not (n771,n772);
and (n772,n89,n287);
and (n773,n88,n289);
nand (n774,n775,n780);
or (n775,n26,n776);
not (n776,n777);
nor (n777,n778,n779);
and (n778,n47,n29);
and (n779,n50,n35);
or (n780,n712,n27);
and (n781,n755,n761);
and (n782,n750,n751);
and (n783,n702,n746);
or (n784,n785,n867);
and (n785,n786,n789);
xor (n786,n787,n788);
xor (n787,n618,n644);
xor (n788,n654,n657);
or (n789,n790,n866);
and (n790,n791,n865);
xor (n791,n792,n864);
or (n792,n793,n863);
and (n793,n794,n841);
xor (n794,n795,n818);
or (n795,n796,n817);
and (n796,n797,n811);
xor (n797,n798,n805);
nand (n798,n799,n804);
or (n799,n800,n383);
not (n800,n801);
nor (n801,n802,n803);
and (n802,n422,n106);
and (n803,n424,n105);
nand (n804,n111,n718);
nand (n805,n806,n810);
or (n806,n807,n129);
nor (n807,n808,n809);
and (n808,n297,n135);
and (n809,n298,n137);
or (n810,n138,n675);
nand (n811,n812,n816);
or (n812,n157,n813);
nor (n813,n814,n815);
and (n814,n165,n197);
and (n815,n166,n199);
or (n816,n158,n681);
and (n817,n798,n805);
or (n818,n819,n840);
and (n819,n820,n834);
xor (n820,n821,n828);
nand (n821,n822,n826);
or (n822,n52,n823);
nor (n823,n824,n825);
and (n824,n227,n48);
and (n825,n225,n51);
nand (n826,n827,n54);
not (n827,n738);
nand (n828,n829,n833);
or (n829,n202,n830);
nor (n830,n831,n832);
and (n831,n206,n146);
and (n832,n207,n148);
or (n833,n212,n757);
nand (n834,n835,n839);
or (n835,n428,n836);
nor (n836,n837,n838);
and (n837,n141,n170);
and (n838,n142,n172);
or (n839,n429,n763);
and (n840,n821,n828);
or (n841,n842,n862);
and (n842,n843,n856);
xor (n843,n844,n850);
nand (n844,n845,n849);
or (n845,n377,n846);
nor (n846,n847,n848);
and (n847,n57,n119);
and (n848,n58,n121);
or (n849,n366,n687);
nand (n850,n851,n855);
or (n851,n281,n852);
nor (n852,n853,n854);
and (n853,n88,n286);
and (n854,n89,n285);
or (n855,n290,n726);
nand (n856,n857,n861);
or (n857,n251,n858);
nor (n858,n859,n860);
and (n859,n214,n395);
and (n860,n215,n397);
or (n861,n252,n732);
and (n862,n844,n850);
and (n863,n795,n818);
xor (n864,n659,n670);
xor (n865,n704,n744);
and (n866,n792,n864);
and (n867,n787,n788);
xor (n868,n650,n694);
and (n869,n699,n784);
nand (n870,n15,n696);
nand (n871,n872,n1519);
nor (n872,n873,n1505);
and (n873,n874,n1190);
and (n874,n875,n1173);
nor (n875,n876,n1088);
nor (n876,n877,n976);
xor (n877,n878,n969);
xor (n878,n879,n958);
or (n879,n880,n957);
and (n880,n881,n928);
xor (n881,n882,n883);
xor (n882,n754,n767);
or (n883,n884,n927);
and (n884,n885,n905);
xor (n885,n886,n887);
xor (n886,n768,n774);
or (n887,n888,n904);
and (n888,n889,n898);
xor (n889,n890,n891);
and (n890,n291,n89);
nand (n891,n892,n897);
or (n892,n26,n893);
not (n893,n894);
nor (n894,n895,n896);
and (n895,n107,n29);
and (n896,n109,n35);
nand (n897,n777,n28);
nand (n898,n899,n903);
or (n899,n383,n900);
nor (n900,n901,n902);
and (n901,n105,n444);
and (n902,n106,n446);
or (n903,n110,n800);
and (n904,n890,n891);
or (n905,n906,n926);
and (n906,n907,n920);
xor (n907,n908,n914);
nand (n908,n909,n913);
or (n909,n129,n910);
nor (n910,n911,n912);
and (n911,n137,n323);
and (n912,n135,n325);
or (n913,n138,n807);
nand (n914,n915,n919);
or (n915,n157,n916);
nor (n916,n917,n918);
and (n917,n165,n94);
and (n918,n166,n96);
or (n919,n158,n813);
nand (n920,n921,n925);
or (n921,n377,n922);
nor (n922,n923,n924);
and (n923,n57,n276);
and (n924,n58,n278);
or (n925,n366,n846);
and (n926,n908,n914);
and (n927,n886,n887);
or (n928,n929,n956);
and (n929,n930,n955);
xor (n930,n931,n954);
or (n931,n932,n953);
and (n932,n933,n947);
xor (n933,n934,n940);
nand (n934,n935,n939);
or (n935,n936,n251);
nor (n936,n937,n938);
and (n937,n214,n152);
and (n938,n215,n154);
or (n939,n252,n858);
nand (n940,n941,n945);
or (n941,n942,n52);
nor (n942,n943,n944);
and (n943,n51,n219);
and (n944,n48,n221);
nand (n945,n946,n54);
not (n946,n823);
nand (n947,n948,n952);
or (n948,n202,n949);
nor (n949,n950,n951);
and (n950,n206,n176);
and (n951,n207,n178);
or (n952,n212,n830);
and (n953,n934,n940);
xor (n954,n820,n834);
xor (n955,n797,n811);
and (n956,n931,n954);
and (n957,n882,n883);
xor (n958,n959,n968);
xor (n959,n960,n967);
or (n960,n961,n966);
and (n961,n962,n965);
xor (n962,n963,n964);
xor (n963,n707,n715);
xor (n964,n672,n685);
xor (n965,n723,n736);
and (n966,n963,n964);
xor (n967,n749,n752);
xor (n968,n791,n865);
or (n969,n970,n975);
and (n970,n971,n974);
xor (n971,n972,n973);
xor (n972,n794,n841);
xor (n973,n962,n965);
xor (n974,n881,n928);
and (n975,n972,n973);
or (n976,n977,n1087);
and (n977,n978,n1086);
xor (n978,n979,n1030);
or (n979,n980,n1029);
and (n980,n981,n1028);
xor (n981,n982,n983);
xor (n982,n843,n856);
or (n983,n984,n1027);
and (n984,n985,n1005);
xor (n985,n986,n992);
nand (n986,n987,n991);
or (n987,n428,n988);
nor (n988,n989,n990);
and (n989,n141,n246);
and (n990,n142,n245);
or (n991,n429,n836);
and (n992,n993,n999);
nor (n993,n994,n165);
nor (n994,n995,n998);
and (n995,n996,n137);
not (n996,n997);
and (n997,n89,n161);
and (n998,n88,n160);
nand (n999,n1000,n1001);
or (n1000,n27,n893);
or (n1001,n26,n1002);
nor (n1002,n1003,n1004);
and (n1003,n35,n119);
and (n1004,n29,n121);
or (n1005,n1006,n1026);
and (n1006,n1007,n1020);
xor (n1007,n1008,n1014);
nand (n1008,n1009,n1013);
or (n1009,n383,n1010);
nor (n1010,n1011,n1012);
and (n1011,n105,n395);
and (n1012,n106,n397);
or (n1013,n110,n900);
nand (n1014,n1015,n1019);
or (n1015,n129,n1016);
nor (n1016,n1017,n1018);
and (n1017,n137,n197);
and (n1018,n135,n199);
or (n1019,n138,n910);
nand (n1020,n1021,n1025);
or (n1021,n157,n1022);
nor (n1022,n1023,n1024);
and (n1023,n88,n166);
and (n1024,n165,n89);
or (n1025,n158,n916);
and (n1026,n1008,n1014);
and (n1027,n986,n992);
xor (n1028,n885,n905);
and (n1029,n982,n983);
or (n1030,n1031,n1085);
and (n1031,n1032,n1062);
xor (n1032,n1033,n1061);
or (n1033,n1034,n1060);
and (n1034,n1035,n1059);
xor (n1035,n1036,n1058);
or (n1036,n1037,n1057);
and (n1037,n1038,n1051);
xor (n1038,n1039,n1045);
nand (n1039,n1040,n1044);
or (n1040,n377,n1041);
nor (n1041,n1042,n1043);
and (n1042,n57,n225);
and (n1043,n58,n227);
or (n1044,n366,n922);
nand (n1045,n1046,n1050);
or (n1046,n251,n1047);
nor (n1047,n1048,n1049);
and (n1048,n214,n146);
and (n1049,n215,n148);
or (n1050,n252,n936);
nand (n1051,n1052,n1056);
or (n1052,n52,n1053);
nor (n1053,n1054,n1055);
and (n1054,n51,n422);
and (n1055,n48,n424);
or (n1056,n742,n942);
and (n1057,n1039,n1045);
xor (n1058,n933,n947);
xor (n1059,n889,n898);
and (n1060,n1036,n1058);
xor (n1061,n930,n955);
or (n1062,n1063,n1084);
and (n1063,n1064,n1083);
xor (n1064,n1065,n1066);
xor (n1065,n907,n920);
or (n1066,n1067,n1082);
and (n1067,n1068,n1081);
xor (n1068,n1069,n1075);
nand (n1069,n1070,n1074);
or (n1070,n202,n1071);
nor (n1071,n1072,n1073);
and (n1072,n206,n170);
and (n1073,n207,n172);
or (n1074,n212,n949);
nand (n1075,n1076,n1080);
or (n1076,n428,n1077);
nor (n1077,n1078,n1079);
and (n1078,n141,n298);
and (n1079,n142,n297);
or (n1080,n429,n988);
xor (n1081,n993,n999);
and (n1082,n1069,n1075);
xor (n1083,n985,n1005);
and (n1084,n1065,n1066);
and (n1085,n1033,n1061);
xor (n1086,n971,n974);
and (n1087,n979,n1030);
nor (n1088,n1089,n1090);
xor (n1089,n978,n1086);
or (n1090,n1091,n1172);
and (n1091,n1092,n1171);
xor (n1092,n1093,n1094);
xor (n1093,n981,n1028);
or (n1094,n1095,n1170);
and (n1095,n1096,n1169);
xor (n1096,n1097,n1162);
or (n1097,n1098,n1161);
and (n1098,n1099,n1139);
xor (n1099,n1100,n1117);
or (n1100,n1101,n1116);
and (n1101,n1102,n1110);
xor (n1102,n1103,n1104);
nor (n1103,n158,n88);
nand (n1104,n1105,n1109);
or (n1105,n26,n1106);
nor (n1106,n1107,n1108);
and (n1107,n35,n276);
and (n1108,n29,n278);
or (n1109,n1002,n27);
nand (n1110,n1111,n1115);
or (n1111,n377,n1112);
nor (n1112,n1113,n1114);
and (n1113,n57,n219);
and (n1114,n58,n221);
or (n1115,n366,n1041);
and (n1116,n1103,n1104);
or (n1117,n1118,n1138);
and (n1118,n1119,n1132);
xor (n1119,n1120,n1126);
nand (n1120,n1121,n1125);
or (n1121,n52,n1122);
nor (n1122,n1123,n1124);
and (n1123,n51,n444);
and (n1124,n48,n446);
or (n1125,n742,n1053);
nand (n1126,n1127,n1131);
or (n1127,n202,n1128);
nor (n1128,n1129,n1130);
and (n1129,n206,n246);
and (n1130,n207,n245);
or (n1131,n1071,n212);
nand (n1132,n1133,n1137);
or (n1133,n428,n1134);
nor (n1134,n1135,n1136);
and (n1135,n141,n323);
and (n1136,n142,n325);
or (n1137,n429,n1077);
and (n1138,n1120,n1126);
or (n1139,n1140,n1160);
and (n1140,n1141,n1154);
xor (n1141,n1142,n1148);
nand (n1142,n1143,n1147);
or (n1143,n129,n1144);
nor (n1144,n1145,n1146);
and (n1145,n137,n94);
and (n1146,n135,n96);
or (n1147,n1016,n138);
nand (n1148,n1149,n1153);
or (n1149,n383,n1150);
nor (n1150,n1151,n1152);
and (n1151,n105,n152);
and (n1152,n106,n154);
or (n1153,n110,n1010);
nand (n1154,n1155,n1159);
or (n1155,n251,n1156);
nor (n1156,n1157,n1158);
and (n1157,n214,n176);
and (n1158,n215,n178);
or (n1159,n252,n1047);
and (n1160,n1142,n1148);
and (n1161,n1100,n1117);
or (n1162,n1163,n1168);
and (n1163,n1164,n1167);
xor (n1164,n1165,n1166);
xor (n1165,n1007,n1020);
xor (n1166,n1038,n1051);
xor (n1167,n1068,n1081);
and (n1168,n1165,n1166);
xor (n1169,n1035,n1059);
and (n1170,n1097,n1162);
xor (n1171,n1032,n1062);
and (n1172,n1093,n1094);
nor (n1173,n1174,n1185);
nor (n1174,n1175,n1182);
xor (n1175,n1176,n1179);
xor (n1176,n1177,n1178);
xor (n1177,n701,n747);
xor (n1178,n786,n789);
or (n1179,n1180,n1181);
and (n1180,n959,n968);
and (n1181,n960,n967);
or (n1182,n1183,n1184);
and (n1183,n878,n969);
and (n1184,n879,n958);
nor (n1185,n1186,n1189);
or (n1186,n1187,n1188);
and (n1187,n1176,n1179);
and (n1188,n1177,n1178);
xor (n1189,n698,n868);
nand (n1190,n1191,n1504);
or (n1191,n1192,n1274);
not (n1192,n1193);
or (n1193,n1194,n1195);
xor (n1194,n1092,n1171);
or (n1195,n1196,n1273);
and (n1196,n1197,n1272);
xor (n1197,n1198,n1199);
xor (n1198,n1064,n1083);
or (n1199,n1200,n1271);
and (n1200,n1201,n1264);
xor (n1201,n1202,n1263);
or (n1202,n1203,n1262);
and (n1203,n1204,n1240);
xor (n1204,n1205,n1218);
and (n1205,n1206,n1212);
nor (n1206,n1207,n137);
nor (n1207,n1208,n1211);
and (n1208,n1209,n141);
not (n1209,n1210);
and (n1210,n89,n134);
and (n1211,n88,n133);
nand (n1212,n1213,n1217);
or (n1213,n26,n1214);
nor (n1214,n1215,n1216);
and (n1215,n35,n225);
and (n1216,n29,n227);
or (n1217,n1106,n27);
or (n1218,n1219,n1239);
and (n1219,n1220,n1233);
xor (n1220,n1221,n1227);
nand (n1221,n1222,n1226);
or (n1222,n377,n1223);
nor (n1223,n1224,n1225);
and (n1224,n57,n422);
and (n1225,n58,n424);
or (n1226,n366,n1112);
nand (n1227,n1228,n1232);
or (n1228,n129,n1229);
nor (n1229,n1230,n1231);
and (n1230,n88,n135);
and (n1231,n137,n89);
or (n1232,n138,n1144);
nand (n1233,n1234,n1238);
or (n1234,n383,n1235);
nor (n1235,n1236,n1237);
and (n1236,n105,n146);
and (n1237,n106,n148);
or (n1238,n110,n1150);
and (n1239,n1221,n1227);
or (n1240,n1241,n1261);
and (n1241,n1242,n1255);
xor (n1242,n1243,n1249);
nand (n1243,n1244,n1248);
or (n1244,n251,n1245);
nor (n1245,n1246,n1247);
and (n1246,n214,n170);
and (n1247,n215,n172);
or (n1248,n252,n1156);
nand (n1249,n1250,n1254);
or (n1250,n52,n1251);
nor (n1251,n1252,n1253);
and (n1252,n51,n395);
and (n1253,n48,n397);
or (n1254,n742,n1122);
nand (n1255,n1256,n1260);
or (n1256,n202,n1257);
nor (n1257,n1258,n1259);
and (n1258,n206,n298);
and (n1259,n207,n297);
or (n1260,n212,n1128);
and (n1261,n1243,n1249);
and (n1262,n1205,n1218);
xor (n1263,n1099,n1139);
or (n1264,n1265,n1270);
and (n1265,n1266,n1269);
xor (n1266,n1267,n1268);
xor (n1267,n1119,n1132);
xor (n1268,n1102,n1110);
xor (n1269,n1141,n1154);
and (n1270,n1267,n1268);
and (n1271,n1202,n1263);
xor (n1272,n1096,n1169);
and (n1273,n1198,n1199);
not (n1274,n1275);
nand (n1275,n1276,n1503);
or (n1276,n1277,n1350);
not (n1277,n1278);
nand (n1278,n1279,n1281);
not (n1279,n1280);
xor (n1280,n1197,n1272);
not (n1281,n1282);
or (n1282,n1283,n1349);
and (n1283,n1284,n1348);
xor (n1284,n1285,n1286);
xor (n1285,n1164,n1167);
or (n1286,n1287,n1347);
and (n1287,n1288,n1319);
xor (n1288,n1289,n1318);
or (n1289,n1290,n1317);
and (n1290,n1291,n1299);
xor (n1291,n1292,n1298);
nand (n1292,n1293,n1297);
or (n1293,n428,n1294);
nor (n1294,n1295,n1296);
and (n1295,n141,n197);
and (n1296,n142,n199);
or (n1297,n429,n1134);
xor (n1298,n1206,n1212);
or (n1299,n1300,n1316);
and (n1300,n1301,n1310);
xor (n1301,n1302,n1303);
nor (n1302,n138,n88);
nand (n1303,n1304,n1309);
or (n1304,n1305,n26);
not (n1305,n1306);
nor (n1306,n1307,n1308);
and (n1307,n219,n29);
and (n1308,n221,n35);
or (n1309,n1214,n27);
nand (n1310,n1311,n1315);
or (n1311,n377,n1312);
nor (n1312,n1313,n1314);
and (n1313,n57,n444);
and (n1314,n58,n446);
or (n1315,n366,n1223);
and (n1316,n1302,n1303);
and (n1317,n1292,n1298);
xor (n1318,n1204,n1240);
or (n1319,n1320,n1346);
and (n1320,n1321,n1345);
xor (n1321,n1322,n1344);
or (n1322,n1323,n1343);
and (n1323,n1324,n1337);
xor (n1324,n1325,n1331);
nand (n1325,n1326,n1330);
or (n1326,n383,n1327);
nor (n1327,n1328,n1329);
and (n1328,n105,n176);
and (n1329,n106,n178);
or (n1330,n110,n1235);
nand (n1331,n1332,n1336);
or (n1332,n251,n1333);
nor (n1333,n1334,n1335);
and (n1334,n214,n246);
and (n1335,n215,n245);
or (n1336,n252,n1245);
nand (n1337,n1338,n1342);
or (n1338,n52,n1339);
nor (n1339,n1340,n1341);
and (n1340,n51,n152);
and (n1341,n48,n154);
or (n1342,n742,n1251);
and (n1343,n1325,n1331);
xor (n1344,n1242,n1255);
xor (n1345,n1220,n1233);
and (n1346,n1322,n1344);
and (n1347,n1289,n1318);
xor (n1348,n1201,n1264);
and (n1349,n1285,n1286);
not (n1350,n1351);
nand (n1351,n1352,n1502);
or (n1352,n1353,n1444);
nor (n1353,n1354,n1355);
xor (n1354,n1284,n1348);
or (n1355,n1356,n1443);
and (n1356,n1357,n1442);
xor (n1357,n1358,n1359);
xor (n1358,n1266,n1269);
or (n1359,n1360,n1441);
and (n1360,n1361,n1392);
xor (n1361,n1362,n1391);
or (n1362,n1363,n1390);
and (n1363,n1364,n1377);
xor (n1364,n1365,n1371);
nand (n1365,n1366,n1370);
or (n1366,n202,n1367);
nor (n1367,n1368,n1369);
and (n1368,n206,n323);
and (n1369,n207,n325);
or (n1370,n212,n1257);
nand (n1371,n1372,n1376);
or (n1372,n428,n1373);
nor (n1373,n1374,n1375);
and (n1374,n141,n94);
and (n1375,n142,n96);
or (n1376,n429,n1294);
and (n1377,n1378,n1384);
nor (n1378,n1379,n141);
nor (n1379,n1380,n1383);
and (n1380,n1381,n206);
not (n1381,n1382);
and (n1382,n89,n432);
and (n1383,n88,n436);
nand (n1384,n1385,n1386);
or (n1385,n27,n1305);
or (n1386,n1387,n26);
nor (n1387,n1388,n1389);
and (n1388,n35,n422);
and (n1389,n29,n424);
and (n1390,n1365,n1371);
xor (n1391,n1291,n1299);
or (n1392,n1393,n1440);
and (n1393,n1394,n1439);
xor (n1394,n1395,n1417);
or (n1395,n1396,n1416);
and (n1396,n1397,n1410);
xor (n1397,n1398,n1404);
nand (n1398,n1399,n1403);
or (n1399,n377,n1400);
nor (n1400,n1401,n1402);
and (n1401,n57,n395);
and (n1402,n58,n397);
or (n1403,n366,n1312);
nand (n1404,n1405,n1409);
or (n1405,n383,n1406);
nor (n1406,n1407,n1408);
and (n1407,n105,n170);
and (n1408,n106,n172);
or (n1409,n110,n1327);
nand (n1410,n1411,n1415);
or (n1411,n251,n1412);
nor (n1412,n1413,n1414);
and (n1413,n214,n298);
and (n1414,n215,n297);
or (n1415,n252,n1333);
and (n1416,n1398,n1404);
or (n1417,n1418,n1438);
and (n1418,n1419,n1432);
xor (n1419,n1420,n1426);
nand (n1420,n1421,n1425);
or (n1421,n52,n1422);
nor (n1422,n1423,n1424);
and (n1423,n51,n146);
and (n1424,n48,n148);
or (n1425,n742,n1339);
nand (n1426,n1427,n1431);
or (n1427,n202,n1428);
nor (n1428,n1429,n1430);
and (n1429,n206,n197);
and (n1430,n207,n199);
or (n1431,n212,n1367);
nand (n1432,n1433,n1437);
or (n1433,n428,n1434);
nor (n1434,n1435,n1436);
and (n1435,n88,n142);
and (n1436,n141,n89);
or (n1437,n429,n1373);
and (n1438,n1420,n1426);
xor (n1439,n1301,n1310);
and (n1440,n1395,n1417);
and (n1441,n1362,n1391);
xor (n1442,n1288,n1319);
and (n1443,n1358,n1359);
nand (n1444,n1445,n1446);
xor (n1445,n1357,n1442);
or (n1446,n1447,n1501);
and (n1447,n1448,n1500);
xor (n1448,n1449,n1450);
xor (n1449,n1321,n1345);
or (n1450,n1451,n1499);
and (n1451,n1452,n1455);
xor (n1452,n1453,n1454);
xor (n1453,n1324,n1337);
xor (n1454,n1364,n1377);
or (n1455,n1456,n1498);
and (n1456,n1457,n1476);
xor (n1457,n1458,n1459);
xor (n1458,n1378,n1384);
or (n1459,n1460,n1475);
and (n1460,n1461,n1469);
xor (n1461,n1462,n1463);
nor (n1462,n429,n88);
nand (n1463,n1464,n1468);
or (n1464,n377,n1465);
nor (n1465,n1466,n1467);
and (n1466,n57,n152);
and (n1467,n58,n154);
or (n1468,n366,n1400);
nand (n1469,n1470,n1474);
or (n1470,n383,n1471);
nor (n1471,n1472,n1473);
and (n1472,n105,n246);
and (n1473,n106,n245);
or (n1474,n110,n1406);
and (n1475,n1462,n1463);
or (n1476,n1477,n1497);
and (n1477,n1478,n1491);
xor (n1478,n1479,n1485);
nand (n1479,n1480,n1484);
or (n1480,n251,n1481);
nor (n1481,n1482,n1483);
and (n1482,n214,n323);
and (n1483,n215,n325);
or (n1484,n252,n1412);
nand (n1485,n1486,n1490);
or (n1486,n26,n1487);
nor (n1487,n1488,n1489);
and (n1488,n35,n444);
and (n1489,n29,n446);
or (n1490,n1387,n27);
nand (n1491,n1492,n1496);
or (n1492,n202,n1493);
nor (n1493,n1494,n1495);
and (n1494,n206,n94);
and (n1495,n207,n96);
or (n1496,n212,n1428);
and (n1497,n1479,n1485);
and (n1498,n1458,n1459);
and (n1499,n1453,n1454);
xor (n1500,n1361,n1392);
and (n1501,n1449,n1450);
nand (n1502,n1354,n1355);
nand (n1503,n1280,n1282);
nand (n1504,n1194,n1195);
nand (n1505,n1506,n1513);
or (n1506,n1507,n1508);
not (n1507,n1173);
not (n1508,n1509);
nand (n1509,n1510,n1512);
or (n1510,n876,n1511);
nand (n1511,n1089,n1090);
nand (n1512,n877,n976);
nor (n1513,n1514,n1518);
and (n1514,n1515,n1517);
not (n1515,n1516);
nand (n1516,n1175,n1182);
not (n1517,n1185);
and (n1518,n1186,n1189);
nand (n1519,n874,n1520,n2035);
or (n1520,n1521,n2034);
and (n1521,n1522,n1584);
xor (n1522,n1523,n1583);
or (n1523,n1524,n1582);
and (n1524,n1525,n1528);
xor (n1525,n1526,n1527);
xor (n1526,n1394,n1439);
xor (n1527,n1452,n1455);
or (n1528,n1529,n1581);
and (n1529,n1530,n1533);
xor (n1530,n1531,n1532);
xor (n1531,n1419,n1432);
xor (n1532,n1397,n1410);
or (n1533,n1534,n1580);
and (n1534,n1535,n1558);
xor (n1535,n1536,n1542);
nand (n1536,n1537,n1541);
or (n1537,n52,n1538);
nor (n1538,n1539,n1540);
and (n1539,n51,n176);
and (n1540,n48,n178);
or (n1541,n742,n1422);
nor (n1542,n1543,n1552);
not (n1543,n1544);
nand (n1544,n1545,n1550);
or (n1545,n1546,n377);
not (n1546,n1547);
nand (n1547,n1548,n1549);
or (n1548,n58,n148);
or (n1549,n57,n146);
nand (n1550,n1551,n471);
not (n1551,n1465);
nand (n1552,n207,n1553);
nand (n1553,n1554,n1555);
or (n1554,n89,n208);
nand (n1555,n1556,n214);
not (n1556,n1557);
and (n1557,n89,n208);
or (n1558,n1559,n1579);
and (n1559,n1560,n1573);
xor (n1560,n1561,n1567);
nand (n1561,n1562,n1566);
or (n1562,n383,n1563);
nor (n1563,n1564,n1565);
and (n1564,n105,n298);
and (n1565,n106,n297);
or (n1566,n110,n1471);
nand (n1567,n1568,n1572);
or (n1568,n251,n1569);
nor (n1569,n1570,n1571);
and (n1570,n214,n197);
and (n1571,n215,n199);
or (n1572,n252,n1481);
nand (n1573,n1574,n1578);
or (n1574,n26,n1575);
nor (n1575,n1576,n1577);
and (n1576,n35,n395);
and (n1577,n29,n397);
or (n1578,n1487,n27);
and (n1579,n1561,n1567);
and (n1580,n1536,n1542);
and (n1581,n1531,n1532);
and (n1582,n1526,n1527);
xor (n1583,n1448,n1500);
or (n1584,n1585,n2033);
and (n1585,n1586,n1620);
xor (n1586,n1587,n1619);
or (n1587,n1588,n1618);
and (n1588,n1589,n1617);
xor (n1589,n1590,n1591);
xor (n1590,n1457,n1476);
or (n1591,n1592,n1616);
and (n1592,n1593,n1596);
xor (n1593,n1594,n1595);
xor (n1594,n1478,n1491);
xor (n1595,n1461,n1469);
or (n1596,n1597,n1615);
and (n1597,n1598,n1611);
xor (n1598,n1599,n1605);
nand (n1599,n1600,n1604);
or (n1600,n1601,n202);
nor (n1601,n1602,n1603);
and (n1602,n88,n207);
and (n1603,n206,n89);
or (n1604,n212,n1493);
nand (n1605,n1606,n1610);
or (n1606,n52,n1607);
nor (n1607,n1608,n1609);
and (n1608,n51,n170);
and (n1609,n48,n172);
or (n1610,n742,n1538);
nand (n1611,n1612,n1614);
or (n1612,n1613,n1543);
not (n1613,n1552);
nand (n1614,n1613,n1543);
and (n1615,n1599,n1605);
and (n1616,n1594,n1595);
xor (n1617,n1530,n1533);
and (n1618,n1590,n1591);
xor (n1619,n1525,n1528);
nand (n1620,n1621,n2027);
or (n1621,n1622,n1732);
not (n1622,n1623);
nor (n1623,n1624,n1682);
nor (n1624,n1625,n1626);
xor (n1625,n1589,n1617);
or (n1626,n1627,n1681);
and (n1627,n1628,n1680);
xor (n1628,n1629,n1630);
xor (n1629,n1535,n1558);
or (n1630,n1631,n1679);
and (n1631,n1632,n1678);
xor (n1632,n1633,n1653);
or (n1633,n1634,n1652);
and (n1634,n1635,n1644);
xor (n1635,n1636,n1637);
nor (n1636,n212,n88);
nand (n1637,n1638,n1643);
or (n1638,n1639,n377);
not (n1639,n1640);
nand (n1640,n1641,n1642);
or (n1641,n58,n178);
or (n1642,n57,n176);
nand (n1643,n471,n1547);
nand (n1644,n1645,n1650);
or (n1645,n1646,n383);
not (n1646,n1647);
nor (n1647,n1648,n1649);
and (n1648,n325,n105);
and (n1649,n323,n106);
nand (n1650,n1651,n111);
not (n1651,n1563);
and (n1652,n1636,n1637);
or (n1653,n1654,n1677);
and (n1654,n1655,n1671);
xor (n1655,n1656,n1665);
nand (n1656,n1657,n1662);
or (n1657,n1658,n251);
not (n1658,n1659);
nand (n1659,n1660,n1661);
or (n1660,n215,n96);
or (n1661,n214,n94);
nand (n1662,n1663,n1664);
not (n1663,n1569);
not (n1664,n252);
nand (n1665,n1666,n1670);
or (n1666,n26,n1667);
nor (n1667,n1668,n1669);
and (n1668,n35,n152);
and (n1669,n29,n154);
or (n1670,n1575,n27);
nand (n1671,n1672,n1676);
or (n1672,n52,n1673);
nor (n1673,n1674,n1675);
and (n1674,n51,n246);
and (n1675,n48,n245);
or (n1676,n742,n1607);
and (n1677,n1656,n1665);
xor (n1678,n1560,n1573);
and (n1679,n1633,n1653);
xor (n1680,n1593,n1596);
and (n1681,n1629,n1630);
nor (n1682,n1683,n1684);
xor (n1683,n1628,n1680);
or (n1684,n1685,n1731);
and (n1685,n1686,n1689);
xor (n1686,n1687,n1688);
xor (n1687,n1598,n1611);
xor (n1688,n1632,n1678);
or (n1689,n1690,n1730);
and (n1690,n1691,n1729);
xor (n1691,n1692,n1706);
and (n1692,n1693,n1699);
and (n1693,n1694,n215);
nand (n1694,n1695,n1696);
or (n1695,n89,n255);
nand (n1696,n1697,n105);
not (n1697,n1698);
and (n1698,n89,n255);
nand (n1699,n1700,n1705);
or (n1700,n1701,n377);
not (n1701,n1702);
nand (n1702,n1703,n1704);
or (n1703,n58,n172);
or (n1704,n57,n170);
nand (n1705,n471,n1640);
or (n1706,n1707,n1728);
and (n1707,n1708,n1722);
xor (n1708,n1709,n1715);
nand (n1709,n1710,n1714);
or (n1710,n1711,n383);
nor (n1711,n1712,n1713);
and (n1712,n105,n197);
and (n1713,n106,n199);
nand (n1714,n111,n1647);
nand (n1715,n1716,n1721);
or (n1716,n1717,n251);
not (n1717,n1718);
nand (n1718,n1719,n1720);
or (n1719,n89,n214);
or (n1720,n88,n215);
nand (n1721,n1664,n1659);
nand (n1722,n1723,n1727);
or (n1723,n26,n1724);
nor (n1724,n1725,n1726);
and (n1725,n35,n146);
and (n1726,n29,n148);
or (n1727,n1667,n27);
and (n1728,n1709,n1715);
xor (n1729,n1635,n1644);
and (n1730,n1692,n1706);
and (n1731,n1687,n1688);
not (n1732,n1733);
or (n1733,n1734,n2026);
and (n1734,n1735,n1772);
xor (n1735,n1736,n1771);
or (n1736,n1737,n1770);
and (n1737,n1738,n1769);
xor (n1738,n1739,n1740);
xor (n1739,n1655,n1671);
or (n1740,n1741,n1768);
and (n1741,n1742,n1750);
xor (n1742,n1743,n1749);
nand (n1743,n1744,n1748);
or (n1744,n52,n1745);
nor (n1745,n1746,n1747);
and (n1746,n51,n298);
and (n1747,n48,n297);
or (n1748,n742,n1673);
xor (n1749,n1693,n1699);
or (n1750,n1751,n1767);
and (n1751,n1752,n1762);
xor (n1752,n1753,n1754);
and (n1753,n1664,n89);
nand (n1754,n1755,n1756);
or (n1755,n1724,n27);
nand (n1756,n1757,n1761);
not (n1757,n1758);
nor (n1758,n1759,n1760);
and (n1759,n35,n176);
and (n1760,n29,n178);
not (n1761,n26);
nand (n1762,n1763,n1766);
or (n1763,n383,n1764);
not (n1764,n1765);
xor (n1765,n96,n105);
or (n1766,n110,n1711);
and (n1767,n1753,n1754);
and (n1768,n1743,n1749);
xor (n1769,n1691,n1729);
and (n1770,n1739,n1740);
xor (n1771,n1686,n1689);
or (n1772,n1773,n2025);
and (n1773,n1774,n1814);
xor (n1774,n1775,n1813);
or (n1775,n1776,n1812);
and (n1776,n1777,n1811);
xor (n1777,n1778,n1779);
xor (n1778,n1708,n1722);
or (n1779,n1780,n1810);
and (n1780,n1781,n1797);
xor (n1781,n1782,n1789);
nand (n1782,n1783,n1788);
or (n1783,n1784,n377);
not (n1784,n1785);
nor (n1785,n1786,n1787);
and (n1786,n246,n58);
and (n1787,n245,n57);
nand (n1788,n471,n1702);
nand (n1789,n1790,n1795);
or (n1790,n1791,n52);
not (n1791,n1792);
nand (n1792,n1793,n1794);
or (n1793,n48,n325);
or (n1794,n51,n323);
nand (n1795,n1796,n54);
not (n1796,n1745);
and (n1797,n1798,n1804);
nor (n1798,n1799,n105);
nor (n1799,n1800,n1803);
and (n1800,n1801,n51);
not (n1801,n1802);
and (n1802,n89,n113);
and (n1803,n88,n126);
nand (n1804,n1805,n1809);
or (n1805,n26,n1806);
nor (n1806,n1807,n1808);
and (n1807,n35,n170);
and (n1808,n29,n172);
or (n1809,n1758,n27);
and (n1810,n1782,n1789);
xor (n1811,n1742,n1750);
and (n1812,n1778,n1779);
xor (n1813,n1738,n1769);
nand (n1814,n1815,n2022,n2024);
nand (n1815,n1816,n1851,n2015);
nand (n1816,n1817,n1819);
not (n1817,n1818);
xor (n1818,n1777,n1811);
not (n1819,n1820);
or (n1820,n1821,n1850);
and (n1821,n1822,n1849);
xor (n1822,n1823,n1848);
or (n1823,n1824,n1847);
and (n1824,n1825,n1840);
xor (n1825,n1826,n1833);
nand (n1826,n1827,n1832);
or (n1827,n1828,n383);
not (n1828,n1829);
nand (n1829,n1830,n1831);
or (n1830,n105,n89);
or (n1831,n88,n106);
nand (n1832,n111,n1765);
nand (n1833,n1834,n1839);
or (n1834,n1835,n377);
not (n1835,n1836);
nor (n1836,n1837,n1838);
and (n1837,n297,n57);
and (n1838,n298,n58);
nand (n1839,n471,n1785);
nand (n1840,n1841,n1846);
or (n1841,n1842,n52);
not (n1842,n1843);
nand (n1843,n1844,n1845);
or (n1844,n48,n199);
or (n1845,n51,n197);
nand (n1846,n54,n1792);
and (n1847,n1826,n1833);
xor (n1848,n1752,n1762);
xor (n1849,n1781,n1797);
and (n1850,n1823,n1848);
nand (n1851,n1852,n2014);
or (n1852,n1853,n1907);
not (n1853,n1854);
nand (n1854,n1855,n1880);
not (n1855,n1856);
xor (n1856,n1857,n1879);
xor (n1857,n1858,n1859);
xor (n1858,n1798,n1804);
or (n1859,n1860,n1878);
and (n1860,n1861,n1871);
xor (n1861,n1862,n1863);
and (n1862,n111,n89);
nand (n1863,n1864,n1869);
or (n1864,n26,n1865);
not (n1865,n1866);
nor (n1866,n1867,n1868);
and (n1867,n246,n29);
and (n1868,n245,n35);
nand (n1869,n1870,n28);
not (n1870,n1806);
nand (n1871,n1872,n1877);
or (n1872,n1873,n377);
not (n1873,n1874);
nor (n1874,n1875,n1876);
and (n1875,n325,n57);
and (n1876,n323,n58);
nand (n1877,n471,n1836);
and (n1878,n1862,n1863);
xor (n1879,n1825,n1840);
not (n1880,n1881);
or (n1881,n1882,n1906);
and (n1882,n1883,n1905);
xor (n1883,n1884,n1891);
nand (n1884,n1885,n1890);
or (n1885,n1886,n52);
not (n1886,n1887);
nor (n1887,n1888,n1889);
and (n1888,n96,n51);
and (n1889,n94,n48);
nand (n1890,n54,n1843);
and (n1891,n1892,n1898);
and (n1892,n1893,n48);
nand (n1893,n1894,n1895);
or (n1894,n89,n56);
nand (n1895,n1896,n57);
not (n1896,n1897);
and (n1897,n89,n56);
nand (n1898,n1899,n1900);
or (n1899,n27,n1865);
nand (n1900,n1901,n1761);
not (n1901,n1902);
nor (n1902,n1903,n1904);
and (n1903,n35,n298);
and (n1904,n29,n297);
xor (n1905,n1861,n1871);
and (n1906,n1884,n1891);
not (n1907,n1908);
nand (n1908,n1909,n2013);
or (n1909,n1910,n1934);
not (n1910,n1911);
nand (n1911,n1912,n1914);
not (n1912,n1913);
xor (n1913,n1883,n1905);
not (n1914,n1915);
or (n1915,n1916,n1933);
and (n1916,n1917,n1932);
xor (n1917,n1918,n1925);
nand (n1918,n1919,n1924);
or (n1919,n1920,n377);
not (n1920,n1921);
nor (n1921,n1922,n1923);
and (n1922,n199,n57);
and (n1923,n197,n58);
nand (n1924,n471,n1874);
nand (n1925,n1926,n1931);
or (n1926,n1927,n52);
not (n1927,n1928);
nand (n1928,n1929,n1930);
or (n1929,n89,n51);
or (n1930,n48,n88);
nand (n1931,n54,n1887);
xor (n1932,n1892,n1898);
and (n1933,n1918,n1925);
not (n1934,n1935);
nand (n1935,n1936,n2012);
or (n1936,n1937,n2007);
nor (n1937,n1938,n2006);
and (n1938,n1939,n1972);
nand (n1939,n1940,n1958);
not (n1940,n1941);
xor (n1941,n1942,n1951);
xor (n1942,n1943,n1944);
and (n1943,n54,n89);
nand (n1944,n1945,n1950);
or (n1945,n1946,n377);
not (n1946,n1947);
nor (n1947,n1948,n1949);
and (n1948,n96,n57);
and (n1949,n94,n58);
nand (n1950,n471,n1921);
nand (n1951,n1952,n1957);
or (n1952,n1953,n26);
not (n1953,n1954);
nand (n1954,n1955,n1956);
or (n1955,n323,n35);
nand (n1956,n35,n323);
or (n1957,n1902,n27);
nand (n1958,n1959,n1966);
nand (n1959,n1960,n1965);
or (n1960,n26,n1961);
not (n1961,n1962);
nand (n1962,n1963,n1964);
or (n1963,n197,n35);
nand (n1964,n35,n197);
nand (n1965,n1954,n28);
not (n1966,n1967);
nand (n1967,n1968,n58);
nand (n1968,n1969,n1970);
or (n1969,n89,n369);
or (n1970,n1971,n29);
and (n1971,n89,n369);
or (n1972,n1973,n2005);
and (n1973,n1974,n1984);
xor (n1974,n1975,n1981);
nand (n1975,n1976,n1977);
or (n1976,n1946,n366);
or (n1977,n377,n1978);
nor (n1978,n1979,n1980);
and (n1979,n58,n88);
and (n1980,n89,n57);
nand (n1981,n1982,n1983);
or (n1982,n1967,n1959);
nand (n1983,n1959,n1967);
nand (n1984,n1985,n2004);
or (n1985,n1986,n1994);
nor (n1986,n1987,n1993);
nand (n1987,n1988,n1989);
or (n1988,n27,n1961);
nand (n1989,n1990,n1761);
nor (n1990,n1991,n1992);
and (n1991,n96,n35);
and (n1992,n94,n29);
and (n1993,n471,n89);
nand (n1994,n1995,n2002);
nand (n1995,n1996,n1998);
or (n1996,n27,n1997);
not (n1997,n1990);
nand (n1998,n1999,n1761);
nand (n1999,n2000,n2001);
or (n2000,n35,n89);
or (n2001,n29,n88);
nor (n2002,n2003,n35);
and (n2003,n89,n28);
nand (n2004,n1987,n1993);
and (n2005,n1975,n1981);
nor (n2006,n1940,n1958);
nor (n2007,n2008,n2009);
xor (n2008,n1917,n1932);
or (n2009,n2010,n2011);
and (n2010,n1942,n1951);
and (n2011,n1943,n1944);
nand (n2012,n2008,n2009);
nand (n2013,n1913,n1915);
nand (n2014,n1881,n1856);
nand (n2015,n2016,n2018);
not (n2016,n2017);
xor (n2017,n1822,n1849);
not (n2018,n2019);
or (n2019,n2020,n2021);
and (n2020,n1857,n1879);
and (n2021,n1858,n1859);
nand (n2022,n1816,n2023);
nor (n2023,n2016,n2018);
nand (n2024,n1818,n1820);
and (n2025,n1775,n1813);
and (n2026,n1736,n1771);
nor (n2027,n2028,n2032);
and (n2028,n2029,n2030);
not (n2029,n1624);
not (n2030,n2031);
nand (n2031,n1683,n1684);
and (n2032,n1625,n1626);
and (n2033,n1587,n1619);
and (n2034,n1523,n1583);
and (n2035,n2036,n1193,n1278);
nor (n2036,n1353,n2037);
nor (n2037,n1445,n1446);
or (n2038,n2039,n3674);
and (n2039,n2040,n3673);
wire s0n2040,s1n2040,notn2040;
or (n2040,s0n2040,s1n2040);
not(notn2040,n7);
and (s0n2040,notn2040,n8);
and (s1n2040,n7,n2041);
xor (n2041,n2042,n3672);
xor (n2042,n2043,n3669);
xor (n2043,n2044,n3668);
xor (n2044,n2045,n3660);
xor (n2045,n2046,n3659);
xor (n2046,n2047,n3644);
xor (n2047,n2048,n3643);
xor (n2048,n2049,n3623);
xor (n2049,n2050,n3622);
xor (n2050,n2051,n3596);
xor (n2051,n2052,n3595);
xor (n2052,n2053,n3563);
xor (n2053,n2054,n3562);
xor (n2054,n2055,n3523);
xor (n2055,n2056,n3522);
xor (n2056,n2057,n3478);
xor (n2057,n2058,n3477);
xor (n2058,n2059,n3426);
xor (n2059,n2060,n3425);
xor (n2060,n2061,n3369);
xor (n2061,n2062,n3368);
xor (n2062,n2063,n3305);
xor (n2063,n2064,n3304);
xor (n2064,n2065,n3236);
xor (n2065,n2066,n3235);
xor (n2066,n2067,n3160);
xor (n2067,n2068,n3159);
xor (n2068,n2069,n3079);
xor (n2069,n2070,n3078);
xor (n2070,n2071,n2991);
xor (n2071,n2072,n2990);
xor (n2072,n2073,n2898);
xor (n2073,n2074,n2897);
xor (n2074,n2075,n2800);
xor (n2075,n2076,n2799);
xor (n2076,n2077,n2695);
xor (n2077,n2078,n2694);
xor (n2078,n2079,n2585);
xor (n2079,n2080,n2584);
xor (n2080,n2081,n2468);
xor (n2081,n2082,n2467);
xor (n2082,n2083,n2349);
xor (n2083,n2084,n2348);
xor (n2084,n2085,n2220);
xor (n2085,n2086,n2219);
xor (n2086,n2087,n2090);
xor (n2087,n2088,n2089);
and (n2088,n348,n28);
and (n2089,n40,n29);
or (n2090,n2091,n2094);
and (n2091,n2092,n2093);
and (n2092,n40,n28);
and (n2093,n33,n29);
and (n2094,n2095,n2096);
xor (n2095,n2092,n2093);
or (n2096,n2097,n2100);
and (n2097,n2098,n2099);
and (n2098,n33,n28);
and (n2099,n374,n29);
and (n2100,n2101,n2102);
xor (n2101,n2098,n2099);
or (n2102,n2103,n2105);
and (n2103,n2104,n489);
and (n2104,n374,n28);
and (n2105,n2106,n2107);
xor (n2106,n2104,n489);
or (n2107,n2108,n2111);
and (n2108,n2109,n2110);
and (n2109,n189,n28);
and (n2110,n68,n29);
and (n2111,n2112,n2113);
xor (n2112,n2109,n2110);
or (n2113,n2114,n2116);
and (n2114,n2115,n778);
and (n2115,n68,n28);
and (n2116,n2117,n2118);
xor (n2117,n2115,n778);
or (n2118,n2119,n2121);
and (n2119,n2120,n895);
and (n2120,n47,n28);
and (n2121,n2122,n2123);
xor (n2122,n2120,n895);
or (n2123,n2124,n2127);
and (n2124,n2125,n2126);
and (n2125,n107,n28);
and (n2126,n119,n29);
and (n2127,n2128,n2129);
xor (n2128,n2125,n2126);
or (n2129,n2130,n2133);
and (n2130,n2131,n2132);
and (n2131,n119,n28);
and (n2132,n276,n29);
and (n2133,n2134,n2135);
xor (n2134,n2131,n2132);
or (n2135,n2136,n2139);
and (n2136,n2137,n2138);
and (n2137,n276,n28);
and (n2138,n225,n29);
and (n2139,n2140,n2141);
xor (n2140,n2137,n2138);
or (n2141,n2142,n2144);
and (n2142,n2143,n1307);
and (n2143,n225,n28);
and (n2144,n2145,n2146);
xor (n2145,n2143,n1307);
or (n2146,n2147,n2150);
and (n2147,n2148,n2149);
and (n2148,n219,n28);
and (n2149,n422,n29);
and (n2150,n2151,n2152);
xor (n2151,n2148,n2149);
or (n2152,n2153,n2156);
and (n2153,n2154,n2155);
and (n2154,n422,n28);
and (n2155,n444,n29);
and (n2156,n2157,n2158);
xor (n2157,n2154,n2155);
or (n2158,n2159,n2162);
and (n2159,n2160,n2161);
and (n2160,n444,n28);
and (n2161,n395,n29);
and (n2162,n2163,n2164);
xor (n2163,n2160,n2161);
or (n2164,n2165,n2168);
and (n2165,n2166,n2167);
and (n2166,n395,n28);
and (n2167,n152,n29);
and (n2168,n2169,n2170);
xor (n2169,n2166,n2167);
or (n2170,n2171,n2174);
and (n2171,n2172,n2173);
and (n2172,n152,n28);
and (n2173,n146,n29);
and (n2174,n2175,n2176);
xor (n2175,n2172,n2173);
or (n2176,n2177,n2180);
and (n2177,n2178,n2179);
and (n2178,n146,n28);
and (n2179,n176,n29);
and (n2180,n2181,n2182);
xor (n2181,n2178,n2179);
or (n2182,n2183,n2186);
and (n2183,n2184,n2185);
and (n2184,n176,n28);
and (n2185,n170,n29);
and (n2186,n2187,n2188);
xor (n2187,n2184,n2185);
or (n2188,n2189,n2191);
and (n2189,n2190,n1867);
and (n2190,n170,n28);
and (n2191,n2192,n2193);
xor (n2192,n2190,n1867);
or (n2193,n2194,n2197);
and (n2194,n2195,n2196);
and (n2195,n246,n28);
and (n2196,n298,n29);
and (n2197,n2198,n2199);
xor (n2198,n2195,n2196);
or (n2199,n2200,n2203);
and (n2200,n2201,n2202);
and (n2201,n298,n28);
and (n2202,n323,n29);
and (n2203,n2204,n2205);
xor (n2204,n2201,n2202);
or (n2205,n2206,n2209);
and (n2206,n2207,n2208);
and (n2207,n323,n28);
and (n2208,n197,n29);
and (n2209,n2210,n2211);
xor (n2210,n2207,n2208);
or (n2211,n2212,n2214);
and (n2212,n2213,n1992);
and (n2213,n197,n28);
and (n2214,n2215,n2216);
xor (n2215,n2213,n1992);
and (n2216,n2217,n2218);
and (n2217,n94,n28);
and (n2218,n89,n29);
and (n2219,n33,n369);
or (n2220,n2221,n2224);
and (n2221,n2222,n2223);
xor (n2222,n2095,n2096);
and (n2223,n374,n369);
and (n2224,n2225,n2226);
xor (n2225,n2222,n2223);
or (n2226,n2227,n2230);
and (n2227,n2228,n2229);
xor (n2228,n2101,n2102);
and (n2229,n189,n369);
and (n2230,n2231,n2232);
xor (n2231,n2228,n2229);
or (n2232,n2233,n2236);
and (n2233,n2234,n2235);
xor (n2234,n2106,n2107);
and (n2235,n68,n369);
and (n2236,n2237,n2238);
xor (n2237,n2234,n2235);
or (n2238,n2239,n2242);
and (n2239,n2240,n2241);
xor (n2240,n2112,n2113);
and (n2241,n47,n369);
and (n2242,n2243,n2244);
xor (n2243,n2240,n2241);
or (n2244,n2245,n2248);
and (n2245,n2246,n2247);
xor (n2246,n2117,n2118);
and (n2247,n107,n369);
and (n2248,n2249,n2250);
xor (n2249,n2246,n2247);
or (n2250,n2251,n2254);
and (n2251,n2252,n2253);
xor (n2252,n2122,n2123);
and (n2253,n119,n369);
and (n2254,n2255,n2256);
xor (n2255,n2252,n2253);
or (n2256,n2257,n2260);
and (n2257,n2258,n2259);
xor (n2258,n2128,n2129);
and (n2259,n276,n369);
and (n2260,n2261,n2262);
xor (n2261,n2258,n2259);
or (n2262,n2263,n2266);
and (n2263,n2264,n2265);
xor (n2264,n2134,n2135);
and (n2265,n225,n369);
and (n2266,n2267,n2268);
xor (n2267,n2264,n2265);
or (n2268,n2269,n2272);
and (n2269,n2270,n2271);
xor (n2270,n2140,n2141);
and (n2271,n219,n369);
and (n2272,n2273,n2274);
xor (n2273,n2270,n2271);
or (n2274,n2275,n2278);
and (n2275,n2276,n2277);
xor (n2276,n2145,n2146);
and (n2277,n422,n369);
and (n2278,n2279,n2280);
xor (n2279,n2276,n2277);
or (n2280,n2281,n2284);
and (n2281,n2282,n2283);
xor (n2282,n2151,n2152);
and (n2283,n444,n369);
and (n2284,n2285,n2286);
xor (n2285,n2282,n2283);
or (n2286,n2287,n2290);
and (n2287,n2288,n2289);
xor (n2288,n2157,n2158);
and (n2289,n395,n369);
and (n2290,n2291,n2292);
xor (n2291,n2288,n2289);
or (n2292,n2293,n2296);
and (n2293,n2294,n2295);
xor (n2294,n2163,n2164);
and (n2295,n152,n369);
and (n2296,n2297,n2298);
xor (n2297,n2294,n2295);
or (n2298,n2299,n2302);
and (n2299,n2300,n2301);
xor (n2300,n2169,n2170);
and (n2301,n146,n369);
and (n2302,n2303,n2304);
xor (n2303,n2300,n2301);
or (n2304,n2305,n2308);
and (n2305,n2306,n2307);
xor (n2306,n2175,n2176);
and (n2307,n176,n369);
and (n2308,n2309,n2310);
xor (n2309,n2306,n2307);
or (n2310,n2311,n2314);
and (n2311,n2312,n2313);
xor (n2312,n2181,n2182);
and (n2313,n170,n369);
and (n2314,n2315,n2316);
xor (n2315,n2312,n2313);
or (n2316,n2317,n2320);
and (n2317,n2318,n2319);
xor (n2318,n2187,n2188);
and (n2319,n246,n369);
and (n2320,n2321,n2322);
xor (n2321,n2318,n2319);
or (n2322,n2323,n2326);
and (n2323,n2324,n2325);
xor (n2324,n2192,n2193);
and (n2325,n298,n369);
and (n2326,n2327,n2328);
xor (n2327,n2324,n2325);
or (n2328,n2329,n2332);
and (n2329,n2330,n2331);
xor (n2330,n2198,n2199);
and (n2331,n323,n369);
and (n2332,n2333,n2334);
xor (n2333,n2330,n2331);
or (n2334,n2335,n2338);
and (n2335,n2336,n2337);
xor (n2336,n2204,n2205);
and (n2337,n197,n369);
and (n2338,n2339,n2340);
xor (n2339,n2336,n2337);
or (n2340,n2341,n2344);
and (n2341,n2342,n2343);
xor (n2342,n2210,n2211);
and (n2343,n94,n369);
and (n2344,n2345,n2346);
xor (n2345,n2342,n2343);
and (n2346,n2347,n1971);
xor (n2347,n2215,n2216);
and (n2348,n374,n58);
or (n2349,n2350,n2353);
and (n2350,n2351,n2352);
xor (n2351,n2225,n2226);
and (n2352,n189,n58);
and (n2353,n2354,n2355);
xor (n2354,n2351,n2352);
or (n2355,n2356,n2359);
and (n2356,n2357,n2358);
xor (n2357,n2231,n2232);
and (n2358,n68,n58);
and (n2359,n2360,n2361);
xor (n2360,n2357,n2358);
or (n2361,n2362,n2365);
and (n2362,n2363,n2364);
xor (n2363,n2237,n2238);
and (n2364,n47,n58);
and (n2365,n2366,n2367);
xor (n2366,n2363,n2364);
or (n2367,n2368,n2371);
and (n2368,n2369,n2370);
xor (n2369,n2243,n2244);
and (n2370,n107,n58);
and (n2371,n2372,n2373);
xor (n2372,n2369,n2370);
or (n2373,n2374,n2377);
and (n2374,n2375,n2376);
xor (n2375,n2249,n2250);
and (n2376,n119,n58);
and (n2377,n2378,n2379);
xor (n2378,n2375,n2376);
or (n2379,n2380,n2383);
and (n2380,n2381,n2382);
xor (n2381,n2255,n2256);
and (n2382,n276,n58);
and (n2383,n2384,n2385);
xor (n2384,n2381,n2382);
or (n2385,n2386,n2389);
and (n2386,n2387,n2388);
xor (n2387,n2261,n2262);
and (n2388,n225,n58);
and (n2389,n2390,n2391);
xor (n2390,n2387,n2388);
or (n2391,n2392,n2395);
and (n2392,n2393,n2394);
xor (n2393,n2267,n2268);
and (n2394,n219,n58);
and (n2395,n2396,n2397);
xor (n2396,n2393,n2394);
or (n2397,n2398,n2401);
and (n2398,n2399,n2400);
xor (n2399,n2273,n2274);
and (n2400,n422,n58);
and (n2401,n2402,n2403);
xor (n2402,n2399,n2400);
or (n2403,n2404,n2407);
and (n2404,n2405,n2406);
xor (n2405,n2279,n2280);
and (n2406,n444,n58);
and (n2407,n2408,n2409);
xor (n2408,n2405,n2406);
or (n2409,n2410,n2413);
and (n2410,n2411,n2412);
xor (n2411,n2285,n2286);
and (n2412,n395,n58);
and (n2413,n2414,n2415);
xor (n2414,n2411,n2412);
or (n2415,n2416,n2419);
and (n2416,n2417,n2418);
xor (n2417,n2291,n2292);
and (n2418,n152,n58);
and (n2419,n2420,n2421);
xor (n2420,n2417,n2418);
or (n2421,n2422,n2425);
and (n2422,n2423,n2424);
xor (n2423,n2297,n2298);
and (n2424,n146,n58);
and (n2425,n2426,n2427);
xor (n2426,n2423,n2424);
or (n2427,n2428,n2431);
and (n2428,n2429,n2430);
xor (n2429,n2303,n2304);
and (n2430,n176,n58);
and (n2431,n2432,n2433);
xor (n2432,n2429,n2430);
or (n2433,n2434,n2437);
and (n2434,n2435,n2436);
xor (n2435,n2309,n2310);
and (n2436,n170,n58);
and (n2437,n2438,n2439);
xor (n2438,n2435,n2436);
or (n2439,n2440,n2442);
and (n2440,n2441,n1786);
xor (n2441,n2315,n2316);
and (n2442,n2443,n2444);
xor (n2443,n2441,n1786);
or (n2444,n2445,n2447);
and (n2445,n2446,n1838);
xor (n2446,n2321,n2322);
and (n2447,n2448,n2449);
xor (n2448,n2446,n1838);
or (n2449,n2450,n2452);
and (n2450,n2451,n1876);
xor (n2451,n2327,n2328);
and (n2452,n2453,n2454);
xor (n2453,n2451,n1876);
or (n2454,n2455,n2457);
and (n2455,n2456,n1923);
xor (n2456,n2333,n2334);
and (n2457,n2458,n2459);
xor (n2458,n2456,n1923);
or (n2459,n2460,n2462);
and (n2460,n2461,n1949);
xor (n2461,n2339,n2340);
and (n2462,n2463,n2464);
xor (n2463,n2461,n1949);
and (n2464,n2465,n2466);
xor (n2465,n2345,n2346);
and (n2466,n89,n58);
and (n2467,n189,n56);
or (n2468,n2469,n2472);
and (n2469,n2470,n2471);
xor (n2470,n2354,n2355);
and (n2471,n68,n56);
and (n2472,n2473,n2474);
xor (n2473,n2470,n2471);
or (n2474,n2475,n2478);
and (n2475,n2476,n2477);
xor (n2476,n2360,n2361);
and (n2477,n47,n56);
and (n2478,n2479,n2480);
xor (n2479,n2476,n2477);
or (n2480,n2481,n2484);
and (n2481,n2482,n2483);
xor (n2482,n2366,n2367);
and (n2483,n107,n56);
and (n2484,n2485,n2486);
xor (n2485,n2482,n2483);
or (n2486,n2487,n2490);
and (n2487,n2488,n2489);
xor (n2488,n2372,n2373);
and (n2489,n119,n56);
and (n2490,n2491,n2492);
xor (n2491,n2488,n2489);
or (n2492,n2493,n2496);
and (n2493,n2494,n2495);
xor (n2494,n2378,n2379);
and (n2495,n276,n56);
and (n2496,n2497,n2498);
xor (n2497,n2494,n2495);
or (n2498,n2499,n2502);
and (n2499,n2500,n2501);
xor (n2500,n2384,n2385);
and (n2501,n225,n56);
and (n2502,n2503,n2504);
xor (n2503,n2500,n2501);
or (n2504,n2505,n2508);
and (n2505,n2506,n2507);
xor (n2506,n2390,n2391);
and (n2507,n219,n56);
and (n2508,n2509,n2510);
xor (n2509,n2506,n2507);
or (n2510,n2511,n2514);
and (n2511,n2512,n2513);
xor (n2512,n2396,n2397);
and (n2513,n422,n56);
and (n2514,n2515,n2516);
xor (n2515,n2512,n2513);
or (n2516,n2517,n2520);
and (n2517,n2518,n2519);
xor (n2518,n2402,n2403);
and (n2519,n444,n56);
and (n2520,n2521,n2522);
xor (n2521,n2518,n2519);
or (n2522,n2523,n2526);
and (n2523,n2524,n2525);
xor (n2524,n2408,n2409);
and (n2525,n395,n56);
and (n2526,n2527,n2528);
xor (n2527,n2524,n2525);
or (n2528,n2529,n2532);
and (n2529,n2530,n2531);
xor (n2530,n2414,n2415);
and (n2531,n152,n56);
and (n2532,n2533,n2534);
xor (n2533,n2530,n2531);
or (n2534,n2535,n2538);
and (n2535,n2536,n2537);
xor (n2536,n2420,n2421);
and (n2537,n146,n56);
and (n2538,n2539,n2540);
xor (n2539,n2536,n2537);
or (n2540,n2541,n2544);
and (n2541,n2542,n2543);
xor (n2542,n2426,n2427);
and (n2543,n176,n56);
and (n2544,n2545,n2546);
xor (n2545,n2542,n2543);
or (n2546,n2547,n2550);
and (n2547,n2548,n2549);
xor (n2548,n2432,n2433);
and (n2549,n170,n56);
and (n2550,n2551,n2552);
xor (n2551,n2548,n2549);
or (n2552,n2553,n2556);
and (n2553,n2554,n2555);
xor (n2554,n2438,n2439);
and (n2555,n246,n56);
and (n2556,n2557,n2558);
xor (n2557,n2554,n2555);
or (n2558,n2559,n2562);
and (n2559,n2560,n2561);
xor (n2560,n2443,n2444);
and (n2561,n298,n56);
and (n2562,n2563,n2564);
xor (n2563,n2560,n2561);
or (n2564,n2565,n2568);
and (n2565,n2566,n2567);
xor (n2566,n2448,n2449);
and (n2567,n323,n56);
and (n2568,n2569,n2570);
xor (n2569,n2566,n2567);
or (n2570,n2571,n2574);
and (n2571,n2572,n2573);
xor (n2572,n2453,n2454);
and (n2573,n197,n56);
and (n2574,n2575,n2576);
xor (n2575,n2572,n2573);
or (n2576,n2577,n2580);
and (n2577,n2578,n2579);
xor (n2578,n2458,n2459);
and (n2579,n94,n56);
and (n2580,n2581,n2582);
xor (n2581,n2578,n2579);
and (n2582,n2583,n1897);
xor (n2583,n2463,n2464);
and (n2584,n68,n48);
or (n2585,n2586,n2588);
and (n2586,n2587,n46);
xor (n2587,n2473,n2474);
and (n2588,n2589,n2590);
xor (n2589,n2587,n46);
or (n2590,n2591,n2594);
and (n2591,n2592,n2593);
xor (n2592,n2479,n2480);
and (n2593,n107,n48);
and (n2594,n2595,n2596);
xor (n2595,n2592,n2593);
or (n2596,n2597,n2600);
and (n2597,n2598,n2599);
xor (n2598,n2485,n2486);
and (n2599,n119,n48);
and (n2600,n2601,n2602);
xor (n2601,n2598,n2599);
or (n2602,n2603,n2606);
and (n2603,n2604,n2605);
xor (n2604,n2491,n2492);
and (n2605,n276,n48);
and (n2606,n2607,n2608);
xor (n2607,n2604,n2605);
or (n2608,n2609,n2612);
and (n2609,n2610,n2611);
xor (n2610,n2497,n2498);
and (n2611,n225,n48);
and (n2612,n2613,n2614);
xor (n2613,n2610,n2611);
or (n2614,n2615,n2618);
and (n2615,n2616,n2617);
xor (n2616,n2503,n2504);
and (n2617,n219,n48);
and (n2618,n2619,n2620);
xor (n2619,n2616,n2617);
or (n2620,n2621,n2624);
and (n2621,n2622,n2623);
xor (n2622,n2509,n2510);
and (n2623,n422,n48);
and (n2624,n2625,n2626);
xor (n2625,n2622,n2623);
or (n2626,n2627,n2630);
and (n2627,n2628,n2629);
xor (n2628,n2515,n2516);
and (n2629,n444,n48);
and (n2630,n2631,n2632);
xor (n2631,n2628,n2629);
or (n2632,n2633,n2636);
and (n2633,n2634,n2635);
xor (n2634,n2521,n2522);
and (n2635,n395,n48);
and (n2636,n2637,n2638);
xor (n2637,n2634,n2635);
or (n2638,n2639,n2642);
and (n2639,n2640,n2641);
xor (n2640,n2527,n2528);
and (n2641,n152,n48);
and (n2642,n2643,n2644);
xor (n2643,n2640,n2641);
or (n2644,n2645,n2648);
and (n2645,n2646,n2647);
xor (n2646,n2533,n2534);
and (n2647,n146,n48);
and (n2648,n2649,n2650);
xor (n2649,n2646,n2647);
or (n2650,n2651,n2654);
and (n2651,n2652,n2653);
xor (n2652,n2539,n2540);
and (n2653,n176,n48);
and (n2654,n2655,n2656);
xor (n2655,n2652,n2653);
or (n2656,n2657,n2660);
and (n2657,n2658,n2659);
xor (n2658,n2545,n2546);
and (n2659,n170,n48);
and (n2660,n2661,n2662);
xor (n2661,n2658,n2659);
or (n2662,n2663,n2666);
and (n2663,n2664,n2665);
xor (n2664,n2551,n2552);
and (n2665,n246,n48);
and (n2666,n2667,n2668);
xor (n2667,n2664,n2665);
or (n2668,n2669,n2672);
and (n2669,n2670,n2671);
xor (n2670,n2557,n2558);
and (n2671,n298,n48);
and (n2672,n2673,n2674);
xor (n2673,n2670,n2671);
or (n2674,n2675,n2678);
and (n2675,n2676,n2677);
xor (n2676,n2563,n2564);
and (n2677,n323,n48);
and (n2678,n2679,n2680);
xor (n2679,n2676,n2677);
or (n2680,n2681,n2684);
and (n2681,n2682,n2683);
xor (n2682,n2569,n2570);
and (n2683,n197,n48);
and (n2684,n2685,n2686);
xor (n2685,n2682,n2683);
or (n2686,n2687,n2689);
and (n2687,n2688,n1889);
xor (n2688,n2575,n2576);
and (n2689,n2690,n2691);
xor (n2690,n2688,n1889);
and (n2691,n2692,n2693);
xor (n2692,n2581,n2582);
and (n2693,n89,n48);
and (n2694,n47,n113);
or (n2695,n2696,n2699);
and (n2696,n2697,n2698);
xor (n2697,n2589,n2590);
and (n2698,n107,n113);
and (n2699,n2700,n2701);
xor (n2700,n2697,n2698);
or (n2701,n2702,n2705);
and (n2702,n2703,n2704);
xor (n2703,n2595,n2596);
and (n2704,n119,n113);
and (n2705,n2706,n2707);
xor (n2706,n2703,n2704);
or (n2707,n2708,n2711);
and (n2708,n2709,n2710);
xor (n2709,n2601,n2602);
and (n2710,n276,n113);
and (n2711,n2712,n2713);
xor (n2712,n2709,n2710);
or (n2713,n2714,n2717);
and (n2714,n2715,n2716);
xor (n2715,n2607,n2608);
and (n2716,n225,n113);
and (n2717,n2718,n2719);
xor (n2718,n2715,n2716);
or (n2719,n2720,n2723);
and (n2720,n2721,n2722);
xor (n2721,n2613,n2614);
and (n2722,n219,n113);
and (n2723,n2724,n2725);
xor (n2724,n2721,n2722);
or (n2725,n2726,n2729);
and (n2726,n2727,n2728);
xor (n2727,n2619,n2620);
and (n2728,n422,n113);
and (n2729,n2730,n2731);
xor (n2730,n2727,n2728);
or (n2731,n2732,n2735);
and (n2732,n2733,n2734);
xor (n2733,n2625,n2626);
and (n2734,n444,n113);
and (n2735,n2736,n2737);
xor (n2736,n2733,n2734);
or (n2737,n2738,n2741);
and (n2738,n2739,n2740);
xor (n2739,n2631,n2632);
and (n2740,n395,n113);
and (n2741,n2742,n2743);
xor (n2742,n2739,n2740);
or (n2743,n2744,n2747);
and (n2744,n2745,n2746);
xor (n2745,n2637,n2638);
and (n2746,n152,n113);
and (n2747,n2748,n2749);
xor (n2748,n2745,n2746);
or (n2749,n2750,n2753);
and (n2750,n2751,n2752);
xor (n2751,n2643,n2644);
and (n2752,n146,n113);
and (n2753,n2754,n2755);
xor (n2754,n2751,n2752);
or (n2755,n2756,n2759);
and (n2756,n2757,n2758);
xor (n2757,n2649,n2650);
and (n2758,n176,n113);
and (n2759,n2760,n2761);
xor (n2760,n2757,n2758);
or (n2761,n2762,n2765);
and (n2762,n2763,n2764);
xor (n2763,n2655,n2656);
and (n2764,n170,n113);
and (n2765,n2766,n2767);
xor (n2766,n2763,n2764);
or (n2767,n2768,n2771);
and (n2768,n2769,n2770);
xor (n2769,n2661,n2662);
and (n2770,n246,n113);
and (n2771,n2772,n2773);
xor (n2772,n2769,n2770);
or (n2773,n2774,n2777);
and (n2774,n2775,n2776);
xor (n2775,n2667,n2668);
and (n2776,n298,n113);
and (n2777,n2778,n2779);
xor (n2778,n2775,n2776);
or (n2779,n2780,n2783);
and (n2780,n2781,n2782);
xor (n2781,n2673,n2674);
and (n2782,n323,n113);
and (n2783,n2784,n2785);
xor (n2784,n2781,n2782);
or (n2785,n2786,n2789);
and (n2786,n2787,n2788);
xor (n2787,n2679,n2680);
and (n2788,n197,n113);
and (n2789,n2790,n2791);
xor (n2790,n2787,n2788);
or (n2791,n2792,n2795);
and (n2792,n2793,n2794);
xor (n2793,n2685,n2686);
and (n2794,n94,n113);
and (n2795,n2796,n2797);
xor (n2796,n2793,n2794);
and (n2797,n2798,n1802);
xor (n2798,n2690,n2691);
and (n2799,n107,n106);
or (n2800,n2801,n2804);
and (n2801,n2802,n2803);
xor (n2802,n2700,n2701);
and (n2803,n119,n106);
and (n2804,n2805,n2806);
xor (n2805,n2802,n2803);
or (n2806,n2807,n2810);
and (n2807,n2808,n2809);
xor (n2808,n2706,n2707);
and (n2809,n276,n106);
and (n2810,n2811,n2812);
xor (n2811,n2808,n2809);
or (n2812,n2813,n2816);
and (n2813,n2814,n2815);
xor (n2814,n2712,n2713);
and (n2815,n225,n106);
and (n2816,n2817,n2818);
xor (n2817,n2814,n2815);
or (n2818,n2819,n2822);
and (n2819,n2820,n2821);
xor (n2820,n2718,n2719);
and (n2821,n219,n106);
and (n2822,n2823,n2824);
xor (n2823,n2820,n2821);
or (n2824,n2825,n2827);
and (n2825,n2826,n802);
xor (n2826,n2724,n2725);
and (n2827,n2828,n2829);
xor (n2828,n2826,n802);
or (n2829,n2830,n2833);
and (n2830,n2831,n2832);
xor (n2831,n2730,n2731);
and (n2832,n444,n106);
and (n2833,n2834,n2835);
xor (n2834,n2831,n2832);
or (n2835,n2836,n2839);
and (n2836,n2837,n2838);
xor (n2837,n2736,n2737);
and (n2838,n395,n106);
and (n2839,n2840,n2841);
xor (n2840,n2837,n2838);
or (n2841,n2842,n2845);
and (n2842,n2843,n2844);
xor (n2843,n2742,n2743);
and (n2844,n152,n106);
and (n2845,n2846,n2847);
xor (n2846,n2843,n2844);
or (n2847,n2848,n2851);
and (n2848,n2849,n2850);
xor (n2849,n2748,n2749);
and (n2850,n146,n106);
and (n2851,n2852,n2853);
xor (n2852,n2849,n2850);
or (n2853,n2854,n2857);
and (n2854,n2855,n2856);
xor (n2855,n2754,n2755);
and (n2856,n176,n106);
and (n2857,n2858,n2859);
xor (n2858,n2855,n2856);
or (n2859,n2860,n2863);
and (n2860,n2861,n2862);
xor (n2861,n2760,n2761);
and (n2862,n170,n106);
and (n2863,n2864,n2865);
xor (n2864,n2861,n2862);
or (n2865,n2866,n2869);
and (n2866,n2867,n2868);
xor (n2867,n2766,n2767);
and (n2868,n246,n106);
and (n2869,n2870,n2871);
xor (n2870,n2867,n2868);
or (n2871,n2872,n2875);
and (n2872,n2873,n2874);
xor (n2873,n2772,n2773);
and (n2874,n298,n106);
and (n2875,n2876,n2877);
xor (n2876,n2873,n2874);
or (n2877,n2878,n2880);
and (n2878,n2879,n1649);
xor (n2879,n2778,n2779);
and (n2880,n2881,n2882);
xor (n2881,n2879,n1649);
or (n2882,n2883,n2886);
and (n2883,n2884,n2885);
xor (n2884,n2784,n2785);
and (n2885,n197,n106);
and (n2886,n2887,n2888);
xor (n2887,n2884,n2885);
or (n2888,n2889,n2892);
and (n2889,n2890,n2891);
xor (n2890,n2790,n2791);
and (n2891,n94,n106);
and (n2892,n2893,n2894);
xor (n2893,n2890,n2891);
and (n2894,n2895,n2896);
xor (n2895,n2796,n2797);
and (n2896,n89,n106);
and (n2897,n119,n255);
or (n2898,n2899,n2902);
and (n2899,n2900,n2901);
xor (n2900,n2805,n2806);
and (n2901,n276,n255);
and (n2902,n2903,n2904);
xor (n2903,n2900,n2901);
or (n2904,n2905,n2908);
and (n2905,n2906,n2907);
xor (n2906,n2811,n2812);
and (n2907,n225,n255);
and (n2908,n2909,n2910);
xor (n2909,n2906,n2907);
or (n2910,n2911,n2914);
and (n2911,n2912,n2913);
xor (n2912,n2817,n2818);
and (n2913,n219,n255);
and (n2914,n2915,n2916);
xor (n2915,n2912,n2913);
or (n2916,n2917,n2920);
and (n2917,n2918,n2919);
xor (n2918,n2823,n2824);
and (n2919,n422,n255);
and (n2920,n2921,n2922);
xor (n2921,n2918,n2919);
or (n2922,n2923,n2926);
and (n2923,n2924,n2925);
xor (n2924,n2828,n2829);
and (n2925,n444,n255);
and (n2926,n2927,n2928);
xor (n2927,n2924,n2925);
or (n2928,n2929,n2932);
and (n2929,n2930,n2931);
xor (n2930,n2834,n2835);
and (n2931,n395,n255);
and (n2932,n2933,n2934);
xor (n2933,n2930,n2931);
or (n2934,n2935,n2938);
and (n2935,n2936,n2937);
xor (n2936,n2840,n2841);
and (n2937,n152,n255);
and (n2938,n2939,n2940);
xor (n2939,n2936,n2937);
or (n2940,n2941,n2944);
and (n2941,n2942,n2943);
xor (n2942,n2846,n2847);
and (n2943,n146,n255);
and (n2944,n2945,n2946);
xor (n2945,n2942,n2943);
or (n2946,n2947,n2950);
and (n2947,n2948,n2949);
xor (n2948,n2852,n2853);
and (n2949,n176,n255);
and (n2950,n2951,n2952);
xor (n2951,n2948,n2949);
or (n2952,n2953,n2956);
and (n2953,n2954,n2955);
xor (n2954,n2858,n2859);
and (n2955,n170,n255);
and (n2956,n2957,n2958);
xor (n2957,n2954,n2955);
or (n2958,n2959,n2962);
and (n2959,n2960,n2961);
xor (n2960,n2864,n2865);
and (n2961,n246,n255);
and (n2962,n2963,n2964);
xor (n2963,n2960,n2961);
or (n2964,n2965,n2968);
and (n2965,n2966,n2967);
xor (n2966,n2870,n2871);
and (n2967,n298,n255);
and (n2968,n2969,n2970);
xor (n2969,n2966,n2967);
or (n2970,n2971,n2974);
and (n2971,n2972,n2973);
xor (n2972,n2876,n2877);
and (n2973,n323,n255);
and (n2974,n2975,n2976);
xor (n2975,n2972,n2973);
or (n2976,n2977,n2980);
and (n2977,n2978,n2979);
xor (n2978,n2881,n2882);
and (n2979,n197,n255);
and (n2980,n2981,n2982);
xor (n2981,n2978,n2979);
or (n2982,n2983,n2986);
and (n2983,n2984,n2985);
xor (n2984,n2887,n2888);
and (n2985,n94,n255);
and (n2986,n2987,n2988);
xor (n2987,n2984,n2985);
and (n2988,n2989,n1698);
xor (n2989,n2893,n2894);
and (n2990,n276,n215);
or (n2991,n2992,n2995);
and (n2992,n2993,n2994);
xor (n2993,n2903,n2904);
and (n2994,n225,n215);
and (n2995,n2996,n2997);
xor (n2996,n2993,n2994);
or (n2997,n2998,n3001);
and (n2998,n2999,n3000);
xor (n2999,n2909,n2910);
and (n3000,n219,n215);
and (n3001,n3002,n3003);
xor (n3002,n2999,n3000);
or (n3003,n3004,n3007);
and (n3004,n3005,n3006);
xor (n3005,n2915,n2916);
and (n3006,n422,n215);
and (n3007,n3008,n3009);
xor (n3008,n3005,n3006);
or (n3009,n3010,n3013);
and (n3010,n3011,n3012);
xor (n3011,n2921,n2922);
and (n3012,n444,n215);
and (n3013,n3014,n3015);
xor (n3014,n3011,n3012);
or (n3015,n3016,n3019);
and (n3016,n3017,n3018);
xor (n3017,n2927,n2928);
and (n3018,n395,n215);
and (n3019,n3020,n3021);
xor (n3020,n3017,n3018);
or (n3021,n3022,n3025);
and (n3022,n3023,n3024);
xor (n3023,n2933,n2934);
and (n3024,n152,n215);
and (n3025,n3026,n3027);
xor (n3026,n3023,n3024);
or (n3027,n3028,n3031);
and (n3028,n3029,n3030);
xor (n3029,n2939,n2940);
and (n3030,n146,n215);
and (n3031,n3032,n3033);
xor (n3032,n3029,n3030);
or (n3033,n3034,n3037);
and (n3034,n3035,n3036);
xor (n3035,n2945,n2946);
and (n3036,n176,n215);
and (n3037,n3038,n3039);
xor (n3038,n3035,n3036);
or (n3039,n3040,n3043);
and (n3040,n3041,n3042);
xor (n3041,n2951,n2952);
and (n3042,n170,n215);
and (n3043,n3044,n3045);
xor (n3044,n3041,n3042);
or (n3045,n3046,n3049);
and (n3046,n3047,n3048);
xor (n3047,n2957,n2958);
and (n3048,n246,n215);
and (n3049,n3050,n3051);
xor (n3050,n3047,n3048);
or (n3051,n3052,n3055);
and (n3052,n3053,n3054);
xor (n3053,n2963,n2964);
and (n3054,n298,n215);
and (n3055,n3056,n3057);
xor (n3056,n3053,n3054);
or (n3057,n3058,n3061);
and (n3058,n3059,n3060);
xor (n3059,n2969,n2970);
and (n3060,n323,n215);
and (n3061,n3062,n3063);
xor (n3062,n3059,n3060);
or (n3063,n3064,n3067);
and (n3064,n3065,n3066);
xor (n3065,n2975,n2976);
and (n3066,n197,n215);
and (n3067,n3068,n3069);
xor (n3068,n3065,n3066);
or (n3069,n3070,n3073);
and (n3070,n3071,n3072);
xor (n3071,n2981,n2982);
and (n3072,n94,n215);
and (n3073,n3074,n3075);
xor (n3074,n3071,n3072);
and (n3075,n3076,n3077);
xor (n3076,n2987,n2988);
and (n3077,n89,n215);
and (n3078,n225,n208);
or (n3079,n3080,n3083);
and (n3080,n3081,n3082);
xor (n3081,n2996,n2997);
and (n3082,n219,n208);
and (n3083,n3084,n3085);
xor (n3084,n3081,n3082);
or (n3085,n3086,n3089);
and (n3086,n3087,n3088);
xor (n3087,n3002,n3003);
and (n3088,n422,n208);
and (n3089,n3090,n3091);
xor (n3090,n3087,n3088);
or (n3091,n3092,n3095);
and (n3092,n3093,n3094);
xor (n3093,n3008,n3009);
and (n3094,n444,n208);
and (n3095,n3096,n3097);
xor (n3096,n3093,n3094);
or (n3097,n3098,n3101);
and (n3098,n3099,n3100);
xor (n3099,n3014,n3015);
and (n3100,n395,n208);
and (n3101,n3102,n3103);
xor (n3102,n3099,n3100);
or (n3103,n3104,n3107);
and (n3104,n3105,n3106);
xor (n3105,n3020,n3021);
and (n3106,n152,n208);
and (n3107,n3108,n3109);
xor (n3108,n3105,n3106);
or (n3109,n3110,n3113);
and (n3110,n3111,n3112);
xor (n3111,n3026,n3027);
and (n3112,n146,n208);
and (n3113,n3114,n3115);
xor (n3114,n3111,n3112);
or (n3115,n3116,n3119);
and (n3116,n3117,n3118);
xor (n3117,n3032,n3033);
and (n3118,n176,n208);
and (n3119,n3120,n3121);
xor (n3120,n3117,n3118);
or (n3121,n3122,n3125);
and (n3122,n3123,n3124);
xor (n3123,n3038,n3039);
and (n3124,n170,n208);
and (n3125,n3126,n3127);
xor (n3126,n3123,n3124);
or (n3127,n3128,n3131);
and (n3128,n3129,n3130);
xor (n3129,n3044,n3045);
and (n3130,n246,n208);
and (n3131,n3132,n3133);
xor (n3132,n3129,n3130);
or (n3133,n3134,n3137);
and (n3134,n3135,n3136);
xor (n3135,n3050,n3051);
and (n3136,n298,n208);
and (n3137,n3138,n3139);
xor (n3138,n3135,n3136);
or (n3139,n3140,n3143);
and (n3140,n3141,n3142);
xor (n3141,n3056,n3057);
and (n3142,n323,n208);
and (n3143,n3144,n3145);
xor (n3144,n3141,n3142);
or (n3145,n3146,n3149);
and (n3146,n3147,n3148);
xor (n3147,n3062,n3063);
and (n3148,n197,n208);
and (n3149,n3150,n3151);
xor (n3150,n3147,n3148);
or (n3151,n3152,n3155);
and (n3152,n3153,n3154);
xor (n3153,n3068,n3069);
and (n3154,n94,n208);
and (n3155,n3156,n3157);
xor (n3156,n3153,n3154);
and (n3157,n3158,n1557);
xor (n3158,n3074,n3075);
and (n3159,n219,n207);
or (n3160,n3161,n3164);
and (n3161,n3162,n3163);
xor (n3162,n3084,n3085);
and (n3163,n422,n207);
and (n3164,n3165,n3166);
xor (n3165,n3162,n3163);
or (n3166,n3167,n3170);
and (n3167,n3168,n3169);
xor (n3168,n3090,n3091);
and (n3169,n444,n207);
and (n3170,n3171,n3172);
xor (n3171,n3168,n3169);
or (n3172,n3173,n3176);
and (n3173,n3174,n3175);
xor (n3174,n3096,n3097);
and (n3175,n395,n207);
and (n3176,n3177,n3178);
xor (n3177,n3174,n3175);
or (n3178,n3179,n3182);
and (n3179,n3180,n3181);
xor (n3180,n3102,n3103);
and (n3181,n152,n207);
and (n3182,n3183,n3184);
xor (n3183,n3180,n3181);
or (n3184,n3185,n3188);
and (n3185,n3186,n3187);
xor (n3186,n3108,n3109);
and (n3187,n146,n207);
and (n3188,n3189,n3190);
xor (n3189,n3186,n3187);
or (n3190,n3191,n3194);
and (n3191,n3192,n3193);
xor (n3192,n3114,n3115);
and (n3193,n176,n207);
and (n3194,n3195,n3196);
xor (n3195,n3192,n3193);
or (n3196,n3197,n3200);
and (n3197,n3198,n3199);
xor (n3198,n3120,n3121);
and (n3199,n170,n207);
and (n3200,n3201,n3202);
xor (n3201,n3198,n3199);
or (n3202,n3203,n3206);
and (n3203,n3204,n3205);
xor (n3204,n3126,n3127);
and (n3205,n246,n207);
and (n3206,n3207,n3208);
xor (n3207,n3204,n3205);
or (n3208,n3209,n3212);
and (n3209,n3210,n3211);
xor (n3210,n3132,n3133);
and (n3211,n298,n207);
and (n3212,n3213,n3214);
xor (n3213,n3210,n3211);
or (n3214,n3215,n3218);
and (n3215,n3216,n3217);
xor (n3216,n3138,n3139);
and (n3217,n323,n207);
and (n3218,n3219,n3220);
xor (n3219,n3216,n3217);
or (n3220,n3221,n3224);
and (n3221,n3222,n3223);
xor (n3222,n3144,n3145);
and (n3223,n197,n207);
and (n3224,n3225,n3226);
xor (n3225,n3222,n3223);
or (n3226,n3227,n3230);
and (n3227,n3228,n3229);
xor (n3228,n3150,n3151);
and (n3229,n94,n207);
and (n3230,n3231,n3232);
xor (n3231,n3228,n3229);
and (n3232,n3233,n3234);
xor (n3233,n3156,n3157);
and (n3234,n89,n207);
and (n3235,n422,n432);
or (n3236,n3237,n3240);
and (n3237,n3238,n3239);
xor (n3238,n3165,n3166);
and (n3239,n444,n432);
and (n3240,n3241,n3242);
xor (n3241,n3238,n3239);
or (n3242,n3243,n3246);
and (n3243,n3244,n3245);
xor (n3244,n3171,n3172);
and (n3245,n395,n432);
and (n3246,n3247,n3248);
xor (n3247,n3244,n3245);
or (n3248,n3249,n3252);
and (n3249,n3250,n3251);
xor (n3250,n3177,n3178);
and (n3251,n152,n432);
and (n3252,n3253,n3254);
xor (n3253,n3250,n3251);
or (n3254,n3255,n3258);
and (n3255,n3256,n3257);
xor (n3256,n3183,n3184);
and (n3257,n146,n432);
and (n3258,n3259,n3260);
xor (n3259,n3256,n3257);
or (n3260,n3261,n3264);
and (n3261,n3262,n3263);
xor (n3262,n3189,n3190);
and (n3263,n176,n432);
and (n3264,n3265,n3266);
xor (n3265,n3262,n3263);
or (n3266,n3267,n3270);
and (n3267,n3268,n3269);
xor (n3268,n3195,n3196);
and (n3269,n170,n432);
and (n3270,n3271,n3272);
xor (n3271,n3268,n3269);
or (n3272,n3273,n3276);
and (n3273,n3274,n3275);
xor (n3274,n3201,n3202);
and (n3275,n246,n432);
and (n3276,n3277,n3278);
xor (n3277,n3274,n3275);
or (n3278,n3279,n3282);
and (n3279,n3280,n3281);
xor (n3280,n3207,n3208);
and (n3281,n298,n432);
and (n3282,n3283,n3284);
xor (n3283,n3280,n3281);
or (n3284,n3285,n3288);
and (n3285,n3286,n3287);
xor (n3286,n3213,n3214);
and (n3287,n323,n432);
and (n3288,n3289,n3290);
xor (n3289,n3286,n3287);
or (n3290,n3291,n3294);
and (n3291,n3292,n3293);
xor (n3292,n3219,n3220);
and (n3293,n197,n432);
and (n3294,n3295,n3296);
xor (n3295,n3292,n3293);
or (n3296,n3297,n3300);
and (n3297,n3298,n3299);
xor (n3298,n3225,n3226);
and (n3299,n94,n432);
and (n3300,n3301,n3302);
xor (n3301,n3298,n3299);
and (n3302,n3303,n1382);
xor (n3303,n3231,n3232);
and (n3304,n444,n142);
or (n3305,n3306,n3309);
and (n3306,n3307,n3308);
xor (n3307,n3241,n3242);
and (n3308,n395,n142);
and (n3309,n3310,n3311);
xor (n3310,n3307,n3308);
or (n3311,n3312,n3315);
and (n3312,n3313,n3314);
xor (n3313,n3247,n3248);
and (n3314,n152,n142);
and (n3315,n3316,n3317);
xor (n3316,n3313,n3314);
or (n3317,n3318,n3321);
and (n3318,n3319,n3320);
xor (n3319,n3253,n3254);
and (n3320,n146,n142);
and (n3321,n3322,n3323);
xor (n3322,n3319,n3320);
or (n3323,n3324,n3327);
and (n3324,n3325,n3326);
xor (n3325,n3259,n3260);
and (n3326,n176,n142);
and (n3327,n3328,n3329);
xor (n3328,n3325,n3326);
or (n3329,n3330,n3333);
and (n3330,n3331,n3332);
xor (n3331,n3265,n3266);
and (n3332,n170,n142);
and (n3333,n3334,n3335);
xor (n3334,n3331,n3332);
or (n3335,n3336,n3339);
and (n3336,n3337,n3338);
xor (n3337,n3271,n3272);
and (n3338,n246,n142);
and (n3339,n3340,n3341);
xor (n3340,n3337,n3338);
or (n3341,n3342,n3345);
and (n3342,n3343,n3344);
xor (n3343,n3277,n3278);
and (n3344,n298,n142);
and (n3345,n3346,n3347);
xor (n3346,n3343,n3344);
or (n3347,n3348,n3351);
and (n3348,n3349,n3350);
xor (n3349,n3283,n3284);
and (n3350,n323,n142);
and (n3351,n3352,n3353);
xor (n3352,n3349,n3350);
or (n3353,n3354,n3357);
and (n3354,n3355,n3356);
xor (n3355,n3289,n3290);
and (n3356,n197,n142);
and (n3357,n3358,n3359);
xor (n3358,n3355,n3356);
or (n3359,n3360,n3363);
and (n3360,n3361,n3362);
xor (n3361,n3295,n3296);
and (n3362,n94,n142);
and (n3363,n3364,n3365);
xor (n3364,n3361,n3362);
and (n3365,n3366,n3367);
xor (n3366,n3301,n3302);
and (n3367,n89,n142);
and (n3368,n395,n134);
or (n3369,n3370,n3373);
and (n3370,n3371,n3372);
xor (n3371,n3310,n3311);
and (n3372,n152,n134);
and (n3373,n3374,n3375);
xor (n3374,n3371,n3372);
or (n3375,n3376,n3379);
and (n3376,n3377,n3378);
xor (n3377,n3316,n3317);
and (n3378,n146,n134);
and (n3379,n3380,n3381);
xor (n3380,n3377,n3378);
or (n3381,n3382,n3385);
and (n3382,n3383,n3384);
xor (n3383,n3322,n3323);
and (n3384,n176,n134);
and (n3385,n3386,n3387);
xor (n3386,n3383,n3384);
or (n3387,n3388,n3391);
and (n3388,n3389,n3390);
xor (n3389,n3328,n3329);
and (n3390,n170,n134);
and (n3391,n3392,n3393);
xor (n3392,n3389,n3390);
or (n3393,n3394,n3397);
and (n3394,n3395,n3396);
xor (n3395,n3334,n3335);
and (n3396,n246,n134);
and (n3397,n3398,n3399);
xor (n3398,n3395,n3396);
or (n3399,n3400,n3403);
and (n3400,n3401,n3402);
xor (n3401,n3340,n3341);
and (n3402,n298,n134);
and (n3403,n3404,n3405);
xor (n3404,n3401,n3402);
or (n3405,n3406,n3409);
and (n3406,n3407,n3408);
xor (n3407,n3346,n3347);
and (n3408,n323,n134);
and (n3409,n3410,n3411);
xor (n3410,n3407,n3408);
or (n3411,n3412,n3415);
and (n3412,n3413,n3414);
xor (n3413,n3352,n3353);
and (n3414,n197,n134);
and (n3415,n3416,n3417);
xor (n3416,n3413,n3414);
or (n3417,n3418,n3421);
and (n3418,n3419,n3420);
xor (n3419,n3358,n3359);
and (n3420,n94,n134);
and (n3421,n3422,n3423);
xor (n3422,n3419,n3420);
and (n3423,n3424,n1210);
xor (n3424,n3364,n3365);
and (n3425,n152,n135);
or (n3426,n3427,n3430);
and (n3427,n3428,n3429);
xor (n3428,n3374,n3375);
and (n3429,n146,n135);
and (n3430,n3431,n3432);
xor (n3431,n3428,n3429);
or (n3432,n3433,n3436);
and (n3433,n3434,n3435);
xor (n3434,n3380,n3381);
and (n3435,n176,n135);
and (n3436,n3437,n3438);
xor (n3437,n3434,n3435);
or (n3438,n3439,n3442);
and (n3439,n3440,n3441);
xor (n3440,n3386,n3387);
and (n3441,n170,n135);
and (n3442,n3443,n3444);
xor (n3443,n3440,n3441);
or (n3444,n3445,n3448);
and (n3445,n3446,n3447);
xor (n3446,n3392,n3393);
and (n3447,n246,n135);
and (n3448,n3449,n3450);
xor (n3449,n3446,n3447);
or (n3450,n3451,n3454);
and (n3451,n3452,n3453);
xor (n3452,n3398,n3399);
and (n3453,n298,n135);
and (n3454,n3455,n3456);
xor (n3455,n3452,n3453);
or (n3456,n3457,n3460);
and (n3457,n3458,n3459);
xor (n3458,n3404,n3405);
and (n3459,n323,n135);
and (n3460,n3461,n3462);
xor (n3461,n3458,n3459);
or (n3462,n3463,n3466);
and (n3463,n3464,n3465);
xor (n3464,n3410,n3411);
and (n3465,n197,n135);
and (n3466,n3467,n3468);
xor (n3467,n3464,n3465);
or (n3468,n3469,n3472);
and (n3469,n3470,n3471);
xor (n3470,n3416,n3417);
and (n3471,n94,n135);
and (n3472,n3473,n3474);
xor (n3473,n3470,n3471);
and (n3474,n3475,n3476);
xor (n3475,n3422,n3423);
and (n3476,n89,n135);
and (n3477,n146,n161);
or (n3478,n3479,n3482);
and (n3479,n3480,n3481);
xor (n3480,n3431,n3432);
and (n3481,n176,n161);
and (n3482,n3483,n3484);
xor (n3483,n3480,n3481);
or (n3484,n3485,n3488);
and (n3485,n3486,n3487);
xor (n3486,n3437,n3438);
and (n3487,n170,n161);
and (n3488,n3489,n3490);
xor (n3489,n3486,n3487);
or (n3490,n3491,n3494);
and (n3491,n3492,n3493);
xor (n3492,n3443,n3444);
and (n3493,n246,n161);
and (n3494,n3495,n3496);
xor (n3495,n3492,n3493);
or (n3496,n3497,n3500);
and (n3497,n3498,n3499);
xor (n3498,n3449,n3450);
and (n3499,n298,n161);
and (n3500,n3501,n3502);
xor (n3501,n3498,n3499);
or (n3502,n3503,n3506);
and (n3503,n3504,n3505);
xor (n3504,n3455,n3456);
and (n3505,n323,n161);
and (n3506,n3507,n3508);
xor (n3507,n3504,n3505);
or (n3508,n3509,n3512);
and (n3509,n3510,n3511);
xor (n3510,n3461,n3462);
and (n3511,n197,n161);
and (n3512,n3513,n3514);
xor (n3513,n3510,n3511);
or (n3514,n3515,n3518);
and (n3515,n3516,n3517);
xor (n3516,n3467,n3468);
and (n3517,n94,n161);
and (n3518,n3519,n3520);
xor (n3519,n3516,n3517);
and (n3520,n3521,n997);
xor (n3521,n3473,n3474);
and (n3522,n176,n166);
or (n3523,n3524,n3527);
and (n3524,n3525,n3526);
xor (n3525,n3483,n3484);
and (n3526,n170,n166);
and (n3527,n3528,n3529);
xor (n3528,n3525,n3526);
or (n3529,n3530,n3533);
and (n3530,n3531,n3532);
xor (n3531,n3489,n3490);
and (n3532,n246,n166);
and (n3533,n3534,n3535);
xor (n3534,n3531,n3532);
or (n3535,n3536,n3539);
and (n3536,n3537,n3538);
xor (n3537,n3495,n3496);
and (n3538,n298,n166);
and (n3539,n3540,n3541);
xor (n3540,n3537,n3538);
or (n3541,n3542,n3545);
and (n3542,n3543,n3544);
xor (n3543,n3501,n3502);
and (n3544,n323,n166);
and (n3545,n3546,n3547);
xor (n3546,n3543,n3544);
or (n3547,n3548,n3551);
and (n3548,n3549,n3550);
xor (n3549,n3507,n3508);
and (n3550,n197,n166);
and (n3551,n3552,n3553);
xor (n3552,n3549,n3550);
or (n3553,n3554,n3557);
and (n3554,n3555,n3556);
xor (n3555,n3513,n3514);
and (n3556,n94,n166);
and (n3557,n3558,n3559);
xor (n3558,n3555,n3556);
and (n3559,n3560,n3561);
xor (n3560,n3519,n3520);
and (n3561,n89,n166);
and (n3562,n170,n287);
or (n3563,n3564,n3567);
and (n3564,n3565,n3566);
xor (n3565,n3528,n3529);
and (n3566,n246,n287);
and (n3567,n3568,n3569);
xor (n3568,n3565,n3566);
or (n3569,n3570,n3573);
and (n3570,n3571,n3572);
xor (n3571,n3534,n3535);
and (n3572,n298,n287);
and (n3573,n3574,n3575);
xor (n3574,n3571,n3572);
or (n3575,n3576,n3579);
and (n3576,n3577,n3578);
xor (n3577,n3540,n3541);
and (n3578,n323,n287);
and (n3579,n3580,n3581);
xor (n3580,n3577,n3578);
or (n3581,n3582,n3585);
and (n3582,n3583,n3584);
xor (n3583,n3546,n3547);
and (n3584,n197,n287);
and (n3585,n3586,n3587);
xor (n3586,n3583,n3584);
or (n3587,n3588,n3591);
and (n3588,n3589,n3590);
xor (n3589,n3552,n3553);
and (n3590,n94,n287);
and (n3591,n3592,n3593);
xor (n3592,n3589,n3590);
and (n3593,n3594,n772);
xor (n3594,n3558,n3559);
and (n3595,n246,n286);
or (n3596,n3597,n3599);
and (n3597,n3598,n299);
xor (n3598,n3568,n3569);
and (n3599,n3600,n3601);
xor (n3600,n3598,n299);
or (n3601,n3602,n3605);
and (n3602,n3603,n3604);
xor (n3603,n3574,n3575);
and (n3604,n323,n286);
and (n3605,n3606,n3607);
xor (n3606,n3603,n3604);
or (n3607,n3608,n3611);
and (n3608,n3609,n3610);
xor (n3609,n3580,n3581);
and (n3610,n197,n286);
and (n3611,n3612,n3613);
xor (n3612,n3609,n3610);
or (n3613,n3614,n3617);
and (n3614,n3615,n3616);
xor (n3615,n3586,n3587);
and (n3616,n94,n286);
and (n3617,n3618,n3619);
xor (n3618,n3615,n3616);
and (n3619,n3620,n3621);
xor (n3620,n3592,n3593);
and (n3621,n89,n286);
and (n3622,n298,n311);
or (n3623,n3624,n3627);
and (n3624,n3625,n3626);
xor (n3625,n3600,n3601);
and (n3626,n323,n311);
and (n3627,n3628,n3629);
xor (n3628,n3625,n3626);
or (n3629,n3630,n3633);
and (n3630,n3631,n3632);
xor (n3631,n3606,n3607);
and (n3632,n197,n311);
and (n3633,n3634,n3635);
xor (n3634,n3631,n3632);
or (n3635,n3636,n3639);
and (n3636,n3637,n3638);
xor (n3637,n3612,n3613);
and (n3638,n94,n311);
and (n3639,n3640,n3641);
xor (n3640,n3637,n3638);
and (n3641,n3642,n480);
xor (n3642,n3618,n3619);
and (n3643,n323,n76);
or (n3644,n3645,n3648);
and (n3645,n3646,n3647);
xor (n3646,n3628,n3629);
and (n3647,n197,n76);
and (n3648,n3649,n3650);
xor (n3649,n3646,n3647);
or (n3650,n3651,n3654);
and (n3651,n3652,n3653);
xor (n3652,n3634,n3635);
and (n3653,n94,n76);
and (n3654,n3655,n3656);
xor (n3655,n3652,n3653);
and (n3656,n3657,n3658);
xor (n3657,n3640,n3641);
and (n3658,n89,n76);
and (n3659,n197,n78);
or (n3660,n3661,n3664);
and (n3661,n3662,n3663);
xor (n3662,n3649,n3650);
and (n3663,n94,n78);
and (n3664,n3665,n3666);
xor (n3665,n3662,n3663);
and (n3666,n3667,n453);
xor (n3667,n3655,n3656);
and (n3668,n94,n84);
and (n3669,n3670,n3671);
xor (n3670,n3665,n3666);
and (n3671,n89,n84);
and (n3672,n89,n358);
nor (n3673,n6,n4);
and (n3674,n8,n3675);
not (n3675,n3673);
endmodule
