module top (out,n12,n17,n19,n20,n22,n26,n29,n35,n53
        ,n67,n68,n69,n70,n71,n72,n73,n74,n78,n79
        ,n80,n84,n86,n88,n125,n127,n128,n129,n140,n141
        ,n142,n143,n155,n156,n157,n158,n171,n172,n173,n174
        ,n180,n182,n183,n186,n188,n191,n193,n194,n195,n275
        ,n381,n384,n386,n540,n542,n543,n546,n549,n550,n551
        ,n552,n555,n557,n561,n572,n573,n590,n593,n595,n596
        ,n598,n602,n608,n611,n613,n615,n619,n622,n624,n626
        ,n630,n633,n635,n637,n639,n647,n650,n652,n654,n658
        ,n661,n663,n665,n669,n672,n674,n676,n680,n683,n685
        ,n687,n695,n698,n700,n702,n706,n709,n711,n713,n717
        ,n720,n722,n724,n728,n731,n733,n735,n743,n746,n748
        ,n750,n767,n770,n772,n774,n783,n786,n788,n790,n799
        ,n802,n804,n806,n815,n818,n820,n822,n831,n834,n836
        ,n838,n846,n849,n851,n853,n926,n929,n931,n933,n937
        ,n940,n942,n944,n948,n951,n953,n955,n959,n962,n964
        ,n966,n975,n978,n980,n982,n986,n989,n991,n993,n997
        ,n1000,n1002,n1004,n1008,n1011,n1013,n1015,n1023,n1026,n1028
        ,n1030,n1034,n1037,n1039,n1041,n1045,n1048,n1050,n1052,n1056
        ,n1059,n1061,n1063,n1239,n1242,n1244,n1246,n1255,n1258,n1260
        ,n1262,n1271,n1274,n1276,n1278,n1287,n1290,n1292,n1294,n1303
        ,n1306,n1308,n1310,n1319,n1322,n1324,n1326,n1335,n1338,n1340
        ,n1342,n1350,n1353,n1355,n1357,n1681,n1684,n1686,n1688,n1696
        ,n1699,n1701,n1703,n1718,n1721,n1723,n1725,n1734,n1737,n1739
        ,n1741,n1750,n1753,n1755,n1757,n1766,n1769,n1771,n1773,n1782
        ,n1785,n1787,n1789,n1797,n1800,n1802,n1804,n2020,n2023,n2025
        ,n2027,n2036,n2039,n2041,n2043,n2052,n2055,n2057,n2059,n2068
        ,n2071,n2073,n2075,n2084,n2087,n2089,n2091,n2100,n2103,n2105
        ,n2107,n2116,n2119,n2121,n2123,n2131,n2134,n2136,n2138);
output out;
input n12;
input n17;
input n19;
input n20;
input n22;
input n26;
input n29;
input n35;
input n53;
input n67;
input n68;
input n69;
input n70;
input n71;
input n72;
input n73;
input n74;
input n78;
input n79;
input n80;
input n84;
input n86;
input n88;
input n125;
input n127;
input n128;
input n129;
input n140;
input n141;
input n142;
input n143;
input n155;
input n156;
input n157;
input n158;
input n171;
input n172;
input n173;
input n174;
input n180;
input n182;
input n183;
input n186;
input n188;
input n191;
input n193;
input n194;
input n195;
input n275;
input n381;
input n384;
input n386;
input n540;
input n542;
input n543;
input n546;
input n549;
input n550;
input n551;
input n552;
input n555;
input n557;
input n561;
input n572;
input n573;
input n590;
input n593;
input n595;
input n596;
input n598;
input n602;
input n608;
input n611;
input n613;
input n615;
input n619;
input n622;
input n624;
input n626;
input n630;
input n633;
input n635;
input n637;
input n639;
input n647;
input n650;
input n652;
input n654;
input n658;
input n661;
input n663;
input n665;
input n669;
input n672;
input n674;
input n676;
input n680;
input n683;
input n685;
input n687;
input n695;
input n698;
input n700;
input n702;
input n706;
input n709;
input n711;
input n713;
input n717;
input n720;
input n722;
input n724;
input n728;
input n731;
input n733;
input n735;
input n743;
input n746;
input n748;
input n750;
input n767;
input n770;
input n772;
input n774;
input n783;
input n786;
input n788;
input n790;
input n799;
input n802;
input n804;
input n806;
input n815;
input n818;
input n820;
input n822;
input n831;
input n834;
input n836;
input n838;
input n846;
input n849;
input n851;
input n853;
input n926;
input n929;
input n931;
input n933;
input n937;
input n940;
input n942;
input n944;
input n948;
input n951;
input n953;
input n955;
input n959;
input n962;
input n964;
input n966;
input n975;
input n978;
input n980;
input n982;
input n986;
input n989;
input n991;
input n993;
input n997;
input n1000;
input n1002;
input n1004;
input n1008;
input n1011;
input n1013;
input n1015;
input n1023;
input n1026;
input n1028;
input n1030;
input n1034;
input n1037;
input n1039;
input n1041;
input n1045;
input n1048;
input n1050;
input n1052;
input n1056;
input n1059;
input n1061;
input n1063;
input n1239;
input n1242;
input n1244;
input n1246;
input n1255;
input n1258;
input n1260;
input n1262;
input n1271;
input n1274;
input n1276;
input n1278;
input n1287;
input n1290;
input n1292;
input n1294;
input n1303;
input n1306;
input n1308;
input n1310;
input n1319;
input n1322;
input n1324;
input n1326;
input n1335;
input n1338;
input n1340;
input n1342;
input n1350;
input n1353;
input n1355;
input n1357;
input n1681;
input n1684;
input n1686;
input n1688;
input n1696;
input n1699;
input n1701;
input n1703;
input n1718;
input n1721;
input n1723;
input n1725;
input n1734;
input n1737;
input n1739;
input n1741;
input n1750;
input n1753;
input n1755;
input n1757;
input n1766;
input n1769;
input n1771;
input n1773;
input n1782;
input n1785;
input n1787;
input n1789;
input n1797;
input n1800;
input n1802;
input n1804;
input n2020;
input n2023;
input n2025;
input n2027;
input n2036;
input n2039;
input n2041;
input n2043;
input n2052;
input n2055;
input n2057;
input n2059;
input n2068;
input n2071;
input n2073;
input n2075;
input n2084;
input n2087;
input n2089;
input n2091;
input n2100;
input n2103;
input n2105;
input n2107;
input n2116;
input n2119;
input n2121;
input n2123;
input n2131;
input n2134;
input n2136;
input n2138;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n8;
wire n9;
wire n10;
wire n11;
wire n13;
wire n14;
wire n15;
wire n16;
wire n18;
wire n21;
wire n23;
wire n24;
wire n25;
wire n27;
wire n28;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n75;
wire n76;
wire n77;
wire n81;
wire n82;
wire n83;
wire n85;
wire n87;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n126;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n181;
wire n184;
wire n185;
wire n187;
wire n189;
wire n190;
wire n192;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n382;
wire n383;
wire n385;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n541;
wire n544;
wire n545;
wire n547;
wire n548;
wire n553;
wire n554;
wire n556;
wire n558;
wire n559;
wire n560;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n591;
wire n592;
wire n594;
wire n597;
wire n599;
wire n600;
wire n601;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n609;
wire n610;
wire n612;
wire n614;
wire n616;
wire n617;
wire n618;
wire n620;
wire n621;
wire n623;
wire n625;
wire n627;
wire n628;
wire n629;
wire n631;
wire n632;
wire n634;
wire n636;
wire n638;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n648;
wire n649;
wire n651;
wire n653;
wire n655;
wire n656;
wire n657;
wire n659;
wire n660;
wire n662;
wire n664;
wire n666;
wire n667;
wire n668;
wire n670;
wire n671;
wire n673;
wire n675;
wire n677;
wire n678;
wire n679;
wire n681;
wire n682;
wire n684;
wire n686;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n696;
wire n697;
wire n699;
wire n701;
wire n703;
wire n704;
wire n705;
wire n707;
wire n708;
wire n710;
wire n712;
wire n714;
wire n715;
wire n716;
wire n718;
wire n719;
wire n721;
wire n723;
wire n725;
wire n726;
wire n727;
wire n729;
wire n730;
wire n732;
wire n734;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n744;
wire n745;
wire n747;
wire n749;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n768;
wire n769;
wire n771;
wire n773;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n784;
wire n785;
wire n787;
wire n789;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n800;
wire n801;
wire n803;
wire n805;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n816;
wire n817;
wire n819;
wire n821;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n832;
wire n833;
wire n835;
wire n837;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n847;
wire n848;
wire n850;
wire n852;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n927;
wire n928;
wire n930;
wire n932;
wire n934;
wire n935;
wire n936;
wire n938;
wire n939;
wire n941;
wire n943;
wire n945;
wire n946;
wire n947;
wire n949;
wire n950;
wire n952;
wire n954;
wire n956;
wire n957;
wire n958;
wire n960;
wire n961;
wire n963;
wire n965;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n976;
wire n977;
wire n979;
wire n981;
wire n983;
wire n984;
wire n985;
wire n987;
wire n988;
wire n990;
wire n992;
wire n994;
wire n995;
wire n996;
wire n998;
wire n999;
wire n1001;
wire n1003;
wire n1005;
wire n1006;
wire n1007;
wire n1009;
wire n1010;
wire n1012;
wire n1014;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1024;
wire n1025;
wire n1027;
wire n1029;
wire n1031;
wire n1032;
wire n1033;
wire n1035;
wire n1036;
wire n1038;
wire n1040;
wire n1042;
wire n1043;
wire n1044;
wire n1046;
wire n1047;
wire n1049;
wire n1051;
wire n1053;
wire n1054;
wire n1055;
wire n1057;
wire n1058;
wire n1060;
wire n1062;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1240;
wire n1241;
wire n1243;
wire n1245;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1256;
wire n1257;
wire n1259;
wire n1261;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1272;
wire n1273;
wire n1275;
wire n1277;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1288;
wire n1289;
wire n1291;
wire n1293;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1304;
wire n1305;
wire n1307;
wire n1309;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1320;
wire n1321;
wire n1323;
wire n1325;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1336;
wire n1337;
wire n1339;
wire n1341;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1351;
wire n1352;
wire n1354;
wire n1356;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1682;
wire n1683;
wire n1685;
wire n1687;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1697;
wire n1698;
wire n1700;
wire n1702;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1719;
wire n1720;
wire n1722;
wire n1724;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1735;
wire n1736;
wire n1738;
wire n1740;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1751;
wire n1752;
wire n1754;
wire n1756;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1767;
wire n1768;
wire n1770;
wire n1772;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1783;
wire n1784;
wire n1786;
wire n1788;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1798;
wire n1799;
wire n1801;
wire n1803;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2021;
wire n2022;
wire n2024;
wire n2026;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2037;
wire n2038;
wire n2040;
wire n2042;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2053;
wire n2054;
wire n2056;
wire n2058;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2069;
wire n2070;
wire n2072;
wire n2074;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2085;
wire n2086;
wire n2088;
wire n2090;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2101;
wire n2102;
wire n2104;
wire n2106;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2117;
wire n2118;
wire n2120;
wire n2122;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2132;
wire n2133;
wire n2135;
wire n2137;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2988;
wire n2989;
wire n2990;
wire n2991;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2996;
wire n2997;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3003;
wire n3004;
wire n3005;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3010;
wire n3011;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3038;
wire n3039;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
wire n3056;
wire n3057;
wire n3058;
wire n3059;
wire n3060;
wire n3061;
wire n3062;
wire n3063;
wire n3064;
wire n3065;
wire n3066;
wire n3067;
wire n3068;
wire n3069;
wire n3070;
wire n3071;
wire n3072;
wire n3073;
wire n3074;
wire n3075;
wire n3076;
wire n3077;
wire n3078;
wire n3079;
wire n3080;
wire n3081;
wire n3082;
wire n3083;
wire n3084;
wire n3085;
wire n3086;
wire n3087;
wire n3088;
wire n3089;
wire n3090;
wire n3091;
wire n3092;
wire n3093;
wire n3094;
wire n3095;
wire n3096;
wire n3097;
wire n3098;
wire n3099;
wire n3100;
wire n3101;
wire n3102;
wire n3103;
wire n3104;
wire n3105;
wire n3106;
wire n3107;
wire n3108;
wire n3109;
wire n3110;
wire n3111;
wire n3112;
wire n3113;
wire n3114;
wire n3115;
wire n3116;
wire n3117;
wire n3118;
wire n3119;
wire n3120;
wire n3121;
wire n3122;
wire n3123;
wire n3124;
wire n3125;
wire n3126;
wire n3127;
wire n3128;
wire n3129;
wire n3130;
wire n3131;
wire n3132;
wire n3133;
wire n3134;
wire n3135;
wire n3136;
wire n3137;
wire n3138;
wire n3139;
wire n3140;
wire n3141;
wire n3142;
wire n3143;
wire n3144;
wire n3145;
wire n3146;
wire n3147;
wire n3148;
wire n3149;
wire n3150;
wire n3151;
wire n3152;
wire n3153;
wire n3154;
wire n3155;
wire n3156;
wire n3157;
wire n3158;
wire n3159;
wire n3160;
wire n3161;
wire n3162;
wire n3163;
wire n3164;
wire n3165;
wire n3166;
wire n3167;
wire n3168;
wire n3169;
wire n3170;
wire n3171;
wire n3172;
wire n3173;
wire n3174;
wire n3175;
wire n3176;
wire n3177;
wire n3178;
wire n3179;
wire n3180;
wire n3181;
wire n3182;
wire n3183;
wire n3184;
wire n3185;
wire n3186;
wire n3187;
wire n3188;
wire n3189;
wire n3190;
wire n3191;
wire n3192;
wire n3193;
wire n3194;
wire n3195;
wire n3196;
wire n3197;
wire n3198;
wire n3199;
wire n3200;
wire n3201;
wire n3202;
wire n3203;
wire n3204;
wire n3205;
wire n3206;
wire n3207;
wire n3208;
wire n3209;
wire n3210;
wire n3211;
wire n3212;
wire n3213;
wire n3214;
wire n3215;
wire n3216;
wire n3217;
wire n3218;
wire n3219;
wire n3220;
wire n3221;
wire n3222;
wire n3223;
wire n3224;
wire n3225;
wire n3226;
wire n3227;
wire n3228;
wire n3229;
wire n3230;
wire n3231;
wire n3232;
wire n3233;
wire n3234;
wire n3235;
wire n3236;
wire n3237;
wire n3238;
wire n3239;
wire n3240;
wire n3241;
wire n3242;
wire n3243;
wire n3244;
wire n3245;
wire n3246;
wire n3247;
wire n3248;
wire n3249;
wire n3250;
wire n3251;
wire n3252;
wire n3253;
wire n3254;
wire n3255;
wire n3256;
wire n3257;
wire n3258;
wire n3259;
wire n3260;
wire n3261;
wire n3262;
wire n3263;
wire n3264;
wire n3265;
wire n3266;
wire n3267;
wire n3268;
wire n3269;
wire n3270;
wire n3271;
wire n3272;
wire n3273;
wire n3274;
wire n3275;
wire n3276;
wire n3277;
wire n3278;
wire n3279;
wire n3280;
wire n3281;
wire n3282;
wire n3283;
wire n3284;
wire n3285;
wire n3286;
wire n3287;
wire n3288;
wire n3289;
wire n3290;
wire n3291;
wire n3292;
wire n3293;
wire n3294;
wire n3295;
wire n3296;
wire n3297;
wire n3298;
wire n3299;
wire n3300;
wire n3301;
wire n3302;
wire n3303;
wire n3304;
wire n3305;
wire n3306;
wire n3307;
wire n3308;
wire n3309;
wire n3310;
wire n3311;
wire n3312;
wire n3313;
wire n3314;
wire n3315;
wire n3316;
wire n3317;
wire n3318;
wire n3319;
wire n3320;
wire n3321;
wire n3322;
wire n3323;
wire n3324;
wire n3325;
wire n3326;
wire n3327;
wire n3328;
wire n3329;
wire n3330;
wire n3331;
wire n3332;
wire n3333;
wire n3334;
wire n3335;
wire n3336;
wire n3337;
wire n3338;
wire n3339;
wire n3340;
wire n3341;
wire n3342;
wire n3343;
wire n3344;
wire n3345;
wire n3346;
wire n3347;
wire n3348;
wire n3349;
wire n3350;
wire n3351;
wire n3352;
wire n3353;
wire n3354;
wire n3355;
wire n3356;
wire n3357;
wire n3358;
wire n3359;
wire n3360;
wire n3361;
wire n3362;
wire n3363;
wire n3364;
wire n3365;
wire n3366;
wire n3367;
wire n3368;
wire n3369;
wire n3370;
wire n3371;
wire n3372;
wire n3373;
wire n3374;
wire n3375;
wire n3376;
wire n3377;
wire n3378;
wire n3379;
wire n3380;
wire n3381;
wire n3382;
wire n3383;
wire n3384;
wire n3385;
wire n3386;
wire n3387;
wire n3388;
wire n3389;
wire n3390;
wire n3391;
wire n3392;
wire n3393;
wire n3394;
wire n3395;
wire n3396;
wire n3397;
wire n3398;
wire n3399;
wire n3400;
wire n3401;
wire n3402;
wire n3403;
wire n3404;
wire n3405;
wire n3406;
wire n3407;
wire n3408;
wire n3409;
wire n3410;
wire n3411;
wire n3412;
wire n3413;
wire n3414;
wire n3415;
wire n3416;
wire n3417;
wire n3418;
wire n3419;
wire n3420;
wire n3421;
wire n3422;
wire n3423;
wire n3424;
wire n3425;
wire n3426;
wire n3427;
wire n3428;
xor (out,n0,n2551);
xor (n0,n1,n2528);
xor (n1,n2,n2429);
xor (n2,n3,n1672);
xor (n3,n4,n1577);
xor (n4,n5,n1232);
xor (n5,n6,n1065);
wire s0n6,s1n6,notn6;
or (n6,s0n6,s1n6);
not(notn6,n919);
and (s0n6,notn6,1'b0);
and (s1n6,n919,n8);
xor (n8,n9,n737);
wire s0n9,s1n9,notn9;
or (n9,s0n9,s1n9);
not(notn9,n583);
and (s0n9,notn9,1'b0);
and (s1n9,n583,n10);
wire s0n10,s1n10,notn10;
or (n10,s0n10,s1n10);
not(notn10,n566);
and (s0n10,notn10,n11);
and (s1n10,n566,n553);
wire s0n11,s1n11,notn11;
or (n11,s0n11,s1n11);
not(notn11,n13);
and (s0n11,notn11,1'b0);
and (s1n11,n13,n12);
and (n13,n14,n547);
and (n14,n15,n31);
or (n15,n16,n21,n25,n28);
and (n16,n17,n18);
and (n18,n19,n20);
and (n21,n22,n23);
and (n23,n24,n20);
not (n24,n19);
and (n25,n26,n27);
nor (n27,n24,n20);
and (n28,n29,n30);
nor (n30,n19,n20);
and (n31,n32,n546);
not (n32,n33);
wire s0n33,s1n33,notn33;
or (n33,s0n33,s1n33);
not(notn33,n545);
and (s0n33,notn33,n34);
and (s1n33,n545,1'b0);
wire s0n34,s1n34,notn34;
or (n34,s0n34,s1n34);
not(notn34,n175);
and (s0n34,notn34,n35);
and (s1n34,n175,n36);
wire s0n36,s1n36,notn36;
or (n36,s0n36,s1n36);
not(notn36,n538);
and (s0n36,notn36,n37);
and (s1n36,n538,n512);
or (n37,n38,n480,n511,1'b0,1'b0,1'b0,1'b0,1'b0);
or (n38,n39,n479);
or (n39,n40,n478);
or (n40,n41,n477);
or (n41,n42,n475);
or (n42,n43,n474);
or (n43,n44,n472);
or (n44,n45,n470);
nor (n45,n46,n395,n404,n416,n428,n439,n450,n461);
or (n46,1'b0,n47,n389,n393);
and (n47,n48,n388);
wire s0n48,s1n48,notn48;
or (n48,s0n48,s1n48);
not(notn48,n379);
and (s0n48,notn48,n49);
and (s1n48,n379,n287);
wire s0n49,s1n49,notn49;
or (n49,s0n49,s1n49);
not(notn49,n246);
and (s0n49,notn49,1'b0);
and (s1n49,n246,n50);
or (n50,n51,n227,n231,n235,n238,n241,n243,1'b0);
and (n51,n52,n54);
not (n52,n53);
and (n54,n55,n200,n211,n221);
wire s0n55,s1n55,notn55;
or (n55,s0n55,s1n55);
not(notn55,n89);
and (s0n55,notn55,n56);
and (s1n55,n89,1'b0);
wire s0n56,s1n56,notn56;
or (n56,s0n56,s1n56);
not(notn56,n87);
and (s0n56,notn56,n57);
and (s1n56,n87,n85);
wire s0n57,s1n57,notn57;
or (n57,s0n57,s1n57);
not(notn57,n81);
and (s0n57,notn57,n58);
and (s1n57,n81,n75);
wire s0n58,s1n58,notn58;
or (n58,s0n58,s1n58);
not(notn58,n74);
and (s0n58,notn58,n59);
and (s1n58,n74,1'b0);
wire s0n59,s1n59,notn59;
or (n59,s0n59,s1n59);
not(notn59,n73);
and (s0n59,notn59,n60);
and (s1n59,n73,1'b1);
wire s0n60,s1n60,notn60;
or (n60,s0n60,s1n60);
not(notn60,n72);
and (s0n60,notn60,n61);
and (s1n60,n72,1'b0);
wire s0n61,s1n61,notn61;
or (n61,s0n61,s1n61);
not(notn61,n71);
and (s0n61,notn61,n62);
and (s1n61,n71,1'b1);
wire s0n62,s1n62,notn62;
or (n62,s0n62,s1n62);
not(notn62,n70);
and (s0n62,notn62,n63);
and (s1n62,n70,1'b0);
wire s0n63,s1n63,notn63;
or (n63,s0n63,s1n63);
not(notn63,n69);
and (s0n63,notn63,n64);
and (s1n63,n69,1'b1);
wire s0n64,s1n64,notn64;
or (n64,s0n64,s1n64);
not(notn64,n68);
and (s0n64,notn64,n65);
and (s1n64,n68,1'b0);
wire s0n65,s1n65,notn65;
or (n65,s0n65,s1n65);
not(notn65,n67);
and (s0n65,notn65,n52);
and (s1n65,n67,1'b1);
wire s0n75,s1n75,notn75;
or (n75,s0n75,s1n75);
not(notn75,n80);
and (s0n75,notn75,n76);
and (s1n75,n80,1'b0);
wire s0n76,s1n76,notn76;
or (n76,s0n76,s1n76);
not(notn76,n79);
and (s0n76,notn76,n77);
and (s1n76,n79,1'b1);
not (n77,n78);
or (n81,n82,n84);
or (n82,n83,n78);
or (n83,n80,n79);
not (n85,n86);
or (n87,n86,n88);
not (n89,n90);
or (n90,n91,n198);
or (n91,n92,n196);
or (n92,n93,n190);
or (n93,n94,n189);
or (n94,n95,n185);
or (n95,n96,n184);
or (n96,n97,n179);
or (n97,n98,n178);
or (n98,n99,n177);
or (n99,n100,n175);
or (n100,n101,n169);
or (n101,n102,n168);
or (n102,n103,n167);
or (n103,n104,n166);
or (n104,n105,n165);
or (n105,n106,n164);
or (n106,n107,n163);
or (n107,n108,n162);
or (n108,n109,n159);
or (n109,n110,n153);
or (n110,n111,n152);
or (n111,n112,n151);
or (n112,n113,n150);
or (n113,n114,n149);
or (n114,n115,n148);
or (n115,n116,n146);
or (n116,n117,n144);
or (n117,n118,n138);
or (n118,n119,n137);
or (n119,n120,n136);
or (n120,n121,n135);
or (n121,n122,n134);
or (n122,n123,n132);
or (n123,n124,n130);
nor (n124,n125,n126,n128,n129);
not (n126,n127);
nor (n130,n125,n126,n131,n129);
not (n131,n128);
and (n132,n125,n127,n128,n133);
not (n133,n129);
and (n134,n125,n126,n128,n133);
nor (n135,n125,n127,n131,n129);
and (n136,n125,n126,n128,n129);
and (n137,n125,n127,n128,n129);
nor (n138,n139,n141,n142,n143);
not (n139,n140);
nor (n144,n139,n145,n142,n143);
not (n145,n141);
and (n146,n139,n141,n142,n147);
not (n147,n143);
and (n148,n140,n141,n142,n147);
and (n149,n140,n145,n142,n147);
and (n150,n139,n145,n142,n143);
and (n151,n140,n145,n142,n143);
and (n152,n140,n141,n142,n143);
nor (n153,n154,n156,n157,n158);
not (n154,n155);
and (n159,n155,n156,n160,n161);
not (n160,n157);
not (n161,n158);
and (n162,n154,n156,n160,n161);
and (n163,n155,n156,n157,n161);
nor (n164,n155,n156,n160,n161);
and (n165,n154,n156,n157,n158);
and (n166,n154,n156,n160,n158);
and (n167,n155,n156,n160,n158);
nor (n168,n154,n156,n157,n161);
nor (n169,n170,n172,n173,n174);
not (n170,n171);
nor (n175,n171,n176,n173,n174);
not (n176,n172);
and (n177,n170,n176,n173,n174);
and (n178,n171,n176,n173,n174);
nor (n179,n180,n181,n183);
not (n181,n182);
and (n184,n180,n182,n183);
and (n185,n186,n187);
not (n187,n188);
nor (n189,n186,n187);
nor (n190,n191,n192,n194,n195);
not (n192,n193);
and (n196,n191,n193,n194,n197);
not (n197,n195);
and (n198,n199,n192,n194,n197);
not (n199,n191);
wire s0n200,s1n200,notn200;
or (n200,s0n200,s1n200);
not(notn200,n89);
and (s0n200,notn200,n201);
and (s1n200,n89,1'b0);
wire s0n201,s1n201,notn201;
or (n201,s0n201,s1n201);
not(notn201,n87);
and (s0n201,notn201,n202);
and (s1n201,n87,1'b0);
wire s0n202,s1n202,notn202;
or (n202,s0n202,s1n202);
not(notn202,n81);
and (s0n202,notn202,n203);
and (s1n202,n81,n83);
wire s0n203,s1n203,notn203;
or (n203,s0n203,s1n203);
not(notn203,n74);
and (s0n203,notn203,n204);
and (s1n203,n74,1'b1);
wire s0n204,s1n204,notn204;
or (n204,s0n204,s1n204);
not(notn204,n73);
and (s0n204,notn204,n205);
and (s1n204,n73,1'b1);
wire s0n205,s1n205,notn205;
or (n205,s0n205,s1n205);
not(notn205,n72);
and (s0n205,notn205,n206);
and (s1n205,n72,1'b0);
wire s0n206,s1n206,notn206;
or (n206,s0n206,s1n206);
not(notn206,n71);
and (s0n206,notn206,n207);
and (s1n206,n71,1'b0);
wire s0n207,s1n207,notn207;
or (n207,s0n207,s1n207);
not(notn207,n70);
and (s0n207,notn207,n208);
and (s1n207,n70,1'b1);
wire s0n208,s1n208,notn208;
or (n208,s0n208,s1n208);
not(notn208,n69);
and (s0n208,notn208,n209);
and (s1n208,n69,1'b1);
wire s0n209,s1n209,notn209;
or (n209,s0n209,s1n209);
not(notn209,n68);
and (s0n209,notn209,n210);
and (s1n209,n68,1'b0);
not (n210,n67);
wire s0n211,s1n211,notn211;
or (n211,s0n211,s1n211);
not(notn211,n89);
and (s0n211,notn211,n212);
and (s1n211,n89,1'b0);
wire s0n212,s1n212,notn212;
or (n212,s0n212,s1n212);
not(notn212,n87);
and (s0n212,notn212,n213);
and (s1n212,n87,1'b0);
wire s0n213,s1n213,notn213;
or (n213,s0n213,s1n213);
not(notn213,n81);
and (s0n213,notn213,n214);
and (s1n213,n81,n220);
wire s0n214,s1n214,notn214;
or (n214,s0n214,s1n214);
not(notn214,n74);
and (s0n214,notn214,n215);
and (s1n214,n74,1'b1);
wire s0n215,s1n215,notn215;
or (n215,s0n215,s1n215);
not(notn215,n73);
and (s0n215,notn215,n216);
and (s1n215,n73,1'b1);
wire s0n216,s1n216,notn216;
or (n216,s0n216,s1n216);
not(notn216,n72);
and (s0n216,notn216,n217);
and (s1n216,n72,1'b0);
wire s0n217,s1n217,notn217;
or (n217,s0n217,s1n217);
not(notn217,n71);
and (s0n217,notn217,n218);
and (s1n217,n71,1'b0);
wire s0n218,s1n218,notn218;
or (n218,s0n218,s1n218);
not(notn218,n70);
and (s0n218,notn218,n219);
and (s1n218,n70,1'b0);
not (n219,n69);
not (n220,n83);
not (n221,n222);
wire s0n222,s1n222,notn222;
or (n222,s0n222,s1n222);
not(notn222,n89);
and (s0n222,notn222,n223);
and (s1n222,n89,1'b0);
wire s0n223,s1n223,notn223;
or (n223,s0n223,s1n223);
not(notn223,n87);
and (s0n223,notn223,n224);
and (s1n223,n87,1'b0);
wire s0n224,s1n224,notn224;
or (n224,s0n224,s1n224);
not(notn224,n81);
and (s0n224,notn224,n225);
and (s1n224,n81,1'b0);
wire s0n225,s1n225,notn225;
or (n225,s0n225,s1n225);
not(notn225,n74);
and (s0n225,notn225,n226);
and (s1n225,n74,1'b0);
not (n226,n73);
and (n227,n228,n229);
not (n228,n68);
and (n229,n230,n200,n211,n221);
not (n230,n55);
and (n231,n232,n233);
not (n232,n70);
and (n233,n55,n234,n211,n221);
not (n234,n200);
and (n235,n236,n237);
not (n236,n72);
and (n237,n230,n234,n211,n221);
and (n238,n239,n240);
not (n239,n74);
nor (n240,n230,n234,n211,n222);
and (n241,n77,n242);
nor (n242,n55,n234,n211,n222);
and (n243,n244,n245);
not (n244,n80);
nor (n245,n230,n200,n211,n222);
or (n246,n247,n276);
wire s0n247,s1n247,notn247;
or (n247,s0n247,s1n247);
not(notn247,n274);
and (s0n247,notn247,n248);
and (s1n247,n274,1'b0);
wire s0n248,s1n248,notn248;
or (n248,s0n248,s1n248);
not(notn248,n273);
and (s0n248,notn248,n249);
and (s1n248,n273,n268);
wire s0n249,s1n249,notn249;
or (n249,s0n249,s1n249);
not(notn249,n267);
and (s0n249,notn249,n250);
and (s1n249,n267,n256);
wire s0n250,s1n250,notn250;
or (n250,s0n250,s1n250);
not(notn250,n255);
and (s0n250,notn250,n251);
and (s1n250,n255,n118);
or (n251,n252,n149);
or (n252,n253,n148);
or (n253,n254,n146);
or (n254,n138,n144);
or (n255,n125,n127,n128,n129);
or (n256,1'b0,1'b0,n257,n263,n265);
and (n257,n258,n261);
or (n258,1'b0,1'b0,n259,n179);
and (n259,n260,n182,n183);
not (n260,n180);
and (n261,n170,n176,n173,n262);
not (n262,n174);
and (n263,n186,n264);
and (n264,n171,n176,n173,n262);
or (n265,n266,n177);
or (n266,n169,n175);
or (n267,n171,n172,n173,n174);
or (n268,n269,n168);
or (n269,n270,n166);
or (n270,n271,n163);
or (n271,n272,n162);
or (n272,n153,n159);
or (n273,n155,n156,n157,n158);
not (n274,n275);
wire s0n276,s1n276,notn276;
or (n276,s0n276,s1n276);
not(notn276,n274);
and (s0n276,notn276,n277);
and (s1n276,n274,1'b0);
wire s0n277,s1n277,notn277;
or (n277,s0n277,s1n277);
not(notn277,n273);
and (s0n277,notn277,n278);
and (s1n277,n273,n286);
wire s0n278,s1n278,notn278;
or (n278,s0n278,s1n278);
not(notn278,n267);
and (s0n278,notn278,n279);
and (s1n278,n267,n282);
wire s0n279,s1n279,notn279;
or (n279,s0n279,s1n279);
not(notn279,n255);
and (s0n279,notn279,n280);
and (s1n279,n255,1'b0);
or (n280,n281,n152);
or (n281,n150,n151);
or (n282,1'b0,n178,n283,n285,1'b0);
and (n283,n284,n261);
or (n284,1'b0,n184,n259,1'b0);
and (n285,n188,n264);
or (n286,n165,n167);
not (n287,n288);
nor (n288,n49,n289,n305,n325,n342,n356,n367,n375);
wire s0n289,s1n289,notn289;
or (n289,s0n289,s1n289);
not(notn289,n246);
and (s0n289,notn289,1'b0);
and (s1n289,n246,n290);
or (n290,n291,n293,n295,n297,n299,n301,n303,1'b0);
and (n291,n292,n54);
xnor (n292,n67,n53);
and (n293,n294,n229);
xnor (n294,n69,n68);
and (n295,n296,n233);
xnor (n296,n71,n70);
and (n297,n298,n237);
xnor (n298,n73,n72);
and (n299,n300,n240);
xnor (n300,n84,n74);
and (n301,n302,n242);
xnor (n302,n79,n78);
and (n303,n304,n245);
xnor (n304,n88,n80);
wire s0n305,s1n305,notn305;
or (n305,s0n305,s1n305);
not(notn305,n246);
and (s0n305,notn305,1'b0);
and (s1n305,n246,n306);
or (n306,n307,n310,n313,n316,n319,n322,1'b0,1'b0);
and (n307,n308,n54);
xnor (n308,n68,n309);
or (n309,n67,n53);
and (n310,n311,n229);
xnor (n311,n70,n312);
or (n312,n69,n68);
and (n313,n314,n233);
xnor (n314,n72,n315);
or (n315,n71,n70);
and (n316,n317,n237);
xnor (n317,n74,n318);
or (n318,n73,n72);
and (n319,n320,n240);
xnor (n320,n78,n321);
or (n321,n84,n74);
and (n322,n323,n242);
xnor (n323,n80,n324);
or (n324,n79,n78);
wire s0n325,s1n325,notn325;
or (n325,s0n325,s1n325);
not(notn325,n246);
and (s0n325,notn325,1'b0);
and (s1n325,n246,n326);
or (n326,n327,n330,n333,n336,n339,1'b0,1'b0,1'b0);
and (n327,n328,n54);
xnor (n328,n69,n329);
or (n329,n68,n309);
and (n330,n331,n229);
xnor (n331,n71,n332);
or (n332,n70,n312);
and (n333,n334,n233);
xnor (n334,n73,n335);
or (n335,n72,n315);
and (n336,n337,n237);
xnor (n337,n84,n338);
or (n338,n74,n318);
and (n339,n340,n240);
xnor (n340,n79,n341);
or (n341,n78,n321);
wire s0n342,s1n342,notn342;
or (n342,s0n342,s1n342);
not(notn342,n246);
and (s0n342,notn342,1'b0);
and (s1n342,n246,n343);
or (n343,n344,n347,n350,n353,1'b0,1'b0,1'b0,1'b0);
and (n344,n345,n54);
xnor (n345,n70,n346);
or (n346,n69,n329);
and (n347,n348,n229);
xnor (n348,n72,n349);
or (n349,n71,n332);
and (n350,n351,n233);
xnor (n351,n74,n352);
or (n352,n73,n335);
and (n353,n354,n237);
xnor (n354,n78,n355);
or (n355,n84,n338);
wire s0n356,s1n356,notn356;
or (n356,s0n356,s1n356);
not(notn356,n246);
and (s0n356,notn356,1'b0);
and (s1n356,n246,n357);
or (n357,n358,n361,n364,1'b0,1'b0,1'b0,1'b0,1'b0);
and (n358,n359,n54);
xnor (n359,n71,n360);
or (n360,n70,n346);
and (n361,n362,n229);
xnor (n362,n73,n363);
or (n363,n72,n349);
and (n364,n365,n233);
xnor (n365,n84,n366);
or (n366,n74,n352);
wire s0n367,s1n367,notn367;
or (n367,s0n367,s1n367);
not(notn367,n246);
and (s0n367,notn367,1'b0);
and (s1n367,n246,n368);
or (n368,n369,n372,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0);
and (n369,n370,n54);
xnor (n370,n72,n371);
or (n371,n71,n360);
and (n372,n373,n229);
xnor (n373,n74,n374);
or (n374,n73,n363);
wire s0n375,s1n375,notn375;
or (n375,s0n375,s1n375);
not(notn375,n246);
and (s0n375,notn375,1'b0);
and (s1n375,n246,n376);
and (n376,n377,n54);
xnor (n377,n73,n378);
or (n378,n72,n371);
nor (n379,n380,n382,n385);
not (n380,n381);
not (n382,n383);
xor (n383,n384,n381);
xor (n385,n386,n387);
and (n387,n384,n381);
and (n388,n247,n276);
and (n389,n390,n391);
xor (n390,n289,n49);
nor (n391,n247,n392);
not (n392,n276);
and (n393,n49,n394);
and (n394,n247,n392);
not (n395,n396);
or (n396,1'b0,n397,n399,n403);
and (n397,n398,n388);
wire s0n398,s1n398,notn398;
or (n398,s0n398,s1n398);
not(notn398,n379);
and (s0n398,notn398,n289);
and (s1n398,n379,1'b0);
and (n399,n400,n391);
xor (n400,n401,n402);
not (n401,n305);
not (n402,n289);
and (n403,n289,n394);
or (n404,1'b0,n405,n407,n415);
and (n405,n406,n388);
wire s0n406,s1n406,notn406;
or (n406,s0n406,s1n406);
not(notn406,n379);
and (s0n406,notn406,n305);
and (s1n406,n379,1'b0);
and (n407,n408,n391);
wire s0n408,s1n408,notn408;
or (n408,s0n408,s1n408);
not(notn408,n49);
and (s0n408,notn408,n409);
and (s1n408,n49,n412);
xor (n409,n410,n411);
not (n410,n325);
and (n411,n401,n402);
xor (n412,n325,n413);
and (n413,n305,n414);
and (n414,n289,n49);
and (n415,n305,n394);
not (n416,n417);
or (n417,1'b0,n418,n420,n427);
and (n418,n419,n388);
wire s0n419,s1n419,notn419;
or (n419,s0n419,s1n419);
not(notn419,n379);
and (s0n419,notn419,n325);
and (s1n419,n379,1'b0);
and (n420,n421,n391);
wire s0n421,s1n421,notn421;
or (n421,s0n421,s1n421);
not(notn421,n49);
and (s0n421,notn421,n422);
and (s1n421,n49,n425);
xor (n422,n423,n424);
not (n423,n342);
and (n424,n410,n411);
xor (n425,n342,n426);
and (n426,n325,n413);
and (n427,n325,n394);
or (n428,1'b0,n429,n431,n438);
and (n429,n430,n388);
wire s0n430,s1n430,notn430;
or (n430,s0n430,s1n430);
not(notn430,n379);
and (s0n430,notn430,n342);
and (s1n430,n379,1'b0);
and (n431,n432,n391);
wire s0n432,s1n432,notn432;
or (n432,s0n432,s1n432);
not(notn432,n49);
and (s0n432,notn432,n433);
and (s1n432,n49,n436);
xor (n433,n434,n435);
not (n434,n356);
and (n435,n423,n424);
xor (n436,n356,n437);
and (n437,n342,n426);
and (n438,n342,n394);
or (n439,1'b0,n440,n442,n449);
and (n440,n441,n388);
wire s0n441,s1n441,notn441;
or (n441,s0n441,s1n441);
not(notn441,n379);
and (s0n441,notn441,n356);
and (s1n441,n379,1'b0);
and (n442,n443,n391);
wire s0n443,s1n443,notn443;
or (n443,s0n443,s1n443);
not(notn443,n49);
and (s0n443,notn443,n444);
and (s1n443,n49,n447);
xor (n444,n445,n446);
not (n445,n367);
and (n446,n434,n435);
xor (n447,n367,n448);
and (n448,n356,n437);
and (n449,n356,n394);
or (n450,1'b0,n451,n453,n460);
and (n451,n452,n388);
wire s0n452,s1n452,notn452;
or (n452,s0n452,s1n452);
not(notn452,n379);
and (s0n452,notn452,n367);
and (s1n452,n379,1'b0);
and (n453,n454,n391);
wire s0n454,s1n454,notn454;
or (n454,s0n454,s1n454);
not(notn454,n49);
and (s0n454,notn454,n455);
and (s1n454,n49,n458);
xor (n455,n456,n457);
not (n456,n375);
and (n457,n445,n446);
xor (n458,n375,n459);
and (n459,n367,n448);
and (n460,n367,n394);
or (n461,1'b0,n462,n464,n469);
and (n462,n463,n388);
wire s0n463,s1n463,notn463;
or (n463,s0n463,s1n463);
not(notn463,n379);
and (s0n463,notn463,n375);
and (s1n463,n379,1'b0);
and (n464,n465,n391);
wire s0n465,s1n465,notn465;
or (n465,s0n465,s1n465);
not(notn465,n49);
and (s0n465,notn465,n466);
and (s1n465,n49,n468);
not (n466,n467);
and (n467,n456,n457);
and (n468,n375,n459);
and (n469,n375,n394);
nor (n470,n471,n395,n404,n416,n428,n439,n450,n461);
not (n471,n46);
nor (n472,n46,n396,n473,n416,n428,n439,n450,n461);
not (n473,n404);
nor (n474,n471,n396,n473,n416,n428,n439,n450,n461);
nor (n475,n46,n395,n473,n417,n476,n439,n450,n461);
not (n476,n428);
nor (n477,n471,n395,n473,n417,n476,n439,n450,n461);
nor (n478,n46,n396,n404,n416,n476,n439,n450,n461);
nor (n479,n471,n396,n404,n416,n476,n439,n450,n461);
or (n480,n481,n496);
or (n481,n482,n495);
or (n482,n483,n494);
or (n483,n484,n493);
or (n484,n485,n492);
or (n485,n486,n491);
or (n486,n487,n490);
or (n487,n488,n489);
nor (n488,n46,n395,n473,n417,n428,n439,n450,n461);
nor (n489,n471,n395,n473,n417,n428,n439,n450,n461);
nor (n490,n46,n396,n404,n416,n428,n439,n450,n461);
nor (n491,n471,n396,n404,n416,n428,n439,n450,n461);
nor (n492,n46,n395,n404,n417,n476,n439,n450,n461);
nor (n493,n471,n395,n404,n417,n476,n439,n450,n461);
nor (n494,n46,n396,n473,n417,n476,n439,n450,n461);
nor (n495,n471,n396,n473,n417,n476,n439,n450,n461);
or (n496,n497,n510);
or (n497,n498,n509);
or (n498,n499,n508);
or (n499,n500,n507);
or (n500,n501,n506);
or (n501,n502,n505);
or (n502,n503,n504);
nor (n503,n46,n395,n473,n416,n428,n439,n450,n461);
nor (n504,n471,n395,n473,n416,n428,n439,n450,n461);
nor (n505,n46,n396,n404,n417,n476,n439,n450,n461);
nor (n506,n471,n396,n404,n417,n476,n439,n450,n461);
nor (n507,n46,n395,n404,n416,n476,n439,n450,n461);
nor (n508,n471,n395,n404,n416,n476,n439,n450,n461);
nor (n509,n46,n396,n473,n416,n476,n439,n450,n461);
nor (n510,n471,n396,n473,n416,n476,n439,n450,n461);
nor (n511,n471,n396,n473,n417,n428,n439,n450,n461);
or (n512,1'b0,n513,n520,n527,n288);
or (n513,n514,n478);
or (n514,n515,n477);
or (n515,n516,n475);
or (n516,n517,n495);
or (n517,n518,n472);
or (n518,n519,n470);
or (n519,n491,n45);
or (n520,n521,n494);
or (n521,n522,n493);
or (n522,n523,n492);
or (n523,n524,n506);
or (n524,n525,n490);
or (n525,n526,n489);
or (n526,n511,n488);
or (n527,n528,n505);
or (n528,n529,n504);
or (n529,n530,n503);
or (n530,n531,n474);
or (n531,n532,n537);
or (n532,n533,n536);
or (n533,n534,n535);
nor (n534,n471,n396,n404,n417,n428,n439,n450,n461);
nor (n535,n46,n395,n404,n417,n428,n439,n450,n461);
nor (n536,n471,n395,n404,n417,n428,n439,n450,n461);
nor (n537,n46,n396,n473,n417,n428,n439,n450,n461);
or (n538,n539,n544);
nor (n539,n540,n541,n543);
not (n541,n542);
and (n544,n540,n542,n543);
nor (n545,n170,n176,n173,n174);
nor (n547,n548,n550,n551,n552);
not (n548,n549);
or (n553,1'b0,n554,n556,n560,n563);
and (n554,n555,n547);
and (n556,n557,n558);
nor (n558,n549,n559,n551,n552);
not (n559,n550);
and (n560,n561,n562);
nor (n562,n548,n559,n551,n552);
and (n563,n12,n564);
and (n564,n548,n559,n551,n565);
not (n565,n552);
and (n566,n31,n567);
not (n567,n568);
wire s0n568,s1n568,notn568;
or (n568,s0n568,s1n568);
not(notn568,n581);
and (s0n568,notn568,n14);
and (s1n568,n581,n569);
or (n569,n570,n574,n577,n579);
and (n570,n17,n571);
and (n571,n572,n573);
and (n574,n22,n575);
and (n575,n576,n573);
not (n576,n572);
and (n577,n26,n578);
nor (n578,n576,n573);
and (n579,n29,n580);
nor (n580,n572,n573);
and (n581,n32,n582);
not (n582,n546);
and (n583,n584,n640);
not (n584,n585);
wire s0n585,s1n585,notn585;
or (n585,s0n585,s1n585);
not(notn585,n31);
and (s0n585,notn585,1'b0);
and (s1n585,n31,n586);
wire s0n586,s1n586,notn586;
or (n586,s0n586,s1n586);
not(notn586,n639);
and (s0n586,notn586,n587);
and (s1n586,n639,n630);
or (n587,n588,n606,n617,n628);
and (n588,n589,n18);
wire s0n589,s1n589,notn589;
or (n589,s0n589,s1n589);
not(notn589,n568);
and (s0n589,notn589,n590);
and (s1n589,n568,n591);
or (n591,n592,n597,n601,n604);
and (n592,n593,n594);
nor (n594,n595,n596);
and (n597,n598,n599);
and (n599,n595,n600);
not (n600,n596);
and (n601,n602,n603);
nor (n603,n595,n600);
and (n604,n590,n605);
and (n605,n595,n596);
and (n606,n607,n23);
wire s0n607,s1n607,notn607;
or (n607,s0n607,s1n607);
not(notn607,n568);
and (s0n607,notn607,n608);
and (s1n607,n568,n609);
or (n609,n610,n612,n614,n616);
and (n610,n611,n594);
and (n612,n613,n599);
and (n614,n615,n603);
and (n616,n608,n605);
and (n617,n618,n27);
wire s0n618,s1n618,notn618;
or (n618,s0n618,s1n618);
not(notn618,n568);
and (s0n618,notn618,n619);
and (s1n618,n568,n620);
or (n620,n621,n623,n625,n627);
and (n621,n622,n594);
and (n623,n624,n599);
and (n625,n626,n603);
and (n627,n619,n605);
and (n628,n629,n30);
wire s0n629,s1n629,notn629;
or (n629,s0n629,s1n629);
not(notn629,n568);
and (s0n629,notn629,n630);
and (s1n629,n568,n631);
or (n631,n632,n634,n636,n638);
and (n632,n633,n594);
and (n634,n635,n599);
and (n636,n637,n603);
and (n638,n630,n605);
and (n640,n641,n689);
not (n641,n642);
wire s0n642,s1n642,notn642;
or (n642,s0n642,s1n642);
not(notn642,n31);
and (s0n642,notn642,1'b0);
and (s1n642,n31,n643);
wire s0n643,s1n643,notn643;
or (n643,s0n643,s1n643);
not(notn643,n639);
and (s0n643,notn643,n644);
and (s1n643,n639,n680);
or (n644,n645,n656,n667,n678);
and (n645,n646,n18);
wire s0n646,s1n646,notn646;
or (n646,s0n646,s1n646);
not(notn646,n568);
and (s0n646,notn646,n647);
and (s1n646,n568,n648);
or (n648,n649,n651,n653,n655);
and (n649,n650,n594);
and (n651,n652,n599);
and (n653,n654,n603);
and (n655,n647,n605);
and (n656,n657,n23);
wire s0n657,s1n657,notn657;
or (n657,s0n657,s1n657);
not(notn657,n568);
and (s0n657,notn657,n658);
and (s1n657,n568,n659);
or (n659,n660,n662,n664,n666);
and (n660,n661,n594);
and (n662,n663,n599);
and (n664,n665,n603);
and (n666,n658,n605);
and (n667,n668,n27);
wire s0n668,s1n668,notn668;
or (n668,s0n668,s1n668);
not(notn668,n568);
and (s0n668,notn668,n669);
and (s1n668,n568,n670);
or (n670,n671,n673,n675,n677);
and (n671,n672,n594);
and (n673,n674,n599);
and (n675,n676,n603);
and (n677,n669,n605);
and (n678,n679,n30);
wire s0n679,s1n679,notn679;
or (n679,s0n679,s1n679);
not(notn679,n568);
and (s0n679,notn679,n680);
and (s1n679,n568,n681);
or (n681,n682,n684,n686,n688);
and (n682,n683,n594);
and (n684,n685,n599);
and (n686,n687,n603);
and (n688,n680,n605);
not (n689,n690);
wire s0n690,s1n690,notn690;
or (n690,s0n690,s1n690);
not(notn690,n31);
and (s0n690,notn690,1'b0);
and (s1n690,n31,n691);
wire s0n691,s1n691,notn691;
or (n691,s0n691,s1n691);
not(notn691,n639);
and (s0n691,notn691,n692);
and (s1n691,n639,n728);
or (n692,n693,n704,n715,n726);
and (n693,n694,n18);
wire s0n694,s1n694,notn694;
or (n694,s0n694,s1n694);
not(notn694,n568);
and (s0n694,notn694,n695);
and (s1n694,n568,n696);
or (n696,n697,n699,n701,n703);
and (n697,n698,n594);
and (n699,n700,n599);
and (n701,n702,n603);
and (n703,n695,n605);
and (n704,n705,n23);
wire s0n705,s1n705,notn705;
or (n705,s0n705,s1n705);
not(notn705,n568);
and (s0n705,notn705,n706);
and (s1n705,n568,n707);
or (n707,n708,n710,n712,n714);
and (n708,n709,n594);
and (n710,n711,n599);
and (n712,n713,n603);
and (n714,n706,n605);
and (n715,n716,n27);
wire s0n716,s1n716,notn716;
or (n716,s0n716,s1n716);
not(notn716,n568);
and (s0n716,notn716,n717);
and (s1n716,n568,n718);
or (n718,n719,n721,n723,n725);
and (n719,n720,n594);
and (n721,n722,n599);
and (n723,n724,n603);
and (n725,n717,n605);
and (n726,n727,n30);
wire s0n727,s1n727,notn727;
or (n727,s0n727,s1n727);
not(notn727,n568);
and (s0n727,notn727,n728);
and (s1n727,n568,n729);
or (n729,n730,n732,n734,n736);
and (n730,n731,n594);
and (n732,n733,n599);
and (n734,n735,n603);
and (n736,n728,n605);
or (n737,n738,n860,n918);
and (n738,n739,n754);
xor (n739,n740,n752);
wire s0n740,s1n740,notn740;
or (n740,s0n740,s1n740);
not(notn740,n583);
and (s0n740,notn740,1'b0);
and (s1n740,n583,n741);
wire s0n741,s1n741,notn741;
or (n741,s0n741,s1n741);
not(notn741,n566);
and (s0n741,notn741,n742);
and (s1n741,n566,n744);
wire s0n742,s1n742,notn742;
or (n742,s0n742,s1n742);
not(notn742,n13);
and (s0n742,notn742,1'b0);
and (s1n742,n13,n743);
or (n744,1'b0,n745,n747,n749,n751);
and (n745,n746,n547);
and (n747,n748,n558);
and (n749,n750,n562);
and (n751,n743,n564);
wire s0n752,s1n752,notn752;
or (n752,s0n752,s1n752);
not(notn752,n753);
and (s0n752,notn752,1'b0);
and (s1n752,n753,n10);
xor (n753,n584,n640);
and (n754,n755,n757);
wire s0n755,s1n755,notn755;
or (n755,s0n755,s1n755);
not(notn755,n756);
and (s0n755,notn755,1'b0);
and (s1n755,n756,n10);
xor (n756,n641,n689);
or (n757,n758,n761,n859);
and (n758,n759,n760);
wire s0n759,s1n759,notn759;
or (n759,s0n759,s1n759);
not(notn759,n756);
and (s0n759,notn759,1'b0);
and (s1n759,n756,n741);
wire s0n760,s1n760,notn760;
or (n760,s0n760,s1n760);
not(notn760,n690);
and (s0n760,notn760,1'b0);
and (s1n760,n690,n10);
and (n761,n760,n762);
or (n762,n763,n777,n858);
and (n763,n764,n776);
wire s0n764,s1n764,notn764;
or (n764,s0n764,s1n764);
not(notn764,n756);
and (s0n764,notn764,1'b0);
and (s1n764,n756,n765);
wire s0n765,s1n765,notn765;
or (n765,s0n765,s1n765);
not(notn765,n566);
and (s0n765,notn765,n766);
and (s1n765,n566,n768);
wire s0n766,s1n766,notn766;
or (n766,s0n766,s1n766);
not(notn766,n13);
and (s0n766,notn766,1'b0);
and (s1n766,n13,n767);
or (n768,1'b0,n769,n771,n773,n775);
and (n769,n770,n547);
and (n771,n772,n558);
and (n773,n774,n562);
and (n775,n767,n564);
wire s0n776,s1n776,notn776;
or (n776,s0n776,s1n776);
not(notn776,n690);
and (s0n776,notn776,1'b0);
and (s1n776,n690,n741);
and (n777,n776,n778);
or (n778,n779,n793,n857);
and (n779,n780,n792);
wire s0n780,s1n780,notn780;
or (n780,s0n780,s1n780);
not(notn780,n756);
and (s0n780,notn780,1'b0);
and (s1n780,n756,n781);
wire s0n781,s1n781,notn781;
or (n781,s0n781,s1n781);
not(notn781,n566);
and (s0n781,notn781,n782);
and (s1n781,n566,n784);
wire s0n782,s1n782,notn782;
or (n782,s0n782,s1n782);
not(notn782,n13);
and (s0n782,notn782,1'b0);
and (s1n782,n13,n783);
or (n784,1'b0,n785,n787,n789,n791);
and (n785,n786,n547);
and (n787,n788,n558);
and (n789,n790,n562);
and (n791,n783,n564);
wire s0n792,s1n792,notn792;
or (n792,s0n792,s1n792);
not(notn792,n690);
and (s0n792,notn792,1'b0);
and (s1n792,n690,n765);
and (n793,n792,n794);
or (n794,n795,n809,n856);
and (n795,n796,n808);
wire s0n796,s1n796,notn796;
or (n796,s0n796,s1n796);
not(notn796,n756);
and (s0n796,notn796,1'b0);
and (s1n796,n756,n797);
wire s0n797,s1n797,notn797;
or (n797,s0n797,s1n797);
not(notn797,n566);
and (s0n797,notn797,n798);
and (s1n797,n566,n800);
wire s0n798,s1n798,notn798;
or (n798,s0n798,s1n798);
not(notn798,n13);
and (s0n798,notn798,1'b0);
and (s1n798,n13,n799);
or (n800,1'b0,n801,n803,n805,n807);
and (n801,n802,n547);
and (n803,n804,n558);
and (n805,n806,n562);
and (n807,n799,n564);
wire s0n808,s1n808,notn808;
or (n808,s0n808,s1n808);
not(notn808,n690);
and (s0n808,notn808,1'b0);
and (s1n808,n690,n781);
and (n809,n808,n810);
or (n810,n811,n825,n827);
and (n811,n812,n824);
wire s0n812,s1n812,notn812;
or (n812,s0n812,s1n812);
not(notn812,n756);
and (s0n812,notn812,1'b0);
and (s1n812,n756,n813);
wire s0n813,s1n813,notn813;
or (n813,s0n813,s1n813);
not(notn813,n566);
and (s0n813,notn813,n814);
and (s1n813,n566,n816);
wire s0n814,s1n814,notn814;
or (n814,s0n814,s1n814);
not(notn814,n13);
and (s0n814,notn814,1'b0);
and (s1n814,n13,n815);
or (n816,1'b0,n817,n819,n821,n823);
and (n817,n818,n547);
and (n819,n820,n558);
and (n821,n822,n562);
and (n823,n815,n564);
wire s0n824,s1n824,notn824;
or (n824,s0n824,s1n824);
not(notn824,n690);
and (s0n824,notn824,1'b0);
and (s1n824,n690,n797);
and (n825,n824,n826);
or (n826,n827,n841,n842);
and (n827,n828,n840);
wire s0n828,s1n828,notn828;
or (n828,s0n828,s1n828);
not(notn828,n756);
and (s0n828,notn828,1'b0);
and (s1n828,n756,n829);
wire s0n829,s1n829,notn829;
or (n829,s0n829,s1n829);
not(notn829,n566);
and (s0n829,notn829,n830);
and (s1n829,n566,n832);
wire s0n830,s1n830,notn830;
or (n830,s0n830,s1n830);
not(notn830,n13);
and (s0n830,notn830,1'b0);
and (s1n830,n13,n831);
or (n832,1'b0,n833,n835,n837,n839);
and (n833,n834,n547);
and (n835,n836,n558);
and (n837,n838,n562);
and (n839,n831,n564);
wire s0n840,s1n840,notn840;
or (n840,s0n840,s1n840);
not(notn840,n690);
and (s0n840,notn840,1'b0);
and (s1n840,n690,n813);
and (n841,n840,n842);
and (n842,n843,n855);
wire s0n843,s1n843,notn843;
or (n843,s0n843,s1n843);
not(notn843,n756);
and (s0n843,notn843,1'b0);
and (s1n843,n756,n844);
wire s0n844,s1n844,notn844;
or (n844,s0n844,s1n844);
not(notn844,n566);
and (s0n844,notn844,n845);
and (s1n844,n566,n847);
wire s0n845,s1n845,notn845;
or (n845,s0n845,s1n845);
not(notn845,n13);
and (s0n845,notn845,1'b0);
and (s1n845,n13,n846);
or (n847,1'b0,n848,n850,n852,n854);
and (n848,n849,n547);
and (n850,n851,n558);
and (n852,n853,n562);
and (n854,n846,n564);
wire s0n855,s1n855,notn855;
or (n855,s0n855,s1n855);
not(notn855,n690);
and (s0n855,notn855,1'b0);
and (s1n855,n690,n829);
and (n856,n796,n810);
and (n857,n780,n794);
and (n858,n764,n778);
and (n859,n759,n762);
and (n860,n754,n861);
or (n861,n862,n867,n917);
and (n862,n863,n866);
xor (n863,n864,n865);
wire s0n864,s1n864,notn864;
or (n864,s0n864,s1n864);
not(notn864,n583);
and (s0n864,notn864,1'b0);
and (s1n864,n583,n765);
wire s0n865,s1n865,notn865;
or (n865,s0n865,s1n865);
not(notn865,n753);
and (s0n865,notn865,1'b0);
and (s1n865,n753,n741);
xor (n866,n755,n757);
and (n867,n866,n868);
or (n868,n869,n875,n916);
and (n869,n870,n873);
xor (n870,n871,n872);
wire s0n871,s1n871,notn871;
or (n871,s0n871,s1n871);
not(notn871,n583);
and (s0n871,notn871,1'b0);
and (s1n871,n583,n781);
wire s0n872,s1n872,notn872;
or (n872,s0n872,s1n872);
not(notn872,n753);
and (s0n872,notn872,1'b0);
and (s1n872,n753,n765);
xor (n873,n874,n762);
xor (n874,n759,n760);
and (n875,n873,n876);
or (n876,n877,n883,n915);
and (n877,n878,n881);
xor (n878,n879,n880);
wire s0n879,s1n879,notn879;
or (n879,s0n879,s1n879);
not(notn879,n583);
and (s0n879,notn879,1'b0);
and (s1n879,n583,n797);
wire s0n880,s1n880,notn880;
or (n880,s0n880,s1n880);
not(notn880,n753);
and (s0n880,notn880,1'b0);
and (s1n880,n753,n781);
xor (n881,n882,n778);
xor (n882,n764,n776);
and (n883,n881,n884);
or (n884,n885,n891,n914);
and (n885,n886,n889);
xor (n886,n887,n888);
wire s0n887,s1n887,notn887;
or (n887,s0n887,s1n887);
not(notn887,n583);
and (s0n887,notn887,1'b0);
and (s1n887,n583,n813);
wire s0n888,s1n888,notn888;
or (n888,s0n888,s1n888);
not(notn888,n753);
and (s0n888,notn888,1'b0);
and (s1n888,n753,n797);
xor (n889,n890,n794);
xor (n890,n780,n792);
and (n891,n889,n892);
or (n892,n893,n899,n913);
and (n893,n894,n897);
xor (n894,n895,n896);
wire s0n895,s1n895,notn895;
or (n895,s0n895,s1n895);
not(notn895,n583);
and (s0n895,notn895,1'b0);
and (s1n895,n583,n829);
wire s0n896,s1n896,notn896;
or (n896,s0n896,s1n896);
not(notn896,n753);
and (s0n896,notn896,1'b0);
and (s1n896,n753,n813);
xor (n897,n898,n810);
xor (n898,n796,n808);
and (n899,n897,n900);
or (n900,n901,n907,n912);
and (n901,n902,n905);
xor (n902,n903,n904);
wire s0n903,s1n903,notn903;
or (n903,s0n903,s1n903);
not(notn903,n583);
and (s0n903,notn903,1'b0);
and (s1n903,n583,n844);
wire s0n904,s1n904,notn904;
or (n904,s0n904,s1n904);
not(notn904,n753);
and (s0n904,notn904,1'b0);
and (s1n904,n753,n829);
xor (n905,n906,n826);
xor (n906,n812,n824);
and (n907,n905,n908);
and (n908,n909,n910);
wire s0n909,s1n909,notn909;
or (n909,s0n909,s1n909);
not(notn909,n753);
and (s0n909,notn909,1'b0);
and (s1n909,n753,n844);
xor (n910,n911,n842);
xor (n911,n828,n840);
and (n912,n902,n908);
and (n913,n894,n900);
and (n914,n886,n892);
and (n915,n878,n884);
and (n916,n870,n876);
and (n917,n863,n868);
and (n918,n739,n861);
and (n919,n920,n968);
not (n920,n921);
wire s0n921,s1n921,notn921;
or (n921,s0n921,s1n921);
not(notn921,n31);
and (s0n921,notn921,1'b0);
and (s1n921,n31,n922);
wire s0n922,s1n922,notn922;
or (n922,s0n922,s1n922);
not(notn922,n639);
and (s0n922,notn922,n923);
and (s1n922,n639,n959);
or (n923,n924,n935,n946,n957);
and (n924,n925,n18);
wire s0n925,s1n925,notn925;
or (n925,s0n925,s1n925);
not(notn925,n568);
and (s0n925,notn925,n926);
and (s1n925,n568,n927);
or (n927,n928,n930,n932,n934);
and (n928,n929,n594);
and (n930,n931,n599);
and (n932,n933,n603);
and (n934,n926,n605);
and (n935,n936,n23);
wire s0n936,s1n936,notn936;
or (n936,s0n936,s1n936);
not(notn936,n568);
and (s0n936,notn936,n937);
and (s1n936,n568,n938);
or (n938,n939,n941,n943,n945);
and (n939,n940,n594);
and (n941,n942,n599);
and (n943,n944,n603);
and (n945,n937,n605);
and (n946,n947,n27);
wire s0n947,s1n947,notn947;
or (n947,s0n947,s1n947);
not(notn947,n568);
and (s0n947,notn947,n948);
and (s1n947,n568,n949);
or (n949,n950,n952,n954,n956);
and (n950,n951,n594);
and (n952,n953,n599);
and (n954,n955,n603);
and (n956,n948,n605);
and (n957,n958,n30);
wire s0n958,s1n958,notn958;
or (n958,s0n958,s1n958);
not(notn958,n568);
and (s0n958,notn958,n959);
and (s1n958,n568,n960);
or (n960,n961,n963,n965,n967);
and (n961,n962,n594);
and (n963,n964,n599);
and (n965,n966,n603);
and (n967,n959,n605);
and (n968,n969,n1017);
not (n969,n970);
wire s0n970,s1n970,notn970;
or (n970,s0n970,s1n970);
not(notn970,n31);
and (s0n970,notn970,1'b0);
and (s1n970,n31,n971);
wire s0n971,s1n971,notn971;
or (n971,s0n971,s1n971);
not(notn971,n639);
and (s0n971,notn971,n972);
and (s1n971,n639,n1008);
or (n972,n973,n984,n995,n1006);
and (n973,n974,n18);
wire s0n974,s1n974,notn974;
or (n974,s0n974,s1n974);
not(notn974,n568);
and (s0n974,notn974,n975);
and (s1n974,n568,n976);
or (n976,n977,n979,n981,n983);
and (n977,n978,n594);
and (n979,n980,n599);
and (n981,n982,n603);
and (n983,n975,n605);
and (n984,n985,n23);
wire s0n985,s1n985,notn985;
or (n985,s0n985,s1n985);
not(notn985,n568);
and (s0n985,notn985,n986);
and (s1n985,n568,n987);
or (n987,n988,n990,n992,n994);
and (n988,n989,n594);
and (n990,n991,n599);
and (n992,n993,n603);
and (n994,n986,n605);
and (n995,n996,n27);
wire s0n996,s1n996,notn996;
or (n996,s0n996,s1n996);
not(notn996,n568);
and (s0n996,notn996,n997);
and (s1n996,n568,n998);
or (n998,n999,n1001,n1003,n1005);
and (n999,n1000,n594);
and (n1001,n1002,n599);
and (n1003,n1004,n603);
and (n1005,n997,n605);
and (n1006,n1007,n30);
wire s0n1007,s1n1007,notn1007;
or (n1007,s0n1007,s1n1007);
not(notn1007,n568);
and (s0n1007,notn1007,n1008);
and (s1n1007,n568,n1009);
or (n1009,n1010,n1012,n1014,n1016);
and (n1010,n1011,n594);
and (n1012,n1013,n599);
and (n1014,n1015,n603);
and (n1016,n1008,n605);
not (n1017,n1018);
wire s0n1018,s1n1018,notn1018;
or (n1018,s0n1018,s1n1018);
not(notn1018,n31);
and (s0n1018,notn1018,1'b0);
and (s1n1018,n31,n1019);
wire s0n1019,s1n1019,notn1019;
or (n1019,s0n1019,s1n1019);
not(notn1019,n639);
and (s0n1019,notn1019,n1020);
and (s1n1019,n639,n1056);
or (n1020,n1021,n1032,n1043,n1054);
and (n1021,n1022,n18);
wire s0n1022,s1n1022,notn1022;
or (n1022,s0n1022,s1n1022);
not(notn1022,n568);
and (s0n1022,notn1022,n1023);
and (s1n1022,n568,n1024);
or (n1024,n1025,n1027,n1029,n1031);
and (n1025,n1026,n594);
and (n1027,n1028,n599);
and (n1029,n1030,n603);
and (n1031,n1023,n605);
and (n1032,n1033,n23);
wire s0n1033,s1n1033,notn1033;
or (n1033,s0n1033,s1n1033);
not(notn1033,n568);
and (s0n1033,notn1033,n1034);
and (s1n1033,n568,n1035);
or (n1035,n1036,n1038,n1040,n1042);
and (n1036,n1037,n594);
and (n1038,n1039,n599);
and (n1040,n1041,n603);
and (n1042,n1034,n605);
and (n1043,n1044,n27);
wire s0n1044,s1n1044,notn1044;
or (n1044,s0n1044,s1n1044);
not(notn1044,n568);
and (s0n1044,notn1044,n1045);
and (s1n1044,n568,n1046);
or (n1046,n1047,n1049,n1051,n1053);
and (n1047,n1048,n594);
and (n1049,n1050,n599);
and (n1051,n1052,n603);
and (n1053,n1045,n605);
and (n1054,n1055,n30);
wire s0n1055,s1n1055,notn1055;
or (n1055,s0n1055,s1n1055);
not(notn1055,n568);
and (s0n1055,notn1055,n1056);
and (s1n1055,n568,n1057);
or (n1057,n1058,n1060,n1062,n1064);
and (n1058,n1059,n594);
and (n1060,n1061,n599);
and (n1062,n1063,n603);
and (n1064,n1056,n605);
or (n1065,n1066,n1146,n1231);
and (n1066,n1067,n1073);
xor (n1067,n1068,n1071);
wire s0n1068,s1n1068,notn1068;
or (n1068,s0n1068,s1n1068);
not(notn1068,n919);
and (s0n1068,notn1068,1'b0);
and (s1n1068,n919,n1069);
xor (n1069,n1070,n861);
xor (n1070,n739,n754);
wire s0n1071,s1n1071,notn1071;
or (n1071,s0n1071,s1n1071);
not(notn1071,n1072);
and (s0n1071,notn1071,1'b0);
and (s1n1071,n1072,n8);
xor (n1072,n920,n968);
and (n1073,n1074,n1076);
wire s0n1074,s1n1074,notn1074;
or (n1074,s0n1074,s1n1074);
not(notn1074,n1075);
and (s0n1074,notn1074,1'b0);
and (s1n1074,n1075,n8);
xor (n1075,n969,n1017);
or (n1076,n1077,n1080,n1145);
and (n1077,n1078,n1079);
wire s0n1078,s1n1078,notn1078;
or (n1078,s0n1078,s1n1078);
not(notn1078,n1075);
and (s0n1078,notn1078,1'b0);
and (s1n1078,n1075,n1069);
wire s0n1079,s1n1079,notn1079;
or (n1079,s0n1079,s1n1079);
not(notn1079,n1018);
and (s0n1079,notn1079,1'b0);
and (s1n1079,n1018,n8);
and (n1080,n1079,n1081);
or (n1081,n1082,n1087,n1144);
and (n1082,n1083,n1086);
wire s0n1083,s1n1083,notn1083;
or (n1083,s0n1083,s1n1083);
not(notn1083,n1075);
and (s0n1083,notn1083,1'b0);
and (s1n1083,n1075,n1084);
xor (n1084,n1085,n868);
xor (n1085,n863,n866);
wire s0n1086,s1n1086,notn1086;
or (n1086,s0n1086,s1n1086);
not(notn1086,n1018);
and (s0n1086,notn1086,1'b0);
and (s1n1086,n1018,n1069);
and (n1087,n1086,n1088);
or (n1088,n1089,n1094,n1143);
and (n1089,n1090,n1093);
wire s0n1090,s1n1090,notn1090;
or (n1090,s0n1090,s1n1090);
not(notn1090,n1075);
and (s0n1090,notn1090,1'b0);
and (s1n1090,n1075,n1091);
xor (n1091,n1092,n876);
xor (n1092,n870,n873);
wire s0n1093,s1n1093,notn1093;
or (n1093,s0n1093,s1n1093);
not(notn1093,n1018);
and (s0n1093,notn1093,1'b0);
and (s1n1093,n1018,n1084);
and (n1094,n1093,n1095);
or (n1095,n1096,n1101,n1142);
and (n1096,n1097,n1100);
wire s0n1097,s1n1097,notn1097;
or (n1097,s0n1097,s1n1097);
not(notn1097,n1075);
and (s0n1097,notn1097,1'b0);
and (s1n1097,n1075,n1098);
xor (n1098,n1099,n884);
xor (n1099,n878,n881);
wire s0n1100,s1n1100,notn1100;
or (n1100,s0n1100,s1n1100);
not(notn1100,n1018);
and (s0n1100,notn1100,1'b0);
and (s1n1100,n1018,n1091);
and (n1101,n1100,n1102);
or (n1102,n1103,n1108,n1141);
and (n1103,n1104,n1107);
wire s0n1104,s1n1104,notn1104;
or (n1104,s0n1104,s1n1104);
not(notn1104,n1075);
and (s0n1104,notn1104,1'b0);
and (s1n1104,n1075,n1105);
xor (n1105,n1106,n892);
xor (n1106,n886,n889);
wire s0n1107,s1n1107,notn1107;
or (n1107,s0n1107,s1n1107);
not(notn1107,n1018);
and (s0n1107,notn1107,1'b0);
and (s1n1107,n1018,n1098);
and (n1108,n1107,n1109);
or (n1109,n1110,n1115,n1140);
and (n1110,n1111,n1114);
wire s0n1111,s1n1111,notn1111;
or (n1111,s0n1111,s1n1111);
not(notn1111,n1075);
and (s0n1111,notn1111,1'b0);
and (s1n1111,n1075,n1112);
xor (n1112,n1113,n900);
xor (n1113,n894,n897);
wire s0n1114,s1n1114,notn1114;
or (n1114,s0n1114,s1n1114);
not(notn1114,n1018);
and (s0n1114,notn1114,1'b0);
and (s1n1114,n1018,n1105);
and (n1115,n1114,n1116);
or (n1116,n1117,n1122,n1139);
and (n1117,n1118,n1121);
wire s0n1118,s1n1118,notn1118;
or (n1118,s0n1118,s1n1118);
not(notn1118,n1075);
and (s0n1118,notn1118,1'b0);
and (s1n1118,n1075,n1119);
xor (n1119,n1120,n908);
xor (n1120,n902,n905);
wire s0n1121,s1n1121,notn1121;
or (n1121,s0n1121,s1n1121);
not(notn1121,n1018);
and (s0n1121,notn1121,1'b0);
and (s1n1121,n1018,n1112);
and (n1122,n1121,n1123);
or (n1123,n1124,n1128,n1130);
and (n1124,n1125,n1127);
wire s0n1125,s1n1125,notn1125;
or (n1125,s0n1125,s1n1125);
not(notn1125,n1075);
and (s0n1125,notn1125,1'b0);
and (s1n1125,n1075,n1126);
xor (n1126,n909,n910);
wire s0n1127,s1n1127,notn1127;
or (n1127,s0n1127,s1n1127);
not(notn1127,n1018);
and (s0n1127,notn1127,1'b0);
and (s1n1127,n1018,n1119);
and (n1128,n1127,n1129);
or (n1129,n1130,n1134,n1135);
and (n1130,n1131,n1133);
wire s0n1131,s1n1131,notn1131;
or (n1131,s0n1131,s1n1131);
not(notn1131,n1075);
and (s0n1131,notn1131,1'b0);
and (s1n1131,n1075,n1132);
xor (n1132,n843,n855);
wire s0n1133,s1n1133,notn1133;
or (n1133,s0n1133,s1n1133);
not(notn1133,n1018);
and (s0n1133,notn1133,1'b0);
and (s1n1133,n1018,n1126);
and (n1134,n1133,n1135);
and (n1135,n1136,n1138);
wire s0n1136,s1n1136,notn1136;
or (n1136,s0n1136,s1n1136);
not(notn1136,n1075);
and (s0n1136,notn1136,1'b0);
and (s1n1136,n1075,n1137);
wire s0n1137,s1n1137,notn1137;
or (n1137,s0n1137,s1n1137);
not(notn1137,n690);
and (s0n1137,notn1137,1'b0);
and (s1n1137,n690,n844);
wire s0n1138,s1n1138,notn1138;
or (n1138,s0n1138,s1n1138);
not(notn1138,n1018);
and (s0n1138,notn1138,1'b0);
and (s1n1138,n1018,n1132);
and (n1139,n1118,n1123);
and (n1140,n1111,n1116);
and (n1141,n1104,n1109);
and (n1142,n1097,n1102);
and (n1143,n1090,n1095);
and (n1144,n1083,n1088);
and (n1145,n1078,n1081);
and (n1146,n1073,n1147);
or (n1147,n1148,n1153,n1230);
and (n1148,n1149,n1152);
xor (n1149,n1150,n1151);
wire s0n1150,s1n1150,notn1150;
or (n1150,s0n1150,s1n1150);
not(notn1150,n919);
and (s0n1150,notn1150,1'b0);
and (s1n1150,n919,n1084);
wire s0n1151,s1n1151,notn1151;
or (n1151,s0n1151,s1n1151);
not(notn1151,n1072);
and (s0n1151,notn1151,1'b0);
and (s1n1151,n1072,n1069);
xor (n1152,n1074,n1076);
and (n1153,n1152,n1154);
or (n1154,n1155,n1161,n1229);
and (n1155,n1156,n1159);
xor (n1156,n1157,n1158);
wire s0n1157,s1n1157,notn1157;
or (n1157,s0n1157,s1n1157);
not(notn1157,n919);
and (s0n1157,notn1157,1'b0);
and (s1n1157,n919,n1091);
wire s0n1158,s1n1158,notn1158;
or (n1158,s0n1158,s1n1158);
not(notn1158,n1072);
and (s0n1158,notn1158,1'b0);
and (s1n1158,n1072,n1084);
xor (n1159,n1160,n1081);
xor (n1160,n1078,n1079);
and (n1161,n1159,n1162);
or (n1162,n1163,n1169,n1228);
and (n1163,n1164,n1167);
xor (n1164,n1165,n1166);
wire s0n1165,s1n1165,notn1165;
or (n1165,s0n1165,s1n1165);
not(notn1165,n919);
and (s0n1165,notn1165,1'b0);
and (s1n1165,n919,n1098);
wire s0n1166,s1n1166,notn1166;
or (n1166,s0n1166,s1n1166);
not(notn1166,n1072);
and (s0n1166,notn1166,1'b0);
and (s1n1166,n1072,n1091);
xor (n1167,n1168,n1088);
xor (n1168,n1083,n1086);
and (n1169,n1167,n1170);
or (n1170,n1171,n1177,n1227);
and (n1171,n1172,n1175);
xor (n1172,n1173,n1174);
wire s0n1173,s1n1173,notn1173;
or (n1173,s0n1173,s1n1173);
not(notn1173,n919);
and (s0n1173,notn1173,1'b0);
and (s1n1173,n919,n1105);
wire s0n1174,s1n1174,notn1174;
or (n1174,s0n1174,s1n1174);
not(notn1174,n1072);
and (s0n1174,notn1174,1'b0);
and (s1n1174,n1072,n1098);
xor (n1175,n1176,n1095);
xor (n1176,n1090,n1093);
and (n1177,n1175,n1178);
or (n1178,n1179,n1185,n1226);
and (n1179,n1180,n1183);
xor (n1180,n1181,n1182);
wire s0n1181,s1n1181,notn1181;
or (n1181,s0n1181,s1n1181);
not(notn1181,n919);
and (s0n1181,notn1181,1'b0);
and (s1n1181,n919,n1112);
wire s0n1182,s1n1182,notn1182;
or (n1182,s0n1182,s1n1182);
not(notn1182,n1072);
and (s0n1182,notn1182,1'b0);
and (s1n1182,n1072,n1105);
xor (n1183,n1184,n1102);
xor (n1184,n1097,n1100);
and (n1185,n1183,n1186);
or (n1186,n1187,n1193,n1225);
and (n1187,n1188,n1191);
xor (n1188,n1189,n1190);
wire s0n1189,s1n1189,notn1189;
or (n1189,s0n1189,s1n1189);
not(notn1189,n919);
and (s0n1189,notn1189,1'b0);
and (s1n1189,n919,n1119);
wire s0n1190,s1n1190,notn1190;
or (n1190,s0n1190,s1n1190);
not(notn1190,n1072);
and (s0n1190,notn1190,1'b0);
and (s1n1190,n1072,n1112);
xor (n1191,n1192,n1109);
xor (n1192,n1104,n1107);
and (n1193,n1191,n1194);
or (n1194,n1195,n1201,n1224);
and (n1195,n1196,n1199);
xor (n1196,n1197,n1198);
wire s0n1197,s1n1197,notn1197;
or (n1197,s0n1197,s1n1197);
not(notn1197,n919);
and (s0n1197,notn1197,1'b0);
and (s1n1197,n919,n1126);
wire s0n1198,s1n1198,notn1198;
or (n1198,s0n1198,s1n1198);
not(notn1198,n1072);
and (s0n1198,notn1198,1'b0);
and (s1n1198,n1072,n1119);
xor (n1199,n1200,n1116);
xor (n1200,n1111,n1114);
and (n1201,n1199,n1202);
or (n1202,n1203,n1209,n1223);
and (n1203,n1204,n1207);
xor (n1204,n1205,n1206);
wire s0n1205,s1n1205,notn1205;
or (n1205,s0n1205,s1n1205);
not(notn1205,n919);
and (s0n1205,notn1205,1'b0);
and (s1n1205,n919,n1132);
wire s0n1206,s1n1206,notn1206;
or (n1206,s0n1206,s1n1206);
not(notn1206,n1072);
and (s0n1206,notn1206,1'b0);
and (s1n1206,n1072,n1126);
xor (n1207,n1208,n1123);
xor (n1208,n1118,n1121);
and (n1209,n1207,n1210);
or (n1210,n1211,n1217,n1222);
and (n1211,n1212,n1215);
xor (n1212,n1213,n1214);
wire s0n1213,s1n1213,notn1213;
or (n1213,s0n1213,s1n1213);
not(notn1213,n919);
and (s0n1213,notn1213,1'b0);
and (s1n1213,n919,n1137);
wire s0n1214,s1n1214,notn1214;
or (n1214,s0n1214,s1n1214);
not(notn1214,n1072);
and (s0n1214,notn1214,1'b0);
and (s1n1214,n1072,n1132);
xor (n1215,n1216,n1129);
xor (n1216,n1125,n1127);
and (n1217,n1215,n1218);
and (n1218,n1219,n1220);
wire s0n1219,s1n1219,notn1219;
or (n1219,s0n1219,s1n1219);
not(notn1219,n1072);
and (s0n1219,notn1219,1'b0);
and (s1n1219,n1072,n1137);
xor (n1220,n1221,n1135);
xor (n1221,n1131,n1133);
and (n1222,n1212,n1218);
and (n1223,n1204,n1210);
and (n1224,n1196,n1202);
and (n1225,n1188,n1194);
and (n1226,n1180,n1186);
and (n1227,n1172,n1178);
and (n1228,n1164,n1170);
and (n1229,n1156,n1162);
and (n1230,n1149,n1154);
and (n1231,n1067,n1147);
xor (n1232,n1233,n1411);
wire s0n1233,s1n1233,notn1233;
or (n1233,s0n1233,s1n1233);
not(notn1233,n919);
and (s0n1233,notn1233,1'b0);
and (s1n1233,n919,n1234);
or (n1234,n1235,n1364,n1410);
and (n1235,n1236,n1248);
wire s0n1236,s1n1236,notn1236;
or (n1236,s0n1236,s1n1236);
not(notn1236,n585);
and (s0n1236,notn1236,1'b0);
and (s1n1236,n585,n1237);
wire s0n1237,s1n1237,notn1237;
or (n1237,s0n1237,s1n1237);
not(notn1237,n566);
and (s0n1237,notn1237,n1238);
and (s1n1237,n566,n1240);
wire s0n1238,s1n1238,notn1238;
or (n1238,s0n1238,s1n1238);
not(notn1238,n13);
and (s0n1238,notn1238,1'b0);
and (s1n1238,n13,n1239);
or (n1240,1'b0,n1241,n1243,n1245,n1247);
and (n1241,n1242,n547);
and (n1243,n1244,n558);
and (n1245,n1246,n562);
and (n1247,n1239,n564);
and (n1248,n1249,n1250);
wire s0n1249,s1n1249,notn1249;
or (n1249,s0n1249,s1n1249);
not(notn1249,n642);
and (s0n1249,notn1249,1'b0);
and (s1n1249,n642,n1237);
or (n1250,n1251,n1265,n1363);
and (n1251,n1252,n1264);
wire s0n1252,s1n1252,notn1252;
or (n1252,s0n1252,s1n1252);
not(notn1252,n642);
and (s0n1252,notn1252,1'b0);
and (s1n1252,n642,n1253);
wire s0n1253,s1n1253,notn1253;
or (n1253,s0n1253,s1n1253);
not(notn1253,n566);
and (s0n1253,notn1253,n1254);
and (s1n1253,n566,n1256);
wire s0n1254,s1n1254,notn1254;
or (n1254,s0n1254,s1n1254);
not(notn1254,n13);
and (s0n1254,notn1254,1'b0);
and (s1n1254,n13,n1255);
or (n1256,1'b0,n1257,n1259,n1261,n1263);
and (n1257,n1258,n547);
and (n1259,n1260,n558);
and (n1261,n1262,n562);
and (n1263,n1255,n564);
wire s0n1264,s1n1264,notn1264;
or (n1264,s0n1264,s1n1264);
not(notn1264,n690);
and (s0n1264,notn1264,1'b0);
and (s1n1264,n690,n1237);
and (n1265,n1264,n1266);
or (n1266,n1267,n1281,n1362);
and (n1267,n1268,n1280);
wire s0n1268,s1n1268,notn1268;
or (n1268,s0n1268,s1n1268);
not(notn1268,n642);
and (s0n1268,notn1268,1'b0);
and (s1n1268,n642,n1269);
wire s0n1269,s1n1269,notn1269;
or (n1269,s0n1269,s1n1269);
not(notn1269,n566);
and (s0n1269,notn1269,n1270);
and (s1n1269,n566,n1272);
wire s0n1270,s1n1270,notn1270;
or (n1270,s0n1270,s1n1270);
not(notn1270,n13);
and (s0n1270,notn1270,1'b0);
and (s1n1270,n13,n1271);
or (n1272,1'b0,n1273,n1275,n1277,n1279);
and (n1273,n1274,n547);
and (n1275,n1276,n558);
and (n1277,n1278,n562);
and (n1279,n1271,n564);
wire s0n1280,s1n1280,notn1280;
or (n1280,s0n1280,s1n1280);
not(notn1280,n690);
and (s0n1280,notn1280,1'b0);
and (s1n1280,n690,n1253);
and (n1281,n1280,n1282);
or (n1282,n1283,n1297,n1361);
and (n1283,n1284,n1296);
wire s0n1284,s1n1284,notn1284;
or (n1284,s0n1284,s1n1284);
not(notn1284,n642);
and (s0n1284,notn1284,1'b0);
and (s1n1284,n642,n1285);
wire s0n1285,s1n1285,notn1285;
or (n1285,s0n1285,s1n1285);
not(notn1285,n566);
and (s0n1285,notn1285,n1286);
and (s1n1285,n566,n1288);
wire s0n1286,s1n1286,notn1286;
or (n1286,s0n1286,s1n1286);
not(notn1286,n13);
and (s0n1286,notn1286,1'b0);
and (s1n1286,n13,n1287);
or (n1288,1'b0,n1289,n1291,n1293,n1295);
and (n1289,n1290,n547);
and (n1291,n1292,n558);
and (n1293,n1294,n562);
and (n1295,n1287,n564);
wire s0n1296,s1n1296,notn1296;
or (n1296,s0n1296,s1n1296);
not(notn1296,n690);
and (s0n1296,notn1296,1'b0);
and (s1n1296,n690,n1269);
and (n1297,n1296,n1298);
or (n1298,n1299,n1313,n1360);
and (n1299,n1300,n1312);
wire s0n1300,s1n1300,notn1300;
or (n1300,s0n1300,s1n1300);
not(notn1300,n642);
and (s0n1300,notn1300,1'b0);
and (s1n1300,n642,n1301);
wire s0n1301,s1n1301,notn1301;
or (n1301,s0n1301,s1n1301);
not(notn1301,n566);
and (s0n1301,notn1301,n1302);
and (s1n1301,n566,n1304);
wire s0n1302,s1n1302,notn1302;
or (n1302,s0n1302,s1n1302);
not(notn1302,n13);
and (s0n1302,notn1302,1'b0);
and (s1n1302,n13,n1303);
or (n1304,1'b0,n1305,n1307,n1309,n1311);
and (n1305,n1306,n547);
and (n1307,n1308,n558);
and (n1309,n1310,n562);
and (n1311,n1303,n564);
wire s0n1312,s1n1312,notn1312;
or (n1312,s0n1312,s1n1312);
not(notn1312,n690);
and (s0n1312,notn1312,1'b0);
and (s1n1312,n690,n1285);
and (n1313,n1312,n1314);
or (n1314,n1315,n1329,n1331);
and (n1315,n1316,n1328);
wire s0n1316,s1n1316,notn1316;
or (n1316,s0n1316,s1n1316);
not(notn1316,n642);
and (s0n1316,notn1316,1'b0);
and (s1n1316,n642,n1317);
wire s0n1317,s1n1317,notn1317;
or (n1317,s0n1317,s1n1317);
not(notn1317,n566);
and (s0n1317,notn1317,n1318);
and (s1n1317,n566,n1320);
wire s0n1318,s1n1318,notn1318;
or (n1318,s0n1318,s1n1318);
not(notn1318,n13);
and (s0n1318,notn1318,1'b0);
and (s1n1318,n13,n1319);
or (n1320,1'b0,n1321,n1323,n1325,n1327);
and (n1321,n1322,n547);
and (n1323,n1324,n558);
and (n1325,n1326,n562);
and (n1327,n1319,n564);
wire s0n1328,s1n1328,notn1328;
or (n1328,s0n1328,s1n1328);
not(notn1328,n690);
and (s0n1328,notn1328,1'b0);
and (s1n1328,n690,n1301);
and (n1329,n1328,n1330);
or (n1330,n1331,n1345,n1346);
and (n1331,n1332,n1344);
wire s0n1332,s1n1332,notn1332;
or (n1332,s0n1332,s1n1332);
not(notn1332,n642);
and (s0n1332,notn1332,1'b0);
and (s1n1332,n642,n1333);
wire s0n1333,s1n1333,notn1333;
or (n1333,s0n1333,s1n1333);
not(notn1333,n566);
and (s0n1333,notn1333,n1334);
and (s1n1333,n566,n1336);
wire s0n1334,s1n1334,notn1334;
or (n1334,s0n1334,s1n1334);
not(notn1334,n13);
and (s0n1334,notn1334,1'b0);
and (s1n1334,n13,n1335);
or (n1336,1'b0,n1337,n1339,n1341,n1343);
and (n1337,n1338,n547);
and (n1339,n1340,n558);
and (n1341,n1342,n562);
and (n1343,n1335,n564);
wire s0n1344,s1n1344,notn1344;
or (n1344,s0n1344,s1n1344);
not(notn1344,n690);
and (s0n1344,notn1344,1'b0);
and (s1n1344,n690,n1317);
and (n1345,n1344,n1346);
and (n1346,n1347,n1359);
wire s0n1347,s1n1347,notn1347;
or (n1347,s0n1347,s1n1347);
not(notn1347,n642);
and (s0n1347,notn1347,1'b0);
and (s1n1347,n642,n1348);
wire s0n1348,s1n1348,notn1348;
or (n1348,s0n1348,s1n1348);
not(notn1348,n566);
and (s0n1348,notn1348,n1349);
and (s1n1348,n566,n1351);
wire s0n1349,s1n1349,notn1349;
or (n1349,s0n1349,s1n1349);
not(notn1349,n13);
and (s0n1349,notn1349,1'b0);
and (s1n1349,n13,n1350);
or (n1351,1'b0,n1352,n1354,n1356,n1358);
and (n1352,n1353,n547);
and (n1354,n1355,n558);
and (n1356,n1357,n562);
and (n1358,n1350,n564);
wire s0n1359,s1n1359,notn1359;
or (n1359,s0n1359,s1n1359);
not(notn1359,n690);
and (s0n1359,notn1359,1'b0);
and (s1n1359,n690,n1333);
and (n1360,n1300,n1314);
and (n1361,n1284,n1298);
and (n1362,n1268,n1282);
and (n1363,n1252,n1266);
and (n1364,n1248,n1365);
or (n1365,n1366,n1369,n1409);
and (n1366,n1367,n1368);
wire s0n1367,s1n1367,notn1367;
or (n1367,s0n1367,s1n1367);
not(notn1367,n585);
and (s0n1367,notn1367,1'b0);
and (s1n1367,n585,n1253);
xor (n1368,n1249,n1250);
and (n1369,n1368,n1370);
or (n1370,n1371,n1375,n1408);
and (n1371,n1372,n1373);
wire s0n1372,s1n1372,notn1372;
or (n1372,s0n1372,s1n1372);
not(notn1372,n585);
and (s0n1372,notn1372,1'b0);
and (s1n1372,n585,n1269);
xor (n1373,n1374,n1266);
xor (n1374,n1252,n1264);
and (n1375,n1373,n1376);
or (n1376,n1377,n1381,n1407);
and (n1377,n1378,n1379);
wire s0n1378,s1n1378,notn1378;
or (n1378,s0n1378,s1n1378);
not(notn1378,n585);
and (s0n1378,notn1378,1'b0);
and (s1n1378,n585,n1285);
xor (n1379,n1380,n1282);
xor (n1380,n1268,n1280);
and (n1381,n1379,n1382);
or (n1382,n1383,n1387,n1406);
and (n1383,n1384,n1385);
wire s0n1384,s1n1384,notn1384;
or (n1384,s0n1384,s1n1384);
not(notn1384,n585);
and (s0n1384,notn1384,1'b0);
and (s1n1384,n585,n1301);
xor (n1385,n1386,n1298);
xor (n1386,n1284,n1296);
and (n1387,n1385,n1388);
or (n1388,n1389,n1393,n1405);
and (n1389,n1390,n1391);
wire s0n1390,s1n1390,notn1390;
or (n1390,s0n1390,s1n1390);
not(notn1390,n585);
and (s0n1390,notn1390,1'b0);
and (s1n1390,n585,n1317);
xor (n1391,n1392,n1314);
xor (n1392,n1300,n1312);
and (n1393,n1391,n1394);
or (n1394,n1395,n1399,n1404);
and (n1395,n1396,n1397);
wire s0n1396,s1n1396,notn1396;
or (n1396,s0n1396,s1n1396);
not(notn1396,n585);
and (s0n1396,notn1396,1'b0);
and (s1n1396,n585,n1333);
xor (n1397,n1398,n1330);
xor (n1398,n1316,n1328);
and (n1399,n1397,n1400);
and (n1400,n1401,n1402);
wire s0n1401,s1n1401,notn1401;
or (n1401,s0n1401,s1n1401);
not(notn1401,n585);
and (s0n1401,notn1401,1'b0);
and (s1n1401,n585,n1348);
xor (n1402,n1403,n1346);
xor (n1403,n1332,n1344);
and (n1404,n1396,n1400);
and (n1405,n1390,n1394);
and (n1406,n1384,n1388);
and (n1407,n1378,n1382);
and (n1408,n1372,n1376);
and (n1409,n1367,n1370);
and (n1410,n1236,n1365);
or (n1411,n1412,n1491,n1576);
and (n1412,n1413,n1418);
xor (n1413,n1414,n1417);
wire s0n1414,s1n1414,notn1414;
or (n1414,s0n1414,s1n1414);
not(notn1414,n919);
and (s0n1414,notn1414,1'b0);
and (s1n1414,n919,n1415);
xor (n1415,n1416,n1365);
xor (n1416,n1236,n1248);
wire s0n1417,s1n1417,notn1417;
or (n1417,s0n1417,s1n1417);
not(notn1417,n1072);
and (s0n1417,notn1417,1'b0);
and (s1n1417,n1072,n1234);
and (n1418,n1419,n1420);
wire s0n1419,s1n1419,notn1419;
or (n1419,s0n1419,s1n1419);
not(notn1419,n1075);
and (s0n1419,notn1419,1'b0);
and (s1n1419,n1075,n1234);
or (n1420,n1421,n1424,n1490);
and (n1421,n1422,n1423);
wire s0n1422,s1n1422,notn1422;
or (n1422,s0n1422,s1n1422);
not(notn1422,n1075);
and (s0n1422,notn1422,1'b0);
and (s1n1422,n1075,n1415);
wire s0n1423,s1n1423,notn1423;
or (n1423,s0n1423,s1n1423);
not(notn1423,n1018);
and (s0n1423,notn1423,1'b0);
and (s1n1423,n1018,n1234);
and (n1424,n1423,n1425);
or (n1425,n1426,n1431,n1489);
and (n1426,n1427,n1430);
wire s0n1427,s1n1427,notn1427;
or (n1427,s0n1427,s1n1427);
not(notn1427,n1075);
and (s0n1427,notn1427,1'b0);
and (s1n1427,n1075,n1428);
xor (n1428,n1429,n1370);
xor (n1429,n1367,n1368);
wire s0n1430,s1n1430,notn1430;
or (n1430,s0n1430,s1n1430);
not(notn1430,n1018);
and (s0n1430,notn1430,1'b0);
and (s1n1430,n1018,n1415);
and (n1431,n1430,n1432);
or (n1432,n1433,n1438,n1488);
and (n1433,n1434,n1437);
wire s0n1434,s1n1434,notn1434;
or (n1434,s0n1434,s1n1434);
not(notn1434,n1075);
and (s0n1434,notn1434,1'b0);
and (s1n1434,n1075,n1435);
xor (n1435,n1436,n1376);
xor (n1436,n1372,n1373);
wire s0n1437,s1n1437,notn1437;
or (n1437,s0n1437,s1n1437);
not(notn1437,n1018);
and (s0n1437,notn1437,1'b0);
and (s1n1437,n1018,n1428);
and (n1438,n1437,n1439);
or (n1439,n1440,n1445,n1487);
and (n1440,n1441,n1444);
wire s0n1441,s1n1441,notn1441;
or (n1441,s0n1441,s1n1441);
not(notn1441,n1075);
and (s0n1441,notn1441,1'b0);
and (s1n1441,n1075,n1442);
xor (n1442,n1443,n1382);
xor (n1443,n1378,n1379);
wire s0n1444,s1n1444,notn1444;
or (n1444,s0n1444,s1n1444);
not(notn1444,n1018);
and (s0n1444,notn1444,1'b0);
and (s1n1444,n1018,n1435);
and (n1445,n1444,n1446);
or (n1446,n1447,n1452,n1486);
and (n1447,n1448,n1451);
wire s0n1448,s1n1448,notn1448;
or (n1448,s0n1448,s1n1448);
not(notn1448,n1075);
and (s0n1448,notn1448,1'b0);
and (s1n1448,n1075,n1449);
xor (n1449,n1450,n1388);
xor (n1450,n1384,n1385);
wire s0n1451,s1n1451,notn1451;
or (n1451,s0n1451,s1n1451);
not(notn1451,n1018);
and (s0n1451,notn1451,1'b0);
and (s1n1451,n1018,n1442);
and (n1452,n1451,n1453);
or (n1453,n1454,n1459,n1485);
and (n1454,n1455,n1458);
wire s0n1455,s1n1455,notn1455;
or (n1455,s0n1455,s1n1455);
not(notn1455,n1075);
and (s0n1455,notn1455,1'b0);
and (s1n1455,n1075,n1456);
xor (n1456,n1457,n1394);
xor (n1457,n1390,n1391);
wire s0n1458,s1n1458,notn1458;
or (n1458,s0n1458,s1n1458);
not(notn1458,n1018);
and (s0n1458,notn1458,1'b0);
and (s1n1458,n1018,n1449);
and (n1459,n1458,n1460);
or (n1460,n1461,n1466,n1484);
and (n1461,n1462,n1465);
wire s0n1462,s1n1462,notn1462;
or (n1462,s0n1462,s1n1462);
not(notn1462,n1075);
and (s0n1462,notn1462,1'b0);
and (s1n1462,n1075,n1463);
xor (n1463,n1464,n1400);
xor (n1464,n1396,n1397);
wire s0n1465,s1n1465,notn1465;
or (n1465,s0n1465,s1n1465);
not(notn1465,n1018);
and (s0n1465,notn1465,1'b0);
and (s1n1465,n1018,n1456);
and (n1466,n1465,n1467);
or (n1467,n1468,n1472,n1474);
and (n1468,n1469,n1471);
wire s0n1469,s1n1469,notn1469;
or (n1469,s0n1469,s1n1469);
not(notn1469,n1075);
and (s0n1469,notn1469,1'b0);
and (s1n1469,n1075,n1470);
xor (n1470,n1401,n1402);
wire s0n1471,s1n1471,notn1471;
or (n1471,s0n1471,s1n1471);
not(notn1471,n1018);
and (s0n1471,notn1471,1'b0);
and (s1n1471,n1018,n1463);
and (n1472,n1471,n1473);
or (n1473,n1474,n1478,n1479);
and (n1474,n1475,n1477);
wire s0n1475,s1n1475,notn1475;
or (n1475,s0n1475,s1n1475);
not(notn1475,n1075);
and (s0n1475,notn1475,1'b0);
and (s1n1475,n1075,n1476);
xor (n1476,n1347,n1359);
wire s0n1477,s1n1477,notn1477;
or (n1477,s0n1477,s1n1477);
not(notn1477,n1018);
and (s0n1477,notn1477,1'b0);
and (s1n1477,n1018,n1470);
and (n1478,n1477,n1479);
and (n1479,n1480,n1483);
wire s0n1480,s1n1480,notn1480;
or (n1480,s0n1480,s1n1480);
not(notn1480,n1075);
and (s0n1480,notn1480,1'b0);
and (s1n1480,n1075,n1481);
not (n1481,n1482);
nand (n1482,n690,n1348);
wire s0n1483,s1n1483,notn1483;
or (n1483,s0n1483,s1n1483);
not(notn1483,n1018);
and (s0n1483,notn1483,1'b0);
and (s1n1483,n1018,n1476);
and (n1484,n1462,n1467);
and (n1485,n1455,n1460);
and (n1486,n1448,n1453);
and (n1487,n1441,n1446);
and (n1488,n1434,n1439);
and (n1489,n1427,n1432);
and (n1490,n1422,n1425);
and (n1491,n1418,n1492);
or (n1492,n1493,n1498,n1575);
and (n1493,n1494,n1497);
xor (n1494,n1495,n1496);
wire s0n1495,s1n1495,notn1495;
or (n1495,s0n1495,s1n1495);
not(notn1495,n919);
and (s0n1495,notn1495,1'b0);
and (s1n1495,n919,n1428);
wire s0n1496,s1n1496,notn1496;
or (n1496,s0n1496,s1n1496);
not(notn1496,n1072);
and (s0n1496,notn1496,1'b0);
and (s1n1496,n1072,n1415);
xor (n1497,n1419,n1420);
and (n1498,n1497,n1499);
or (n1499,n1500,n1506,n1574);
and (n1500,n1501,n1504);
xor (n1501,n1502,n1503);
wire s0n1502,s1n1502,notn1502;
or (n1502,s0n1502,s1n1502);
not(notn1502,n919);
and (s0n1502,notn1502,1'b0);
and (s1n1502,n919,n1435);
wire s0n1503,s1n1503,notn1503;
or (n1503,s0n1503,s1n1503);
not(notn1503,n1072);
and (s0n1503,notn1503,1'b0);
and (s1n1503,n1072,n1428);
xor (n1504,n1505,n1425);
xor (n1505,n1422,n1423);
and (n1506,n1504,n1507);
or (n1507,n1508,n1514,n1573);
and (n1508,n1509,n1512);
xor (n1509,n1510,n1511);
wire s0n1510,s1n1510,notn1510;
or (n1510,s0n1510,s1n1510);
not(notn1510,n919);
and (s0n1510,notn1510,1'b0);
and (s1n1510,n919,n1442);
wire s0n1511,s1n1511,notn1511;
or (n1511,s0n1511,s1n1511);
not(notn1511,n1072);
and (s0n1511,notn1511,1'b0);
and (s1n1511,n1072,n1435);
xor (n1512,n1513,n1432);
xor (n1513,n1427,n1430);
and (n1514,n1512,n1515);
or (n1515,n1516,n1522,n1572);
and (n1516,n1517,n1520);
xor (n1517,n1518,n1519);
wire s0n1518,s1n1518,notn1518;
or (n1518,s0n1518,s1n1518);
not(notn1518,n919);
and (s0n1518,notn1518,1'b0);
and (s1n1518,n919,n1449);
wire s0n1519,s1n1519,notn1519;
or (n1519,s0n1519,s1n1519);
not(notn1519,n1072);
and (s0n1519,notn1519,1'b0);
and (s1n1519,n1072,n1442);
xor (n1520,n1521,n1439);
xor (n1521,n1434,n1437);
and (n1522,n1520,n1523);
or (n1523,n1524,n1530,n1571);
and (n1524,n1525,n1528);
xor (n1525,n1526,n1527);
wire s0n1526,s1n1526,notn1526;
or (n1526,s0n1526,s1n1526);
not(notn1526,n919);
and (s0n1526,notn1526,1'b0);
and (s1n1526,n919,n1456);
wire s0n1527,s1n1527,notn1527;
or (n1527,s0n1527,s1n1527);
not(notn1527,n1072);
and (s0n1527,notn1527,1'b0);
and (s1n1527,n1072,n1449);
xor (n1528,n1529,n1446);
xor (n1529,n1441,n1444);
and (n1530,n1528,n1531);
or (n1531,n1532,n1538,n1570);
and (n1532,n1533,n1536);
xor (n1533,n1534,n1535);
wire s0n1534,s1n1534,notn1534;
or (n1534,s0n1534,s1n1534);
not(notn1534,n919);
and (s0n1534,notn1534,1'b0);
and (s1n1534,n919,n1463);
wire s0n1535,s1n1535,notn1535;
or (n1535,s0n1535,s1n1535);
not(notn1535,n1072);
and (s0n1535,notn1535,1'b0);
and (s1n1535,n1072,n1456);
xor (n1536,n1537,n1453);
xor (n1537,n1448,n1451);
and (n1538,n1536,n1539);
or (n1539,n1540,n1546,n1569);
and (n1540,n1541,n1544);
xor (n1541,n1542,n1543);
wire s0n1542,s1n1542,notn1542;
or (n1542,s0n1542,s1n1542);
not(notn1542,n919);
and (s0n1542,notn1542,1'b0);
and (s1n1542,n919,n1470);
wire s0n1543,s1n1543,notn1543;
or (n1543,s0n1543,s1n1543);
not(notn1543,n1072);
and (s0n1543,notn1543,1'b0);
and (s1n1543,n1072,n1463);
xor (n1544,n1545,n1460);
xor (n1545,n1455,n1458);
and (n1546,n1544,n1547);
or (n1547,n1548,n1554,n1568);
and (n1548,n1549,n1552);
xor (n1549,n1550,n1551);
wire s0n1550,s1n1550,notn1550;
or (n1550,s0n1550,s1n1550);
not(notn1550,n919);
and (s0n1550,notn1550,1'b0);
and (s1n1550,n919,n1476);
wire s0n1551,s1n1551,notn1551;
or (n1551,s0n1551,s1n1551);
not(notn1551,n1072);
and (s0n1551,notn1551,1'b0);
and (s1n1551,n1072,n1470);
xor (n1552,n1553,n1467);
xor (n1553,n1462,n1465);
and (n1554,n1552,n1555);
or (n1555,n1556,n1562,n1567);
and (n1556,n1557,n1560);
xor (n1557,n1558,n1559);
wire s0n1558,s1n1558,notn1558;
or (n1558,s0n1558,s1n1558);
not(notn1558,n919);
and (s0n1558,notn1558,1'b0);
and (s1n1558,n919,n1481);
wire s0n1559,s1n1559,notn1559;
or (n1559,s0n1559,s1n1559);
not(notn1559,n1072);
and (s0n1559,notn1559,1'b0);
and (s1n1559,n1072,n1476);
xor (n1560,n1561,n1473);
xor (n1561,n1469,n1471);
and (n1562,n1560,n1563);
and (n1563,n1564,n1565);
wire s0n1564,s1n1564,notn1564;
or (n1564,s0n1564,s1n1564);
not(notn1564,n1072);
and (s0n1564,notn1564,1'b0);
and (s1n1564,n1072,n1481);
xor (n1565,n1566,n1479);
xor (n1566,n1475,n1477);
and (n1567,n1557,n1563);
and (n1568,n1549,n1555);
and (n1569,n1541,n1547);
and (n1570,n1533,n1539);
and (n1571,n1525,n1531);
and (n1572,n1517,n1523);
and (n1573,n1509,n1515);
and (n1574,n1501,n1507);
and (n1575,n1494,n1499);
and (n1576,n1413,n1492);
or (n1577,n1578,n1583,n1671);
and (n1578,n1579,n1581);
xor (n1579,n1580,n1147);
xor (n1580,n1067,n1073);
xor (n1581,n1582,n1492);
xor (n1582,n1413,n1418);
and (n1583,n1581,n1584);
or (n1584,n1585,n1590,n1670);
and (n1585,n1586,n1588);
xor (n1586,n1587,n1154);
xor (n1587,n1149,n1152);
xor (n1588,n1589,n1499);
xor (n1589,n1494,n1497);
and (n1590,n1588,n1591);
or (n1591,n1592,n1597,n1669);
and (n1592,n1593,n1595);
xor (n1593,n1594,n1162);
xor (n1594,n1156,n1159);
xor (n1595,n1596,n1507);
xor (n1596,n1501,n1504);
and (n1597,n1595,n1598);
or (n1598,n1599,n1604,n1668);
and (n1599,n1600,n1602);
xor (n1600,n1601,n1170);
xor (n1601,n1164,n1167);
xor (n1602,n1603,n1515);
xor (n1603,n1509,n1512);
and (n1604,n1602,n1605);
or (n1605,n1606,n1611,n1667);
and (n1606,n1607,n1609);
xor (n1607,n1608,n1178);
xor (n1608,n1172,n1175);
xor (n1609,n1610,n1523);
xor (n1610,n1517,n1520);
and (n1611,n1609,n1612);
or (n1612,n1613,n1618,n1666);
and (n1613,n1614,n1616);
xor (n1614,n1615,n1186);
xor (n1615,n1180,n1183);
xor (n1616,n1617,n1531);
xor (n1617,n1525,n1528);
and (n1618,n1616,n1619);
or (n1619,n1620,n1625,n1665);
and (n1620,n1621,n1623);
xor (n1621,n1622,n1194);
xor (n1622,n1188,n1191);
xor (n1623,n1624,n1539);
xor (n1624,n1533,n1536);
and (n1625,n1623,n1626);
or (n1626,n1627,n1632,n1664);
and (n1627,n1628,n1630);
xor (n1628,n1629,n1202);
xor (n1629,n1196,n1199);
xor (n1630,n1631,n1547);
xor (n1631,n1541,n1544);
and (n1632,n1630,n1633);
or (n1633,n1634,n1639,n1663);
and (n1634,n1635,n1637);
xor (n1635,n1636,n1210);
xor (n1636,n1204,n1207);
xor (n1637,n1638,n1555);
xor (n1638,n1549,n1552);
and (n1639,n1637,n1640);
or (n1640,n1641,n1646,n1662);
and (n1641,n1642,n1644);
xor (n1642,n1643,n1218);
xor (n1643,n1212,n1215);
xor (n1644,n1645,n1563);
xor (n1645,n1557,n1560);
and (n1646,n1644,n1647);
or (n1647,n1648,n1651,n1661);
and (n1648,n1649,n1650);
xor (n1649,n1219,n1220);
xor (n1650,n1564,n1565);
and (n1651,n1650,n1652);
or (n1652,n1653,n1656,n1660);
and (n1653,n1654,n1655);
xor (n1654,n1136,n1138);
xor (n1655,n1480,n1483);
and (n1656,n1655,n1657);
and (n1657,n1658,n1659);
wire s0n1658,s1n1658,notn1658;
or (n1658,s0n1658,s1n1658);
not(notn1658,n1018);
and (s0n1658,notn1658,1'b0);
and (s1n1658,n1018,n1137);
wire s0n1659,s1n1659,notn1659;
or (n1659,s0n1659,s1n1659);
not(notn1659,n1018);
and (s0n1659,notn1659,1'b0);
and (s1n1659,n1018,n1481);
and (n1660,n1654,n1657);
and (n1661,n1649,n1652);
and (n1662,n1642,n1647);
and (n1663,n1635,n1640);
and (n1664,n1628,n1633);
and (n1665,n1621,n1626);
and (n1666,n1614,n1619);
and (n1667,n1607,n1612);
and (n1668,n1600,n1605);
and (n1669,n1593,n1598);
and (n1670,n1586,n1591);
and (n1671,n1579,n1584);
xor (n1672,n1673,n2334);
xor (n1673,n1674,n2012);
or (n1674,n1675,n1944,n2011);
and (n1675,n1676,n1870);
wire s0n1676,s1n1676,notn1676;
or (n1676,s0n1676,s1n1676);
not(notn1676,n921);
and (s0n1676,notn1676,1'b0);
and (s1n1676,n921,n1677);
xor (n1677,n1678,n1690);
wire s0n1678,s1n1678,notn1678;
or (n1678,s0n1678,s1n1678);
not(notn1678,n583);
and (s0n1678,notn1678,1'b0);
and (s1n1678,n583,n1679);
wire s0n1679,s1n1679,notn1679;
or (n1679,s0n1679,s1n1679);
not(notn1679,n566);
and (s0n1679,notn1679,n1680);
and (s1n1679,n566,n1682);
wire s0n1680,s1n1680,notn1680;
or (n1680,s0n1680,s1n1680);
not(notn1680,n13);
and (s0n1680,notn1680,1'b0);
and (s1n1680,n13,n1681);
or (n1682,1'b0,n1683,n1685,n1687,n1689);
and (n1683,n1684,n547);
and (n1685,n1686,n558);
and (n1687,n1688,n562);
and (n1689,n1681,n564);
or (n1690,n1691,n1811,n1869);
and (n1691,n1692,n1706);
xor (n1692,n1693,n1705);
wire s0n1693,s1n1693,notn1693;
or (n1693,s0n1693,s1n1693);
not(notn1693,n583);
and (s0n1693,notn1693,1'b0);
and (s1n1693,n583,n1694);
wire s0n1694,s1n1694,notn1694;
or (n1694,s0n1694,s1n1694);
not(notn1694,n566);
and (s0n1694,notn1694,n1695);
and (s1n1694,n566,n1697);
wire s0n1695,s1n1695,notn1695;
or (n1695,s0n1695,s1n1695);
not(notn1695,n13);
and (s0n1695,notn1695,1'b0);
and (s1n1695,n13,n1696);
or (n1697,1'b0,n1698,n1700,n1702,n1704);
and (n1698,n1699,n547);
and (n1700,n1701,n558);
and (n1702,n1703,n562);
and (n1704,n1696,n564);
wire s0n1705,s1n1705,notn1705;
or (n1705,s0n1705,s1n1705);
not(notn1705,n753);
and (s0n1705,notn1705,1'b0);
and (s1n1705,n753,n1679);
and (n1706,n1707,n1708);
wire s0n1707,s1n1707,notn1707;
or (n1707,s0n1707,s1n1707);
not(notn1707,n756);
and (s0n1707,notn1707,1'b0);
and (s1n1707,n756,n1679);
or (n1708,n1709,n1712,n1810);
and (n1709,n1710,n1711);
wire s0n1710,s1n1710,notn1710;
or (n1710,s0n1710,s1n1710);
not(notn1710,n756);
and (s0n1710,notn1710,1'b0);
and (s1n1710,n756,n1694);
wire s0n1711,s1n1711,notn1711;
or (n1711,s0n1711,s1n1711);
not(notn1711,n690);
and (s0n1711,notn1711,1'b0);
and (s1n1711,n690,n1679);
and (n1712,n1711,n1713);
or (n1713,n1714,n1728,n1809);
and (n1714,n1715,n1727);
wire s0n1715,s1n1715,notn1715;
or (n1715,s0n1715,s1n1715);
not(notn1715,n756);
and (s0n1715,notn1715,1'b0);
and (s1n1715,n756,n1716);
wire s0n1716,s1n1716,notn1716;
or (n1716,s0n1716,s1n1716);
not(notn1716,n566);
and (s0n1716,notn1716,n1717);
and (s1n1716,n566,n1719);
wire s0n1717,s1n1717,notn1717;
or (n1717,s0n1717,s1n1717);
not(notn1717,n13);
and (s0n1717,notn1717,1'b0);
and (s1n1717,n13,n1718);
or (n1719,1'b0,n1720,n1722,n1724,n1726);
and (n1720,n1721,n547);
and (n1722,n1723,n558);
and (n1724,n1725,n562);
and (n1726,n1718,n564);
wire s0n1727,s1n1727,notn1727;
or (n1727,s0n1727,s1n1727);
not(notn1727,n690);
and (s0n1727,notn1727,1'b0);
and (s1n1727,n690,n1694);
and (n1728,n1727,n1729);
or (n1729,n1730,n1744,n1808);
and (n1730,n1731,n1743);
wire s0n1731,s1n1731,notn1731;
or (n1731,s0n1731,s1n1731);
not(notn1731,n756);
and (s0n1731,notn1731,1'b0);
and (s1n1731,n756,n1732);
wire s0n1732,s1n1732,notn1732;
or (n1732,s0n1732,s1n1732);
not(notn1732,n566);
and (s0n1732,notn1732,n1733);
and (s1n1732,n566,n1735);
wire s0n1733,s1n1733,notn1733;
or (n1733,s0n1733,s1n1733);
not(notn1733,n13);
and (s0n1733,notn1733,1'b0);
and (s1n1733,n13,n1734);
or (n1735,1'b0,n1736,n1738,n1740,n1742);
and (n1736,n1737,n547);
and (n1738,n1739,n558);
and (n1740,n1741,n562);
and (n1742,n1734,n564);
wire s0n1743,s1n1743,notn1743;
or (n1743,s0n1743,s1n1743);
not(notn1743,n690);
and (s0n1743,notn1743,1'b0);
and (s1n1743,n690,n1716);
and (n1744,n1743,n1745);
or (n1745,n1746,n1760,n1807);
and (n1746,n1747,n1759);
wire s0n1747,s1n1747,notn1747;
or (n1747,s0n1747,s1n1747);
not(notn1747,n756);
and (s0n1747,notn1747,1'b0);
and (s1n1747,n756,n1748);
wire s0n1748,s1n1748,notn1748;
or (n1748,s0n1748,s1n1748);
not(notn1748,n566);
and (s0n1748,notn1748,n1749);
and (s1n1748,n566,n1751);
wire s0n1749,s1n1749,notn1749;
or (n1749,s0n1749,s1n1749);
not(notn1749,n13);
and (s0n1749,notn1749,1'b0);
and (s1n1749,n13,n1750);
or (n1751,1'b0,n1752,n1754,n1756,n1758);
and (n1752,n1753,n547);
and (n1754,n1755,n558);
and (n1756,n1757,n562);
and (n1758,n1750,n564);
wire s0n1759,s1n1759,notn1759;
or (n1759,s0n1759,s1n1759);
not(notn1759,n690);
and (s0n1759,notn1759,1'b0);
and (s1n1759,n690,n1732);
and (n1760,n1759,n1761);
or (n1761,n1762,n1776,n1778);
and (n1762,n1763,n1775);
wire s0n1763,s1n1763,notn1763;
or (n1763,s0n1763,s1n1763);
not(notn1763,n756);
and (s0n1763,notn1763,1'b0);
and (s1n1763,n756,n1764);
wire s0n1764,s1n1764,notn1764;
or (n1764,s0n1764,s1n1764);
not(notn1764,n566);
and (s0n1764,notn1764,n1765);
and (s1n1764,n566,n1767);
wire s0n1765,s1n1765,notn1765;
or (n1765,s0n1765,s1n1765);
not(notn1765,n13);
and (s0n1765,notn1765,1'b0);
and (s1n1765,n13,n1766);
or (n1767,1'b0,n1768,n1770,n1772,n1774);
and (n1768,n1769,n547);
and (n1770,n1771,n558);
and (n1772,n1773,n562);
and (n1774,n1766,n564);
wire s0n1775,s1n1775,notn1775;
or (n1775,s0n1775,s1n1775);
not(notn1775,n690);
and (s0n1775,notn1775,1'b0);
and (s1n1775,n690,n1748);
and (n1776,n1775,n1777);
or (n1777,n1778,n1792,n1793);
and (n1778,n1779,n1791);
wire s0n1779,s1n1779,notn1779;
or (n1779,s0n1779,s1n1779);
not(notn1779,n756);
and (s0n1779,notn1779,1'b0);
and (s1n1779,n756,n1780);
wire s0n1780,s1n1780,notn1780;
or (n1780,s0n1780,s1n1780);
not(notn1780,n566);
and (s0n1780,notn1780,n1781);
and (s1n1780,n566,n1783);
wire s0n1781,s1n1781,notn1781;
or (n1781,s0n1781,s1n1781);
not(notn1781,n13);
and (s0n1781,notn1781,1'b0);
and (s1n1781,n13,n1782);
or (n1783,1'b0,n1784,n1786,n1788,n1790);
and (n1784,n1785,n547);
and (n1786,n1787,n558);
and (n1788,n1789,n562);
and (n1790,n1782,n564);
wire s0n1791,s1n1791,notn1791;
or (n1791,s0n1791,s1n1791);
not(notn1791,n690);
and (s0n1791,notn1791,1'b0);
and (s1n1791,n690,n1764);
and (n1792,n1791,n1793);
and (n1793,n1794,n1806);
wire s0n1794,s1n1794,notn1794;
or (n1794,s0n1794,s1n1794);
not(notn1794,n756);
and (s0n1794,notn1794,1'b0);
and (s1n1794,n756,n1795);
wire s0n1795,s1n1795,notn1795;
or (n1795,s0n1795,s1n1795);
not(notn1795,n566);
and (s0n1795,notn1795,n1796);
and (s1n1795,n566,n1798);
wire s0n1796,s1n1796,notn1796;
or (n1796,s0n1796,s1n1796);
not(notn1796,n13);
and (s0n1796,notn1796,1'b0);
and (s1n1796,n13,n1797);
or (n1798,1'b0,n1799,n1801,n1803,n1805);
and (n1799,n1800,n547);
and (n1801,n1802,n558);
and (n1803,n1804,n562);
and (n1805,n1797,n564);
wire s0n1806,s1n1806,notn1806;
or (n1806,s0n1806,s1n1806);
not(notn1806,n690);
and (s0n1806,notn1806,1'b0);
and (s1n1806,n690,n1780);
and (n1807,n1747,n1761);
and (n1808,n1731,n1745);
and (n1809,n1715,n1729);
and (n1810,n1710,n1713);
and (n1811,n1706,n1812);
or (n1812,n1813,n1818,n1868);
and (n1813,n1814,n1817);
xor (n1814,n1815,n1816);
wire s0n1815,s1n1815,notn1815;
or (n1815,s0n1815,s1n1815);
not(notn1815,n583);
and (s0n1815,notn1815,1'b0);
and (s1n1815,n583,n1716);
wire s0n1816,s1n1816,notn1816;
or (n1816,s0n1816,s1n1816);
not(notn1816,n753);
and (s0n1816,notn1816,1'b0);
and (s1n1816,n753,n1694);
xor (n1817,n1707,n1708);
and (n1818,n1817,n1819);
or (n1819,n1820,n1826,n1867);
and (n1820,n1821,n1824);
xor (n1821,n1822,n1823);
wire s0n1822,s1n1822,notn1822;
or (n1822,s0n1822,s1n1822);
not(notn1822,n583);
and (s0n1822,notn1822,1'b0);
and (s1n1822,n583,n1732);
wire s0n1823,s1n1823,notn1823;
or (n1823,s0n1823,s1n1823);
not(notn1823,n753);
and (s0n1823,notn1823,1'b0);
and (s1n1823,n753,n1716);
xor (n1824,n1825,n1713);
xor (n1825,n1710,n1711);
and (n1826,n1824,n1827);
or (n1827,n1828,n1834,n1866);
and (n1828,n1829,n1832);
xor (n1829,n1830,n1831);
wire s0n1830,s1n1830,notn1830;
or (n1830,s0n1830,s1n1830);
not(notn1830,n583);
and (s0n1830,notn1830,1'b0);
and (s1n1830,n583,n1748);
wire s0n1831,s1n1831,notn1831;
or (n1831,s0n1831,s1n1831);
not(notn1831,n753);
and (s0n1831,notn1831,1'b0);
and (s1n1831,n753,n1732);
xor (n1832,n1833,n1729);
xor (n1833,n1715,n1727);
and (n1834,n1832,n1835);
or (n1835,n1836,n1842,n1865);
and (n1836,n1837,n1840);
xor (n1837,n1838,n1839);
wire s0n1838,s1n1838,notn1838;
or (n1838,s0n1838,s1n1838);
not(notn1838,n583);
and (s0n1838,notn1838,1'b0);
and (s1n1838,n583,n1764);
wire s0n1839,s1n1839,notn1839;
or (n1839,s0n1839,s1n1839);
not(notn1839,n753);
and (s0n1839,notn1839,1'b0);
and (s1n1839,n753,n1748);
xor (n1840,n1841,n1745);
xor (n1841,n1731,n1743);
and (n1842,n1840,n1843);
or (n1843,n1844,n1850,n1864);
and (n1844,n1845,n1848);
xor (n1845,n1846,n1847);
wire s0n1846,s1n1846,notn1846;
or (n1846,s0n1846,s1n1846);
not(notn1846,n583);
and (s0n1846,notn1846,1'b0);
and (s1n1846,n583,n1780);
wire s0n1847,s1n1847,notn1847;
or (n1847,s0n1847,s1n1847);
not(notn1847,n753);
and (s0n1847,notn1847,1'b0);
and (s1n1847,n753,n1764);
xor (n1848,n1849,n1761);
xor (n1849,n1747,n1759);
and (n1850,n1848,n1851);
or (n1851,n1852,n1858,n1863);
and (n1852,n1853,n1856);
xor (n1853,n1854,n1855);
wire s0n1854,s1n1854,notn1854;
or (n1854,s0n1854,s1n1854);
not(notn1854,n583);
and (s0n1854,notn1854,1'b0);
and (s1n1854,n583,n1795);
wire s0n1855,s1n1855,notn1855;
or (n1855,s0n1855,s1n1855);
not(notn1855,n753);
and (s0n1855,notn1855,1'b0);
and (s1n1855,n753,n1780);
xor (n1856,n1857,n1777);
xor (n1857,n1763,n1775);
and (n1858,n1856,n1859);
and (n1859,n1860,n1861);
wire s0n1860,s1n1860,notn1860;
or (n1860,s0n1860,s1n1860);
not(notn1860,n753);
and (s0n1860,notn1860,1'b0);
and (s1n1860,n753,n1795);
xor (n1861,n1862,n1793);
xor (n1862,n1779,n1791);
and (n1863,n1853,n1859);
and (n1864,n1845,n1851);
and (n1865,n1837,n1843);
and (n1866,n1829,n1835);
and (n1867,n1821,n1827);
and (n1868,n1814,n1819);
and (n1869,n1692,n1812);
and (n1870,n1871,n1872);
wire s0n1871,s1n1871,notn1871;
or (n1871,s0n1871,s1n1871);
not(notn1871,n970);
and (s0n1871,notn1871,1'b0);
and (s1n1871,n970,n1677);
or (n1872,n1873,n1878,n1943);
and (n1873,n1874,n1877);
wire s0n1874,s1n1874,notn1874;
or (n1874,s0n1874,s1n1874);
not(notn1874,n970);
and (s0n1874,notn1874,1'b0);
and (s1n1874,n970,n1875);
xor (n1875,n1876,n1812);
xor (n1876,n1692,n1706);
wire s0n1877,s1n1877,notn1877;
or (n1877,s0n1877,s1n1877);
not(notn1877,n1018);
and (s0n1877,notn1877,1'b0);
and (s1n1877,n1018,n1677);
and (n1878,n1877,n1879);
or (n1879,n1880,n1885,n1942);
and (n1880,n1881,n1884);
wire s0n1881,s1n1881,notn1881;
or (n1881,s0n1881,s1n1881);
not(notn1881,n970);
and (s0n1881,notn1881,1'b0);
and (s1n1881,n970,n1882);
xor (n1882,n1883,n1819);
xor (n1883,n1814,n1817);
wire s0n1884,s1n1884,notn1884;
or (n1884,s0n1884,s1n1884);
not(notn1884,n1018);
and (s0n1884,notn1884,1'b0);
and (s1n1884,n1018,n1875);
and (n1885,n1884,n1886);
or (n1886,n1887,n1892,n1941);
and (n1887,n1888,n1891);
wire s0n1888,s1n1888,notn1888;
or (n1888,s0n1888,s1n1888);
not(notn1888,n970);
and (s0n1888,notn1888,1'b0);
and (s1n1888,n970,n1889);
xor (n1889,n1890,n1827);
xor (n1890,n1821,n1824);
wire s0n1891,s1n1891,notn1891;
or (n1891,s0n1891,s1n1891);
not(notn1891,n1018);
and (s0n1891,notn1891,1'b0);
and (s1n1891,n1018,n1882);
and (n1892,n1891,n1893);
or (n1893,n1894,n1899,n1940);
and (n1894,n1895,n1898);
wire s0n1895,s1n1895,notn1895;
or (n1895,s0n1895,s1n1895);
not(notn1895,n970);
and (s0n1895,notn1895,1'b0);
and (s1n1895,n970,n1896);
xor (n1896,n1897,n1835);
xor (n1897,n1829,n1832);
wire s0n1898,s1n1898,notn1898;
or (n1898,s0n1898,s1n1898);
not(notn1898,n1018);
and (s0n1898,notn1898,1'b0);
and (s1n1898,n1018,n1889);
and (n1899,n1898,n1900);
or (n1900,n1901,n1906,n1939);
and (n1901,n1902,n1905);
wire s0n1902,s1n1902,notn1902;
or (n1902,s0n1902,s1n1902);
not(notn1902,n970);
and (s0n1902,notn1902,1'b0);
and (s1n1902,n970,n1903);
xor (n1903,n1904,n1843);
xor (n1904,n1837,n1840);
wire s0n1905,s1n1905,notn1905;
or (n1905,s0n1905,s1n1905);
not(notn1905,n1018);
and (s0n1905,notn1905,1'b0);
and (s1n1905,n1018,n1896);
and (n1906,n1905,n1907);
or (n1907,n1908,n1913,n1938);
and (n1908,n1909,n1912);
wire s0n1909,s1n1909,notn1909;
or (n1909,s0n1909,s1n1909);
not(notn1909,n970);
and (s0n1909,notn1909,1'b0);
and (s1n1909,n970,n1910);
xor (n1910,n1911,n1851);
xor (n1911,n1845,n1848);
wire s0n1912,s1n1912,notn1912;
or (n1912,s0n1912,s1n1912);
not(notn1912,n1018);
and (s0n1912,notn1912,1'b0);
and (s1n1912,n1018,n1903);
and (n1913,n1912,n1914);
or (n1914,n1915,n1920,n1937);
and (n1915,n1916,n1919);
wire s0n1916,s1n1916,notn1916;
or (n1916,s0n1916,s1n1916);
not(notn1916,n970);
and (s0n1916,notn1916,1'b0);
and (s1n1916,n970,n1917);
xor (n1917,n1918,n1859);
xor (n1918,n1853,n1856);
wire s0n1919,s1n1919,notn1919;
or (n1919,s0n1919,s1n1919);
not(notn1919,n1018);
and (s0n1919,notn1919,1'b0);
and (s1n1919,n1018,n1910);
and (n1920,n1919,n1921);
or (n1921,n1922,n1926,n1928);
and (n1922,n1923,n1925);
wire s0n1923,s1n1923,notn1923;
or (n1923,s0n1923,s1n1923);
not(notn1923,n970);
and (s0n1923,notn1923,1'b0);
and (s1n1923,n970,n1924);
xor (n1924,n1860,n1861);
wire s0n1925,s1n1925,notn1925;
or (n1925,s0n1925,s1n1925);
not(notn1925,n1018);
and (s0n1925,notn1925,1'b0);
and (s1n1925,n1018,n1917);
and (n1926,n1925,n1927);
or (n1927,n1928,n1932,n1933);
and (n1928,n1929,n1931);
wire s0n1929,s1n1929,notn1929;
or (n1929,s0n1929,s1n1929);
not(notn1929,n970);
and (s0n1929,notn1929,1'b0);
and (s1n1929,n970,n1930);
xor (n1930,n1794,n1806);
wire s0n1931,s1n1931,notn1931;
or (n1931,s0n1931,s1n1931);
not(notn1931,n1018);
and (s0n1931,notn1931,1'b0);
and (s1n1931,n1018,n1924);
and (n1932,n1931,n1933);
and (n1933,n1934,n1936);
wire s0n1934,s1n1934,notn1934;
or (n1934,s0n1934,s1n1934);
not(notn1934,n970);
and (s0n1934,notn1934,1'b0);
and (s1n1934,n970,n1935);
wire s0n1935,s1n1935,notn1935;
or (n1935,s0n1935,s1n1935);
not(notn1935,n690);
and (s0n1935,notn1935,1'b0);
and (s1n1935,n690,n1795);
wire s0n1936,s1n1936,notn1936;
or (n1936,s0n1936,s1n1936);
not(notn1936,n1018);
and (s0n1936,notn1936,1'b0);
and (s1n1936,n1018,n1930);
and (n1937,n1916,n1921);
and (n1938,n1909,n1914);
and (n1939,n1902,n1907);
and (n1940,n1895,n1900);
and (n1941,n1888,n1893);
and (n1942,n1881,n1886);
and (n1943,n1874,n1879);
and (n1944,n1870,n1945);
or (n1945,n1946,n1949,n2010);
and (n1946,n1947,n1948);
wire s0n1947,s1n1947,notn1947;
or (n1947,s0n1947,s1n1947);
not(notn1947,n921);
and (s0n1947,notn1947,1'b0);
and (s1n1947,n921,n1875);
xor (n1948,n1871,n1872);
and (n1949,n1948,n1950);
or (n1950,n1951,n1955,n2009);
and (n1951,n1952,n1953);
wire s0n1952,s1n1952,notn1952;
or (n1952,s0n1952,s1n1952);
not(notn1952,n921);
and (s0n1952,notn1952,1'b0);
and (s1n1952,n921,n1882);
xor (n1953,n1954,n1879);
xor (n1954,n1874,n1877);
and (n1955,n1953,n1956);
or (n1956,n1957,n1961,n2008);
and (n1957,n1958,n1959);
wire s0n1958,s1n1958,notn1958;
or (n1958,s0n1958,s1n1958);
not(notn1958,n921);
and (s0n1958,notn1958,1'b0);
and (s1n1958,n921,n1889);
xor (n1959,n1960,n1886);
xor (n1960,n1881,n1884);
and (n1961,n1959,n1962);
or (n1962,n1963,n1967,n2007);
and (n1963,n1964,n1965);
wire s0n1964,s1n1964,notn1964;
or (n1964,s0n1964,s1n1964);
not(notn1964,n921);
and (s0n1964,notn1964,1'b0);
and (s1n1964,n921,n1896);
xor (n1965,n1966,n1893);
xor (n1966,n1888,n1891);
and (n1967,n1965,n1968);
or (n1968,n1969,n1973,n2006);
and (n1969,n1970,n1971);
wire s0n1970,s1n1970,notn1970;
or (n1970,s0n1970,s1n1970);
not(notn1970,n921);
and (s0n1970,notn1970,1'b0);
and (s1n1970,n921,n1903);
xor (n1971,n1972,n1900);
xor (n1972,n1895,n1898);
and (n1973,n1971,n1974);
or (n1974,n1975,n1979,n2005);
and (n1975,n1976,n1977);
wire s0n1976,s1n1976,notn1976;
or (n1976,s0n1976,s1n1976);
not(notn1976,n921);
and (s0n1976,notn1976,1'b0);
and (s1n1976,n921,n1910);
xor (n1977,n1978,n1907);
xor (n1978,n1902,n1905);
and (n1979,n1977,n1980);
or (n1980,n1981,n1985,n2004);
and (n1981,n1982,n1983);
wire s0n1982,s1n1982,notn1982;
or (n1982,s0n1982,s1n1982);
not(notn1982,n921);
and (s0n1982,notn1982,1'b0);
and (s1n1982,n921,n1917);
xor (n1983,n1984,n1914);
xor (n1984,n1909,n1912);
and (n1985,n1983,n1986);
or (n1986,n1987,n1991,n2003);
and (n1987,n1988,n1989);
wire s0n1988,s1n1988,notn1988;
or (n1988,s0n1988,s1n1988);
not(notn1988,n921);
and (s0n1988,notn1988,1'b0);
and (s1n1988,n921,n1924);
xor (n1989,n1990,n1921);
xor (n1990,n1916,n1919);
and (n1991,n1989,n1992);
or (n1992,n1993,n1997,n2002);
and (n1993,n1994,n1995);
wire s0n1994,s1n1994,notn1994;
or (n1994,s0n1994,s1n1994);
not(notn1994,n921);
and (s0n1994,notn1994,1'b0);
and (s1n1994,n921,n1930);
xor (n1995,n1996,n1927);
xor (n1996,n1923,n1925);
and (n1997,n1995,n1998);
and (n1998,n1999,n2000);
wire s0n1999,s1n1999,notn1999;
or (n1999,s0n1999,s1n1999);
not(notn1999,n921);
and (s0n1999,notn1999,1'b0);
and (s1n1999,n921,n1935);
xor (n2000,n2001,n1933);
xor (n2001,n1929,n1931);
and (n2002,n1994,n1998);
and (n2003,n1988,n1992);
and (n2004,n1982,n1986);
and (n2005,n1976,n1980);
and (n2006,n1970,n1974);
and (n2007,n1964,n1968);
and (n2008,n1958,n1962);
and (n2009,n1952,n1956);
and (n2010,n1947,n1950);
and (n2011,n1676,n1945);
or (n2012,n2013,n2266,n2333);
and (n2013,n2014,n2192);
wire s0n2014,s1n2014,notn2014;
or (n2014,s0n2014,s1n2014);
not(notn2014,n921);
and (s0n2014,notn2014,1'b0);
and (s1n2014,n921,n2015);
or (n2015,n2016,n2145,n2191);
and (n2016,n2017,n2029);
wire s0n2017,s1n2017,notn2017;
or (n2017,s0n2017,s1n2017);
not(notn2017,n585);
and (s0n2017,notn2017,1'b0);
and (s1n2017,n585,n2018);
wire s0n2018,s1n2018,notn2018;
or (n2018,s0n2018,s1n2018);
not(notn2018,n566);
and (s0n2018,notn2018,n2019);
and (s1n2018,n566,n2021);
wire s0n2019,s1n2019,notn2019;
or (n2019,s0n2019,s1n2019);
not(notn2019,n13);
and (s0n2019,notn2019,1'b0);
and (s1n2019,n13,n2020);
or (n2021,1'b0,n2022,n2024,n2026,n2028);
and (n2022,n2023,n547);
and (n2024,n2025,n558);
and (n2026,n2027,n562);
and (n2028,n2020,n564);
and (n2029,n2030,n2031);
wire s0n2030,s1n2030,notn2030;
or (n2030,s0n2030,s1n2030);
not(notn2030,n642);
and (s0n2030,notn2030,1'b0);
and (s1n2030,n642,n2018);
or (n2031,n2032,n2046,n2144);
and (n2032,n2033,n2045);
wire s0n2033,s1n2033,notn2033;
or (n2033,s0n2033,s1n2033);
not(notn2033,n642);
and (s0n2033,notn2033,1'b0);
and (s1n2033,n642,n2034);
wire s0n2034,s1n2034,notn2034;
or (n2034,s0n2034,s1n2034);
not(notn2034,n566);
and (s0n2034,notn2034,n2035);
and (s1n2034,n566,n2037);
wire s0n2035,s1n2035,notn2035;
or (n2035,s0n2035,s1n2035);
not(notn2035,n13);
and (s0n2035,notn2035,1'b0);
and (s1n2035,n13,n2036);
or (n2037,1'b0,n2038,n2040,n2042,n2044);
and (n2038,n2039,n547);
and (n2040,n2041,n558);
and (n2042,n2043,n562);
and (n2044,n2036,n564);
wire s0n2045,s1n2045,notn2045;
or (n2045,s0n2045,s1n2045);
not(notn2045,n690);
and (s0n2045,notn2045,1'b0);
and (s1n2045,n690,n2018);
and (n2046,n2045,n2047);
or (n2047,n2048,n2062,n2143);
and (n2048,n2049,n2061);
wire s0n2049,s1n2049,notn2049;
or (n2049,s0n2049,s1n2049);
not(notn2049,n642);
and (s0n2049,notn2049,1'b0);
and (s1n2049,n642,n2050);
wire s0n2050,s1n2050,notn2050;
or (n2050,s0n2050,s1n2050);
not(notn2050,n566);
and (s0n2050,notn2050,n2051);
and (s1n2050,n566,n2053);
wire s0n2051,s1n2051,notn2051;
or (n2051,s0n2051,s1n2051);
not(notn2051,n13);
and (s0n2051,notn2051,1'b0);
and (s1n2051,n13,n2052);
or (n2053,1'b0,n2054,n2056,n2058,n2060);
and (n2054,n2055,n547);
and (n2056,n2057,n558);
and (n2058,n2059,n562);
and (n2060,n2052,n564);
wire s0n2061,s1n2061,notn2061;
or (n2061,s0n2061,s1n2061);
not(notn2061,n690);
and (s0n2061,notn2061,1'b0);
and (s1n2061,n690,n2034);
and (n2062,n2061,n2063);
or (n2063,n2064,n2078,n2142);
and (n2064,n2065,n2077);
wire s0n2065,s1n2065,notn2065;
or (n2065,s0n2065,s1n2065);
not(notn2065,n642);
and (s0n2065,notn2065,1'b0);
and (s1n2065,n642,n2066);
wire s0n2066,s1n2066,notn2066;
or (n2066,s0n2066,s1n2066);
not(notn2066,n566);
and (s0n2066,notn2066,n2067);
and (s1n2066,n566,n2069);
wire s0n2067,s1n2067,notn2067;
or (n2067,s0n2067,s1n2067);
not(notn2067,n13);
and (s0n2067,notn2067,1'b0);
and (s1n2067,n13,n2068);
or (n2069,1'b0,n2070,n2072,n2074,n2076);
and (n2070,n2071,n547);
and (n2072,n2073,n558);
and (n2074,n2075,n562);
and (n2076,n2068,n564);
wire s0n2077,s1n2077,notn2077;
or (n2077,s0n2077,s1n2077);
not(notn2077,n690);
and (s0n2077,notn2077,1'b0);
and (s1n2077,n690,n2050);
and (n2078,n2077,n2079);
or (n2079,n2080,n2094,n2141);
and (n2080,n2081,n2093);
wire s0n2081,s1n2081,notn2081;
or (n2081,s0n2081,s1n2081);
not(notn2081,n642);
and (s0n2081,notn2081,1'b0);
and (s1n2081,n642,n2082);
wire s0n2082,s1n2082,notn2082;
or (n2082,s0n2082,s1n2082);
not(notn2082,n566);
and (s0n2082,notn2082,n2083);
and (s1n2082,n566,n2085);
wire s0n2083,s1n2083,notn2083;
or (n2083,s0n2083,s1n2083);
not(notn2083,n13);
and (s0n2083,notn2083,1'b0);
and (s1n2083,n13,n2084);
or (n2085,1'b0,n2086,n2088,n2090,n2092);
and (n2086,n2087,n547);
and (n2088,n2089,n558);
and (n2090,n2091,n562);
and (n2092,n2084,n564);
wire s0n2093,s1n2093,notn2093;
or (n2093,s0n2093,s1n2093);
not(notn2093,n690);
and (s0n2093,notn2093,1'b0);
and (s1n2093,n690,n2066);
and (n2094,n2093,n2095);
or (n2095,n2096,n2110,n2112);
and (n2096,n2097,n2109);
wire s0n2097,s1n2097,notn2097;
or (n2097,s0n2097,s1n2097);
not(notn2097,n642);
and (s0n2097,notn2097,1'b0);
and (s1n2097,n642,n2098);
wire s0n2098,s1n2098,notn2098;
or (n2098,s0n2098,s1n2098);
not(notn2098,n566);
and (s0n2098,notn2098,n2099);
and (s1n2098,n566,n2101);
wire s0n2099,s1n2099,notn2099;
or (n2099,s0n2099,s1n2099);
not(notn2099,n13);
and (s0n2099,notn2099,1'b0);
and (s1n2099,n13,n2100);
or (n2101,1'b0,n2102,n2104,n2106,n2108);
and (n2102,n2103,n547);
and (n2104,n2105,n558);
and (n2106,n2107,n562);
and (n2108,n2100,n564);
wire s0n2109,s1n2109,notn2109;
or (n2109,s0n2109,s1n2109);
not(notn2109,n690);
and (s0n2109,notn2109,1'b0);
and (s1n2109,n690,n2082);
and (n2110,n2109,n2111);
or (n2111,n2112,n2126,n2127);
and (n2112,n2113,n2125);
wire s0n2113,s1n2113,notn2113;
or (n2113,s0n2113,s1n2113);
not(notn2113,n642);
and (s0n2113,notn2113,1'b0);
and (s1n2113,n642,n2114);
wire s0n2114,s1n2114,notn2114;
or (n2114,s0n2114,s1n2114);
not(notn2114,n566);
and (s0n2114,notn2114,n2115);
and (s1n2114,n566,n2117);
wire s0n2115,s1n2115,notn2115;
or (n2115,s0n2115,s1n2115);
not(notn2115,n13);
and (s0n2115,notn2115,1'b0);
and (s1n2115,n13,n2116);
or (n2117,1'b0,n2118,n2120,n2122,n2124);
and (n2118,n2119,n547);
and (n2120,n2121,n558);
and (n2122,n2123,n562);
and (n2124,n2116,n564);
wire s0n2125,s1n2125,notn2125;
or (n2125,s0n2125,s1n2125);
not(notn2125,n690);
and (s0n2125,notn2125,1'b0);
and (s1n2125,n690,n2098);
and (n2126,n2125,n2127);
and (n2127,n2128,n2140);
wire s0n2128,s1n2128,notn2128;
or (n2128,s0n2128,s1n2128);
not(notn2128,n642);
and (s0n2128,notn2128,1'b0);
and (s1n2128,n642,n2129);
wire s0n2129,s1n2129,notn2129;
or (n2129,s0n2129,s1n2129);
not(notn2129,n566);
and (s0n2129,notn2129,n2130);
and (s1n2129,n566,n2132);
wire s0n2130,s1n2130,notn2130;
or (n2130,s0n2130,s1n2130);
not(notn2130,n13);
and (s0n2130,notn2130,1'b0);
and (s1n2130,n13,n2131);
or (n2132,1'b0,n2133,n2135,n2137,n2139);
and (n2133,n2134,n547);
and (n2135,n2136,n558);
and (n2137,n2138,n562);
and (n2139,n2131,n564);
wire s0n2140,s1n2140,notn2140;
or (n2140,s0n2140,s1n2140);
not(notn2140,n690);
and (s0n2140,notn2140,1'b0);
and (s1n2140,n690,n2114);
and (n2141,n2081,n2095);
and (n2142,n2065,n2079);
and (n2143,n2049,n2063);
and (n2144,n2033,n2047);
and (n2145,n2029,n2146);
or (n2146,n2147,n2150,n2190);
and (n2147,n2148,n2149);
wire s0n2148,s1n2148,notn2148;
or (n2148,s0n2148,s1n2148);
not(notn2148,n585);
and (s0n2148,notn2148,1'b0);
and (s1n2148,n585,n2034);
xor (n2149,n2030,n2031);
and (n2150,n2149,n2151);
or (n2151,n2152,n2156,n2189);
and (n2152,n2153,n2154);
wire s0n2153,s1n2153,notn2153;
or (n2153,s0n2153,s1n2153);
not(notn2153,n585);
and (s0n2153,notn2153,1'b0);
and (s1n2153,n585,n2050);
xor (n2154,n2155,n2047);
xor (n2155,n2033,n2045);
and (n2156,n2154,n2157);
or (n2157,n2158,n2162,n2188);
and (n2158,n2159,n2160);
wire s0n2159,s1n2159,notn2159;
or (n2159,s0n2159,s1n2159);
not(notn2159,n585);
and (s0n2159,notn2159,1'b0);
and (s1n2159,n585,n2066);
xor (n2160,n2161,n2063);
xor (n2161,n2049,n2061);
and (n2162,n2160,n2163);
or (n2163,n2164,n2168,n2187);
and (n2164,n2165,n2166);
wire s0n2165,s1n2165,notn2165;
or (n2165,s0n2165,s1n2165);
not(notn2165,n585);
and (s0n2165,notn2165,1'b0);
and (s1n2165,n585,n2082);
xor (n2166,n2167,n2079);
xor (n2167,n2065,n2077);
and (n2168,n2166,n2169);
or (n2169,n2170,n2174,n2186);
and (n2170,n2171,n2172);
wire s0n2171,s1n2171,notn2171;
or (n2171,s0n2171,s1n2171);
not(notn2171,n585);
and (s0n2171,notn2171,1'b0);
and (s1n2171,n585,n2098);
xor (n2172,n2173,n2095);
xor (n2173,n2081,n2093);
and (n2174,n2172,n2175);
or (n2175,n2176,n2180,n2185);
and (n2176,n2177,n2178);
wire s0n2177,s1n2177,notn2177;
or (n2177,s0n2177,s1n2177);
not(notn2177,n585);
and (s0n2177,notn2177,1'b0);
and (s1n2177,n585,n2114);
xor (n2178,n2179,n2111);
xor (n2179,n2097,n2109);
and (n2180,n2178,n2181);
and (n2181,n2182,n2183);
wire s0n2182,s1n2182,notn2182;
or (n2182,s0n2182,s1n2182);
not(notn2182,n585);
and (s0n2182,notn2182,1'b0);
and (s1n2182,n585,n2129);
xor (n2183,n2184,n2127);
xor (n2184,n2113,n2125);
and (n2185,n2177,n2181);
and (n2186,n2171,n2175);
and (n2187,n2165,n2169);
and (n2188,n2159,n2163);
and (n2189,n2153,n2157);
and (n2190,n2148,n2151);
and (n2191,n2017,n2146);
and (n2192,n2193,n2194);
wire s0n2193,s1n2193,notn2193;
or (n2193,s0n2193,s1n2193);
not(notn2193,n970);
and (s0n2193,notn2193,1'b0);
and (s1n2193,n970,n2015);
or (n2194,n2195,n2200,n2265);
and (n2195,n2196,n2199);
wire s0n2196,s1n2196,notn2196;
or (n2196,s0n2196,s1n2196);
not(notn2196,n970);
and (s0n2196,notn2196,1'b0);
and (s1n2196,n970,n2197);
xor (n2197,n2198,n2146);
xor (n2198,n2017,n2029);
wire s0n2199,s1n2199,notn2199;
or (n2199,s0n2199,s1n2199);
not(notn2199,n1018);
and (s0n2199,notn2199,1'b0);
and (s1n2199,n1018,n2015);
and (n2200,n2199,n2201);
or (n2201,n2202,n2207,n2264);
and (n2202,n2203,n2206);
wire s0n2203,s1n2203,notn2203;
or (n2203,s0n2203,s1n2203);
not(notn2203,n970);
and (s0n2203,notn2203,1'b0);
and (s1n2203,n970,n2204);
xor (n2204,n2205,n2151);
xor (n2205,n2148,n2149);
wire s0n2206,s1n2206,notn2206;
or (n2206,s0n2206,s1n2206);
not(notn2206,n1018);
and (s0n2206,notn2206,1'b0);
and (s1n2206,n1018,n2197);
and (n2207,n2206,n2208);
or (n2208,n2209,n2214,n2263);
and (n2209,n2210,n2213);
wire s0n2210,s1n2210,notn2210;
or (n2210,s0n2210,s1n2210);
not(notn2210,n970);
and (s0n2210,notn2210,1'b0);
and (s1n2210,n970,n2211);
xor (n2211,n2212,n2157);
xor (n2212,n2153,n2154);
wire s0n2213,s1n2213,notn2213;
or (n2213,s0n2213,s1n2213);
not(notn2213,n1018);
and (s0n2213,notn2213,1'b0);
and (s1n2213,n1018,n2204);
and (n2214,n2213,n2215);
or (n2215,n2216,n2221,n2262);
and (n2216,n2217,n2220);
wire s0n2217,s1n2217,notn2217;
or (n2217,s0n2217,s1n2217);
not(notn2217,n970);
and (s0n2217,notn2217,1'b0);
and (s1n2217,n970,n2218);
xor (n2218,n2219,n2163);
xor (n2219,n2159,n2160);
wire s0n2220,s1n2220,notn2220;
or (n2220,s0n2220,s1n2220);
not(notn2220,n1018);
and (s0n2220,notn2220,1'b0);
and (s1n2220,n1018,n2211);
and (n2221,n2220,n2222);
or (n2222,n2223,n2228,n2261);
and (n2223,n2224,n2227);
wire s0n2224,s1n2224,notn2224;
or (n2224,s0n2224,s1n2224);
not(notn2224,n970);
and (s0n2224,notn2224,1'b0);
and (s1n2224,n970,n2225);
xor (n2225,n2226,n2169);
xor (n2226,n2165,n2166);
wire s0n2227,s1n2227,notn2227;
or (n2227,s0n2227,s1n2227);
not(notn2227,n1018);
and (s0n2227,notn2227,1'b0);
and (s1n2227,n1018,n2218);
and (n2228,n2227,n2229);
or (n2229,n2230,n2235,n2260);
and (n2230,n2231,n2234);
wire s0n2231,s1n2231,notn2231;
or (n2231,s0n2231,s1n2231);
not(notn2231,n970);
and (s0n2231,notn2231,1'b0);
and (s1n2231,n970,n2232);
xor (n2232,n2233,n2175);
xor (n2233,n2171,n2172);
wire s0n2234,s1n2234,notn2234;
or (n2234,s0n2234,s1n2234);
not(notn2234,n1018);
and (s0n2234,notn2234,1'b0);
and (s1n2234,n1018,n2225);
and (n2235,n2234,n2236);
or (n2236,n2237,n2242,n2259);
and (n2237,n2238,n2241);
wire s0n2238,s1n2238,notn2238;
or (n2238,s0n2238,s1n2238);
not(notn2238,n970);
and (s0n2238,notn2238,1'b0);
and (s1n2238,n970,n2239);
xor (n2239,n2240,n2181);
xor (n2240,n2177,n2178);
wire s0n2241,s1n2241,notn2241;
or (n2241,s0n2241,s1n2241);
not(notn2241,n1018);
and (s0n2241,notn2241,1'b0);
and (s1n2241,n1018,n2232);
and (n2242,n2241,n2243);
or (n2243,n2244,n2248,n2250);
and (n2244,n2245,n2247);
wire s0n2245,s1n2245,notn2245;
or (n2245,s0n2245,s1n2245);
not(notn2245,n970);
and (s0n2245,notn2245,1'b0);
and (s1n2245,n970,n2246);
xor (n2246,n2182,n2183);
wire s0n2247,s1n2247,notn2247;
or (n2247,s0n2247,s1n2247);
not(notn2247,n1018);
and (s0n2247,notn2247,1'b0);
and (s1n2247,n1018,n2239);
and (n2248,n2247,n2249);
or (n2249,n2250,n2254,n2255);
and (n2250,n2251,n2253);
wire s0n2251,s1n2251,notn2251;
or (n2251,s0n2251,s1n2251);
not(notn2251,n970);
and (s0n2251,notn2251,1'b0);
and (s1n2251,n970,n2252);
xor (n2252,n2128,n2140);
wire s0n2253,s1n2253,notn2253;
or (n2253,s0n2253,s1n2253);
not(notn2253,n1018);
and (s0n2253,notn2253,1'b0);
and (s1n2253,n1018,n2246);
and (n2254,n2253,n2255);
and (n2255,n2256,n2258);
wire s0n2256,s1n2256,notn2256;
or (n2256,s0n2256,s1n2256);
not(notn2256,n970);
and (s0n2256,notn2256,1'b0);
and (s1n2256,n970,n2257);
wire s0n2257,s1n2257,notn2257;
or (n2257,s0n2257,s1n2257);
not(notn2257,n690);
and (s0n2257,notn2257,1'b0);
and (s1n2257,n690,n2129);
wire s0n2258,s1n2258,notn2258;
or (n2258,s0n2258,s1n2258);
not(notn2258,n1018);
and (s0n2258,notn2258,1'b0);
and (s1n2258,n1018,n2252);
and (n2259,n2238,n2243);
and (n2260,n2231,n2236);
and (n2261,n2224,n2229);
and (n2262,n2217,n2222);
and (n2263,n2210,n2215);
and (n2264,n2203,n2208);
and (n2265,n2196,n2201);
and (n2266,n2192,n2267);
or (n2267,n2268,n2271,n2332);
and (n2268,n2269,n2270);
wire s0n2269,s1n2269,notn2269;
or (n2269,s0n2269,s1n2269);
not(notn2269,n921);
and (s0n2269,notn2269,1'b0);
and (s1n2269,n921,n2197);
xor (n2270,n2193,n2194);
and (n2271,n2270,n2272);
or (n2272,n2273,n2277,n2331);
and (n2273,n2274,n2275);
wire s0n2274,s1n2274,notn2274;
or (n2274,s0n2274,s1n2274);
not(notn2274,n921);
and (s0n2274,notn2274,1'b0);
and (s1n2274,n921,n2204);
xor (n2275,n2276,n2201);
xor (n2276,n2196,n2199);
and (n2277,n2275,n2278);
or (n2278,n2279,n2283,n2330);
and (n2279,n2280,n2281);
wire s0n2280,s1n2280,notn2280;
or (n2280,s0n2280,s1n2280);
not(notn2280,n921);
and (s0n2280,notn2280,1'b0);
and (s1n2280,n921,n2211);
xor (n2281,n2282,n2208);
xor (n2282,n2203,n2206);
and (n2283,n2281,n2284);
or (n2284,n2285,n2289,n2329);
and (n2285,n2286,n2287);
wire s0n2286,s1n2286,notn2286;
or (n2286,s0n2286,s1n2286);
not(notn2286,n921);
and (s0n2286,notn2286,1'b0);
and (s1n2286,n921,n2218);
xor (n2287,n2288,n2215);
xor (n2288,n2210,n2213);
and (n2289,n2287,n2290);
or (n2290,n2291,n2295,n2328);
and (n2291,n2292,n2293);
wire s0n2292,s1n2292,notn2292;
or (n2292,s0n2292,s1n2292);
not(notn2292,n921);
and (s0n2292,notn2292,1'b0);
and (s1n2292,n921,n2225);
xor (n2293,n2294,n2222);
xor (n2294,n2217,n2220);
and (n2295,n2293,n2296);
or (n2296,n2297,n2301,n2327);
and (n2297,n2298,n2299);
wire s0n2298,s1n2298,notn2298;
or (n2298,s0n2298,s1n2298);
not(notn2298,n921);
and (s0n2298,notn2298,1'b0);
and (s1n2298,n921,n2232);
xor (n2299,n2300,n2229);
xor (n2300,n2224,n2227);
and (n2301,n2299,n2302);
or (n2302,n2303,n2307,n2326);
and (n2303,n2304,n2305);
wire s0n2304,s1n2304,notn2304;
or (n2304,s0n2304,s1n2304);
not(notn2304,n921);
and (s0n2304,notn2304,1'b0);
and (s1n2304,n921,n2239);
xor (n2305,n2306,n2236);
xor (n2306,n2231,n2234);
and (n2307,n2305,n2308);
or (n2308,n2309,n2313,n2325);
and (n2309,n2310,n2311);
wire s0n2310,s1n2310,notn2310;
or (n2310,s0n2310,s1n2310);
not(notn2310,n921);
and (s0n2310,notn2310,1'b0);
and (s1n2310,n921,n2246);
xor (n2311,n2312,n2243);
xor (n2312,n2238,n2241);
and (n2313,n2311,n2314);
or (n2314,n2315,n2319,n2324);
and (n2315,n2316,n2317);
wire s0n2316,s1n2316,notn2316;
or (n2316,s0n2316,s1n2316);
not(notn2316,n921);
and (s0n2316,notn2316,1'b0);
and (s1n2316,n921,n2252);
xor (n2317,n2318,n2249);
xor (n2318,n2245,n2247);
and (n2319,n2317,n2320);
and (n2320,n2321,n2322);
wire s0n2321,s1n2321,notn2321;
or (n2321,s0n2321,s1n2321);
not(notn2321,n921);
and (s0n2321,notn2321,1'b0);
and (s1n2321,n921,n2257);
xor (n2322,n2323,n2255);
xor (n2323,n2251,n2253);
and (n2324,n2316,n2320);
and (n2325,n2310,n2314);
and (n2326,n2304,n2308);
and (n2327,n2298,n2302);
and (n2328,n2292,n2296);
and (n2329,n2286,n2290);
and (n2330,n2280,n2284);
and (n2331,n2274,n2278);
and (n2332,n2269,n2272);
and (n2333,n2014,n2267);
or (n2334,n2335,n2340,n2428);
and (n2335,n2336,n2338);
xor (n2336,n2337,n1945);
xor (n2337,n1676,n1870);
xor (n2338,n2339,n2267);
xor (n2339,n2014,n2192);
and (n2340,n2338,n2341);
or (n2341,n2342,n2347,n2427);
and (n2342,n2343,n2345);
xor (n2343,n2344,n1950);
xor (n2344,n1947,n1948);
xor (n2345,n2346,n2272);
xor (n2346,n2269,n2270);
and (n2347,n2345,n2348);
or (n2348,n2349,n2354,n2426);
and (n2349,n2350,n2352);
xor (n2350,n2351,n1956);
xor (n2351,n1952,n1953);
xor (n2352,n2353,n2278);
xor (n2353,n2274,n2275);
and (n2354,n2352,n2355);
or (n2355,n2356,n2361,n2425);
and (n2356,n2357,n2359);
xor (n2357,n2358,n1962);
xor (n2358,n1958,n1959);
xor (n2359,n2360,n2284);
xor (n2360,n2280,n2281);
and (n2361,n2359,n2362);
or (n2362,n2363,n2368,n2424);
and (n2363,n2364,n2366);
xor (n2364,n2365,n1968);
xor (n2365,n1964,n1965);
xor (n2366,n2367,n2290);
xor (n2367,n2286,n2287);
and (n2368,n2366,n2369);
or (n2369,n2370,n2375,n2423);
and (n2370,n2371,n2373);
xor (n2371,n2372,n1974);
xor (n2372,n1970,n1971);
xor (n2373,n2374,n2296);
xor (n2374,n2292,n2293);
and (n2375,n2373,n2376);
or (n2376,n2377,n2382,n2422);
and (n2377,n2378,n2380);
xor (n2378,n2379,n1980);
xor (n2379,n1976,n1977);
xor (n2380,n2381,n2302);
xor (n2381,n2298,n2299);
and (n2382,n2380,n2383);
or (n2383,n2384,n2389,n2421);
and (n2384,n2385,n2387);
xor (n2385,n2386,n1986);
xor (n2386,n1982,n1983);
xor (n2387,n2388,n2308);
xor (n2388,n2304,n2305);
and (n2389,n2387,n2390);
or (n2390,n2391,n2396,n2420);
and (n2391,n2392,n2394);
xor (n2392,n2393,n1992);
xor (n2393,n1988,n1989);
xor (n2394,n2395,n2314);
xor (n2395,n2310,n2311);
and (n2396,n2394,n2397);
or (n2397,n2398,n2403,n2419);
and (n2398,n2399,n2401);
xor (n2399,n2400,n1998);
xor (n2400,n1994,n1995);
xor (n2401,n2402,n2320);
xor (n2402,n2316,n2317);
and (n2403,n2401,n2404);
or (n2404,n2405,n2408,n2418);
and (n2405,n2406,n2407);
xor (n2406,n1999,n2000);
xor (n2407,n2321,n2322);
and (n2408,n2407,n2409);
or (n2409,n2410,n2413,n2417);
and (n2410,n2411,n2412);
xor (n2411,n1934,n1936);
xor (n2412,n2256,n2258);
and (n2413,n2412,n2414);
and (n2414,n2415,n2416);
wire s0n2415,s1n2415,notn2415;
or (n2415,s0n2415,s1n2415);
not(notn2415,n1018);
and (s0n2415,notn2415,1'b0);
and (s1n2415,n1018,n1935);
wire s0n2416,s1n2416,notn2416;
or (n2416,s0n2416,s1n2416);
not(notn2416,n1018);
and (s0n2416,notn2416,1'b0);
and (s1n2416,n1018,n2257);
and (n2417,n2411,n2414);
and (n2418,n2406,n2409);
and (n2419,n2399,n2404);
and (n2420,n2392,n2397);
and (n2421,n2385,n2390);
and (n2422,n2378,n2383);
and (n2423,n2371,n2376);
and (n2424,n2364,n2369);
and (n2425,n2357,n2362);
and (n2426,n2350,n2355);
and (n2427,n2343,n2348);
and (n2428,n2336,n2341);
or (n2429,n2430,n2435,n2527);
and (n2430,n2431,n2433);
xor (n2431,n2432,n1584);
xor (n2432,n1579,n1581);
xor (n2433,n2434,n2341);
xor (n2434,n2336,n2338);
and (n2435,n2433,n2436);
or (n2436,n2437,n2442,n2526);
and (n2437,n2438,n2440);
xor (n2438,n2439,n1591);
xor (n2439,n1586,n1588);
xor (n2440,n2441,n2348);
xor (n2441,n2343,n2345);
and (n2442,n2440,n2443);
or (n2443,n2444,n2449,n2525);
and (n2444,n2445,n2447);
xor (n2445,n2446,n1598);
xor (n2446,n1593,n1595);
xor (n2447,n2448,n2355);
xor (n2448,n2350,n2352);
and (n2449,n2447,n2450);
or (n2450,n2451,n2456,n2524);
and (n2451,n2452,n2454);
xor (n2452,n2453,n1605);
xor (n2453,n1600,n1602);
xor (n2454,n2455,n2362);
xor (n2455,n2357,n2359);
and (n2456,n2454,n2457);
or (n2457,n2458,n2463,n2523);
and (n2458,n2459,n2461);
xor (n2459,n2460,n1612);
xor (n2460,n1607,n1609);
xor (n2461,n2462,n2369);
xor (n2462,n2364,n2366);
and (n2463,n2461,n2464);
or (n2464,n2465,n2470,n2522);
and (n2465,n2466,n2468);
xor (n2466,n2467,n1619);
xor (n2467,n1614,n1616);
xor (n2468,n2469,n2376);
xor (n2469,n2371,n2373);
and (n2470,n2468,n2471);
or (n2471,n2472,n2477,n2521);
and (n2472,n2473,n2475);
xor (n2473,n2474,n1626);
xor (n2474,n1621,n1623);
xor (n2475,n2476,n2383);
xor (n2476,n2378,n2380);
and (n2477,n2475,n2478);
or (n2478,n2479,n2484,n2520);
and (n2479,n2480,n2482);
xor (n2480,n2481,n1633);
xor (n2481,n1628,n1630);
xor (n2482,n2483,n2390);
xor (n2483,n2385,n2387);
and (n2484,n2482,n2485);
or (n2485,n2486,n2491,n2519);
and (n2486,n2487,n2489);
xor (n2487,n2488,n1640);
xor (n2488,n1635,n1637);
xor (n2489,n2490,n2397);
xor (n2490,n2392,n2394);
and (n2491,n2489,n2492);
or (n2492,n2493,n2498,n2518);
and (n2493,n2494,n2496);
xor (n2494,n2495,n1647);
xor (n2495,n1642,n1644);
xor (n2496,n2497,n2404);
xor (n2497,n2399,n2401);
and (n2498,n2496,n2499);
or (n2499,n2500,n2505,n2517);
and (n2500,n2501,n2503);
xor (n2501,n2502,n1652);
xor (n2502,n1649,n1650);
xor (n2503,n2504,n2409);
xor (n2504,n2406,n2407);
and (n2505,n2503,n2506);
or (n2506,n2507,n2512,n2516);
and (n2507,n2508,n2510);
xor (n2508,n2509,n1657);
xor (n2509,n1654,n1655);
xor (n2510,n2511,n2414);
xor (n2511,n2411,n2412);
and (n2512,n2510,n2513);
and (n2513,n2514,n2515);
xor (n2514,n1658,n1659);
xor (n2515,n2415,n2416);
and (n2516,n2508,n2513);
and (n2517,n2501,n2506);
and (n2518,n2494,n2499);
and (n2519,n2487,n2492);
and (n2520,n2480,n2485);
and (n2521,n2473,n2478);
and (n2522,n2466,n2471);
and (n2523,n2459,n2464);
and (n2524,n2452,n2457);
and (n2525,n2445,n2450);
and (n2526,n2438,n2443);
and (n2527,n2431,n2436);
and (n2528,n2529,n2531);
xor (n2529,n2530,n2436);
xor (n2530,n2431,n2433);
and (n2531,n2532,n2534);
xor (n2532,n2533,n2443);
xor (n2533,n2438,n2440);
and (n2534,n2535,n2537);
xor (n2535,n2536,n2450);
xor (n2536,n2445,n2447);
and (n2537,n2538,n2540);
xor (n2538,n2539,n2457);
xor (n2539,n2452,n2454);
and (n2540,n2541,n2543);
xor (n2541,n2542,n2464);
xor (n2542,n2459,n2461);
and (n2543,n2544,n2546);
xor (n2544,n2545,n2471);
xor (n2545,n2466,n2468);
and (n2546,n2547,n2549);
xor (n2547,n2548,n2478);
xor (n2548,n2473,n2475);
xor (n2549,n2550,n2485);
xor (n2550,n2480,n2482);
nand (n2551,n2552,n3401);
not (n2552,n2553);
or (n2553,n2554,n3400);
and (n2554,n2555,n2992);
xor (n2555,n2556,n2934);
xor (n2556,n2557,n2883);
xor (n2557,n2558,n2858);
or (n2558,n2559,n2857);
and (n2559,n2560,n2706);
xor (n2560,n2561,n2681);
xor (n2561,n2562,n2608);
xor (n2562,n2563,n2565);
xor (n2563,n2564,n1151);
xor (n2564,n1074,n1947);
xor (n2565,n2566,n2193);
xor (n2566,n2567,n2606);
or (n2567,n2568,n2605);
and (n2568,n2569,n2274);
xor (n2569,n2570,n1503);
and (n2570,n2571,n1511);
xor (n2571,n1510,n2572);
xor (n2572,n2573,n2582);
xor (n2573,n2574,n2581);
xor (n2574,n2575,n2580);
xor (n2575,n2576,n2578);
nor (n2576,n2577,n1017);
not (n2577,n2017);
nor (n2578,n2579,n1017);
not (n2579,n1236);
and (n2580,n2578,n1252);
and (n2581,n2576,n2033);
or (n2582,n2583,n2604);
and (n2583,n2584,n2595);
xor (n2584,n2585,n2589);
nor (n2585,n2586,n1017);
xnor (n2586,n2587,n2588);
not (n2587,n1367);
not (n2588,n1249);
and (n2589,n2590,n1018);
nand (n2590,n2591,n2593);
or (n2591,n2592,n2148);
not (n2592,n2030);
or (n2593,n2594,n2030);
not (n2594,n2148);
and (n2595,n2596,n1018);
or (n2596,n2597,n2602);
nor (n2597,n2598,n2601);
and (n2598,n2599,n2600);
not (n2599,n2153);
not (n2600,n2045);
not (n2601,n2033);
nor (n2602,n2603,n2577);
not (n2603,n2077);
and (n2604,n2585,n2589);
and (n2605,n2570,n1503);
xor (n2606,n2607,n1496);
xor (n2607,n1419,n1495);
or (n2608,n2609,n2680);
and (n2609,n2610,n2616);
xor (n2610,n2611,n2615);
or (n2611,n2612,n2614);
and (n2612,n2613,n1166);
xor (n2613,n1958,n1881);
and (n2614,n1958,n1881);
xor (n2615,n2569,n2274);
and (n2616,n2617,n1083);
xor (n2617,n1165,n2618);
or (n2618,n2619,n2679);
and (n2619,n2620,n2651);
xor (n2620,n2286,n2621);
and (n2621,n2622,n2645);
or (n2622,n2623,n2644);
and (n2623,n2624,n2642);
xor (n2624,n2625,n2633);
and (n2625,n2626,n1018);
nand (n2626,n2627,n2629,n2632);
or (n2627,n2628,n2599);
not (n2628,n2109);
or (n2629,n2630,n2631);
not (n2630,n2159);
not (n2631,n2081);
not (n2632,n2064);
and (n2633,n2634,n1018);
nand (n2634,n2635,n2638,n2641);
or (n2635,n2636,n2637);
not (n2636,n1328);
not (n2637,n1372);
or (n2638,n2639,n2640);
not (n2639,n1378);
not (n2640,n1300);
not (n2641,n1283);
nor (n2642,n2643,n1017);
xor (n2643,n1380,n2639);
and (n2644,n2625,n2633);
and (n2645,n2646,n1018);
nor (n2646,n2647,n2649);
and (n2647,n2648,n2033);
xor (n2648,n2599,n2600);
and (n2649,n2650,n2601);
not (n2650,n2648);
or (n2651,n2652,n2678);
and (n2652,n2653,n2292);
xor (n2653,n1527,n2654);
xor (n2654,n2655,n2670);
xor (n2655,n2656,n2663);
and (n2656,n2657,n1018);
nand (n2657,n2658,n2662);
or (n2658,n2659,n2639);
and (n2659,n2660,n2661);
not (n2660,n1268);
not (n2661,n1280);
not (n2662,n1267);
and (n2663,n2664,n1018);
nand (n2664,n2665,n2669);
or (n2665,n2666,n2630);
and (n2666,n2667,n2668);
not (n2667,n2049);
not (n2668,n2061);
not (n2669,n2048);
and (n2670,n2671,n1018);
nor (n2671,n2672,n2675);
and (n2672,n2673,n1252);
xor (n2673,n2637,n2674);
not (n2674,n1264);
and (n2675,n2676,n2677);
not (n2676,n2673);
not (n2677,n1252);
and (n2678,n1527,n2654);
and (n2679,n2286,n2621);
and (n2680,n2611,n2615);
xor (n2681,n2682,n2702);
xor (n2682,n2683,n2692);
xor (n2683,n2684,n2269);
xor (n2684,n1150,n2685);
and (n2685,n2686,n2689);
or (n2686,n2687,n2688);
and (n2687,n2573,n2582);
and (n2688,n2574,n2581);
or (n2689,n2690,n2691);
and (n2690,n2575,n2580);
and (n2691,n2576,n2578);
or (n2692,n2693,n2701);
and (n2693,n2694,n1158);
xor (n2694,n2695,n1952);
or (n2695,n2696,n2700);
and (n2696,n2697,n2203);
xor (n2697,n2698,n2699);
xor (n2698,n2571,n1511);
and (n2699,n1517,n1434);
and (n2700,n2698,n2699);
and (n2701,n2695,n1952);
or (n2702,n2703,n2705);
and (n2703,n2704,n1078);
xor (n2704,n1079,n1877);
and (n2705,n1079,n1877);
or (n2706,n2707,n2856);
and (n2707,n2708,n2733);
xor (n2708,n2709,n2710);
xor (n2709,n2610,n2616);
or (n2710,n2711,n2732);
and (n2711,n2712,n2719);
xor (n2712,n2713,n2718);
or (n2713,n2714,n2717);
and (n2714,n2715,n1891);
xor (n2715,n1174,n2716);
xor (n2716,n2620,n2651);
and (n2717,n1174,n2716);
xor (n2718,n2617,n1083);
or (n2719,n2720,n2731);
and (n2720,n2721,n1090);
xor (n2721,n1888,n2722);
or (n2722,n2723,n2730);
and (n2723,n2724,n1181);
xor (n2724,n2725,n2727);
xor (n2725,n2726,n1526);
xor (n2726,n2622,n2645);
and (n2727,n2728,n2298);
xor (n2728,n2729,n1534);
xor (n2729,n2624,n2642);
and (n2730,n2725,n2727);
and (n2731,n1888,n2722);
and (n2732,n2713,n2718);
or (n2733,n2734,n2855);
and (n2734,n2735,n2838);
xor (n2735,n2736,n2837);
or (n2736,n2737,n2836);
and (n2737,n2738,n1093);
xor (n2738,n2739,n2803);
or (n2739,n2740,n2802);
and (n2740,n2741,n1182);
xor (n2741,n2742,n2762);
xor (n2742,n2743,n2217);
xor (n2743,n1441,n2744);
or (n2744,n2745,n2761);
and (n2745,n2746,n1535);
xor (n2746,n2747,n2759);
or (n2747,n2748,n2754);
and (n2748,n2749,n1018);
or (n2749,n2750,n1299);
nor (n2750,n2751,n2753);
and (n2751,n2752,n2640);
not (n2752,n1312);
not (n2753,n1390);
and (n2754,n2755,n1018);
nand (n2755,n2756,n2757);
not (n2756,n2080);
nand (n2757,n2758,n2171);
or (n2758,n2081,n2093);
nor (n2759,n1017,n2760);
xor (n2760,n2161,n2630);
and (n2761,n2747,n2759);
and (n2762,n2763,n2801);
xor (n2763,n2764,n2799);
or (n2764,n2765,n2798);
and (n2765,n2766,n2304);
xor (n2766,n2767,n2776);
and (n2767,n2768,n2772);
xor (n2768,n2769,n1550);
and (n2769,n2770,n1018);
xnor (n2770,n2771,n2173);
not (n2771,n2171);
and (n2772,n2773,n2774);
and (n2773,n2416,n2171);
nor (n2774,n2775,n2753);
not (n2775,n1659);
or (n2776,n2777,n2797);
and (n2777,n2778,n2795);
xor (n2778,n2779,n2787);
and (n2779,n2780,n1018);
not (n2780,n2781);
nor (n2781,n2782,n2783);
and (n2782,n2171,n2113);
and (n2783,n2784,n2109);
nand (n2784,n2785,n2786);
not (n2785,n2177);
not (n2786,n2097);
and (n2787,n2788,n1018);
not (n2788,n2789);
nor (n2789,n2790,n2791);
and (n2790,n1390,n1332);
nor (n2791,n2792,n2636);
and (n2792,n2793,n2794);
not (n2793,n1396);
not (n2794,n1316);
and (n2795,n2796,n1018);
xnor (n2796,n2753,n1392);
and (n2797,n2779,n2787);
and (n2798,n2767,n2776);
and (n2799,n2800,n1455);
xor (n2800,n2231,n1542);
xor (n2801,n2728,n2298);
and (n2802,n2742,n2762);
or (n2803,n2804,n2835);
and (n2804,n2805,n1970);
xor (n2805,n2806,n2807);
xor (n2806,n2653,n2292);
or (n2807,n2808,n2834);
and (n2808,n2809,n2224);
xor (n2809,n1448,n2810);
or (n2810,n2811,n2833);
and (n2811,n2812,n1543);
xor (n2812,n2813,n2822);
and (n2813,n2814,n1018);
not (n2814,n2815);
nor (n2815,n2816,n2820);
and (n2816,n2817,n2065);
not (n2817,n2818);
xor (n2818,n2603,n2819);
not (n2819,n2165);
and (n2820,n2818,n2821);
not (n2821,n2065);
and (n2822,n2823,n1018);
nand (n2823,n2824,n2831);
or (n2824,n1284,n2825);
not (n2825,n2826);
nand (n2826,n2827,n2829);
or (n2827,n1296,n2828);
not (n2828,n1384);
or (n2829,n1384,n2830);
not (n2830,n1296);
or (n2831,n2826,n2832);
not (n2832,n1284);
and (n2833,n2813,n2822);
and (n2834,n1448,n2810);
and (n2835,n2806,n2807);
and (n2836,n2739,n2803);
xor (n2837,n2613,n1166);
xor (n2838,n2839,n1086);
xor (n2839,n1884,n2840);
xor (n2840,n2841,n2280);
xor (n2841,n1427,n2842);
or (n2842,n2843,n2854);
and (n2843,n2844,n2851);
xor (n2844,n2845,n2846);
xor (n2845,n2584,n2595);
and (n2846,n2847,n1018);
or (n2847,n2848,n2850);
nor (n2848,n2849,n2677);
and (n2849,n2637,n2674);
nor (n2850,n2830,n2579);
or (n2851,n2852,n2853);
and (n2852,n2655,n2670);
and (n2853,n2656,n2663);
and (n2854,n2845,n2846);
and (n2855,n2736,n2837);
and (n2856,n2709,n2710);
and (n2857,n2561,n2681);
xor (n2858,n2859,n2880);
xor (n2859,n2860,n2867);
xor (n2860,n2861,n2864);
xor (n2861,n2862,n2863);
and (n2862,n2684,n2269);
and (n2863,n2607,n1496);
or (n2864,n2865,n2866);
and (n2865,n2564,n1151);
and (n2866,n1074,n1947);
and (n2867,n2868,n2875);
xor (n2868,n2869,n1871);
or (n2869,n2870,n2874);
and (n2870,n2871,n1874);
xor (n2871,n1422,n2872);
xor (n2872,n2873,n1502);
xor (n2873,n2686,n2689);
and (n2874,n1422,n2872);
and (n2875,n2876,n2196);
xor (n2876,n1157,n2877);
or (n2877,n2878,n2879);
and (n2878,n2841,n2280);
and (n2879,n1427,n2842);
or (n2880,n2881,n2882);
and (n2881,n2682,n2702);
and (n2882,n2683,n2692);
xor (n2883,n2884,n2896);
xor (n2884,n2885,n2888);
or (n2885,n2886,n2887);
and (n2886,n2562,n2608);
and (n2887,n2563,n2565);
xor (n2888,n2889,n2894);
xor (n2889,n2890,n2893);
or (n2890,n2891,n2892);
and (n2891,n2566,n2193);
and (n2892,n2567,n2606);
xor (n2893,n1413,n1068);
xor (n2894,n2895,n1071);
xor (n2895,n1676,n2014);
or (n2896,n2897,n2933);
and (n2897,n2898,n2909);
xor (n2898,n2899,n2908);
or (n2899,n2900,n2907);
and (n2900,n2901,n2906);
xor (n2901,n2902,n2905);
or (n2902,n2903,n2904);
and (n2903,n2839,n1086);
and (n2904,n1884,n2840);
xor (n2905,n2871,n1874);
xor (n2906,n2694,n1158);
and (n2907,n2902,n2905);
xor (n2908,n2868,n2875);
or (n2909,n2910,n2932);
and (n2910,n2911,n2931);
xor (n2911,n2912,n2913);
xor (n2912,n2876,n2196);
or (n2913,n2914,n2930);
and (n2914,n2915,n2925);
xor (n2915,n2916,n2917);
xor (n2916,n2697,n2203);
or (n2917,n2918,n2924);
and (n2918,n2919,n2210);
xor (n2919,n2920,n2923);
or (n2920,n2921,n2922);
and (n2921,n2743,n2217);
and (n2922,n1441,n2744);
xor (n2923,n2844,n2851);
and (n2924,n2920,n2923);
or (n2925,n2926,n2929);
and (n2926,n2927,n1964);
xor (n2927,n1173,n2928);
xor (n2928,n1517,n1434);
and (n2929,n1173,n2928);
and (n2930,n2916,n2917);
xor (n2931,n2704,n1078);
and (n2932,n2912,n2913);
and (n2933,n2899,n2908);
or (n2934,n2935,n2991);
and (n2935,n2936,n2990);
xor (n2936,n2937,n2989);
or (n2937,n2938,n2988);
and (n2938,n2939,n2942);
xor (n2939,n2940,n2941);
xor (n2940,n2911,n2931);
xor (n2941,n2901,n2906);
or (n2942,n2943,n2987);
and (n2943,n2944,n2977);
xor (n2944,n2945,n2976);
or (n2945,n2946,n2975);
and (n2946,n2947,n2950);
xor (n2947,n2948,n2949);
xor (n2948,n2927,n1964);
xor (n2949,n2919,n2210);
or (n2950,n2951,n2974);
and (n2951,n2952,n1898);
xor (n2952,n2953,n2956);
and (n2953,n2954,n1976);
xor (n2954,n1189,n2955);
xor (n2955,n2746,n1535);
or (n2956,n2957,n2973);
and (n2957,n2958,n1190);
xor (n2958,n2959,n2960);
xor (n2959,n2809,n2224);
or (n2960,n2961,n2972);
and (n2961,n2962,n2968);
xor (n2962,n2963,n2964);
xor (n2963,n2812,n1543);
nand (n2964,n2965,n2747);
or (n2965,n2966,n2967);
not (n2966,n2754);
not (n2967,n2748);
or (n2968,n2969,n2971);
and (n2969,n2970,n1462);
xor (n2970,n1551,n2310);
and (n2971,n1551,n2310);
and (n2972,n2963,n2964);
and (n2973,n2959,n2960);
and (n2974,n2953,n2956);
and (n2975,n2948,n2949);
xor (n2976,n2915,n2925);
or (n2977,n2978,n2986);
and (n2978,n2979,n2985);
xor (n2979,n2980,n2981);
xor (n2980,n2715,n1891);
or (n2981,n2982,n2984);
and (n2982,n2983,n1100);
xor (n2983,n1097,n1895);
and (n2984,n1097,n1895);
xor (n2985,n2721,n1090);
and (n2986,n2980,n2981);
and (n2987,n2945,n2976);
and (n2988,n2940,n2941);
xor (n2989,n2898,n2909);
xor (n2990,n2560,n2706);
and (n2991,n2937,n2989);
or (n2992,n2993,n3399);
and (n2993,n2994,n3070);
xor (n2994,n2995,n2996);
xor (n2995,n2936,n2990);
or (n2996,n2997,n3069);
and (n2997,n2998,n3068);
xor (n2998,n2999,n3067);
or (n2999,n3000,n3066);
and (n3000,n3001,n3065);
xor (n3001,n3002,n3003);
xor (n3002,n2712,n2719);
or (n3003,n3004,n3064);
and (n3004,n3005,n3041);
xor (n3005,n3006,n3007);
xor (n3006,n2738,n1093);
or (n3007,n3008,n3040);
and (n3008,n3009,n3012);
xor (n3009,n3010,n3011);
xor (n3010,n2724,n1181);
xor (n3011,n2805,n1970);
or (n3012,n3013,n3039);
and (n3013,n3014,n1902);
xor (n3014,n3015,n1104);
and (n3015,n3016,n3038);
and (n3016,n3017,n3022);
or (n3017,n3018,n3021);
and (n3018,n3019,n2245);
xor (n3019,n1559,n3020);
xor (n3020,n2773,n2774);
and (n3021,n1559,n3020);
and (n3022,n3023,n3031);
xor (n3023,n3024,n1213);
and (n3024,n3025,n1018);
nand (n3025,n3026,n3030);
or (n3026,n2786,n3027);
nand (n3027,n3028,n3029);
or (n3028,n2177,n2628);
nand (n3029,n2177,n2628);
nand (n3030,n3027,n2786);
and (n3031,n3032,n1018);
nand (n3032,n3033,n3037);
or (n3033,n2794,n3034);
nand (n3034,n3035,n3036);
or (n3035,n1328,n2793);
nand (n3036,n1328,n2793);
nand (n3037,n3034,n2794);
xor (n3038,n2766,n2304);
and (n3039,n3015,n1104);
and (n3040,n3010,n3011);
or (n3041,n3042,n3063);
and (n3042,n3043,n3062);
xor (n3043,n3044,n3061);
or (n3044,n3045,n3060);
and (n3045,n3046,n1107);
xor (n3046,n3047,n3059);
or (n3047,n3048,n3058);
and (n3048,n3049,n1198);
xor (n3049,n3050,n3051);
xor (n3050,n2800,n1455);
or (n3051,n3052,n3057);
and (n3052,n3053,n2238);
xor (n3053,n3054,n3055);
xor (n3054,n2778,n2795);
and (n3055,n2316,n3056);
and (n3056,n2321,n1999);
and (n3057,n3054,n3055);
and (n3058,n3050,n3051);
xor (n3059,n2763,n2801);
and (n3060,n3047,n3059);
xor (n3061,n2741,n1182);
xor (n3062,n2983,n1100);
and (n3063,n3044,n3061);
and (n3064,n3006,n3007);
xor (n3065,n2735,n2838);
and (n3066,n3002,n3003);
xor (n3067,n2708,n2733);
xor (n3068,n2939,n2942);
and (n3069,n2999,n3067);
or (n3070,n3071,n3398);
and (n3071,n3072,n3167);
xor (n3072,n3073,n3074);
xor (n3073,n2998,n3068);
or (n3074,n3075,n3166);
and (n3075,n3076,n3165);
xor (n3076,n3077,n3078);
xor (n3077,n2944,n2977);
or (n3078,n3079,n3164);
and (n3079,n3080,n3163);
xor (n3080,n3081,n3082);
xor (n3081,n2947,n2950);
or (n3082,n3083,n3162);
and (n3083,n3084,n3100);
xor (n3084,n3085,n3099);
or (n3085,n3086,n3098);
and (n3086,n3087,n3089);
xor (n3087,n1905,n3088);
xor (n3088,n2954,n1976);
or (n3089,n3090,n3097);
and (n3090,n3091,n1111);
xor (n3091,n3092,n1982);
or (n3092,n3093,n3096);
and (n3093,n3094,n1206);
xor (n3094,n1988,n3095);
xor (n3095,n2768,n2772);
and (n3096,n1988,n3095);
and (n3097,n3092,n1982);
and (n3098,n1905,n3088);
xor (n3099,n2952,n1898);
or (n3100,n3101,n3161);
and (n3101,n3102,n3160);
xor (n3102,n3103,n3104);
xor (n3103,n2958,n1190);
or (n3104,n3105,n3159);
and (n3105,n3106,n1912);
xor (n3106,n1909,n3107);
or (n3107,n3108,n3158);
and (n3108,n3109,n3135);
xor (n3109,n3110,n3111);
xor (n3110,n2970,n1462);
or (n3111,n3112,n3134);
and (n3112,n3113,n1469);
xor (n3113,n3114,n3124);
or (n3114,n3115,n3123);
and (n3115,n3116,n3118);
xor (n3116,n3117,n2251);
xor (n3117,n2321,n1999);
and (n3118,n3119,n1018);
nand (n3119,n3120,n3122);
or (n3120,n1401,n3121);
not (n3121,n1344);
nand (n3122,n1401,n3121);
and (n3123,n3117,n2251);
or (n3124,n3125,n3133);
and (n3125,n3126,n3129);
xor (n3126,n3127,n3128);
and (n3127,n1332,n1018);
and (n3128,n2113,n1018);
and (n3129,n3130,n1018);
xor (n3130,n3131,n3132);
not (n3131,n2125);
not (n3132,n2182);
and (n3133,n3127,n3128);
and (n3134,n3114,n3124);
or (n3135,n3136,n3157);
and (n3136,n3137,n1994);
xor (n3137,n3138,n3155);
or (n3138,n3139,n3154);
and (n3139,n3140,n1219);
xor (n3140,n3141,n3149);
or (n3141,n3142,n3148);
and (n3142,n3143,n3146);
xor (n3143,n3144,n2256);
nor (n3144,n3145,n1017);
not (n3145,n1359);
nor (n3146,n3147,n1017);
not (n3147,n2140);
and (n3148,n3144,n2256);
and (n3149,n3150,n3152);
nor (n3150,n3151,n1017);
not (n3151,n1347);
nor (n3152,n3153,n1017);
not (n3153,n2128);
and (n3154,n3141,n3149);
xor (n3155,n3156,n1558);
xor (n3156,n2316,n3056);
and (n3157,n3138,n3155);
and (n3158,n3110,n3111);
and (n3159,n1909,n3107);
xor (n3160,n3014,n1902);
and (n3161,n3103,n3104);
and (n3162,n3085,n3099);
xor (n3163,n2979,n2985);
and (n3164,n3081,n3082);
xor (n3165,n3001,n3065);
and (n3166,n3077,n3078);
or (n3167,n3168,n3397);
and (n3168,n3169,n3221);
xor (n3169,n3170,n3220);
or (n3170,n3171,n3219);
and (n3171,n3172,n3218);
xor (n3172,n3173,n3217);
or (n3173,n3174,n3216);
and (n3174,n3175,n3215);
xor (n3175,n3176,n3214);
or (n3176,n3177,n3213);
and (n3177,n3178,n3212);
xor (n3178,n3179,n3206);
or (n3179,n3180,n3205);
and (n3180,n3181,n3200);
xor (n3181,n3182,n3184);
xor (n3182,n3183,n1197);
xor (n3183,n3016,n3038);
or (n3184,n3185,n3199);
and (n3185,n3186,n1118);
xor (n3186,n3187,n3197);
or (n3187,n3188,n3196);
and (n3188,n3189,n3195);
xor (n3189,n1214,n3190);
or (n3190,n3191,n3194);
and (n3191,n3192,n1564);
xor (n3192,n3193,n1475);
xor (n3193,n3126,n3129);
and (n3194,n3193,n1475);
xor (n3195,n3019,n2245);
and (n3196,n1214,n3190);
xor (n3197,n3198,n1205);
xor (n3198,n3017,n3022);
and (n3199,n3187,n3197);
or (n3200,n3201,n3204);
and (n3201,n3202,n1121);
xor (n3202,n1916,n3203);
xor (n3203,n3053,n2238);
and (n3204,n1916,n3203);
and (n3205,n3182,n3184);
or (n3206,n3207,n3211);
and (n3207,n3208,n1114);
xor (n3208,n3209,n3210);
xor (n3209,n2962,n2968);
xor (n3210,n3049,n1198);
and (n3211,n3209,n3210);
xor (n3212,n3046,n1107);
and (n3213,n3179,n3206);
xor (n3214,n3009,n3012);
xor (n3215,n3043,n3062);
and (n3216,n3176,n3214);
xor (n3217,n3005,n3041);
xor (n3218,n3080,n3163);
and (n3219,n3173,n3217);
xor (n3220,n3076,n3165);
or (n3221,n3222,n3396);
and (n3222,n3223,n3288);
xor (n3223,n3224,n3287);
or (n3224,n3225,n3286);
and (n3225,n3226,n3285);
xor (n3226,n3227,n3228);
xor (n3227,n3084,n3100);
or (n3228,n3229,n3284);
and (n3229,n3230,n3283);
xor (n3230,n3231,n3232);
xor (n3231,n3087,n3089);
or (n3232,n3233,n3282);
and (n3233,n3234,n3246);
xor (n3234,n3235,n3236);
xor (n3235,n3091,n1111);
or (n3236,n3237,n3245);
and (n3237,n3238,n1919);
xor (n3238,n3239,n3240);
xor (n3239,n3094,n1206);
or (n3240,n3241,n3244);
and (n3241,n3242,n1125);
xor (n3242,n1923,n3243);
xor (n3243,n3023,n3031);
and (n3244,n1923,n3243);
and (n3245,n3239,n3240);
or (n3246,n3247,n3281);
and (n3247,n3248,n3266);
xor (n3248,n3249,n3250);
xor (n3249,n3109,n3135);
or (n3250,n3251,n3265);
and (n3251,n3252,n1925);
xor (n3252,n3253,n3264);
or (n3253,n3254,n3263);
and (n3254,n3255,n1131);
xor (n3255,n3256,n3257);
xor (n3256,n3116,n3118);
or (n3257,n3258,n3262);
and (n3258,n3259,n3261);
xor (n3259,n3260,n1934);
and (n3260,n1659,n2415);
xor (n3261,n3150,n3152);
and (n3262,n3260,n1934);
and (n3263,n3256,n3257);
xor (n3264,n3113,n1469);
and (n3265,n3253,n3264);
or (n3266,n3267,n3280);
and (n3267,n3268,n1127);
xor (n3268,n3269,n3270);
xor (n3269,n3137,n1994);
or (n3270,n3271,n3279);
and (n3271,n3272,n1929);
xor (n3272,n3273,n3274);
xor (n3273,n3192,n1564);
or (n3274,n3275,n3278);
and (n3275,n3276,n1480);
xor (n3276,n1136,n3277);
xor (n3277,n3143,n3146);
and (n3278,n1136,n3277);
and (n3279,n3273,n3274);
and (n3280,n3269,n3270);
and (n3281,n3249,n3250);
and (n3282,n3235,n3236);
xor (n3283,n3102,n3160);
and (n3284,n3231,n3232);
xor (n3285,n3175,n3215);
and (n3286,n3227,n3228);
xor (n3287,n3172,n3218);
nand (n3288,n3289,n3395);
or (n3289,n3290,n3305);
nor (n3290,n3291,n3292);
xor (n3291,n3226,n3285);
or (n3292,n3293,n3304);
and (n3293,n3294,n3303);
xor (n3294,n3295,n3296);
xor (n3295,n3178,n3212);
or (n3296,n3297,n3302);
and (n3297,n3298,n3301);
xor (n3298,n3299,n3300);
xor (n3299,n3106,n1912);
xor (n3300,n3208,n1114);
xor (n3301,n3181,n3200);
and (n3302,n3299,n3300);
xor (n3303,n3230,n3283);
and (n3304,n3295,n3296);
and (n3305,n3306,n3394);
nand (n3306,n3307,n3322);
or (n3307,n3308,n3309);
xor (n3308,n3294,n3303);
or (n3309,n3310,n3321);
and (n3310,n3311,n3320);
xor (n3311,n3312,n3319);
or (n3312,n3313,n3318);
and (n3313,n3314,n3317);
xor (n3314,n3315,n3316);
xor (n3315,n3202,n1121);
xor (n3316,n3186,n1118);
xor (n3317,n3238,n1919);
and (n3318,n3315,n3316);
xor (n3319,n3234,n3246);
xor (n3320,n3298,n3301);
and (n3321,n3312,n3319);
nand (n3322,n3323,n3387);
nand (n3323,n3324,n3359,n3362);
or (n3324,n3325,n3358);
or (n3325,n3326,n3357);
and (n3326,n3327,n3356);
xor (n3327,n3328,n3345);
or (n3328,n3329,n3344);
and (n3329,n3330,n3343);
xor (n3330,n3331,n3332);
xor (n3331,n3252,n1925);
or (n3332,n3333,n3342);
and (n3333,n3334,n3341);
xor (n3334,n3335,n3336);
xor (n3335,n3255,n1131);
or (n3336,n3337,n3340);
and (n3337,n3338,n1936);
xor (n3338,n3339,n1138);
xor (n3339,n3259,n3261);
and (n3340,n3339,n1138);
xor (n3341,n3272,n1929);
and (n3342,n3335,n3336);
xor (n3343,n3268,n1127);
and (n3344,n3331,n3332);
or (n3345,n3346,n3355);
and (n3346,n3347,n3354);
xor (n3347,n3348,n3353);
or (n3348,n3349,n3352);
and (n3349,n3350,n1133);
xor (n3350,n1931,n3351);
xor (n3351,n3140,n1219);
and (n3352,n1931,n3351);
xor (n3353,n3189,n3195);
xor (n3354,n3242,n1125);
and (n3355,n3348,n3353);
xor (n3356,n3248,n3266);
and (n3357,n3328,n3345);
xor (n3358,n3311,n3320);
or (n3359,n3360,n3361);
xor (n3360,n3327,n3356);
xor (n3361,n3314,n3317);
nand (n3362,n3363,n3383);
or (n3363,n3364,n3367);
nor (n3364,n3365,n3366);
xor (n3365,n3330,n3343);
xor (n3366,n3347,n3354);
nand (n3367,n3368,n3371,n3374);
or (n3368,n3369,n3370);
xor (n3369,n3350,n1133);
xor (n3370,n3334,n3341);
or (n3371,n3372,n3373);
xor (n3372,n3276,n1480);
xor (n3373,n3338,n1936);
nand (n3374,n3375,n3378);
or (n3375,n3376,n3377);
not (n3376,n3372);
not (n3377,n3373);
nor (n3378,n3379,n3382);
and (n3379,n3380,n3381);
xor (n3380,n1659,n2415);
or (n3381,n1658,n2416);
and (n3382,n1658,n2416);
nor (n3383,n3384,n3386);
and (n3384,n3385,n3369,n3370);
not (n3385,n3364);
and (n3386,n3365,n3366);
nor (n3387,n3388,n3392);
and (n3388,n3358,n3389);
nand (n3389,n3390,n3391);
not (n3390,n3325);
nand (n3391,n3360,n3361);
and (n3392,n3393,n3325);
not (n3393,n3391);
nand (n3394,n3308,n3309);
nand (n3395,n3291,n3292);
and (n3396,n3224,n3287);
and (n3397,n3170,n3220);
and (n3398,n3073,n3074);
and (n3399,n2995,n2996);
and (n3400,n2556,n2934);
nand (n3401,n3402,n3428);
or (n3402,n3403,n3424);
not (n3403,n3404);
nand (n3404,n3405,n3409);
not (n3405,n3406);
or (n3406,n3407,n3408);
and (n3407,n2884,n2896);
and (n3408,n2885,n2888);
nor (n3409,n3410,n3423);
not (n3410,n3411);
nor (n3411,n3412,n3420);
not (n3412,n3413);
nor (n3413,n3414,n3415);
and (n3414,n2895,n1071);
not (n3415,n3416);
nor (n3416,n3417,n3418);
and (n3417,n1413,n1068);
not (n3418,n3419);
xnor (n3419,n6,n1233);
or (n3420,n3421,n3422);
and (n3421,n2889,n2894);
and (n3422,n2890,n2893);
and (n3423,n2859,n2880);
not (n3424,n3425);
or (n3425,n3426,n3427);
and (n3426,n2557,n2883);
and (n3427,n2558,n2858);
or (n3428,n3425,n3404);
endmodule
