module top (out,n9,n21,n23,n24,n26,n28,n29,n34,n41
        ,n48,n54,n57,n58,n76,n77,n89,n90,n96,n97
        ,n116,n117,n123,n124,n129,n135,n144,n153,n168,n181
        ,n187,n206,n212,n672,n690,n697,n701,n706,n712,n718
        ,n724,n729,n751,n762,n777,n788,n799);
output out;
input n9;
input n21;
input n23;
input n24;
input n26;
input n28;
input n29;
input n34;
input n41;
input n48;
input n54;
input n57;
input n58;
input n76;
input n77;
input n89;
input n90;
input n96;
input n97;
input n116;
input n117;
input n123;
input n124;
input n129;
input n135;
input n144;
input n153;
input n168;
input n181;
input n187;
input n206;
input n212;
input n672;
input n690;
input n697;
input n701;
input n706;
input n712;
input n718;
input n724;
input n729;
input n751;
input n762;
input n777;
input n788;
input n799;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n22;
wire n25;
wire n27;
wire n30;
wire n31;
wire n32;
wire n33;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n55;
wire n56;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n125;
wire n126;
wire n127;
wire n128;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n143;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n698;
wire n699;
wire n700;
wire n702;
wire n703;
wire n704;
wire n705;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n725;
wire n726;
wire n727;
wire n728;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
xor (out,n0,n813);
nand (n0,n1,n812);
or (n1,n2,n674);
not (n2,n3);
nand (n3,n4,n673);
not (n4,n5);
nor (n5,n6,n672);
nand (n6,n7,n98);
or (n7,n8,n10);
not (n8,n9);
not (n10,n11);
xor (n11,n12,n94);
xor (n12,n13,n91);
xor (n13,n14,n87);
xor (n14,n15,n78);
xor (n15,n16,n74);
xor (n16,n17,n59);
xor (n17,n18,n55);
xor (n18,n19,n30);
xor (n19,n20,n25);
and (n20,n21,n22);
wire s0n22,s1n22,notn22;
or (n22,s0n22,s1n22);
not(notn22,n9);
and (s0n22,notn22,n23);
and (s1n22,n9,n24);
and (n25,n26,n27);
wire s0n27,s1n27,notn27;
or (n27,s0n27,s1n27);
not(notn27,n9);
and (s0n27,notn27,n28);
and (s1n27,n9,n29);
or (n30,n31,n35);
and (n31,n32,n33);
and (n32,n26,n22);
and (n33,n34,n27);
and (n35,n36,n37);
xor (n36,n32,n33);
or (n37,n38,n42);
and (n38,n39,n40);
and (n39,n34,n22);
and (n40,n41,n27);
and (n42,n43,n44);
xor (n43,n39,n40);
or (n44,n45,n49);
and (n45,n46,n47);
and (n46,n41,n22);
and (n47,n48,n27);
and (n49,n50,n51);
xor (n50,n46,n47);
and (n51,n52,n53);
and (n52,n48,n22);
and (n53,n54,n27);
and (n55,n34,n56);
wire s0n56,s1n56,notn56;
or (n56,s0n56,s1n56);
not(notn56,n9);
and (s0n56,notn56,n57);
and (s1n56,n9,n58);
or (n59,n60,n63);
and (n60,n61,n62);
xor (n61,n36,n37);
and (n62,n41,n56);
and (n63,n64,n65);
xor (n64,n61,n62);
or (n65,n66,n69);
and (n66,n67,n68);
xor (n67,n43,n44);
and (n68,n48,n56);
and (n69,n70,n71);
xor (n70,n67,n68);
and (n71,n72,n73);
xor (n72,n50,n51);
and (n73,n54,n56);
and (n74,n41,n75);
wire s0n75,s1n75,notn75;
or (n75,s0n75,s1n75);
not(notn75,n9);
and (s0n75,notn75,n76);
and (s1n75,n9,n77);
or (n78,n79,n82);
and (n79,n80,n81);
xor (n80,n64,n65);
and (n81,n48,n75);
and (n82,n83,n84);
xor (n83,n80,n81);
and (n84,n85,n86);
xor (n85,n70,n71);
and (n86,n54,n75);
and (n87,n48,n88);
wire s0n88,s1n88,notn88;
or (n88,s0n88,s1n88);
not(notn88,n9);
and (s0n88,notn88,n89);
and (s1n88,n9,n90);
and (n91,n92,n93);
xor (n92,n83,n84);
and (n93,n54,n88);
and (n94,n54,n95);
wire s0n95,s1n95,notn95;
or (n95,s0n95,s1n95);
not(notn95,n9);
and (s0n95,notn95,n96);
and (s1n95,n9,n97);
nand (n98,n99,n8);
nand (n99,n100,n671);
or (n100,n101,n339);
not (n101,n102);
nand (n102,n103,n338);
not (n103,n104);
nor (n104,n105,n292);
xor (n105,n106,n252);
xor (n106,n107,n171);
xor (n107,n108,n149);
xor (n108,n109,n138);
nand (n109,n110,n132);
or (n110,n111,n126);
nand (n111,n112,n120);
nor (n112,n113,n118);
and (n113,n114,n95);
not (n114,n115);
wire s0n115,s1n115,notn115;
or (n115,s0n115,s1n115);
not(notn115,n9);
and (s0n115,notn115,n116);
and (s1n115,n9,n117);
and (n118,n115,n119);
not (n119,n95);
nand (n120,n121,n125);
or (n121,n114,n122);
wire s0n122,s1n122,notn122;
or (n122,s0n122,s1n122);
not(notn122,n9);
and (s0n122,notn122,n123);
and (s1n122,n9,n124);
nand (n125,n122,n114);
nor (n126,n127,n130);
and (n127,n128,n129);
not (n128,n122);
and (n130,n122,n131);
not (n131,n129);
or (n132,n112,n133);
nor (n133,n134,n136);
and (n134,n135,n128);
and (n136,n137,n122);
not (n137,n135);
nor (n138,n139,n145);
nand (n139,n122,n140);
not (n140,n141);
wire s0n141,s1n141,notn141;
or (n141,s0n141,s1n141);
not(notn141,n9);
and (s0n141,notn141,1'b0);
and (s1n141,n9,n143);
and (n143,n144,n124);
nor (n145,n146,n148);
and (n146,n141,n147);
not (n147,n21);
and (n148,n140,n21);
nand (n149,n150,n161);
or (n150,n151,n156);
nor (n151,n152,n154);
and (n152,n119,n153);
and (n154,n95,n155);
not (n155,n153);
not (n156,n157);
nand (n157,n158,n160);
or (n158,n159,n75);
not (n159,n88);
nand (n160,n75,n159);
or (n161,n162,n166);
nand (n162,n156,n163);
nand (n163,n164,n165);
or (n164,n159,n95);
nand (n165,n95,n159);
nor (n166,n167,n169);
and (n167,n119,n168);
and (n169,n95,n170);
not (n170,n168);
xor (n171,n172,n228);
xor (n172,n173,n215);
xor (n173,n174,n191);
nand (n174,n175,n184);
or (n175,n176,n179);
not (n176,n177);
nor (n177,n178,n22);
not (n178,n27);
nor (n179,n180,n182);
and (n180,n178,n181);
and (n182,n27,n183);
not (n183,n181);
or (n184,n185,n190);
nor (n185,n186,n188);
and (n186,n178,n187);
and (n188,n27,n189);
not (n189,n187);
not (n190,n22);
nand (n191,n192,n209);
or (n192,n193,n203);
not (n193,n194);
and (n194,n195,n199);
nand (n195,n196,n198);
or (n196,n197,n75);
not (n197,n56);
nand (n198,n75,n197);
not (n199,n200);
nand (n200,n201,n202);
or (n201,n197,n27);
nand (n202,n27,n197);
nor (n203,n204,n207);
and (n204,n205,n206);
not (n205,n75);
and (n207,n75,n208);
not (n208,n206);
or (n209,n210,n199);
nor (n210,n211,n213);
and (n211,n205,n212);
and (n213,n75,n214);
not (n214,n212);
and (n215,n216,n222);
nand (n216,n217,n221);
or (n217,n176,n218);
nor (n218,n219,n220);
and (n219,n178,n212);
and (n220,n27,n214);
or (n221,n179,n190);
nand (n222,n223,n227);
or (n223,n193,n224);
nor (n224,n225,n226);
and (n225,n205,n153);
and (n226,n75,n155);
or (n227,n203,n199);
or (n228,n229,n251);
and (n229,n230,n245);
xor (n230,n231,n240);
nand (n231,n232,n237);
or (n232,n233,n111);
not (n233,n234);
nor (n234,n235,n236);
and (n235,n21,n122);
and (n236,n147,n128);
nand (n237,n238,n239);
not (n238,n126);
not (n239,n112);
nor (n240,n139,n241);
nor (n241,n242,n244);
and (n242,n141,n243);
not (n243,n26);
and (n244,n140,n26);
nand (n245,n246,n250);
or (n246,n162,n247);
nor (n247,n248,n249);
and (n248,n119,n135);
and (n249,n95,n137);
or (n250,n156,n166);
and (n251,n231,n240);
or (n252,n253,n291);
and (n253,n254,n269);
xor (n254,n255,n256);
xor (n255,n216,n222);
and (n256,n257,n263);
nand (n257,n258,n262);
or (n258,n176,n259);
nor (n259,n260,n261);
and (n260,n178,n206);
and (n261,n27,n208);
or (n262,n218,n190);
nand (n263,n264,n268);
or (n264,n193,n265);
nor (n265,n266,n267);
and (n266,n205,n168);
and (n267,n75,n170);
or (n268,n199,n224);
or (n269,n270,n290);
and (n270,n271,n284);
xor (n271,n272,n279);
nand (n272,n273,n278);
or (n273,n274,n111);
not (n274,n275);
nor (n275,n276,n277);
and (n276,n26,n122);
and (n277,n243,n128);
nand (n278,n239,n234);
nor (n279,n139,n280);
nor (n280,n281,n283);
and (n281,n141,n282);
not (n282,n34);
and (n283,n140,n34);
nand (n284,n285,n289);
or (n285,n162,n286);
nor (n286,n287,n288);
and (n287,n119,n129);
and (n288,n95,n131);
or (n289,n156,n247);
and (n290,n272,n279);
and (n291,n255,n256);
or (n292,n293,n337);
and (n293,n294,n297);
xor (n294,n295,n296);
xor (n295,n230,n245);
xor (n296,n254,n269);
or (n297,n298,n336);
and (n298,n299,n314);
xor (n299,n300,n301);
xor (n300,n257,n263);
and (n301,n302,n308);
nand (n302,n303,n307);
or (n303,n176,n304);
nor (n304,n305,n306);
and (n305,n178,n153);
and (n306,n27,n155);
or (n307,n259,n190);
nand (n308,n309,n313);
or (n309,n193,n310);
nor (n310,n311,n312);
and (n311,n205,n135);
and (n312,n75,n137);
or (n313,n265,n199);
or (n314,n315,n335);
and (n315,n316,n329);
xor (n316,n317,n324);
nand (n317,n318,n323);
or (n318,n319,n111);
not (n319,n320);
nor (n320,n321,n322);
and (n321,n34,n122);
and (n322,n282,n128);
nand (n323,n239,n275);
nor (n324,n139,n325);
nor (n325,n326,n328);
and (n326,n141,n327);
not (n327,n41);
and (n328,n140,n41);
nand (n329,n330,n334);
or (n330,n162,n331);
nor (n331,n332,n333);
and (n332,n119,n21);
and (n333,n95,n147);
or (n334,n156,n286);
and (n335,n317,n324);
and (n336,n300,n301);
and (n337,n295,n296);
nand (n338,n105,n292);
not (n339,n340);
nand (n340,n341,n670);
or (n341,n342,n376);
not (n342,n343);
nand (n343,n344,n346);
not (n344,n345);
xor (n345,n294,n297);
not (n346,n347);
or (n347,n348,n375);
and (n348,n349,n352);
xor (n349,n350,n351);
xor (n350,n271,n284);
xor (n351,n299,n314);
and (n352,n353,n354);
xor (n353,n302,n308);
or (n354,n355,n374);
and (n355,n356,n368);
xor (n356,n357,n363);
nand (n357,n358,n362);
or (n358,n359,n111);
nor (n359,n360,n361);
and (n360,n41,n128);
and (n361,n327,n122);
nand (n362,n320,n239);
nor (n363,n139,n364);
nor (n364,n365,n367);
and (n365,n141,n366);
not (n366,n48);
and (n367,n140,n48);
nand (n368,n369,n373);
or (n369,n176,n370);
nor (n370,n371,n372);
and (n371,n178,n168);
and (n372,n27,n170);
or (n373,n304,n190);
and (n374,n357,n363);
and (n375,n350,n351);
not (n376,n377);
nand (n377,n378,n530,n669);
nand (n378,n379,n523);
nand (n379,n380,n522);
or (n380,n381,n511);
nor (n381,n382,n510);
and (n382,n383,n482);
not (n383,n384);
nor (n384,n385,n465);
or (n385,n386,n464);
and (n386,n387,n435);
xor (n387,n388,n422);
or (n388,n389,n421);
and (n389,n390,n412);
xor (n390,n391,n402);
nand (n391,n392,n398);
or (n392,n393,n111);
not (n393,n394);
nand (n394,n395,n396);
or (n395,n128,n54);
or (n396,n122,n397);
not (n397,n54);
or (n398,n112,n399);
nor (n399,n400,n401);
and (n400,n48,n128);
and (n401,n366,n122);
nand (n402,n403,n408);
or (n403,n404,n193);
not (n404,n405);
nand (n405,n406,n407);
or (n406,n75,n243);
or (n407,n205,n26);
nand (n408,n200,n409);
nor (n409,n410,n411);
and (n410,n21,n75);
and (n411,n147,n205);
nand (n412,n413,n417);
or (n413,n162,n414);
nor (n414,n415,n416);
and (n415,n119,n41);
and (n416,n95,n327);
or (n417,n156,n418);
nor (n418,n419,n420);
and (n419,n119,n34);
and (n420,n95,n282);
and (n421,n391,n402);
xor (n422,n423,n432);
xor (n423,n424,n426);
and (n424,n425,n54);
not (n425,n139);
nand (n426,n427,n431);
or (n427,n176,n428);
nor (n428,n429,n430);
and (n429,n137,n27);
and (n430,n135,n178);
or (n431,n370,n190);
nand (n432,n433,n434);
or (n433,n111,n399);
or (n434,n112,n359);
xor (n435,n436,n450);
xor (n436,n437,n444);
nand (n437,n438,n440);
or (n438,n193,n439);
not (n439,n409);
or (n440,n199,n441);
nor (n441,n442,n443);
and (n442,n205,n129);
and (n443,n75,n131);
nand (n444,n445,n446);
or (n445,n162,n418);
or (n446,n156,n447);
nor (n447,n448,n449);
and (n448,n119,n26);
and (n449,n95,n243);
and (n450,n451,n456);
nor (n451,n452,n128);
nor (n452,n453,n455);
and (n453,n119,n454);
nand (n454,n115,n54);
and (n455,n114,n397);
nand (n456,n457,n462);
or (n457,n458,n176);
not (n458,n459);
nor (n459,n460,n461);
and (n460,n129,n27);
and (n461,n131,n178);
nand (n462,n463,n22);
not (n463,n428);
and (n464,n388,n422);
xor (n465,n466,n471);
xor (n466,n467,n468);
xor (n467,n356,n368);
or (n468,n469,n470);
and (n469,n436,n450);
and (n470,n437,n444);
xor (n471,n472,n479);
xor (n472,n473,n476);
nand (n473,n474,n475);
or (n474,n162,n447);
or (n475,n156,n331);
nand (n476,n477,n478);
or (n477,n193,n441);
or (n478,n310,n199);
or (n479,n480,n481);
and (n480,n423,n432);
and (n481,n424,n426);
not (n482,n483);
nand (n483,n484,n485);
xor (n484,n387,n435);
or (n485,n486,n509);
and (n486,n487,n508);
xor (n487,n488,n489);
xor (n488,n451,n456);
or (n489,n490,n507);
and (n490,n491,n500);
xor (n491,n492,n493);
and (n492,n239,n54);
nand (n493,n494,n495);
or (n494,n190,n458);
nand (n495,n496,n177);
not (n496,n497);
nor (n497,n498,n499);
and (n498,n21,n178);
and (n499,n147,n27);
nand (n500,n501,n506);
or (n501,n502,n193);
not (n502,n503);
nor (n503,n504,n505);
and (n504,n34,n75);
and (n505,n205,n282);
nand (n506,n200,n405);
and (n507,n492,n493);
xor (n508,n390,n412);
and (n509,n488,n489);
and (n510,n385,n465);
nor (n511,n512,n519);
xor (n512,n513,n516);
xor (n513,n514,n515);
xor (n514,n316,n329);
xor (n515,n353,n354);
or (n516,n517,n518);
and (n517,n472,n479);
and (n518,n473,n476);
or (n519,n520,n521);
and (n520,n466,n471);
and (n521,n467,n468);
nand (n522,n512,n519);
nand (n523,n524,n526);
not (n524,n525);
xor (n525,n349,n352);
not (n526,n527);
or (n527,n528,n529);
and (n528,n513,n516);
and (n529,n514,n515);
nand (n530,n523,n531,n668);
nor (n531,n532,n665);
nor (n532,n533,n663);
and (n533,n534,n658);
or (n534,n535,n657);
and (n535,n536,n576);
xor (n536,n537,n569);
or (n537,n538,n568);
and (n538,n539,n557);
xor (n539,n540,n546);
nand (n540,n541,n545);
or (n541,n542,n193);
not (n542,n543);
nor (n543,n544,n74);
and (n544,n327,n205);
nand (n545,n200,n503);
nand (n546,n547,n552);
or (n547,n548,n156);
not (n548,n549);
nor (n549,n550,n551);
and (n550,n48,n95);
and (n551,n366,n119);
nand (n552,n553,n554);
not (n553,n162);
nand (n554,n555,n556);
or (n555,n119,n54);
or (n556,n95,n397);
xor (n557,n558,n562);
and (n558,n559,n95);
nand (n559,n560,n561);
or (n560,n75,n93);
or (n561,n88,n54);
nand (n562,n563,n567);
or (n563,n176,n564);
nor (n564,n565,n566);
and (n565,n178,n26);
and (n566,n27,n243);
or (n567,n497,n190);
and (n568,n540,n546);
xor (n569,n570,n575);
xor (n570,n571,n574);
nand (n571,n572,n573);
or (n572,n548,n162);
or (n573,n156,n414);
and (n574,n558,n562);
xor (n575,n491,n500);
or (n576,n577,n656);
and (n577,n578,n597);
xor (n578,n579,n596);
or (n579,n580,n595);
and (n580,n581,n589);
xor (n581,n582,n583);
and (n582,n157,n54);
nand (n583,n584,n588);
or (n584,n585,n193);
not (n585,n586);
nor (n586,n81,n587);
and (n587,n366,n205);
nand (n588,n543,n200);
nand (n589,n590,n594);
or (n590,n176,n591);
not (n591,n592);
nor (n592,n593,n33);
and (n593,n282,n178);
or (n594,n564,n190);
and (n595,n582,n583);
xor (n596,n539,n557);
or (n597,n598,n655);
and (n598,n599,n654);
xor (n599,n600,n613);
nor (n600,n601,n609);
not (n601,n602);
nand (n602,n603,n608);
or (n603,n604,n176);
not (n604,n605);
nand (n605,n606,n607);
or (n606,n327,n27);
nand (n607,n27,n327);
nand (n608,n592,n22);
nand (n609,n610,n75);
nand (n610,n611,n612);
or (n611,n27,n73);
or (n612,n56,n54);
nand (n613,n614,n652);
or (n614,n615,n638);
not (n615,n616);
nand (n616,n617,n637);
or (n617,n618,n627);
nor (n618,n619,n626);
nand (n619,n620,n625);
or (n620,n621,n176);
not (n621,n622);
nand (n622,n623,n624);
or (n623,n366,n27);
nand (n624,n27,n366);
nand (n625,n605,n22);
nor (n626,n199,n397);
nand (n627,n628,n635);
nand (n628,n629,n634);
or (n629,n630,n176);
not (n630,n631);
nand (n631,n632,n633);
or (n632,n178,n54);
or (n633,n27,n397);
nand (n634,n622,n22);
nor (n635,n636,n178);
and (n636,n54,n22);
nand (n637,n619,n626);
not (n638,n639);
nand (n639,n640,n648);
not (n640,n641);
nand (n641,n642,n647);
or (n642,n643,n193);
not (n643,n644);
nand (n644,n645,n646);
or (n645,n205,n54);
or (n646,n75,n397);
nand (n647,n200,n586);
nor (n648,n649,n651);
and (n649,n601,n650);
not (n650,n609);
and (n651,n602,n609);
nand (n652,n653,n641);
not (n653,n648);
xor (n654,n581,n589);
and (n655,n600,n613);
and (n656,n579,n596);
and (n657,n537,n569);
or (n658,n659,n660);
xor (n659,n487,n508);
or (n660,n661,n662);
and (n661,n570,n575);
and (n662,n571,n574);
not (n663,n664);
nand (n664,n659,n660);
nand (n665,n666,n383);
not (n666,n667);
nor (n667,n484,n485);
not (n668,n511);
nand (n669,n525,n527);
nand (n670,n345,n347);
or (n671,n340,n102);
nand (n673,n6,n672);
not (n674,n675);
nand (n675,n676,n800,n811);
or (n676,n677,n789);
nand (n677,n678,n738,n763);
not (n678,n679);
not (n679,n680);
or (n680,n681,n691,n737);
not (n681,n682);
nand (n682,n683,n690);
and (n683,n684,n8);
nand (n684,n685,n689);
or (n685,n686,n687);
not (n686,n534);
not (n687,n688);
nand (n688,n658,n664);
or (n689,n688,n534);
and (n691,n683,n692);
or (n692,n693,n698,n736);
not (n693,n694);
nand (n694,n695,n697);
and (n695,n696,n8);
xor (n696,n536,n576);
and (n698,n695,n699);
or (n699,n700,n703,n735);
and (n700,n701,n702);
wire s0n702,s1n702,notn702;
or (n702,s0n702,s1n702);
not(notn702,n9);
and (s0n702,notn702,n11);
and (s1n702,n9,1'b0);
and (n703,n702,n704);
or (n704,n705,n709,n734);
and (n705,n706,n707);
wire s0n707,s1n707,notn707;
or (n707,s0n707,s1n707);
not(notn707,n9);
and (s0n707,notn707,n708);
and (s1n707,n9,1'b0);
xor (n708,n92,n93);
and (n709,n707,n710);
or (n710,n711,n715,n733);
and (n711,n712,n713);
wire s0n713,s1n713,notn713;
or (n713,s0n713,s1n713);
not(notn713,n9);
and (s0n713,notn713,n714);
and (s1n713,n9,1'b0);
xor (n714,n85,n86);
and (n715,n713,n716);
or (n716,n717,n721,n732);
and (n717,n718,n719);
wire s0n719,s1n719,notn719;
or (n719,s0n719,s1n719);
not(notn719,n9);
and (s0n719,notn719,n720);
and (s1n719,n9,1'b0);
xor (n720,n72,n73);
and (n721,n719,n722);
or (n722,n723,n727,n731);
and (n723,n724,n725);
wire s0n725,s1n725,notn725;
or (n725,s0n725,s1n725);
not(notn725,n9);
and (s0n725,notn725,n726);
and (s1n725,n9,1'b0);
xor (n726,n52,n53);
and (n727,n725,n728);
and (n728,n729,n730);
wire s0n730,s1n730,notn730;
or (n730,s0n730,s1n730);
not(notn730,n9);
and (s0n730,notn730,n636);
and (s1n730,n9,1'b0);
and (n731,n724,n728);
and (n732,n718,n722);
and (n733,n712,n716);
and (n734,n706,n710);
and (n735,n701,n704);
and (n736,n697,n699);
and (n737,n690,n692);
nor (n738,n739,n752);
nor (n739,n740,n751);
nand (n740,n741,n743);
or (n741,n8,n742);
not (n742,n714);
nand (n743,n744,n8);
xnor (n744,n745,n746);
nand (n745,n523,n669);
nand (n746,n747,n522);
or (n747,n511,n748);
not (n748,n749);
nand (n749,n750,n381);
not (n750,n531);
nor (n752,n753,n762);
nand (n753,n754,n756);
or (n754,n8,n755);
not (n755,n720);
nand (n756,n757,n8);
nand (n757,n758,n761);
or (n758,n759,n748);
not (n759,n760);
nand (n760,n668,n522);
or (n761,n749,n760);
nor (n763,n764,n778);
nor (n764,n765,n777);
nand (n765,n766,n768);
or (n766,n8,n767);
not (n767,n726);
nand (n768,n769,n8);
nand (n769,n770,n776);
or (n770,n771,n773);
not (n771,n772);
or (n772,n510,n384);
not (n773,n774);
nand (n774,n775,n483);
or (n775,n532,n667);
or (n776,n774,n772);
nor (n778,n779,n788);
or (n779,n780,n781);
and (n780,n9,n636);
and (n781,n8,n782);
nand (n782,n783,n787);
or (n783,n784,n785);
not (n784,n532);
not (n785,n786);
nor (n786,n482,n667);
or (n787,n786,n532);
nor (n789,n790,n799);
nand (n790,n791,n793);
or (n791,n8,n792);
not (n792,n708);
nand (n793,n794,n8);
nand (n794,n795,n798);
or (n795,n796,n376);
not (n796,n797);
nand (n797,n343,n670);
or (n798,n377,n797);
or (n800,n789,n801);
nor (n801,n802,n807);
and (n802,n738,n803);
nand (n803,n804,n806);
or (n804,n764,n805);
nand (n805,n779,n788);
nand (n806,n765,n777);
nand (n807,n808,n810);
or (n808,n739,n809);
nand (n809,n753,n762);
nand (n810,n740,n751);
nand (n811,n790,n799);
or (n812,n675,n3);
xor (n813,n814,n1203);
xor (n814,n672,n815);
wire s0n815,s1n815,notn815;
or (n815,s0n815,s1n815);
not(notn815,n9);
and (s0n815,notn815,n816);
and (s1n815,n9,n11);
xor (n816,n817,n1164);
xor (n817,n818,n1201);
xor (n818,n819,n1159);
xor (n819,n820,n1194);
xor (n820,n821,n1153);
xor (n821,n822,n1182);
xor (n822,n823,n1147);
xor (n823,n824,n1165);
xor (n824,n825,n1141);
xor (n825,n826,n1138);
xor (n826,n827,n1137);
xor (n827,n828,n1107);
xor (n828,n829,n1106);
xor (n829,n830,n1067);
xor (n830,n831,n1066);
xor (n831,n832,n1024);
xor (n832,n833,n1023);
xor (n833,n834,n978);
xor (n834,n835,n977);
xor (n835,n836,n934);
xor (n836,n837,n933);
xor (n837,n838,n888);
xor (n838,n839,n887);
xor (n839,n840,n843);
xor (n840,n841,n842);
and (n841,n187,n22);
and (n842,n181,n27);
or (n843,n844,n847);
and (n844,n845,n846);
and (n845,n181,n22);
and (n846,n212,n27);
and (n847,n848,n849);
xor (n848,n845,n846);
or (n849,n850,n853);
and (n850,n851,n852);
and (n851,n212,n22);
and (n852,n206,n27);
and (n853,n854,n855);
xor (n854,n851,n852);
or (n855,n856,n859);
and (n856,n857,n858);
and (n857,n206,n22);
and (n858,n153,n27);
and (n859,n860,n861);
xor (n860,n857,n858);
or (n861,n862,n865);
and (n862,n863,n864);
and (n863,n153,n22);
and (n864,n168,n27);
and (n865,n866,n867);
xor (n866,n863,n864);
or (n867,n868,n871);
and (n868,n869,n870);
and (n869,n168,n22);
and (n870,n135,n27);
and (n871,n872,n873);
xor (n872,n869,n870);
or (n873,n874,n876);
and (n874,n875,n460);
and (n875,n135,n22);
and (n876,n877,n878);
xor (n877,n875,n460);
or (n878,n879,n882);
and (n879,n880,n881);
and (n880,n129,n22);
and (n881,n21,n27);
and (n882,n883,n884);
xor (n883,n880,n881);
or (n884,n885,n886);
and (n885,n20,n25);
and (n886,n19,n30);
and (n887,n212,n56);
or (n888,n889,n892);
and (n889,n890,n891);
xor (n890,n848,n849);
and (n891,n206,n56);
and (n892,n893,n894);
xor (n893,n890,n891);
or (n894,n895,n898);
and (n895,n896,n897);
xor (n896,n854,n855);
and (n897,n153,n56);
and (n898,n899,n900);
xor (n899,n896,n897);
or (n900,n901,n904);
and (n901,n902,n903);
xor (n902,n860,n861);
and (n903,n168,n56);
and (n904,n905,n906);
xor (n905,n902,n903);
or (n906,n907,n910);
and (n907,n908,n909);
xor (n908,n866,n867);
and (n909,n135,n56);
and (n910,n911,n912);
xor (n911,n908,n909);
or (n912,n913,n916);
and (n913,n914,n915);
xor (n914,n872,n873);
and (n915,n129,n56);
and (n916,n917,n918);
xor (n917,n914,n915);
or (n918,n919,n922);
and (n919,n920,n921);
xor (n920,n877,n878);
and (n921,n21,n56);
and (n922,n923,n924);
xor (n923,n920,n921);
or (n924,n925,n928);
and (n925,n926,n927);
xor (n926,n883,n884);
and (n927,n26,n56);
and (n928,n929,n930);
xor (n929,n926,n927);
or (n930,n931,n932);
and (n931,n18,n55);
and (n932,n17,n59);
and (n933,n206,n75);
or (n934,n935,n938);
and (n935,n936,n937);
xor (n936,n893,n894);
and (n937,n153,n75);
and (n938,n939,n940);
xor (n939,n936,n937);
or (n940,n941,n944);
and (n941,n942,n943);
xor (n942,n899,n900);
and (n943,n168,n75);
and (n944,n945,n946);
xor (n945,n942,n943);
or (n946,n947,n950);
and (n947,n948,n949);
xor (n948,n905,n906);
and (n949,n135,n75);
and (n950,n951,n952);
xor (n951,n948,n949);
or (n952,n953,n956);
and (n953,n954,n955);
xor (n954,n911,n912);
and (n955,n129,n75);
and (n956,n957,n958);
xor (n957,n954,n955);
or (n958,n959,n961);
and (n959,n960,n410);
xor (n960,n917,n918);
and (n961,n962,n963);
xor (n962,n960,n410);
or (n963,n964,n967);
and (n964,n965,n966);
xor (n965,n923,n924);
and (n966,n26,n75);
and (n967,n968,n969);
xor (n968,n965,n966);
or (n969,n970,n972);
and (n970,n971,n504);
xor (n971,n929,n930);
and (n972,n973,n974);
xor (n973,n971,n504);
or (n974,n975,n976);
and (n975,n16,n74);
and (n976,n15,n78);
and (n977,n153,n88);
or (n978,n979,n982);
and (n979,n980,n981);
xor (n980,n939,n940);
and (n981,n168,n88);
and (n982,n983,n984);
xor (n983,n980,n981);
or (n984,n985,n988);
and (n985,n986,n987);
xor (n986,n945,n946);
and (n987,n135,n88);
and (n988,n989,n990);
xor (n989,n986,n987);
or (n990,n991,n994);
and (n991,n992,n993);
xor (n992,n951,n952);
and (n993,n129,n88);
and (n994,n995,n996);
xor (n995,n992,n993);
or (n996,n997,n1000);
and (n997,n998,n999);
xor (n998,n957,n958);
and (n999,n21,n88);
and (n1000,n1001,n1002);
xor (n1001,n998,n999);
or (n1002,n1003,n1006);
and (n1003,n1004,n1005);
xor (n1004,n962,n963);
and (n1005,n26,n88);
and (n1006,n1007,n1008);
xor (n1007,n1004,n1005);
or (n1008,n1009,n1012);
and (n1009,n1010,n1011);
xor (n1010,n968,n969);
and (n1011,n34,n88);
and (n1012,n1013,n1014);
xor (n1013,n1010,n1011);
or (n1014,n1015,n1018);
and (n1015,n1016,n1017);
xor (n1016,n973,n974);
and (n1017,n41,n88);
and (n1018,n1019,n1020);
xor (n1019,n1016,n1017);
or (n1020,n1021,n1022);
and (n1021,n14,n87);
and (n1022,n13,n91);
and (n1023,n168,n95);
or (n1024,n1025,n1028);
and (n1025,n1026,n1027);
xor (n1026,n983,n984);
and (n1027,n135,n95);
and (n1028,n1029,n1030);
xor (n1029,n1026,n1027);
or (n1030,n1031,n1034);
and (n1031,n1032,n1033);
xor (n1032,n989,n990);
and (n1033,n129,n95);
and (n1034,n1035,n1036);
xor (n1035,n1032,n1033);
or (n1036,n1037,n1040);
and (n1037,n1038,n1039);
xor (n1038,n995,n996);
and (n1039,n21,n95);
and (n1040,n1041,n1042);
xor (n1041,n1038,n1039);
or (n1042,n1043,n1046);
and (n1043,n1044,n1045);
xor (n1044,n1001,n1002);
and (n1045,n26,n95);
and (n1046,n1047,n1048);
xor (n1047,n1044,n1045);
or (n1048,n1049,n1052);
and (n1049,n1050,n1051);
xor (n1050,n1007,n1008);
and (n1051,n34,n95);
and (n1052,n1053,n1054);
xor (n1053,n1050,n1051);
or (n1054,n1055,n1058);
and (n1055,n1056,n1057);
xor (n1056,n1013,n1014);
and (n1057,n41,n95);
and (n1058,n1059,n1060);
xor (n1059,n1056,n1057);
or (n1060,n1061,n1063);
and (n1061,n1062,n550);
xor (n1062,n1019,n1020);
and (n1063,n1064,n1065);
xor (n1064,n1062,n550);
and (n1065,n12,n94);
and (n1066,n135,n115);
or (n1067,n1068,n1071);
and (n1068,n1069,n1070);
xor (n1069,n1029,n1030);
and (n1070,n129,n115);
and (n1071,n1072,n1073);
xor (n1072,n1069,n1070);
or (n1073,n1074,n1077);
and (n1074,n1075,n1076);
xor (n1075,n1035,n1036);
and (n1076,n21,n115);
and (n1077,n1078,n1079);
xor (n1078,n1075,n1076);
or (n1079,n1080,n1083);
and (n1080,n1081,n1082);
xor (n1081,n1041,n1042);
and (n1082,n26,n115);
and (n1083,n1084,n1085);
xor (n1084,n1081,n1082);
or (n1085,n1086,n1089);
and (n1086,n1087,n1088);
xor (n1087,n1047,n1048);
and (n1088,n34,n115);
and (n1089,n1090,n1091);
xor (n1090,n1087,n1088);
or (n1091,n1092,n1095);
and (n1092,n1093,n1094);
xor (n1093,n1053,n1054);
and (n1094,n41,n115);
and (n1095,n1096,n1097);
xor (n1096,n1093,n1094);
or (n1097,n1098,n1101);
and (n1098,n1099,n1100);
xor (n1099,n1059,n1060);
and (n1100,n48,n115);
and (n1101,n1102,n1103);
xor (n1102,n1099,n1100);
and (n1103,n1104,n1105);
xor (n1104,n1064,n1065);
not (n1105,n454);
and (n1106,n129,n122);
or (n1107,n1108,n1110);
and (n1108,n1109,n235);
xor (n1109,n1072,n1073);
and (n1110,n1111,n1112);
xor (n1111,n1109,n235);
or (n1112,n1113,n1115);
and (n1113,n1114,n276);
xor (n1114,n1078,n1079);
and (n1115,n1116,n1117);
xor (n1116,n1114,n276);
or (n1117,n1118,n1120);
and (n1118,n1119,n321);
xor (n1119,n1084,n1085);
and (n1120,n1121,n1122);
xor (n1121,n1119,n321);
or (n1122,n1123,n1126);
and (n1123,n1124,n1125);
xor (n1124,n1090,n1091);
and (n1125,n41,n122);
and (n1126,n1127,n1128);
xor (n1127,n1124,n1125);
or (n1128,n1129,n1132);
and (n1129,n1130,n1131);
xor (n1130,n1096,n1097);
and (n1131,n48,n122);
and (n1132,n1133,n1134);
xor (n1133,n1130,n1131);
and (n1134,n1135,n1136);
xor (n1135,n1102,n1103);
and (n1136,n54,n122);
and (n1137,n21,n141);
or (n1138,n1139,n1142);
and (n1139,n1140,n1141);
xor (n1140,n1111,n1112);
and (n1141,n26,n141);
and (n1142,n1143,n1144);
xor (n1143,n1140,n1141);
or (n1144,n1145,n1148);
and (n1145,n1146,n1147);
xor (n1146,n1116,n1117);
and (n1147,n34,n141);
and (n1148,n1149,n1150);
xor (n1149,n1146,n1147);
or (n1150,n1151,n1154);
and (n1151,n1152,n1153);
xor (n1152,n1121,n1122);
and (n1153,n41,n141);
and (n1154,n1155,n1156);
xor (n1155,n1152,n1153);
or (n1156,n1157,n1160);
and (n1157,n1158,n1159);
xor (n1158,n1127,n1128);
and (n1159,n48,n141);
and (n1160,n1161,n1162);
xor (n1161,n1158,n1159);
and (n1162,n1163,n1164);
xor (n1163,n1133,n1134);
and (n1164,n54,n141);
or (n1165,n1166,n1168);
and (n1166,n1167,n1147);
xor (n1167,n1143,n1144);
and (n1168,n1169,n1170);
xor (n1169,n1167,n1147);
or (n1170,n1171,n1173);
and (n1171,n1172,n1153);
xor (n1172,n1149,n1150);
and (n1173,n1174,n1175);
xor (n1174,n1172,n1153);
or (n1175,n1176,n1178);
and (n1176,n1177,n1159);
xor (n1177,n1155,n1156);
and (n1178,n1179,n1180);
xor (n1179,n1177,n1159);
and (n1180,n1181,n1164);
xor (n1181,n1161,n1162);
or (n1182,n1183,n1185);
and (n1183,n1184,n1153);
xor (n1184,n1169,n1170);
and (n1185,n1186,n1187);
xor (n1186,n1184,n1153);
or (n1187,n1188,n1190);
and (n1188,n1189,n1159);
xor (n1189,n1174,n1175);
and (n1190,n1191,n1192);
xor (n1191,n1189,n1159);
and (n1192,n1193,n1164);
xor (n1193,n1179,n1180);
or (n1194,n1195,n1197);
and (n1195,n1196,n1159);
xor (n1196,n1186,n1187);
and (n1197,n1198,n1199);
xor (n1198,n1196,n1159);
and (n1199,n1200,n1164);
xor (n1200,n1191,n1192);
and (n1201,n1202,n1164);
xor (n1202,n1198,n1199);
or (n1203,n1204,n1207,n1232);
and (n1204,n799,n1205);
wire s0n1205,s1n1205,notn1205;
or (n1205,s0n1205,s1n1205);
not(notn1205,n9);
and (s0n1205,notn1205,n1206);
and (s1n1205,n9,n708);
xor (n1206,n1202,n1164);
and (n1207,n1205,n1208);
or (n1208,n1209,n1212,n1231);
and (n1209,n751,n1210);
wire s0n1210,s1n1210,notn1210;
or (n1210,s0n1210,s1n1210);
not(notn1210,n9);
and (s0n1210,notn1210,n1211);
and (s1n1210,n9,n714);
xor (n1211,n1200,n1164);
and (n1212,n1210,n1213);
or (n1213,n1214,n1217,n1230);
and (n1214,n762,n1215);
wire s0n1215,s1n1215,notn1215;
or (n1215,s0n1215,s1n1215);
not(notn1215,n9);
and (s0n1215,notn1215,n1216);
and (s1n1215,n9,n720);
xor (n1216,n1193,n1164);
and (n1217,n1215,n1218);
or (n1218,n1219,n1222,n1229);
and (n1219,n777,n1220);
wire s0n1220,s1n1220,notn1220;
or (n1220,s0n1220,s1n1220);
not(notn1220,n9);
and (s0n1220,notn1220,n1221);
and (s1n1220,n9,n726);
xor (n1221,n1181,n1164);
and (n1222,n1220,n1223);
or (n1223,n1224,n1227,n1228);
and (n1224,n788,n1225);
wire s0n1225,s1n1225,notn1225;
or (n1225,s0n1225,s1n1225);
not(notn1225,n9);
and (s0n1225,notn1225,n1226);
and (s1n1225,n9,n636);
xor (n1226,n1163,n1164);
and (n1227,n1225,n680);
and (n1228,n788,n680);
and (n1229,n777,n1223);
and (n1230,n762,n1218);
and (n1231,n751,n1213);
and (n1232,n799,n1208);
endmodule
