module top (out,n12,n15,n17,n18,n20,n32,n35,n37,n38
        ,n40,n44,n52,n54,n55,n57,n61,n64,n70,n88
        ,n102,n103,n104,n105,n106,n107,n108,n109,n113,n114
        ,n115,n119,n121,n123,n160,n162,n163,n164,n175,n176
        ,n177,n178,n190,n191,n192,n193,n206,n207,n208,n209
        ,n215,n217,n218,n221,n223,n226,n228,n229,n230,n310
        ,n416,n419,n421,n575,n577,n578,n581,n585,n586,n598
        ,n601,n603,n605,n609,n612,n614,n616,n620,n623,n625
        ,n627,n629,n678,n681,n683,n685,n689,n692,n694,n696
        ,n700,n703,n705,n707,n711,n714,n716,n718,n751,n754
        ,n756,n758,n762,n765,n767,n769,n773,n776,n778,n780
        ,n784,n787,n789,n791,n825,n828,n830,n832,n836,n839
        ,n841,n843,n847,n850,n852,n854,n858,n861,n863,n865
        ,n895,n925,n926,n953,n954,n963,n964,n973,n974,n988
        ,n989,n992,n993,n996,n997,n1000,n1001,n1008,n1009,n1012
        ,n1013,n1016,n1017,n1020,n1021,n1028,n1029,n1032,n1033,n1036
        ,n1037,n1040,n1041,n1050,n1051,n1065,n1066,n1084,n1085,n1088
        ,n1089,n1092,n1093,n1096,n1097,n1102,n1103,n1106,n1107,n1110
        ,n1111,n1114,n1115,n1120,n1121,n1124,n1125,n1128,n1129,n1132
        ,n1133,n1138,n1139,n1142,n1143,n1146,n1147,n1150,n1151,n1157
        ,n1158,n1172,n1173,n1191,n1192,n1195,n1196,n1199,n1200,n1203
        ,n1204,n1209,n1210,n1213,n1214,n1217,n1218,n1221,n1222,n1227
        ,n1228,n1231,n1232,n1235,n1236,n1239,n1240,n1245,n1246,n1249
        ,n1250,n1253,n1254,n1257,n1258,n1264,n1265,n1279,n1280,n1298
        ,n1299,n1302,n1303,n1306,n1307,n1310,n1311,n1316,n1317,n1320
        ,n1321,n1324,n1325,n1328,n1329,n1334,n1335,n1338,n1339,n1342
        ,n1343,n1346,n1347,n1352,n1353,n1356,n1357,n1360,n1361,n1364
        ,n1365,n1371,n1372,n1386,n1387,n1405,n1406,n1409,n1410,n1413
        ,n1414,n1417,n1418,n1423,n1424,n1427,n1428,n1431,n1432,n1435
        ,n1436,n1441,n1442,n1445,n1446,n1449,n1450,n1453,n1454,n1459
        ,n1460,n1463,n1464,n1467,n1468,n1471,n1472,n1478,n1479,n1493
        ,n1494,n1512,n1513,n1516,n1517,n1520,n1521,n1524,n1525,n1530
        ,n1531,n1534,n1535,n1538,n1539,n1542,n1543,n1548,n1549,n1552
        ,n1553,n1556,n1557,n1560,n1561,n1566,n1567,n1570,n1571,n1574
        ,n1575,n1578,n1579,n1585,n1586,n1600,n1601,n1619,n1620,n1623
        ,n1624,n1627,n1628,n1631,n1632,n1637,n1638,n1641,n1642,n1645
        ,n1646,n1649,n1650,n1655,n1656,n1659,n1660,n1663,n1664,n1667
        ,n1668,n1673,n1674,n1677,n1678,n1681,n1682,n1685,n1686,n1692
        ,n1693,n1707,n1708,n1725,n1726,n1729,n1730,n1733,n1734,n1737
        ,n1738,n1743,n1744,n1747,n1748,n1751,n1752,n1755,n1756,n1761
        ,n1762,n1765,n1766,n1769,n1770,n1773,n1774,n1779,n1780,n1783
        ,n1784,n1787,n1788,n1791,n1792,n1798,n1799,n1813,n1814,n1855
        ,n1856,n1870,n1871,n1877,n1878,n1892,n1893,n1920,n1921,n1935
        ,n1936,n1942,n1943,n1957,n1958,n1985,n1986,n2000,n2001,n2007
        ,n2008,n2022,n2023,n2050,n2051,n2065,n2066,n2072,n2073,n2087
        ,n2088,n2115,n2116,n2130,n2131,n2137,n2138,n2152,n2153,n2180
        ,n2181,n2195,n2196,n2202,n2203,n2217,n2218,n2245,n2246,n2260
        ,n2261,n2267,n2268,n2282,n2283,n2309,n2310,n2324,n2325,n2331
        ,n2332,n2346,n2347,n2464,n2465,n2474,n2475,n2481,n2482,n2491
        ,n2492,n2509,n2510,n2519,n2520,n2526,n2527,n2536,n2537,n2554
        ,n2555,n2564,n2565,n2571,n2572,n2581,n2582,n2599,n2600,n2609
        ,n2610,n2616,n2617,n2626,n2627,n2644,n2645,n2654,n2655,n2661
        ,n2662,n2671,n2672,n2689,n2690,n2699,n2700,n2706,n2707,n2716
        ,n2717,n2734,n2735,n2744,n2745,n2751,n2752,n2761,n2762,n2778
        ,n2779,n2788,n2789,n2795,n2796,n2805,n2806,n3073,n3083,n3087
        ,n3089,n3094,n3096,n3101,n3103,n3108,n3110,n3120,n3121,n3135
        ,n3140,n3145,n3152,n3155,n3158,n3161,n3166,n3167,n3170,n3173
        ,n3176,n3181,n3184,n3187,n3190,n3191,n3198,n3199,n3202,n3205
        ,n3208,n3213,n3216,n3219,n3222,n3227,n3228,n3231,n3234,n3237
        ,n3242,n3245,n3248,n3251,n3252,n3262,n3263,n3266,n3269,n3272
        ,n3277,n3280,n3283,n3286,n3291,n3292,n3295,n3298,n3301,n3306
        ,n3309,n3312,n3315,n3316,n3323,n3324,n3327,n3330,n3333,n3338
        ,n3341,n3344,n3347,n3352,n3353,n3356,n3359,n3362,n3367,n3370
        ,n3373,n3376,n3377,n3387,n3388,n3391,n3394,n3397,n3402,n3405
        ,n3408,n3411,n3416,n3417,n3420,n3423,n3426,n3431,n3434,n3437
        ,n3440,n3441,n3448,n3449,n3452,n3455,n3458,n3463,n3466,n3469
        ,n3472,n3477,n3478,n3481,n3484,n3487,n3492,n3495,n3498,n3501
        ,n3502,n3512,n3513,n3516,n3519,n3522,n3527,n3530,n3533,n3536
        ,n3541,n3542,n3545,n3548,n3551,n3556,n3559,n3562,n3565,n3566
        ,n3573,n3574,n3577,n3580,n3583,n3588,n3591,n3594,n3597,n3602
        ,n3603,n3606,n3609,n3612,n3617,n3620,n3623,n3626,n3627,n3637
        ,n3638,n3641,n3644,n3647,n3652,n3655,n3658,n3661,n3666,n3667
        ,n3670,n3673,n3676,n3681,n3684,n3687,n3690,n3691,n3698,n3699
        ,n3702,n3705,n3708,n3713,n3716,n3719,n3722,n3727,n3728,n3731
        ,n3734,n3737,n3742,n3745,n3748,n3751,n3752,n3762,n3763,n3766
        ,n3769,n3772,n3777,n3780,n3783,n3786,n3791,n3792,n3795,n3798
        ,n3801,n3806,n3809,n3812,n3815,n3816,n3823,n3824,n3827,n3830
        ,n3833,n3838,n3841,n3844,n3847,n3852,n3853,n3856,n3859,n3862
        ,n3867,n3870,n3873,n3876,n3877,n3887,n3888,n3891,n3894,n3897
        ,n3902,n3905,n3908,n3911,n3916,n3917,n3920,n3923,n3926,n3931
        ,n3934,n3937,n3940,n3941,n3948,n3949,n3952,n3955,n3958,n3963
        ,n3966,n3969,n3972,n3977,n3978,n3981,n3984,n3987,n3992,n3995
        ,n3998,n4001,n4002,n4011,n4012,n4015,n4018,n4021,n4026,n4029
        ,n4032,n4035,n4040,n4041,n4044,n4047,n4050,n4055,n4058,n4061
        ,n4064,n4065,n4072,n4073,n4076,n4079,n4082,n4087,n4090,n4093
        ,n4096,n4101,n4102,n4105,n4108,n4111,n4116,n4119,n4122,n4125
        ,n4126,n4144,n4146,n4150,n4152,n4157,n4159,n4205,n4248,n4294
        ,n4337,n4383,n4426,n4472,n4515,n4561,n4604,n4650,n4693,n4739
        ,n4782,n4827,n4870,n4884,n4886,n4890,n4892,n4897,n4899,n4904
        ,n4906,n4911,n4913,n4925,n4926,n4929,n4932,n4935,n4940,n4943
        ,n4946,n4949,n4950,n4957,n4958,n4961,n4964,n4967,n4972,n4975
        ,n4978,n4981,n4984,n4996,n4997,n5000,n5003,n5006,n5011,n5014
        ,n5017,n5020,n5021,n5028,n5029,n5032,n5035,n5038,n5043,n5046
        ,n5049,n5052,n5055,n5067,n5068,n5071,n5074,n5077,n5082,n5085
        ,n5088,n5091,n5092,n5099,n5100,n5103,n5106,n5109,n5114,n5117
        ,n5120,n5123,n5126,n5138,n5139,n5142,n5145,n5148,n5153,n5156
        ,n5159,n5162,n5163,n5170,n5171,n5174,n5177,n5180,n5185,n5188
        ,n5191,n5194,n5197,n5209,n5210,n5213,n5216,n5219,n5224,n5227
        ,n5230,n5233,n5234,n5241,n5242,n5245,n5248,n5251,n5256,n5259
        ,n5262,n5265,n5268,n5280,n5281,n5284,n5287,n5290,n5295,n5298
        ,n5301,n5304,n5305,n5312,n5313,n5316,n5319,n5322,n5327,n5330
        ,n5333,n5336,n5339,n5351,n5352,n5355,n5358,n5361,n5366,n5369
        ,n5372,n5375,n5376,n5383,n5384,n5387,n5390,n5393,n5398,n5401
        ,n5404,n5407,n5410,n5421,n5422,n5425,n5428,n5431,n5436,n5439
        ,n5442,n5445,n5446,n5453,n5454,n5457,n5460,n5463,n5468,n5471
        ,n5474,n5477,n5480,n5784,n5786,n5793,n5795,n5809,n5811,n5818
        ,n5820,n5825,n5827,n5832,n5834,n5848,n5850,n5857,n5859,n6025
        ,n6028,n6137,n6140,n6249,n6252,n6361,n6364,n6469,n6472,n6577
        ,n6580,n6684,n6687,n6837,n6848,n6851,n6853,n6855,n6859,n6862
        ,n6864,n6866,n6870,n6873,n6875,n6877,n6881,n6884,n6886,n6888
        ,n6900,n6903,n6905,n6907,n6911,n6914,n6916,n6918,n6922,n6925
        ,n6927,n6929,n6933,n6936,n6938,n6940,n6979,n7000,n7013,n7026
        ,n7039,n7052,n7064,n7142,n7151,n7166,n7189,n7202,n7220,n7247
        ,n7267,n7326,n7337,n7346,n7362,n7375,n7388,n7400,n7442,n7452
        ,n7464,n7497,n7554,n7582,n7605,n7634,n7655);
output out;
input n12;
input n15;
input n17;
input n18;
input n20;
input n32;
input n35;
input n37;
input n38;
input n40;
input n44;
input n52;
input n54;
input n55;
input n57;
input n61;
input n64;
input n70;
input n88;
input n102;
input n103;
input n104;
input n105;
input n106;
input n107;
input n108;
input n109;
input n113;
input n114;
input n115;
input n119;
input n121;
input n123;
input n160;
input n162;
input n163;
input n164;
input n175;
input n176;
input n177;
input n178;
input n190;
input n191;
input n192;
input n193;
input n206;
input n207;
input n208;
input n209;
input n215;
input n217;
input n218;
input n221;
input n223;
input n226;
input n228;
input n229;
input n230;
input n310;
input n416;
input n419;
input n421;
input n575;
input n577;
input n578;
input n581;
input n585;
input n586;
input n598;
input n601;
input n603;
input n605;
input n609;
input n612;
input n614;
input n616;
input n620;
input n623;
input n625;
input n627;
input n629;
input n678;
input n681;
input n683;
input n685;
input n689;
input n692;
input n694;
input n696;
input n700;
input n703;
input n705;
input n707;
input n711;
input n714;
input n716;
input n718;
input n751;
input n754;
input n756;
input n758;
input n762;
input n765;
input n767;
input n769;
input n773;
input n776;
input n778;
input n780;
input n784;
input n787;
input n789;
input n791;
input n825;
input n828;
input n830;
input n832;
input n836;
input n839;
input n841;
input n843;
input n847;
input n850;
input n852;
input n854;
input n858;
input n861;
input n863;
input n865;
input n895;
input n925;
input n926;
input n953;
input n954;
input n963;
input n964;
input n973;
input n974;
input n988;
input n989;
input n992;
input n993;
input n996;
input n997;
input n1000;
input n1001;
input n1008;
input n1009;
input n1012;
input n1013;
input n1016;
input n1017;
input n1020;
input n1021;
input n1028;
input n1029;
input n1032;
input n1033;
input n1036;
input n1037;
input n1040;
input n1041;
input n1050;
input n1051;
input n1065;
input n1066;
input n1084;
input n1085;
input n1088;
input n1089;
input n1092;
input n1093;
input n1096;
input n1097;
input n1102;
input n1103;
input n1106;
input n1107;
input n1110;
input n1111;
input n1114;
input n1115;
input n1120;
input n1121;
input n1124;
input n1125;
input n1128;
input n1129;
input n1132;
input n1133;
input n1138;
input n1139;
input n1142;
input n1143;
input n1146;
input n1147;
input n1150;
input n1151;
input n1157;
input n1158;
input n1172;
input n1173;
input n1191;
input n1192;
input n1195;
input n1196;
input n1199;
input n1200;
input n1203;
input n1204;
input n1209;
input n1210;
input n1213;
input n1214;
input n1217;
input n1218;
input n1221;
input n1222;
input n1227;
input n1228;
input n1231;
input n1232;
input n1235;
input n1236;
input n1239;
input n1240;
input n1245;
input n1246;
input n1249;
input n1250;
input n1253;
input n1254;
input n1257;
input n1258;
input n1264;
input n1265;
input n1279;
input n1280;
input n1298;
input n1299;
input n1302;
input n1303;
input n1306;
input n1307;
input n1310;
input n1311;
input n1316;
input n1317;
input n1320;
input n1321;
input n1324;
input n1325;
input n1328;
input n1329;
input n1334;
input n1335;
input n1338;
input n1339;
input n1342;
input n1343;
input n1346;
input n1347;
input n1352;
input n1353;
input n1356;
input n1357;
input n1360;
input n1361;
input n1364;
input n1365;
input n1371;
input n1372;
input n1386;
input n1387;
input n1405;
input n1406;
input n1409;
input n1410;
input n1413;
input n1414;
input n1417;
input n1418;
input n1423;
input n1424;
input n1427;
input n1428;
input n1431;
input n1432;
input n1435;
input n1436;
input n1441;
input n1442;
input n1445;
input n1446;
input n1449;
input n1450;
input n1453;
input n1454;
input n1459;
input n1460;
input n1463;
input n1464;
input n1467;
input n1468;
input n1471;
input n1472;
input n1478;
input n1479;
input n1493;
input n1494;
input n1512;
input n1513;
input n1516;
input n1517;
input n1520;
input n1521;
input n1524;
input n1525;
input n1530;
input n1531;
input n1534;
input n1535;
input n1538;
input n1539;
input n1542;
input n1543;
input n1548;
input n1549;
input n1552;
input n1553;
input n1556;
input n1557;
input n1560;
input n1561;
input n1566;
input n1567;
input n1570;
input n1571;
input n1574;
input n1575;
input n1578;
input n1579;
input n1585;
input n1586;
input n1600;
input n1601;
input n1619;
input n1620;
input n1623;
input n1624;
input n1627;
input n1628;
input n1631;
input n1632;
input n1637;
input n1638;
input n1641;
input n1642;
input n1645;
input n1646;
input n1649;
input n1650;
input n1655;
input n1656;
input n1659;
input n1660;
input n1663;
input n1664;
input n1667;
input n1668;
input n1673;
input n1674;
input n1677;
input n1678;
input n1681;
input n1682;
input n1685;
input n1686;
input n1692;
input n1693;
input n1707;
input n1708;
input n1725;
input n1726;
input n1729;
input n1730;
input n1733;
input n1734;
input n1737;
input n1738;
input n1743;
input n1744;
input n1747;
input n1748;
input n1751;
input n1752;
input n1755;
input n1756;
input n1761;
input n1762;
input n1765;
input n1766;
input n1769;
input n1770;
input n1773;
input n1774;
input n1779;
input n1780;
input n1783;
input n1784;
input n1787;
input n1788;
input n1791;
input n1792;
input n1798;
input n1799;
input n1813;
input n1814;
input n1855;
input n1856;
input n1870;
input n1871;
input n1877;
input n1878;
input n1892;
input n1893;
input n1920;
input n1921;
input n1935;
input n1936;
input n1942;
input n1943;
input n1957;
input n1958;
input n1985;
input n1986;
input n2000;
input n2001;
input n2007;
input n2008;
input n2022;
input n2023;
input n2050;
input n2051;
input n2065;
input n2066;
input n2072;
input n2073;
input n2087;
input n2088;
input n2115;
input n2116;
input n2130;
input n2131;
input n2137;
input n2138;
input n2152;
input n2153;
input n2180;
input n2181;
input n2195;
input n2196;
input n2202;
input n2203;
input n2217;
input n2218;
input n2245;
input n2246;
input n2260;
input n2261;
input n2267;
input n2268;
input n2282;
input n2283;
input n2309;
input n2310;
input n2324;
input n2325;
input n2331;
input n2332;
input n2346;
input n2347;
input n2464;
input n2465;
input n2474;
input n2475;
input n2481;
input n2482;
input n2491;
input n2492;
input n2509;
input n2510;
input n2519;
input n2520;
input n2526;
input n2527;
input n2536;
input n2537;
input n2554;
input n2555;
input n2564;
input n2565;
input n2571;
input n2572;
input n2581;
input n2582;
input n2599;
input n2600;
input n2609;
input n2610;
input n2616;
input n2617;
input n2626;
input n2627;
input n2644;
input n2645;
input n2654;
input n2655;
input n2661;
input n2662;
input n2671;
input n2672;
input n2689;
input n2690;
input n2699;
input n2700;
input n2706;
input n2707;
input n2716;
input n2717;
input n2734;
input n2735;
input n2744;
input n2745;
input n2751;
input n2752;
input n2761;
input n2762;
input n2778;
input n2779;
input n2788;
input n2789;
input n2795;
input n2796;
input n2805;
input n2806;
input n3073;
input n3083;
input n3087;
input n3089;
input n3094;
input n3096;
input n3101;
input n3103;
input n3108;
input n3110;
input n3120;
input n3121;
input n3135;
input n3140;
input n3145;
input n3152;
input n3155;
input n3158;
input n3161;
input n3166;
input n3167;
input n3170;
input n3173;
input n3176;
input n3181;
input n3184;
input n3187;
input n3190;
input n3191;
input n3198;
input n3199;
input n3202;
input n3205;
input n3208;
input n3213;
input n3216;
input n3219;
input n3222;
input n3227;
input n3228;
input n3231;
input n3234;
input n3237;
input n3242;
input n3245;
input n3248;
input n3251;
input n3252;
input n3262;
input n3263;
input n3266;
input n3269;
input n3272;
input n3277;
input n3280;
input n3283;
input n3286;
input n3291;
input n3292;
input n3295;
input n3298;
input n3301;
input n3306;
input n3309;
input n3312;
input n3315;
input n3316;
input n3323;
input n3324;
input n3327;
input n3330;
input n3333;
input n3338;
input n3341;
input n3344;
input n3347;
input n3352;
input n3353;
input n3356;
input n3359;
input n3362;
input n3367;
input n3370;
input n3373;
input n3376;
input n3377;
input n3387;
input n3388;
input n3391;
input n3394;
input n3397;
input n3402;
input n3405;
input n3408;
input n3411;
input n3416;
input n3417;
input n3420;
input n3423;
input n3426;
input n3431;
input n3434;
input n3437;
input n3440;
input n3441;
input n3448;
input n3449;
input n3452;
input n3455;
input n3458;
input n3463;
input n3466;
input n3469;
input n3472;
input n3477;
input n3478;
input n3481;
input n3484;
input n3487;
input n3492;
input n3495;
input n3498;
input n3501;
input n3502;
input n3512;
input n3513;
input n3516;
input n3519;
input n3522;
input n3527;
input n3530;
input n3533;
input n3536;
input n3541;
input n3542;
input n3545;
input n3548;
input n3551;
input n3556;
input n3559;
input n3562;
input n3565;
input n3566;
input n3573;
input n3574;
input n3577;
input n3580;
input n3583;
input n3588;
input n3591;
input n3594;
input n3597;
input n3602;
input n3603;
input n3606;
input n3609;
input n3612;
input n3617;
input n3620;
input n3623;
input n3626;
input n3627;
input n3637;
input n3638;
input n3641;
input n3644;
input n3647;
input n3652;
input n3655;
input n3658;
input n3661;
input n3666;
input n3667;
input n3670;
input n3673;
input n3676;
input n3681;
input n3684;
input n3687;
input n3690;
input n3691;
input n3698;
input n3699;
input n3702;
input n3705;
input n3708;
input n3713;
input n3716;
input n3719;
input n3722;
input n3727;
input n3728;
input n3731;
input n3734;
input n3737;
input n3742;
input n3745;
input n3748;
input n3751;
input n3752;
input n3762;
input n3763;
input n3766;
input n3769;
input n3772;
input n3777;
input n3780;
input n3783;
input n3786;
input n3791;
input n3792;
input n3795;
input n3798;
input n3801;
input n3806;
input n3809;
input n3812;
input n3815;
input n3816;
input n3823;
input n3824;
input n3827;
input n3830;
input n3833;
input n3838;
input n3841;
input n3844;
input n3847;
input n3852;
input n3853;
input n3856;
input n3859;
input n3862;
input n3867;
input n3870;
input n3873;
input n3876;
input n3877;
input n3887;
input n3888;
input n3891;
input n3894;
input n3897;
input n3902;
input n3905;
input n3908;
input n3911;
input n3916;
input n3917;
input n3920;
input n3923;
input n3926;
input n3931;
input n3934;
input n3937;
input n3940;
input n3941;
input n3948;
input n3949;
input n3952;
input n3955;
input n3958;
input n3963;
input n3966;
input n3969;
input n3972;
input n3977;
input n3978;
input n3981;
input n3984;
input n3987;
input n3992;
input n3995;
input n3998;
input n4001;
input n4002;
input n4011;
input n4012;
input n4015;
input n4018;
input n4021;
input n4026;
input n4029;
input n4032;
input n4035;
input n4040;
input n4041;
input n4044;
input n4047;
input n4050;
input n4055;
input n4058;
input n4061;
input n4064;
input n4065;
input n4072;
input n4073;
input n4076;
input n4079;
input n4082;
input n4087;
input n4090;
input n4093;
input n4096;
input n4101;
input n4102;
input n4105;
input n4108;
input n4111;
input n4116;
input n4119;
input n4122;
input n4125;
input n4126;
input n4144;
input n4146;
input n4150;
input n4152;
input n4157;
input n4159;
input n4205;
input n4248;
input n4294;
input n4337;
input n4383;
input n4426;
input n4472;
input n4515;
input n4561;
input n4604;
input n4650;
input n4693;
input n4739;
input n4782;
input n4827;
input n4870;
input n4884;
input n4886;
input n4890;
input n4892;
input n4897;
input n4899;
input n4904;
input n4906;
input n4911;
input n4913;
input n4925;
input n4926;
input n4929;
input n4932;
input n4935;
input n4940;
input n4943;
input n4946;
input n4949;
input n4950;
input n4957;
input n4958;
input n4961;
input n4964;
input n4967;
input n4972;
input n4975;
input n4978;
input n4981;
input n4984;
input n4996;
input n4997;
input n5000;
input n5003;
input n5006;
input n5011;
input n5014;
input n5017;
input n5020;
input n5021;
input n5028;
input n5029;
input n5032;
input n5035;
input n5038;
input n5043;
input n5046;
input n5049;
input n5052;
input n5055;
input n5067;
input n5068;
input n5071;
input n5074;
input n5077;
input n5082;
input n5085;
input n5088;
input n5091;
input n5092;
input n5099;
input n5100;
input n5103;
input n5106;
input n5109;
input n5114;
input n5117;
input n5120;
input n5123;
input n5126;
input n5138;
input n5139;
input n5142;
input n5145;
input n5148;
input n5153;
input n5156;
input n5159;
input n5162;
input n5163;
input n5170;
input n5171;
input n5174;
input n5177;
input n5180;
input n5185;
input n5188;
input n5191;
input n5194;
input n5197;
input n5209;
input n5210;
input n5213;
input n5216;
input n5219;
input n5224;
input n5227;
input n5230;
input n5233;
input n5234;
input n5241;
input n5242;
input n5245;
input n5248;
input n5251;
input n5256;
input n5259;
input n5262;
input n5265;
input n5268;
input n5280;
input n5281;
input n5284;
input n5287;
input n5290;
input n5295;
input n5298;
input n5301;
input n5304;
input n5305;
input n5312;
input n5313;
input n5316;
input n5319;
input n5322;
input n5327;
input n5330;
input n5333;
input n5336;
input n5339;
input n5351;
input n5352;
input n5355;
input n5358;
input n5361;
input n5366;
input n5369;
input n5372;
input n5375;
input n5376;
input n5383;
input n5384;
input n5387;
input n5390;
input n5393;
input n5398;
input n5401;
input n5404;
input n5407;
input n5410;
input n5421;
input n5422;
input n5425;
input n5428;
input n5431;
input n5436;
input n5439;
input n5442;
input n5445;
input n5446;
input n5453;
input n5454;
input n5457;
input n5460;
input n5463;
input n5468;
input n5471;
input n5474;
input n5477;
input n5480;
input n5784;
input n5786;
input n5793;
input n5795;
input n5809;
input n5811;
input n5818;
input n5820;
input n5825;
input n5827;
input n5832;
input n5834;
input n5848;
input n5850;
input n5857;
input n5859;
input n6025;
input n6028;
input n6137;
input n6140;
input n6249;
input n6252;
input n6361;
input n6364;
input n6469;
input n6472;
input n6577;
input n6580;
input n6684;
input n6687;
input n6837;
input n6848;
input n6851;
input n6853;
input n6855;
input n6859;
input n6862;
input n6864;
input n6866;
input n6870;
input n6873;
input n6875;
input n6877;
input n6881;
input n6884;
input n6886;
input n6888;
input n6900;
input n6903;
input n6905;
input n6907;
input n6911;
input n6914;
input n6916;
input n6918;
input n6922;
input n6925;
input n6927;
input n6929;
input n6933;
input n6936;
input n6938;
input n6940;
input n6979;
input n7000;
input n7013;
input n7026;
input n7039;
input n7052;
input n7064;
input n7142;
input n7151;
input n7166;
input n7189;
input n7202;
input n7220;
input n7247;
input n7267;
input n7326;
input n7337;
input n7346;
input n7362;
input n7375;
input n7388;
input n7400;
input n7442;
input n7452;
input n7464;
input n7497;
input n7554;
input n7582;
input n7605;
input n7634;
input n7655;
wire n0;
wire n1;
wire n2;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n13;
wire n14;
wire n16;
wire n19;
wire n21;
wire n22;
wire n23;
wire n24;
wire n25;
wire n26;
wire n27;
wire n28;
wire n29;
wire n30;
wire n31;
wire n33;
wire n34;
wire n36;
wire n39;
wire n41;
wire n42;
wire n43;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n53;
wire n56;
wire n58;
wire n59;
wire n60;
wire n62;
wire n63;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n110;
wire n111;
wire n112;
wire n116;
wire n117;
wire n118;
wire n120;
wire n122;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n161;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n216;
wire n219;
wire n220;
wire n222;
wire n224;
wire n225;
wire n227;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n417;
wire n418;
wire n420;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n576;
wire n579;
wire n580;
wire n582;
wire n583;
wire n584;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n599;
wire n600;
wire n602;
wire n604;
wire n606;
wire n607;
wire n608;
wire n610;
wire n611;
wire n613;
wire n615;
wire n617;
wire n618;
wire n619;
wire n621;
wire n622;
wire n624;
wire n626;
wire n628;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n679;
wire n680;
wire n682;
wire n684;
wire n686;
wire n687;
wire n688;
wire n690;
wire n691;
wire n693;
wire n695;
wire n697;
wire n698;
wire n699;
wire n701;
wire n702;
wire n704;
wire n706;
wire n708;
wire n709;
wire n710;
wire n712;
wire n713;
wire n715;
wire n717;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n752;
wire n753;
wire n755;
wire n757;
wire n759;
wire n760;
wire n761;
wire n763;
wire n764;
wire n766;
wire n768;
wire n770;
wire n771;
wire n772;
wire n774;
wire n775;
wire n777;
wire n779;
wire n781;
wire n782;
wire n783;
wire n785;
wire n786;
wire n788;
wire n790;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n826;
wire n827;
wire n829;
wire n831;
wire n833;
wire n834;
wire n835;
wire n837;
wire n838;
wire n840;
wire n842;
wire n844;
wire n845;
wire n846;
wire n848;
wire n849;
wire n851;
wire n853;
wire n855;
wire n856;
wire n857;
wire n859;
wire n860;
wire n862;
wire n864;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n990;
wire n991;
wire n994;
wire n995;
wire n998;
wire n999;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1010;
wire n1011;
wire n1014;
wire n1015;
wire n1018;
wire n1019;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1030;
wire n1031;
wire n1034;
wire n1035;
wire n1038;
wire n1039;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1086;
wire n1087;
wire n1090;
wire n1091;
wire n1094;
wire n1095;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1104;
wire n1105;
wire n1108;
wire n1109;
wire n1112;
wire n1113;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1122;
wire n1123;
wire n1126;
wire n1127;
wire n1130;
wire n1131;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1140;
wire n1141;
wire n1144;
wire n1145;
wire n1148;
wire n1149;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1193;
wire n1194;
wire n1197;
wire n1198;
wire n1201;
wire n1202;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1211;
wire n1212;
wire n1215;
wire n1216;
wire n1219;
wire n1220;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1229;
wire n1230;
wire n1233;
wire n1234;
wire n1237;
wire n1238;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1247;
wire n1248;
wire n1251;
wire n1252;
wire n1255;
wire n1256;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1300;
wire n1301;
wire n1304;
wire n1305;
wire n1308;
wire n1309;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1318;
wire n1319;
wire n1322;
wire n1323;
wire n1326;
wire n1327;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1336;
wire n1337;
wire n1340;
wire n1341;
wire n1344;
wire n1345;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1354;
wire n1355;
wire n1358;
wire n1359;
wire n1362;
wire n1363;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1407;
wire n1408;
wire n1411;
wire n1412;
wire n1415;
wire n1416;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1425;
wire n1426;
wire n1429;
wire n1430;
wire n1433;
wire n1434;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1443;
wire n1444;
wire n1447;
wire n1448;
wire n1451;
wire n1452;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1461;
wire n1462;
wire n1465;
wire n1466;
wire n1469;
wire n1470;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1514;
wire n1515;
wire n1518;
wire n1519;
wire n1522;
wire n1523;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1532;
wire n1533;
wire n1536;
wire n1537;
wire n1540;
wire n1541;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1550;
wire n1551;
wire n1554;
wire n1555;
wire n1558;
wire n1559;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1568;
wire n1569;
wire n1572;
wire n1573;
wire n1576;
wire n1577;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1621;
wire n1622;
wire n1625;
wire n1626;
wire n1629;
wire n1630;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1639;
wire n1640;
wire n1643;
wire n1644;
wire n1647;
wire n1648;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1657;
wire n1658;
wire n1661;
wire n1662;
wire n1665;
wire n1666;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1675;
wire n1676;
wire n1679;
wire n1680;
wire n1683;
wire n1684;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1727;
wire n1728;
wire n1731;
wire n1732;
wire n1735;
wire n1736;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1745;
wire n1746;
wire n1749;
wire n1750;
wire n1753;
wire n1754;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1763;
wire n1764;
wire n1767;
wire n1768;
wire n1771;
wire n1772;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1781;
wire n1782;
wire n1785;
wire n1786;
wire n1789;
wire n1790;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2988;
wire n2989;
wire n2990;
wire n2991;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2996;
wire n2997;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3003;
wire n3004;
wire n3005;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3010;
wire n3011;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3038;
wire n3039;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
wire n3056;
wire n3057;
wire n3058;
wire n3059;
wire n3060;
wire n3061;
wire n3062;
wire n3063;
wire n3064;
wire n3065;
wire n3066;
wire n3067;
wire n3068;
wire n3069;
wire n3070;
wire n3071;
wire n3072;
wire n3074;
wire n3075;
wire n3076;
wire n3077;
wire n3078;
wire n3079;
wire n3080;
wire n3081;
wire n3082;
wire n3084;
wire n3085;
wire n3086;
wire n3088;
wire n3090;
wire n3091;
wire n3092;
wire n3093;
wire n3095;
wire n3097;
wire n3098;
wire n3099;
wire n3100;
wire n3102;
wire n3104;
wire n3105;
wire n3106;
wire n3107;
wire n3109;
wire n3111;
wire n3112;
wire n3113;
wire n3114;
wire n3115;
wire n3116;
wire n3117;
wire n3118;
wire n3119;
wire n3122;
wire n3123;
wire n3124;
wire n3125;
wire n3126;
wire n3127;
wire n3128;
wire n3129;
wire n3130;
wire n3131;
wire n3132;
wire n3133;
wire n3134;
wire n3136;
wire n3137;
wire n3138;
wire n3139;
wire n3141;
wire n3142;
wire n3143;
wire n3144;
wire n3146;
wire n3147;
wire n3148;
wire n3149;
wire n3150;
wire n3151;
wire n3153;
wire n3154;
wire n3156;
wire n3157;
wire n3159;
wire n3160;
wire n3162;
wire n3163;
wire n3164;
wire n3165;
wire n3168;
wire n3169;
wire n3171;
wire n3172;
wire n3174;
wire n3175;
wire n3177;
wire n3178;
wire n3179;
wire n3180;
wire n3182;
wire n3183;
wire n3185;
wire n3186;
wire n3188;
wire n3189;
wire n3192;
wire n3193;
wire n3194;
wire n3195;
wire n3196;
wire n3197;
wire n3200;
wire n3201;
wire n3203;
wire n3204;
wire n3206;
wire n3207;
wire n3209;
wire n3210;
wire n3211;
wire n3212;
wire n3214;
wire n3215;
wire n3217;
wire n3218;
wire n3220;
wire n3221;
wire n3223;
wire n3224;
wire n3225;
wire n3226;
wire n3229;
wire n3230;
wire n3232;
wire n3233;
wire n3235;
wire n3236;
wire n3238;
wire n3239;
wire n3240;
wire n3241;
wire n3243;
wire n3244;
wire n3246;
wire n3247;
wire n3249;
wire n3250;
wire n3253;
wire n3254;
wire n3255;
wire n3256;
wire n3257;
wire n3258;
wire n3259;
wire n3260;
wire n3261;
wire n3264;
wire n3265;
wire n3267;
wire n3268;
wire n3270;
wire n3271;
wire n3273;
wire n3274;
wire n3275;
wire n3276;
wire n3278;
wire n3279;
wire n3281;
wire n3282;
wire n3284;
wire n3285;
wire n3287;
wire n3288;
wire n3289;
wire n3290;
wire n3293;
wire n3294;
wire n3296;
wire n3297;
wire n3299;
wire n3300;
wire n3302;
wire n3303;
wire n3304;
wire n3305;
wire n3307;
wire n3308;
wire n3310;
wire n3311;
wire n3313;
wire n3314;
wire n3317;
wire n3318;
wire n3319;
wire n3320;
wire n3321;
wire n3322;
wire n3325;
wire n3326;
wire n3328;
wire n3329;
wire n3331;
wire n3332;
wire n3334;
wire n3335;
wire n3336;
wire n3337;
wire n3339;
wire n3340;
wire n3342;
wire n3343;
wire n3345;
wire n3346;
wire n3348;
wire n3349;
wire n3350;
wire n3351;
wire n3354;
wire n3355;
wire n3357;
wire n3358;
wire n3360;
wire n3361;
wire n3363;
wire n3364;
wire n3365;
wire n3366;
wire n3368;
wire n3369;
wire n3371;
wire n3372;
wire n3374;
wire n3375;
wire n3378;
wire n3379;
wire n3380;
wire n3381;
wire n3382;
wire n3383;
wire n3384;
wire n3385;
wire n3386;
wire n3389;
wire n3390;
wire n3392;
wire n3393;
wire n3395;
wire n3396;
wire n3398;
wire n3399;
wire n3400;
wire n3401;
wire n3403;
wire n3404;
wire n3406;
wire n3407;
wire n3409;
wire n3410;
wire n3412;
wire n3413;
wire n3414;
wire n3415;
wire n3418;
wire n3419;
wire n3421;
wire n3422;
wire n3424;
wire n3425;
wire n3427;
wire n3428;
wire n3429;
wire n3430;
wire n3432;
wire n3433;
wire n3435;
wire n3436;
wire n3438;
wire n3439;
wire n3442;
wire n3443;
wire n3444;
wire n3445;
wire n3446;
wire n3447;
wire n3450;
wire n3451;
wire n3453;
wire n3454;
wire n3456;
wire n3457;
wire n3459;
wire n3460;
wire n3461;
wire n3462;
wire n3464;
wire n3465;
wire n3467;
wire n3468;
wire n3470;
wire n3471;
wire n3473;
wire n3474;
wire n3475;
wire n3476;
wire n3479;
wire n3480;
wire n3482;
wire n3483;
wire n3485;
wire n3486;
wire n3488;
wire n3489;
wire n3490;
wire n3491;
wire n3493;
wire n3494;
wire n3496;
wire n3497;
wire n3499;
wire n3500;
wire n3503;
wire n3504;
wire n3505;
wire n3506;
wire n3507;
wire n3508;
wire n3509;
wire n3510;
wire n3511;
wire n3514;
wire n3515;
wire n3517;
wire n3518;
wire n3520;
wire n3521;
wire n3523;
wire n3524;
wire n3525;
wire n3526;
wire n3528;
wire n3529;
wire n3531;
wire n3532;
wire n3534;
wire n3535;
wire n3537;
wire n3538;
wire n3539;
wire n3540;
wire n3543;
wire n3544;
wire n3546;
wire n3547;
wire n3549;
wire n3550;
wire n3552;
wire n3553;
wire n3554;
wire n3555;
wire n3557;
wire n3558;
wire n3560;
wire n3561;
wire n3563;
wire n3564;
wire n3567;
wire n3568;
wire n3569;
wire n3570;
wire n3571;
wire n3572;
wire n3575;
wire n3576;
wire n3578;
wire n3579;
wire n3581;
wire n3582;
wire n3584;
wire n3585;
wire n3586;
wire n3587;
wire n3589;
wire n3590;
wire n3592;
wire n3593;
wire n3595;
wire n3596;
wire n3598;
wire n3599;
wire n3600;
wire n3601;
wire n3604;
wire n3605;
wire n3607;
wire n3608;
wire n3610;
wire n3611;
wire n3613;
wire n3614;
wire n3615;
wire n3616;
wire n3618;
wire n3619;
wire n3621;
wire n3622;
wire n3624;
wire n3625;
wire n3628;
wire n3629;
wire n3630;
wire n3631;
wire n3632;
wire n3633;
wire n3634;
wire n3635;
wire n3636;
wire n3639;
wire n3640;
wire n3642;
wire n3643;
wire n3645;
wire n3646;
wire n3648;
wire n3649;
wire n3650;
wire n3651;
wire n3653;
wire n3654;
wire n3656;
wire n3657;
wire n3659;
wire n3660;
wire n3662;
wire n3663;
wire n3664;
wire n3665;
wire n3668;
wire n3669;
wire n3671;
wire n3672;
wire n3674;
wire n3675;
wire n3677;
wire n3678;
wire n3679;
wire n3680;
wire n3682;
wire n3683;
wire n3685;
wire n3686;
wire n3688;
wire n3689;
wire n3692;
wire n3693;
wire n3694;
wire n3695;
wire n3696;
wire n3697;
wire n3700;
wire n3701;
wire n3703;
wire n3704;
wire n3706;
wire n3707;
wire n3709;
wire n3710;
wire n3711;
wire n3712;
wire n3714;
wire n3715;
wire n3717;
wire n3718;
wire n3720;
wire n3721;
wire n3723;
wire n3724;
wire n3725;
wire n3726;
wire n3729;
wire n3730;
wire n3732;
wire n3733;
wire n3735;
wire n3736;
wire n3738;
wire n3739;
wire n3740;
wire n3741;
wire n3743;
wire n3744;
wire n3746;
wire n3747;
wire n3749;
wire n3750;
wire n3753;
wire n3754;
wire n3755;
wire n3756;
wire n3757;
wire n3758;
wire n3759;
wire n3760;
wire n3761;
wire n3764;
wire n3765;
wire n3767;
wire n3768;
wire n3770;
wire n3771;
wire n3773;
wire n3774;
wire n3775;
wire n3776;
wire n3778;
wire n3779;
wire n3781;
wire n3782;
wire n3784;
wire n3785;
wire n3787;
wire n3788;
wire n3789;
wire n3790;
wire n3793;
wire n3794;
wire n3796;
wire n3797;
wire n3799;
wire n3800;
wire n3802;
wire n3803;
wire n3804;
wire n3805;
wire n3807;
wire n3808;
wire n3810;
wire n3811;
wire n3813;
wire n3814;
wire n3817;
wire n3818;
wire n3819;
wire n3820;
wire n3821;
wire n3822;
wire n3825;
wire n3826;
wire n3828;
wire n3829;
wire n3831;
wire n3832;
wire n3834;
wire n3835;
wire n3836;
wire n3837;
wire n3839;
wire n3840;
wire n3842;
wire n3843;
wire n3845;
wire n3846;
wire n3848;
wire n3849;
wire n3850;
wire n3851;
wire n3854;
wire n3855;
wire n3857;
wire n3858;
wire n3860;
wire n3861;
wire n3863;
wire n3864;
wire n3865;
wire n3866;
wire n3868;
wire n3869;
wire n3871;
wire n3872;
wire n3874;
wire n3875;
wire n3878;
wire n3879;
wire n3880;
wire n3881;
wire n3882;
wire n3883;
wire n3884;
wire n3885;
wire n3886;
wire n3889;
wire n3890;
wire n3892;
wire n3893;
wire n3895;
wire n3896;
wire n3898;
wire n3899;
wire n3900;
wire n3901;
wire n3903;
wire n3904;
wire n3906;
wire n3907;
wire n3909;
wire n3910;
wire n3912;
wire n3913;
wire n3914;
wire n3915;
wire n3918;
wire n3919;
wire n3921;
wire n3922;
wire n3924;
wire n3925;
wire n3927;
wire n3928;
wire n3929;
wire n3930;
wire n3932;
wire n3933;
wire n3935;
wire n3936;
wire n3938;
wire n3939;
wire n3942;
wire n3943;
wire n3944;
wire n3945;
wire n3946;
wire n3947;
wire n3950;
wire n3951;
wire n3953;
wire n3954;
wire n3956;
wire n3957;
wire n3959;
wire n3960;
wire n3961;
wire n3962;
wire n3964;
wire n3965;
wire n3967;
wire n3968;
wire n3970;
wire n3971;
wire n3973;
wire n3974;
wire n3975;
wire n3976;
wire n3979;
wire n3980;
wire n3982;
wire n3983;
wire n3985;
wire n3986;
wire n3988;
wire n3989;
wire n3990;
wire n3991;
wire n3993;
wire n3994;
wire n3996;
wire n3997;
wire n3999;
wire n4000;
wire n4003;
wire n4004;
wire n4005;
wire n4006;
wire n4007;
wire n4008;
wire n4009;
wire n4010;
wire n4013;
wire n4014;
wire n4016;
wire n4017;
wire n4019;
wire n4020;
wire n4022;
wire n4023;
wire n4024;
wire n4025;
wire n4027;
wire n4028;
wire n4030;
wire n4031;
wire n4033;
wire n4034;
wire n4036;
wire n4037;
wire n4038;
wire n4039;
wire n4042;
wire n4043;
wire n4045;
wire n4046;
wire n4048;
wire n4049;
wire n4051;
wire n4052;
wire n4053;
wire n4054;
wire n4056;
wire n4057;
wire n4059;
wire n4060;
wire n4062;
wire n4063;
wire n4066;
wire n4067;
wire n4068;
wire n4069;
wire n4070;
wire n4071;
wire n4074;
wire n4075;
wire n4077;
wire n4078;
wire n4080;
wire n4081;
wire n4083;
wire n4084;
wire n4085;
wire n4086;
wire n4088;
wire n4089;
wire n4091;
wire n4092;
wire n4094;
wire n4095;
wire n4097;
wire n4098;
wire n4099;
wire n4100;
wire n4103;
wire n4104;
wire n4106;
wire n4107;
wire n4109;
wire n4110;
wire n4112;
wire n4113;
wire n4114;
wire n4115;
wire n4117;
wire n4118;
wire n4120;
wire n4121;
wire n4123;
wire n4124;
wire n4127;
wire n4128;
wire n4129;
wire n4130;
wire n4131;
wire n4132;
wire n4133;
wire n4134;
wire n4135;
wire n4136;
wire n4137;
wire n4138;
wire n4139;
wire n4140;
wire n4141;
wire n4142;
wire n4143;
wire n4145;
wire n4147;
wire n4148;
wire n4149;
wire n4151;
wire n4153;
wire n4154;
wire n4155;
wire n4156;
wire n4158;
wire n4160;
wire n4161;
wire n4162;
wire n4163;
wire n4164;
wire n4165;
wire n4166;
wire n4167;
wire n4168;
wire n4169;
wire n4170;
wire n4171;
wire n4172;
wire n4173;
wire n4174;
wire n4175;
wire n4176;
wire n4177;
wire n4178;
wire n4179;
wire n4180;
wire n4181;
wire n4182;
wire n4183;
wire n4184;
wire n4185;
wire n4186;
wire n4187;
wire n4188;
wire n4189;
wire n4190;
wire n4191;
wire n4192;
wire n4193;
wire n4194;
wire n4195;
wire n4196;
wire n4197;
wire n4198;
wire n4199;
wire n4200;
wire n4201;
wire n4202;
wire n4203;
wire n4204;
wire n4206;
wire n4207;
wire n4208;
wire n4209;
wire n4210;
wire n4211;
wire n4212;
wire n4213;
wire n4214;
wire n4215;
wire n4216;
wire n4217;
wire n4218;
wire n4219;
wire n4220;
wire n4221;
wire n4222;
wire n4223;
wire n4224;
wire n4225;
wire n4226;
wire n4227;
wire n4228;
wire n4229;
wire n4230;
wire n4231;
wire n4232;
wire n4233;
wire n4234;
wire n4235;
wire n4236;
wire n4237;
wire n4238;
wire n4239;
wire n4240;
wire n4241;
wire n4242;
wire n4243;
wire n4244;
wire n4245;
wire n4246;
wire n4247;
wire n4249;
wire n4250;
wire n4251;
wire n4252;
wire n4253;
wire n4254;
wire n4255;
wire n4256;
wire n4257;
wire n4258;
wire n4259;
wire n4260;
wire n4261;
wire n4262;
wire n4263;
wire n4264;
wire n4265;
wire n4266;
wire n4267;
wire n4268;
wire n4269;
wire n4270;
wire n4271;
wire n4272;
wire n4273;
wire n4274;
wire n4275;
wire n4276;
wire n4277;
wire n4278;
wire n4279;
wire n4280;
wire n4281;
wire n4282;
wire n4283;
wire n4284;
wire n4285;
wire n4286;
wire n4287;
wire n4288;
wire n4289;
wire n4290;
wire n4291;
wire n4292;
wire n4293;
wire n4295;
wire n4296;
wire n4297;
wire n4298;
wire n4299;
wire n4300;
wire n4301;
wire n4302;
wire n4303;
wire n4304;
wire n4305;
wire n4306;
wire n4307;
wire n4308;
wire n4309;
wire n4310;
wire n4311;
wire n4312;
wire n4313;
wire n4314;
wire n4315;
wire n4316;
wire n4317;
wire n4318;
wire n4319;
wire n4320;
wire n4321;
wire n4322;
wire n4323;
wire n4324;
wire n4325;
wire n4326;
wire n4327;
wire n4328;
wire n4329;
wire n4330;
wire n4331;
wire n4332;
wire n4333;
wire n4334;
wire n4335;
wire n4336;
wire n4338;
wire n4339;
wire n4340;
wire n4341;
wire n4342;
wire n4343;
wire n4344;
wire n4345;
wire n4346;
wire n4347;
wire n4348;
wire n4349;
wire n4350;
wire n4351;
wire n4352;
wire n4353;
wire n4354;
wire n4355;
wire n4356;
wire n4357;
wire n4358;
wire n4359;
wire n4360;
wire n4361;
wire n4362;
wire n4363;
wire n4364;
wire n4365;
wire n4366;
wire n4367;
wire n4368;
wire n4369;
wire n4370;
wire n4371;
wire n4372;
wire n4373;
wire n4374;
wire n4375;
wire n4376;
wire n4377;
wire n4378;
wire n4379;
wire n4380;
wire n4381;
wire n4382;
wire n4384;
wire n4385;
wire n4386;
wire n4387;
wire n4388;
wire n4389;
wire n4390;
wire n4391;
wire n4392;
wire n4393;
wire n4394;
wire n4395;
wire n4396;
wire n4397;
wire n4398;
wire n4399;
wire n4400;
wire n4401;
wire n4402;
wire n4403;
wire n4404;
wire n4405;
wire n4406;
wire n4407;
wire n4408;
wire n4409;
wire n4410;
wire n4411;
wire n4412;
wire n4413;
wire n4414;
wire n4415;
wire n4416;
wire n4417;
wire n4418;
wire n4419;
wire n4420;
wire n4421;
wire n4422;
wire n4423;
wire n4424;
wire n4425;
wire n4427;
wire n4428;
wire n4429;
wire n4430;
wire n4431;
wire n4432;
wire n4433;
wire n4434;
wire n4435;
wire n4436;
wire n4437;
wire n4438;
wire n4439;
wire n4440;
wire n4441;
wire n4442;
wire n4443;
wire n4444;
wire n4445;
wire n4446;
wire n4447;
wire n4448;
wire n4449;
wire n4450;
wire n4451;
wire n4452;
wire n4453;
wire n4454;
wire n4455;
wire n4456;
wire n4457;
wire n4458;
wire n4459;
wire n4460;
wire n4461;
wire n4462;
wire n4463;
wire n4464;
wire n4465;
wire n4466;
wire n4467;
wire n4468;
wire n4469;
wire n4470;
wire n4471;
wire n4473;
wire n4474;
wire n4475;
wire n4476;
wire n4477;
wire n4478;
wire n4479;
wire n4480;
wire n4481;
wire n4482;
wire n4483;
wire n4484;
wire n4485;
wire n4486;
wire n4487;
wire n4488;
wire n4489;
wire n4490;
wire n4491;
wire n4492;
wire n4493;
wire n4494;
wire n4495;
wire n4496;
wire n4497;
wire n4498;
wire n4499;
wire n4500;
wire n4501;
wire n4502;
wire n4503;
wire n4504;
wire n4505;
wire n4506;
wire n4507;
wire n4508;
wire n4509;
wire n4510;
wire n4511;
wire n4512;
wire n4513;
wire n4514;
wire n4516;
wire n4517;
wire n4518;
wire n4519;
wire n4520;
wire n4521;
wire n4522;
wire n4523;
wire n4524;
wire n4525;
wire n4526;
wire n4527;
wire n4528;
wire n4529;
wire n4530;
wire n4531;
wire n4532;
wire n4533;
wire n4534;
wire n4535;
wire n4536;
wire n4537;
wire n4538;
wire n4539;
wire n4540;
wire n4541;
wire n4542;
wire n4543;
wire n4544;
wire n4545;
wire n4546;
wire n4547;
wire n4548;
wire n4549;
wire n4550;
wire n4551;
wire n4552;
wire n4553;
wire n4554;
wire n4555;
wire n4556;
wire n4557;
wire n4558;
wire n4559;
wire n4560;
wire n4562;
wire n4563;
wire n4564;
wire n4565;
wire n4566;
wire n4567;
wire n4568;
wire n4569;
wire n4570;
wire n4571;
wire n4572;
wire n4573;
wire n4574;
wire n4575;
wire n4576;
wire n4577;
wire n4578;
wire n4579;
wire n4580;
wire n4581;
wire n4582;
wire n4583;
wire n4584;
wire n4585;
wire n4586;
wire n4587;
wire n4588;
wire n4589;
wire n4590;
wire n4591;
wire n4592;
wire n4593;
wire n4594;
wire n4595;
wire n4596;
wire n4597;
wire n4598;
wire n4599;
wire n4600;
wire n4601;
wire n4602;
wire n4603;
wire n4605;
wire n4606;
wire n4607;
wire n4608;
wire n4609;
wire n4610;
wire n4611;
wire n4612;
wire n4613;
wire n4614;
wire n4615;
wire n4616;
wire n4617;
wire n4618;
wire n4619;
wire n4620;
wire n4621;
wire n4622;
wire n4623;
wire n4624;
wire n4625;
wire n4626;
wire n4627;
wire n4628;
wire n4629;
wire n4630;
wire n4631;
wire n4632;
wire n4633;
wire n4634;
wire n4635;
wire n4636;
wire n4637;
wire n4638;
wire n4639;
wire n4640;
wire n4641;
wire n4642;
wire n4643;
wire n4644;
wire n4645;
wire n4646;
wire n4647;
wire n4648;
wire n4649;
wire n4651;
wire n4652;
wire n4653;
wire n4654;
wire n4655;
wire n4656;
wire n4657;
wire n4658;
wire n4659;
wire n4660;
wire n4661;
wire n4662;
wire n4663;
wire n4664;
wire n4665;
wire n4666;
wire n4667;
wire n4668;
wire n4669;
wire n4670;
wire n4671;
wire n4672;
wire n4673;
wire n4674;
wire n4675;
wire n4676;
wire n4677;
wire n4678;
wire n4679;
wire n4680;
wire n4681;
wire n4682;
wire n4683;
wire n4684;
wire n4685;
wire n4686;
wire n4687;
wire n4688;
wire n4689;
wire n4690;
wire n4691;
wire n4692;
wire n4694;
wire n4695;
wire n4696;
wire n4697;
wire n4698;
wire n4699;
wire n4700;
wire n4701;
wire n4702;
wire n4703;
wire n4704;
wire n4705;
wire n4706;
wire n4707;
wire n4708;
wire n4709;
wire n4710;
wire n4711;
wire n4712;
wire n4713;
wire n4714;
wire n4715;
wire n4716;
wire n4717;
wire n4718;
wire n4719;
wire n4720;
wire n4721;
wire n4722;
wire n4723;
wire n4724;
wire n4725;
wire n4726;
wire n4727;
wire n4728;
wire n4729;
wire n4730;
wire n4731;
wire n4732;
wire n4733;
wire n4734;
wire n4735;
wire n4736;
wire n4737;
wire n4738;
wire n4740;
wire n4741;
wire n4742;
wire n4743;
wire n4744;
wire n4745;
wire n4746;
wire n4747;
wire n4748;
wire n4749;
wire n4750;
wire n4751;
wire n4752;
wire n4753;
wire n4754;
wire n4755;
wire n4756;
wire n4757;
wire n4758;
wire n4759;
wire n4760;
wire n4761;
wire n4762;
wire n4763;
wire n4764;
wire n4765;
wire n4766;
wire n4767;
wire n4768;
wire n4769;
wire n4770;
wire n4771;
wire n4772;
wire n4773;
wire n4774;
wire n4775;
wire n4776;
wire n4777;
wire n4778;
wire n4779;
wire n4780;
wire n4781;
wire n4783;
wire n4784;
wire n4785;
wire n4786;
wire n4787;
wire n4788;
wire n4789;
wire n4790;
wire n4791;
wire n4792;
wire n4793;
wire n4794;
wire n4795;
wire n4796;
wire n4797;
wire n4798;
wire n4799;
wire n4800;
wire n4801;
wire n4802;
wire n4803;
wire n4804;
wire n4805;
wire n4806;
wire n4807;
wire n4808;
wire n4809;
wire n4810;
wire n4811;
wire n4812;
wire n4813;
wire n4814;
wire n4815;
wire n4816;
wire n4817;
wire n4818;
wire n4819;
wire n4820;
wire n4821;
wire n4822;
wire n4823;
wire n4824;
wire n4825;
wire n4826;
wire n4828;
wire n4829;
wire n4830;
wire n4831;
wire n4832;
wire n4833;
wire n4834;
wire n4835;
wire n4836;
wire n4837;
wire n4838;
wire n4839;
wire n4840;
wire n4841;
wire n4842;
wire n4843;
wire n4844;
wire n4845;
wire n4846;
wire n4847;
wire n4848;
wire n4849;
wire n4850;
wire n4851;
wire n4852;
wire n4853;
wire n4854;
wire n4855;
wire n4856;
wire n4857;
wire n4858;
wire n4859;
wire n4860;
wire n4861;
wire n4862;
wire n4863;
wire n4864;
wire n4865;
wire n4866;
wire n4867;
wire n4868;
wire n4869;
wire n4871;
wire n4872;
wire n4873;
wire n4874;
wire n4875;
wire n4876;
wire n4877;
wire n4878;
wire n4879;
wire n4880;
wire n4881;
wire n4882;
wire n4883;
wire n4885;
wire n4887;
wire n4888;
wire n4889;
wire n4891;
wire n4893;
wire n4894;
wire n4895;
wire n4896;
wire n4898;
wire n4900;
wire n4901;
wire n4902;
wire n4903;
wire n4905;
wire n4907;
wire n4908;
wire n4909;
wire n4910;
wire n4912;
wire n4914;
wire n4915;
wire n4916;
wire n4917;
wire n4918;
wire n4919;
wire n4920;
wire n4921;
wire n4922;
wire n4923;
wire n4924;
wire n4927;
wire n4928;
wire n4930;
wire n4931;
wire n4933;
wire n4934;
wire n4936;
wire n4937;
wire n4938;
wire n4939;
wire n4941;
wire n4942;
wire n4944;
wire n4945;
wire n4947;
wire n4948;
wire n4951;
wire n4952;
wire n4953;
wire n4954;
wire n4955;
wire n4956;
wire n4959;
wire n4960;
wire n4962;
wire n4963;
wire n4965;
wire n4966;
wire n4968;
wire n4969;
wire n4970;
wire n4971;
wire n4973;
wire n4974;
wire n4976;
wire n4977;
wire n4979;
wire n4980;
wire n4982;
wire n4983;
wire n4985;
wire n4986;
wire n4987;
wire n4988;
wire n4989;
wire n4990;
wire n4991;
wire n4992;
wire n4993;
wire n4994;
wire n4995;
wire n4998;
wire n4999;
wire n5001;
wire n5002;
wire n5004;
wire n5005;
wire n5007;
wire n5008;
wire n5009;
wire n5010;
wire n5012;
wire n5013;
wire n5015;
wire n5016;
wire n5018;
wire n5019;
wire n5022;
wire n5023;
wire n5024;
wire n5025;
wire n5026;
wire n5027;
wire n5030;
wire n5031;
wire n5033;
wire n5034;
wire n5036;
wire n5037;
wire n5039;
wire n5040;
wire n5041;
wire n5042;
wire n5044;
wire n5045;
wire n5047;
wire n5048;
wire n5050;
wire n5051;
wire n5053;
wire n5054;
wire n5056;
wire n5057;
wire n5058;
wire n5059;
wire n5060;
wire n5061;
wire n5062;
wire n5063;
wire n5064;
wire n5065;
wire n5066;
wire n5069;
wire n5070;
wire n5072;
wire n5073;
wire n5075;
wire n5076;
wire n5078;
wire n5079;
wire n5080;
wire n5081;
wire n5083;
wire n5084;
wire n5086;
wire n5087;
wire n5089;
wire n5090;
wire n5093;
wire n5094;
wire n5095;
wire n5096;
wire n5097;
wire n5098;
wire n5101;
wire n5102;
wire n5104;
wire n5105;
wire n5107;
wire n5108;
wire n5110;
wire n5111;
wire n5112;
wire n5113;
wire n5115;
wire n5116;
wire n5118;
wire n5119;
wire n5121;
wire n5122;
wire n5124;
wire n5125;
wire n5127;
wire n5128;
wire n5129;
wire n5130;
wire n5131;
wire n5132;
wire n5133;
wire n5134;
wire n5135;
wire n5136;
wire n5137;
wire n5140;
wire n5141;
wire n5143;
wire n5144;
wire n5146;
wire n5147;
wire n5149;
wire n5150;
wire n5151;
wire n5152;
wire n5154;
wire n5155;
wire n5157;
wire n5158;
wire n5160;
wire n5161;
wire n5164;
wire n5165;
wire n5166;
wire n5167;
wire n5168;
wire n5169;
wire n5172;
wire n5173;
wire n5175;
wire n5176;
wire n5178;
wire n5179;
wire n5181;
wire n5182;
wire n5183;
wire n5184;
wire n5186;
wire n5187;
wire n5189;
wire n5190;
wire n5192;
wire n5193;
wire n5195;
wire n5196;
wire n5198;
wire n5199;
wire n5200;
wire n5201;
wire n5202;
wire n5203;
wire n5204;
wire n5205;
wire n5206;
wire n5207;
wire n5208;
wire n5211;
wire n5212;
wire n5214;
wire n5215;
wire n5217;
wire n5218;
wire n5220;
wire n5221;
wire n5222;
wire n5223;
wire n5225;
wire n5226;
wire n5228;
wire n5229;
wire n5231;
wire n5232;
wire n5235;
wire n5236;
wire n5237;
wire n5238;
wire n5239;
wire n5240;
wire n5243;
wire n5244;
wire n5246;
wire n5247;
wire n5249;
wire n5250;
wire n5252;
wire n5253;
wire n5254;
wire n5255;
wire n5257;
wire n5258;
wire n5260;
wire n5261;
wire n5263;
wire n5264;
wire n5266;
wire n5267;
wire n5269;
wire n5270;
wire n5271;
wire n5272;
wire n5273;
wire n5274;
wire n5275;
wire n5276;
wire n5277;
wire n5278;
wire n5279;
wire n5282;
wire n5283;
wire n5285;
wire n5286;
wire n5288;
wire n5289;
wire n5291;
wire n5292;
wire n5293;
wire n5294;
wire n5296;
wire n5297;
wire n5299;
wire n5300;
wire n5302;
wire n5303;
wire n5306;
wire n5307;
wire n5308;
wire n5309;
wire n5310;
wire n5311;
wire n5314;
wire n5315;
wire n5317;
wire n5318;
wire n5320;
wire n5321;
wire n5323;
wire n5324;
wire n5325;
wire n5326;
wire n5328;
wire n5329;
wire n5331;
wire n5332;
wire n5334;
wire n5335;
wire n5337;
wire n5338;
wire n5340;
wire n5341;
wire n5342;
wire n5343;
wire n5344;
wire n5345;
wire n5346;
wire n5347;
wire n5348;
wire n5349;
wire n5350;
wire n5353;
wire n5354;
wire n5356;
wire n5357;
wire n5359;
wire n5360;
wire n5362;
wire n5363;
wire n5364;
wire n5365;
wire n5367;
wire n5368;
wire n5370;
wire n5371;
wire n5373;
wire n5374;
wire n5377;
wire n5378;
wire n5379;
wire n5380;
wire n5381;
wire n5382;
wire n5385;
wire n5386;
wire n5388;
wire n5389;
wire n5391;
wire n5392;
wire n5394;
wire n5395;
wire n5396;
wire n5397;
wire n5399;
wire n5400;
wire n5402;
wire n5403;
wire n5405;
wire n5406;
wire n5408;
wire n5409;
wire n5411;
wire n5412;
wire n5413;
wire n5414;
wire n5415;
wire n5416;
wire n5417;
wire n5418;
wire n5419;
wire n5420;
wire n5423;
wire n5424;
wire n5426;
wire n5427;
wire n5429;
wire n5430;
wire n5432;
wire n5433;
wire n5434;
wire n5435;
wire n5437;
wire n5438;
wire n5440;
wire n5441;
wire n5443;
wire n5444;
wire n5447;
wire n5448;
wire n5449;
wire n5450;
wire n5451;
wire n5452;
wire n5455;
wire n5456;
wire n5458;
wire n5459;
wire n5461;
wire n5462;
wire n5464;
wire n5465;
wire n5466;
wire n5467;
wire n5469;
wire n5470;
wire n5472;
wire n5473;
wire n5475;
wire n5476;
wire n5478;
wire n5479;
wire n5481;
wire n5482;
wire n5483;
wire n5484;
wire n5485;
wire n5486;
wire n5487;
wire n5488;
wire n5489;
wire n5490;
wire n5491;
wire n5492;
wire n5493;
wire n5494;
wire n5495;
wire n5496;
wire n5497;
wire n5498;
wire n5499;
wire n5500;
wire n5501;
wire n5502;
wire n5503;
wire n5504;
wire n5505;
wire n5506;
wire n5507;
wire n5508;
wire n5509;
wire n5510;
wire n5511;
wire n5512;
wire n5513;
wire n5514;
wire n5515;
wire n5516;
wire n5517;
wire n5518;
wire n5519;
wire n5520;
wire n5521;
wire n5522;
wire n5523;
wire n5524;
wire n5525;
wire n5526;
wire n5527;
wire n5528;
wire n5529;
wire n5530;
wire n5531;
wire n5532;
wire n5533;
wire n5534;
wire n5535;
wire n5536;
wire n5537;
wire n5538;
wire n5539;
wire n5540;
wire n5541;
wire n5542;
wire n5543;
wire n5544;
wire n5545;
wire n5546;
wire n5547;
wire n5548;
wire n5549;
wire n5550;
wire n5551;
wire n5552;
wire n5553;
wire n5554;
wire n5555;
wire n5556;
wire n5557;
wire n5558;
wire n5559;
wire n5560;
wire n5561;
wire n5562;
wire n5563;
wire n5564;
wire n5565;
wire n5566;
wire n5567;
wire n5568;
wire n5569;
wire n5570;
wire n5571;
wire n5572;
wire n5573;
wire n5574;
wire n5575;
wire n5576;
wire n5577;
wire n5578;
wire n5579;
wire n5580;
wire n5581;
wire n5582;
wire n5583;
wire n5584;
wire n5585;
wire n5586;
wire n5587;
wire n5588;
wire n5589;
wire n5590;
wire n5591;
wire n5592;
wire n5593;
wire n5594;
wire n5595;
wire n5596;
wire n5597;
wire n5598;
wire n5599;
wire n5600;
wire n5601;
wire n5602;
wire n5603;
wire n5604;
wire n5605;
wire n5606;
wire n5607;
wire n5608;
wire n5609;
wire n5610;
wire n5611;
wire n5612;
wire n5613;
wire n5614;
wire n5615;
wire n5616;
wire n5617;
wire n5618;
wire n5619;
wire n5620;
wire n5621;
wire n5622;
wire n5623;
wire n5624;
wire n5625;
wire n5626;
wire n5627;
wire n5628;
wire n5629;
wire n5630;
wire n5631;
wire n5632;
wire n5633;
wire n5634;
wire n5635;
wire n5636;
wire n5637;
wire n5638;
wire n5639;
wire n5640;
wire n5641;
wire n5642;
wire n5643;
wire n5644;
wire n5645;
wire n5646;
wire n5647;
wire n5648;
wire n5649;
wire n5650;
wire n5651;
wire n5652;
wire n5653;
wire n5654;
wire n5655;
wire n5656;
wire n5657;
wire n5658;
wire n5659;
wire n5660;
wire n5661;
wire n5662;
wire n5663;
wire n5664;
wire n5665;
wire n5666;
wire n5667;
wire n5668;
wire n5669;
wire n5670;
wire n5671;
wire n5672;
wire n5673;
wire n5674;
wire n5675;
wire n5676;
wire n5677;
wire n5678;
wire n5679;
wire n5680;
wire n5681;
wire n5682;
wire n5683;
wire n5684;
wire n5685;
wire n5686;
wire n5687;
wire n5688;
wire n5689;
wire n5690;
wire n5691;
wire n5692;
wire n5693;
wire n5694;
wire n5695;
wire n5696;
wire n5697;
wire n5698;
wire n5699;
wire n5700;
wire n5701;
wire n5702;
wire n5703;
wire n5704;
wire n5705;
wire n5706;
wire n5707;
wire n5708;
wire n5709;
wire n5710;
wire n5711;
wire n5712;
wire n5713;
wire n5714;
wire n5715;
wire n5716;
wire n5717;
wire n5718;
wire n5719;
wire n5720;
wire n5721;
wire n5722;
wire n5723;
wire n5724;
wire n5725;
wire n5726;
wire n5727;
wire n5728;
wire n5729;
wire n5730;
wire n5731;
wire n5732;
wire n5733;
wire n5734;
wire n5735;
wire n5736;
wire n5737;
wire n5738;
wire n5739;
wire n5740;
wire n5741;
wire n5742;
wire n5743;
wire n5744;
wire n5745;
wire n5746;
wire n5747;
wire n5748;
wire n5749;
wire n5750;
wire n5751;
wire n5752;
wire n5753;
wire n5754;
wire n5755;
wire n5756;
wire n5757;
wire n5758;
wire n5759;
wire n5760;
wire n5761;
wire n5762;
wire n5763;
wire n5764;
wire n5765;
wire n5766;
wire n5767;
wire n5768;
wire n5769;
wire n5770;
wire n5771;
wire n5772;
wire n5773;
wire n5774;
wire n5775;
wire n5776;
wire n5777;
wire n5778;
wire n5779;
wire n5780;
wire n5781;
wire n5782;
wire n5783;
wire n5785;
wire n5787;
wire n5788;
wire n5789;
wire n5790;
wire n5791;
wire n5792;
wire n5794;
wire n5796;
wire n5797;
wire n5798;
wire n5799;
wire n5800;
wire n5801;
wire n5802;
wire n5803;
wire n5804;
wire n5805;
wire n5806;
wire n5807;
wire n5808;
wire n5810;
wire n5812;
wire n5813;
wire n5814;
wire n5815;
wire n5816;
wire n5817;
wire n5819;
wire n5821;
wire n5822;
wire n5823;
wire n5824;
wire n5826;
wire n5828;
wire n5829;
wire n5830;
wire n5831;
wire n5833;
wire n5835;
wire n5836;
wire n5837;
wire n5838;
wire n5839;
wire n5840;
wire n5841;
wire n5842;
wire n5843;
wire n5844;
wire n5845;
wire n5846;
wire n5847;
wire n5849;
wire n5851;
wire n5852;
wire n5853;
wire n5854;
wire n5855;
wire n5856;
wire n5858;
wire n5860;
wire n5861;
wire n5862;
wire n5863;
wire n5864;
wire n5865;
wire n5866;
wire n5867;
wire n5868;
wire n5869;
wire n5870;
wire n5871;
wire n5872;
wire n5873;
wire n5874;
wire n5875;
wire n5876;
wire n5877;
wire n5878;
wire n5879;
wire n5880;
wire n5881;
wire n5882;
wire n5883;
wire n5884;
wire n5885;
wire n5886;
wire n5887;
wire n5888;
wire n5889;
wire n5890;
wire n5891;
wire n5892;
wire n5893;
wire n5894;
wire n5895;
wire n5896;
wire n5897;
wire n5898;
wire n5899;
wire n5900;
wire n5901;
wire n5902;
wire n5903;
wire n5904;
wire n5905;
wire n5906;
wire n5907;
wire n5908;
wire n5909;
wire n5910;
wire n5911;
wire n5912;
wire n5913;
wire n5914;
wire n5915;
wire n5916;
wire n5917;
wire n5918;
wire n5919;
wire n5920;
wire n5921;
wire n5922;
wire n5923;
wire n5924;
wire n5925;
wire n5926;
wire n5927;
wire n5928;
wire n5929;
wire n5930;
wire n5931;
wire n5932;
wire n5933;
wire n5934;
wire n5935;
wire n5936;
wire n5937;
wire n5938;
wire n5939;
wire n5940;
wire n5941;
wire n5942;
wire n5943;
wire n5944;
wire n5945;
wire n5946;
wire n5947;
wire n5948;
wire n5949;
wire n5950;
wire n5951;
wire n5952;
wire n5953;
wire n5954;
wire n5955;
wire n5956;
wire n5957;
wire n5958;
wire n5959;
wire n5960;
wire n5961;
wire n5962;
wire n5963;
wire n5964;
wire n5965;
wire n5966;
wire n5967;
wire n5968;
wire n5969;
wire n5970;
wire n5971;
wire n5972;
wire n5973;
wire n5974;
wire n5975;
wire n5976;
wire n5977;
wire n5978;
wire n5979;
wire n5980;
wire n5981;
wire n5982;
wire n5983;
wire n5984;
wire n5985;
wire n5986;
wire n5987;
wire n5988;
wire n5989;
wire n5990;
wire n5991;
wire n5992;
wire n5993;
wire n5994;
wire n5995;
wire n5996;
wire n5997;
wire n5998;
wire n5999;
wire n6000;
wire n6001;
wire n6002;
wire n6003;
wire n6004;
wire n6005;
wire n6006;
wire n6007;
wire n6008;
wire n6009;
wire n6010;
wire n6011;
wire n6012;
wire n6013;
wire n6014;
wire n6015;
wire n6016;
wire n6017;
wire n6018;
wire n6019;
wire n6020;
wire n6021;
wire n6022;
wire n6023;
wire n6024;
wire n6026;
wire n6027;
wire n6029;
wire n6030;
wire n6031;
wire n6032;
wire n6033;
wire n6034;
wire n6035;
wire n6036;
wire n6037;
wire n6038;
wire n6039;
wire n6040;
wire n6041;
wire n6042;
wire n6043;
wire n6044;
wire n6045;
wire n6046;
wire n6047;
wire n6048;
wire n6049;
wire n6050;
wire n6051;
wire n6052;
wire n6053;
wire n6054;
wire n6055;
wire n6056;
wire n6057;
wire n6058;
wire n6059;
wire n6060;
wire n6061;
wire n6062;
wire n6063;
wire n6064;
wire n6065;
wire n6066;
wire n6067;
wire n6068;
wire n6069;
wire n6070;
wire n6071;
wire n6072;
wire n6073;
wire n6074;
wire n6075;
wire n6076;
wire n6077;
wire n6078;
wire n6079;
wire n6080;
wire n6081;
wire n6082;
wire n6083;
wire n6084;
wire n6085;
wire n6086;
wire n6087;
wire n6088;
wire n6089;
wire n6090;
wire n6091;
wire n6092;
wire n6093;
wire n6094;
wire n6095;
wire n6096;
wire n6097;
wire n6098;
wire n6099;
wire n6100;
wire n6101;
wire n6102;
wire n6103;
wire n6104;
wire n6105;
wire n6106;
wire n6107;
wire n6108;
wire n6109;
wire n6110;
wire n6111;
wire n6112;
wire n6113;
wire n6114;
wire n6115;
wire n6116;
wire n6117;
wire n6118;
wire n6119;
wire n6120;
wire n6121;
wire n6122;
wire n6123;
wire n6124;
wire n6125;
wire n6126;
wire n6127;
wire n6128;
wire n6129;
wire n6130;
wire n6131;
wire n6132;
wire n6133;
wire n6134;
wire n6135;
wire n6136;
wire n6138;
wire n6139;
wire n6141;
wire n6142;
wire n6143;
wire n6144;
wire n6145;
wire n6146;
wire n6147;
wire n6148;
wire n6149;
wire n6150;
wire n6151;
wire n6152;
wire n6153;
wire n6154;
wire n6155;
wire n6156;
wire n6157;
wire n6158;
wire n6159;
wire n6160;
wire n6161;
wire n6162;
wire n6163;
wire n6164;
wire n6165;
wire n6166;
wire n6167;
wire n6168;
wire n6169;
wire n6170;
wire n6171;
wire n6172;
wire n6173;
wire n6174;
wire n6175;
wire n6176;
wire n6177;
wire n6178;
wire n6179;
wire n6180;
wire n6181;
wire n6182;
wire n6183;
wire n6184;
wire n6185;
wire n6186;
wire n6187;
wire n6188;
wire n6189;
wire n6190;
wire n6191;
wire n6192;
wire n6193;
wire n6194;
wire n6195;
wire n6196;
wire n6197;
wire n6198;
wire n6199;
wire n6200;
wire n6201;
wire n6202;
wire n6203;
wire n6204;
wire n6205;
wire n6206;
wire n6207;
wire n6208;
wire n6209;
wire n6210;
wire n6211;
wire n6212;
wire n6213;
wire n6214;
wire n6215;
wire n6216;
wire n6217;
wire n6218;
wire n6219;
wire n6220;
wire n6221;
wire n6222;
wire n6223;
wire n6224;
wire n6225;
wire n6226;
wire n6227;
wire n6228;
wire n6229;
wire n6230;
wire n6231;
wire n6232;
wire n6233;
wire n6234;
wire n6235;
wire n6236;
wire n6237;
wire n6238;
wire n6239;
wire n6240;
wire n6241;
wire n6242;
wire n6243;
wire n6244;
wire n6245;
wire n6246;
wire n6247;
wire n6248;
wire n6250;
wire n6251;
wire n6253;
wire n6254;
wire n6255;
wire n6256;
wire n6257;
wire n6258;
wire n6259;
wire n6260;
wire n6261;
wire n6262;
wire n6263;
wire n6264;
wire n6265;
wire n6266;
wire n6267;
wire n6268;
wire n6269;
wire n6270;
wire n6271;
wire n6272;
wire n6273;
wire n6274;
wire n6275;
wire n6276;
wire n6277;
wire n6278;
wire n6279;
wire n6280;
wire n6281;
wire n6282;
wire n6283;
wire n6284;
wire n6285;
wire n6286;
wire n6287;
wire n6288;
wire n6289;
wire n6290;
wire n6291;
wire n6292;
wire n6293;
wire n6294;
wire n6295;
wire n6296;
wire n6297;
wire n6298;
wire n6299;
wire n6300;
wire n6301;
wire n6302;
wire n6303;
wire n6304;
wire n6305;
wire n6306;
wire n6307;
wire n6308;
wire n6309;
wire n6310;
wire n6311;
wire n6312;
wire n6313;
wire n6314;
wire n6315;
wire n6316;
wire n6317;
wire n6318;
wire n6319;
wire n6320;
wire n6321;
wire n6322;
wire n6323;
wire n6324;
wire n6325;
wire n6326;
wire n6327;
wire n6328;
wire n6329;
wire n6330;
wire n6331;
wire n6332;
wire n6333;
wire n6334;
wire n6335;
wire n6336;
wire n6337;
wire n6338;
wire n6339;
wire n6340;
wire n6341;
wire n6342;
wire n6343;
wire n6344;
wire n6345;
wire n6346;
wire n6347;
wire n6348;
wire n6349;
wire n6350;
wire n6351;
wire n6352;
wire n6353;
wire n6354;
wire n6355;
wire n6356;
wire n6357;
wire n6358;
wire n6359;
wire n6360;
wire n6362;
wire n6363;
wire n6365;
wire n6366;
wire n6367;
wire n6368;
wire n6369;
wire n6370;
wire n6371;
wire n6372;
wire n6373;
wire n6374;
wire n6375;
wire n6376;
wire n6377;
wire n6378;
wire n6379;
wire n6380;
wire n6381;
wire n6382;
wire n6383;
wire n6384;
wire n6385;
wire n6386;
wire n6387;
wire n6388;
wire n6389;
wire n6390;
wire n6391;
wire n6392;
wire n6393;
wire n6394;
wire n6395;
wire n6396;
wire n6397;
wire n6398;
wire n6399;
wire n6400;
wire n6401;
wire n6402;
wire n6403;
wire n6404;
wire n6405;
wire n6406;
wire n6407;
wire n6408;
wire n6409;
wire n6410;
wire n6411;
wire n6412;
wire n6413;
wire n6414;
wire n6415;
wire n6416;
wire n6417;
wire n6418;
wire n6419;
wire n6420;
wire n6421;
wire n6422;
wire n6423;
wire n6424;
wire n6425;
wire n6426;
wire n6427;
wire n6428;
wire n6429;
wire n6430;
wire n6431;
wire n6432;
wire n6433;
wire n6434;
wire n6435;
wire n6436;
wire n6437;
wire n6438;
wire n6439;
wire n6440;
wire n6441;
wire n6442;
wire n6443;
wire n6444;
wire n6445;
wire n6446;
wire n6447;
wire n6448;
wire n6449;
wire n6450;
wire n6451;
wire n6452;
wire n6453;
wire n6454;
wire n6455;
wire n6456;
wire n6457;
wire n6458;
wire n6459;
wire n6460;
wire n6461;
wire n6462;
wire n6463;
wire n6464;
wire n6465;
wire n6466;
wire n6467;
wire n6468;
wire n6470;
wire n6471;
wire n6473;
wire n6474;
wire n6475;
wire n6476;
wire n6477;
wire n6478;
wire n6479;
wire n6480;
wire n6481;
wire n6482;
wire n6483;
wire n6484;
wire n6485;
wire n6486;
wire n6487;
wire n6488;
wire n6489;
wire n6490;
wire n6491;
wire n6492;
wire n6493;
wire n6494;
wire n6495;
wire n6496;
wire n6497;
wire n6498;
wire n6499;
wire n6500;
wire n6501;
wire n6502;
wire n6503;
wire n6504;
wire n6505;
wire n6506;
wire n6507;
wire n6508;
wire n6509;
wire n6510;
wire n6511;
wire n6512;
wire n6513;
wire n6514;
wire n6515;
wire n6516;
wire n6517;
wire n6518;
wire n6519;
wire n6520;
wire n6521;
wire n6522;
wire n6523;
wire n6524;
wire n6525;
wire n6526;
wire n6527;
wire n6528;
wire n6529;
wire n6530;
wire n6531;
wire n6532;
wire n6533;
wire n6534;
wire n6535;
wire n6536;
wire n6537;
wire n6538;
wire n6539;
wire n6540;
wire n6541;
wire n6542;
wire n6543;
wire n6544;
wire n6545;
wire n6546;
wire n6547;
wire n6548;
wire n6549;
wire n6550;
wire n6551;
wire n6552;
wire n6553;
wire n6554;
wire n6555;
wire n6556;
wire n6557;
wire n6558;
wire n6559;
wire n6560;
wire n6561;
wire n6562;
wire n6563;
wire n6564;
wire n6565;
wire n6566;
wire n6567;
wire n6568;
wire n6569;
wire n6570;
wire n6571;
wire n6572;
wire n6573;
wire n6574;
wire n6575;
wire n6576;
wire n6578;
wire n6579;
wire n6581;
wire n6582;
wire n6583;
wire n6584;
wire n6585;
wire n6586;
wire n6587;
wire n6588;
wire n6589;
wire n6590;
wire n6591;
wire n6592;
wire n6593;
wire n6594;
wire n6595;
wire n6596;
wire n6597;
wire n6598;
wire n6599;
wire n6600;
wire n6601;
wire n6602;
wire n6603;
wire n6604;
wire n6605;
wire n6606;
wire n6607;
wire n6608;
wire n6609;
wire n6610;
wire n6611;
wire n6612;
wire n6613;
wire n6614;
wire n6615;
wire n6616;
wire n6617;
wire n6618;
wire n6619;
wire n6620;
wire n6621;
wire n6622;
wire n6623;
wire n6624;
wire n6625;
wire n6626;
wire n6627;
wire n6628;
wire n6629;
wire n6630;
wire n6631;
wire n6632;
wire n6633;
wire n6634;
wire n6635;
wire n6636;
wire n6637;
wire n6638;
wire n6639;
wire n6640;
wire n6641;
wire n6642;
wire n6643;
wire n6644;
wire n6645;
wire n6646;
wire n6647;
wire n6648;
wire n6649;
wire n6650;
wire n6651;
wire n6652;
wire n6653;
wire n6654;
wire n6655;
wire n6656;
wire n6657;
wire n6658;
wire n6659;
wire n6660;
wire n6661;
wire n6662;
wire n6663;
wire n6664;
wire n6665;
wire n6666;
wire n6667;
wire n6668;
wire n6669;
wire n6670;
wire n6671;
wire n6672;
wire n6673;
wire n6674;
wire n6675;
wire n6676;
wire n6677;
wire n6678;
wire n6679;
wire n6680;
wire n6681;
wire n6682;
wire n6683;
wire n6685;
wire n6686;
wire n6688;
wire n6689;
wire n6690;
wire n6691;
wire n6692;
wire n6693;
wire n6694;
wire n6695;
wire n6696;
wire n6697;
wire n6698;
wire n6699;
wire n6700;
wire n6701;
wire n6702;
wire n6703;
wire n6704;
wire n6705;
wire n6706;
wire n6707;
wire n6708;
wire n6709;
wire n6710;
wire n6711;
wire n6712;
wire n6713;
wire n6714;
wire n6715;
wire n6716;
wire n6717;
wire n6718;
wire n6719;
wire n6720;
wire n6721;
wire n6722;
wire n6723;
wire n6724;
wire n6725;
wire n6726;
wire n6727;
wire n6728;
wire n6729;
wire n6730;
wire n6731;
wire n6732;
wire n6733;
wire n6734;
wire n6735;
wire n6736;
wire n6737;
wire n6738;
wire n6739;
wire n6740;
wire n6741;
wire n6742;
wire n6743;
wire n6744;
wire n6745;
wire n6746;
wire n6747;
wire n6748;
wire n6749;
wire n6750;
wire n6751;
wire n6752;
wire n6753;
wire n6754;
wire n6755;
wire n6756;
wire n6757;
wire n6758;
wire n6759;
wire n6760;
wire n6761;
wire n6762;
wire n6763;
wire n6764;
wire n6765;
wire n6766;
wire n6767;
wire n6768;
wire n6769;
wire n6770;
wire n6771;
wire n6772;
wire n6773;
wire n6774;
wire n6775;
wire n6776;
wire n6777;
wire n6778;
wire n6779;
wire n6780;
wire n6781;
wire n6782;
wire n6783;
wire n6784;
wire n6785;
wire n6786;
wire n6787;
wire n6788;
wire n6789;
wire n6790;
wire n6791;
wire n6792;
wire n6793;
wire n6794;
wire n6795;
wire n6796;
wire n6797;
wire n6798;
wire n6799;
wire n6800;
wire n6801;
wire n6802;
wire n6803;
wire n6804;
wire n6805;
wire n6806;
wire n6807;
wire n6808;
wire n6809;
wire n6810;
wire n6811;
wire n6812;
wire n6813;
wire n6814;
wire n6815;
wire n6816;
wire n6817;
wire n6818;
wire n6819;
wire n6820;
wire n6821;
wire n6822;
wire n6823;
wire n6824;
wire n6825;
wire n6826;
wire n6827;
wire n6828;
wire n6829;
wire n6830;
wire n6831;
wire n6832;
wire n6833;
wire n6834;
wire n6835;
wire n6836;
wire n6838;
wire n6839;
wire n6840;
wire n6841;
wire n6842;
wire n6843;
wire n6844;
wire n6845;
wire n6846;
wire n6847;
wire n6849;
wire n6850;
wire n6852;
wire n6854;
wire n6856;
wire n6857;
wire n6858;
wire n6860;
wire n6861;
wire n6863;
wire n6865;
wire n6867;
wire n6868;
wire n6869;
wire n6871;
wire n6872;
wire n6874;
wire n6876;
wire n6878;
wire n6879;
wire n6880;
wire n6882;
wire n6883;
wire n6885;
wire n6887;
wire n6889;
wire n6890;
wire n6891;
wire n6892;
wire n6893;
wire n6894;
wire n6895;
wire n6896;
wire n6897;
wire n6898;
wire n6899;
wire n6901;
wire n6902;
wire n6904;
wire n6906;
wire n6908;
wire n6909;
wire n6910;
wire n6912;
wire n6913;
wire n6915;
wire n6917;
wire n6919;
wire n6920;
wire n6921;
wire n6923;
wire n6924;
wire n6926;
wire n6928;
wire n6930;
wire n6931;
wire n6932;
wire n6934;
wire n6935;
wire n6937;
wire n6939;
wire n6941;
wire n6942;
wire n6943;
wire n6944;
wire n6945;
wire n6946;
wire n6947;
wire n6948;
wire n6949;
wire n6950;
wire n6951;
wire n6952;
wire n6953;
wire n6954;
wire n6955;
wire n6956;
wire n6957;
wire n6958;
wire n6959;
wire n6960;
wire n6961;
wire n6962;
wire n6963;
wire n6964;
wire n6965;
wire n6966;
wire n6967;
wire n6968;
wire n6969;
wire n6970;
wire n6971;
wire n6972;
wire n6973;
wire n6974;
wire n6975;
wire n6976;
wire n6977;
wire n6978;
wire n6980;
wire n6981;
wire n6982;
wire n6983;
wire n6984;
wire n6985;
wire n6986;
wire n6987;
wire n6988;
wire n6989;
wire n6990;
wire n6991;
wire n6992;
wire n6993;
wire n6994;
wire n6995;
wire n6996;
wire n6997;
wire n6998;
wire n6999;
wire n7001;
wire n7002;
wire n7003;
wire n7004;
wire n7005;
wire n7006;
wire n7007;
wire n7008;
wire n7009;
wire n7010;
wire n7011;
wire n7012;
wire n7014;
wire n7015;
wire n7016;
wire n7017;
wire n7018;
wire n7019;
wire n7020;
wire n7021;
wire n7022;
wire n7023;
wire n7024;
wire n7025;
wire n7027;
wire n7028;
wire n7029;
wire n7030;
wire n7031;
wire n7032;
wire n7033;
wire n7034;
wire n7035;
wire n7036;
wire n7037;
wire n7038;
wire n7040;
wire n7041;
wire n7042;
wire n7043;
wire n7044;
wire n7045;
wire n7046;
wire n7047;
wire n7048;
wire n7049;
wire n7050;
wire n7051;
wire n7053;
wire n7054;
wire n7055;
wire n7056;
wire n7057;
wire n7058;
wire n7059;
wire n7060;
wire n7061;
wire n7062;
wire n7063;
wire n7065;
wire n7066;
wire n7067;
wire n7068;
wire n7069;
wire n7070;
wire n7071;
wire n7072;
wire n7073;
wire n7074;
wire n7075;
wire n7076;
wire n7077;
wire n7078;
wire n7079;
wire n7080;
wire n7081;
wire n7082;
wire n7083;
wire n7084;
wire n7085;
wire n7086;
wire n7087;
wire n7088;
wire n7089;
wire n7090;
wire n7091;
wire n7092;
wire n7093;
wire n7094;
wire n7095;
wire n7096;
wire n7097;
wire n7098;
wire n7099;
wire n7100;
wire n7101;
wire n7102;
wire n7103;
wire n7104;
wire n7105;
wire n7106;
wire n7107;
wire n7108;
wire n7109;
wire n7110;
wire n7111;
wire n7112;
wire n7113;
wire n7114;
wire n7115;
wire n7116;
wire n7117;
wire n7118;
wire n7119;
wire n7120;
wire n7121;
wire n7122;
wire n7123;
wire n7124;
wire n7125;
wire n7126;
wire n7127;
wire n7128;
wire n7129;
wire n7130;
wire n7131;
wire n7132;
wire n7133;
wire n7134;
wire n7135;
wire n7136;
wire n7137;
wire n7138;
wire n7139;
wire n7140;
wire n7141;
wire n7143;
wire n7144;
wire n7145;
wire n7146;
wire n7147;
wire n7148;
wire n7149;
wire n7150;
wire n7152;
wire n7153;
wire n7154;
wire n7155;
wire n7156;
wire n7157;
wire n7158;
wire n7159;
wire n7160;
wire n7161;
wire n7162;
wire n7163;
wire n7164;
wire n7165;
wire n7167;
wire n7168;
wire n7169;
wire n7170;
wire n7171;
wire n7172;
wire n7173;
wire n7174;
wire n7175;
wire n7176;
wire n7177;
wire n7178;
wire n7179;
wire n7180;
wire n7181;
wire n7182;
wire n7183;
wire n7184;
wire n7185;
wire n7186;
wire n7187;
wire n7188;
wire n7190;
wire n7191;
wire n7192;
wire n7193;
wire n7194;
wire n7195;
wire n7196;
wire n7197;
wire n7198;
wire n7199;
wire n7200;
wire n7201;
wire n7203;
wire n7204;
wire n7205;
wire n7206;
wire n7207;
wire n7208;
wire n7209;
wire n7210;
wire n7211;
wire n7212;
wire n7213;
wire n7214;
wire n7215;
wire n7216;
wire n7217;
wire n7218;
wire n7219;
wire n7221;
wire n7222;
wire n7223;
wire n7224;
wire n7225;
wire n7226;
wire n7227;
wire n7228;
wire n7229;
wire n7230;
wire n7231;
wire n7232;
wire n7233;
wire n7234;
wire n7235;
wire n7236;
wire n7237;
wire n7238;
wire n7239;
wire n7240;
wire n7241;
wire n7242;
wire n7243;
wire n7244;
wire n7245;
wire n7246;
wire n7248;
wire n7249;
wire n7250;
wire n7251;
wire n7252;
wire n7253;
wire n7254;
wire n7255;
wire n7256;
wire n7257;
wire n7258;
wire n7259;
wire n7260;
wire n7261;
wire n7262;
wire n7263;
wire n7264;
wire n7265;
wire n7266;
wire n7268;
wire n7269;
wire n7270;
wire n7271;
wire n7272;
wire n7273;
wire n7274;
wire n7275;
wire n7276;
wire n7277;
wire n7278;
wire n7279;
wire n7280;
wire n7281;
wire n7282;
wire n7283;
wire n7284;
wire n7285;
wire n7286;
wire n7287;
wire n7288;
wire n7289;
wire n7290;
wire n7291;
wire n7292;
wire n7293;
wire n7294;
wire n7295;
wire n7296;
wire n7297;
wire n7298;
wire n7299;
wire n7300;
wire n7301;
wire n7302;
wire n7303;
wire n7304;
wire n7305;
wire n7306;
wire n7307;
wire n7308;
wire n7309;
wire n7310;
wire n7311;
wire n7312;
wire n7313;
wire n7314;
wire n7315;
wire n7316;
wire n7317;
wire n7318;
wire n7319;
wire n7320;
wire n7321;
wire n7322;
wire n7323;
wire n7324;
wire n7325;
wire n7327;
wire n7328;
wire n7329;
wire n7330;
wire n7331;
wire n7332;
wire n7333;
wire n7334;
wire n7335;
wire n7336;
wire n7338;
wire n7339;
wire n7340;
wire n7341;
wire n7342;
wire n7343;
wire n7344;
wire n7345;
wire n7347;
wire n7348;
wire n7349;
wire n7350;
wire n7351;
wire n7352;
wire n7353;
wire n7354;
wire n7355;
wire n7356;
wire n7357;
wire n7358;
wire n7359;
wire n7360;
wire n7361;
wire n7363;
wire n7364;
wire n7365;
wire n7366;
wire n7367;
wire n7368;
wire n7369;
wire n7370;
wire n7371;
wire n7372;
wire n7373;
wire n7374;
wire n7376;
wire n7377;
wire n7378;
wire n7379;
wire n7380;
wire n7381;
wire n7382;
wire n7383;
wire n7384;
wire n7385;
wire n7386;
wire n7387;
wire n7389;
wire n7390;
wire n7391;
wire n7392;
wire n7393;
wire n7394;
wire n7395;
wire n7396;
wire n7397;
wire n7398;
wire n7399;
wire n7401;
wire n7402;
wire n7403;
wire n7404;
wire n7405;
wire n7406;
wire n7407;
wire n7408;
wire n7409;
wire n7410;
wire n7411;
wire n7412;
wire n7413;
wire n7414;
wire n7415;
wire n7416;
wire n7417;
wire n7418;
wire n7419;
wire n7420;
wire n7421;
wire n7422;
wire n7423;
wire n7424;
wire n7425;
wire n7426;
wire n7427;
wire n7428;
wire n7429;
wire n7430;
wire n7431;
wire n7432;
wire n7433;
wire n7434;
wire n7435;
wire n7436;
wire n7437;
wire n7438;
wire n7439;
wire n7440;
wire n7441;
wire n7443;
wire n7444;
wire n7445;
wire n7446;
wire n7447;
wire n7448;
wire n7449;
wire n7450;
wire n7451;
wire n7453;
wire n7454;
wire n7455;
wire n7456;
wire n7457;
wire n7458;
wire n7459;
wire n7460;
wire n7461;
wire n7462;
wire n7463;
wire n7465;
wire n7466;
wire n7467;
wire n7468;
wire n7469;
wire n7470;
wire n7471;
wire n7472;
wire n7473;
wire n7474;
wire n7475;
wire n7476;
wire n7477;
wire n7478;
wire n7479;
wire n7480;
wire n7481;
wire n7482;
wire n7483;
wire n7484;
wire n7485;
wire n7486;
wire n7487;
wire n7488;
wire n7489;
wire n7490;
wire n7491;
wire n7492;
wire n7493;
wire n7494;
wire n7495;
wire n7496;
wire n7498;
wire n7499;
wire n7500;
wire n7501;
wire n7502;
wire n7503;
wire n7504;
wire n7505;
wire n7506;
wire n7507;
wire n7508;
wire n7509;
wire n7510;
wire n7511;
wire n7512;
wire n7513;
wire n7514;
wire n7515;
wire n7516;
wire n7517;
wire n7518;
wire n7519;
wire n7520;
wire n7521;
wire n7522;
wire n7523;
wire n7524;
wire n7525;
wire n7526;
wire n7527;
wire n7528;
wire n7529;
wire n7530;
wire n7531;
wire n7532;
wire n7533;
wire n7534;
wire n7535;
wire n7536;
wire n7537;
wire n7538;
wire n7539;
wire n7540;
wire n7541;
wire n7542;
wire n7543;
wire n7544;
wire n7545;
wire n7546;
wire n7547;
wire n7548;
wire n7549;
wire n7550;
wire n7551;
wire n7552;
wire n7553;
wire n7555;
wire n7556;
wire n7557;
wire n7558;
wire n7559;
wire n7560;
wire n7561;
wire n7562;
wire n7563;
wire n7564;
wire n7565;
wire n7566;
wire n7567;
wire n7568;
wire n7569;
wire n7570;
wire n7571;
wire n7572;
wire n7573;
wire n7574;
wire n7575;
wire n7576;
wire n7577;
wire n7578;
wire n7579;
wire n7580;
wire n7581;
wire n7583;
wire n7584;
wire n7585;
wire n7586;
wire n7587;
wire n7588;
wire n7589;
wire n7590;
wire n7591;
wire n7592;
wire n7593;
wire n7594;
wire n7595;
wire n7596;
wire n7597;
wire n7598;
wire n7599;
wire n7600;
wire n7601;
wire n7602;
wire n7603;
wire n7604;
wire n7606;
wire n7607;
wire n7608;
wire n7609;
wire n7610;
wire n7611;
wire n7612;
wire n7613;
wire n7614;
wire n7615;
wire n7616;
wire n7617;
wire n7618;
wire n7619;
wire n7620;
wire n7621;
wire n7622;
wire n7623;
wire n7624;
wire n7625;
wire n7626;
wire n7627;
wire n7628;
wire n7629;
wire n7630;
wire n7631;
wire n7632;
wire n7633;
wire n7635;
wire n7636;
wire n7637;
wire n7638;
wire n7639;
wire n7640;
wire n7641;
wire n7642;
wire n7643;
wire n7644;
wire n7645;
wire n7646;
wire n7647;
wire n7648;
wire n7649;
wire n7650;
wire n7651;
wire n7652;
wire n7653;
wire n7654;
wire n7656;
wire n7657;
wire n7658;
wire n7659;
wire n7660;
wire n7661;
wire n7662;
wire n7663;
wire n7664;
wire n7665;
wire n7666;
wire n7667;
wire n7668;
wire n7669;
wire n7670;
wire n7671;
wire n7672;
wire n7673;
wire n7674;
wire n7675;
wire n7676;
wire n7677;
wire n7678;
wire n7679;
wire n7680;
wire n7681;
wire n7682;
wire n7683;
wire n7684;
wire n7685;
wire n7686;
wire n7687;
wire n7688;
wire n7689;
wire n7690;
wire n7691;
wire n7692;
wire n7693;
wire n7694;
wire n7695;
wire n7696;
wire n7697;
wire n7698;
wire n7699;
wire n7700;
wire n7701;
wire n7702;
wire n7703;
wire n7704;
wire n7705;
wire n7706;
wire n7707;
wire n7708;
wire n7709;
wire n7710;
wire n7711;
wire n7712;
wire n7713;
wire n7714;
wire n7715;
wire n7716;
wire n7717;
wire n7718;
wire n7719;
wire n7720;
wire n7721;
wire n7722;
wire n7723;
wire n7724;
wire n7725;
wire n7726;
wire n7727;
wire n7728;
wire n7729;
wire n7730;
wire n7731;
wire n7732;
wire n7733;
wire n7734;
wire n7735;
wire n7736;
wire n7737;
wire n7738;
wire n7739;
wire n7740;
wire n7741;
wire n7742;
wire n7743;
wire n7744;
wire n7745;
wire n7746;
wire n7747;
wire n7748;
wire n7749;
wire n7750;
wire n7751;
wire n7752;
wire n7753;
wire n7754;
wire n7755;
wire n7756;
wire n7757;
wire n7758;
wire n7759;
wire n7760;
wire n7761;
wire n7762;
wire n7763;
wire n7764;
wire n7765;
wire n7766;
wire n7767;
wire n7768;
wire n7769;
wire n7770;
wire n7771;
wire n7772;
wire n7773;
wire n7774;
wire n7775;
wire n7776;
wire n7777;
wire n7778;
wire n7779;
wire n7780;
wire n7781;
wire n7782;
wire n7783;
wire n7784;
wire n7785;
wire n7786;
wire n7787;
wire n7788;
wire n7789;
wire n7790;
wire n7791;
wire n7792;
wire n7793;
wire n7794;
wire n7795;
wire n7796;
wire n7797;
wire n7798;
wire n7799;
wire n7800;
wire n7801;
wire n7802;
wire n7803;
wire n7804;
wire n7805;
wire n7806;
wire n7807;
wire n7808;
wire n7809;
wire n7810;
wire n7811;
wire n7812;
wire n7813;
wire n7814;
wire n7815;
wire n7816;
wire n7817;
wire n7818;
wire n7819;
wire n7820;
wire n7821;
wire n7822;
wire n7823;
wire n7824;
wire n7825;
wire n7826;
wire n7827;
wire n7828;
wire n7829;
wire n7830;
wire n7831;
wire n7832;
wire n7833;
wire n7834;
wire n7835;
wire n7836;
wire n7837;
wire n7838;
wire n7839;
wire n7840;
wire n7841;
wire n7842;
wire n7843;
wire n7844;
wire n7845;
wire n7846;
wire n7847;
wire n7848;
wire n7849;
wire n7850;
wire n7851;
wire n7852;
wire n7853;
wire n7854;
wire n7855;
wire n7856;
wire n7857;
wire n7858;
wire n7859;
wire n7860;
wire n7861;
wire n7862;
wire n7863;
wire n7864;
wire n7865;
wire n7866;
wire n7867;
wire n7868;
wire n7869;
wire n7870;
wire n7871;
wire n7872;
wire n7873;
wire n7874;
wire n7875;
wire n7876;
wire n7877;
wire n7878;
wire n7879;
wire n7880;
wire n7881;
wire n7882;
wire n7883;
wire n7884;
wire n7885;
wire n7886;
wire n7887;
wire n7888;
wire n7889;
wire n7890;
wire n7891;
wire n7892;
wire n7893;
wire n7894;
wire n7895;
wire n7896;
wire n7897;
wire n7898;
wire n7899;
wire n7900;
wire n7901;
wire n7902;
wire n7903;
wire n7904;
wire n7905;
wire n7906;
wire n7907;
wire n7908;
wire n7909;
wire n7910;
wire n7911;
wire n7912;
wire n7913;
wire n7914;
wire n7915;
wire n7916;
wire n7917;
wire n7918;
wire n7919;
wire n7920;
wire n7921;
wire n7922;
wire n7923;
wire n7924;
wire n7925;
wire n7926;
wire n7927;
wire n7928;
wire n7929;
wire n7930;
wire n7931;
wire n7932;
wire n7933;
wire n7934;
wire n7935;
wire n7936;
wire n7937;
wire n7938;
wire n7939;
wire n7940;
wire n7941;
wire n7942;
wire n7943;
wire n7944;
wire n7945;
wire n7946;
wire n7947;
wire n7948;
wire n7949;
wire n7950;
wire n7951;
wire n7952;
wire n7953;
wire n7954;
wire n7955;
wire n7956;
wire n7957;
wire n7958;
wire n7959;
wire n7960;
wire n7961;
wire n7962;
wire n7963;
wire n7964;
wire n7965;
wire n7966;
wire n7967;
wire n7968;
wire n7969;
wire n7970;
wire n7971;
wire n7972;
wire n7973;
wire n7974;
wire n7975;
wire n7976;
wire n7977;
wire n7978;
wire n7979;
wire n7980;
wire n7981;
wire n7982;
wire n7983;
wire n7984;
wire n7985;
wire n7986;
wire n7987;
wire n7988;
wire n7989;
wire n7990;
wire n7991;
wire n7992;
wire n7993;
wire n7994;
wire n7995;
wire n7996;
wire n7997;
wire n7998;
wire n7999;
wire n8000;
wire n8001;
wire n8002;
wire n8003;
wire n8004;
wire n8005;
wire n8006;
wire n8007;
wire n8008;
wire n8009;
wire n8010;
wire n8011;
wire n8012;
wire n8013;
wire n8014;
wire n8015;
wire n8016;
wire n8017;
wire n8018;
wire n8019;
wire n8020;
wire n8021;
wire n8022;
wire n8023;
wire n8024;
wire n8025;
wire n8026;
wire n8027;
wire n8028;
wire n8029;
wire n8030;
wire n8031;
wire n8032;
wire n8033;
wire n8034;
wire n8035;
wire n8036;
wire n8037;
wire n8038;
wire n8039;
wire n8040;
wire n8041;
wire n8042;
wire n8043;
wire n8044;
wire n8045;
wire n8046;
wire n8047;
wire n8048;
wire n8049;
wire n8050;
wire n8051;
wire n8052;
wire n8053;
wire n8054;
wire n8055;
wire n8056;
wire n8057;
wire n8058;
wire n8059;
wire n8060;
wire n8061;
wire n8062;
wire n8063;
wire n8064;
wire n8065;
wire n8066;
wire n8067;
wire n8068;
wire n8069;
wire n8070;
wire n8071;
wire n8072;
wire n8073;
wire n8074;
wire n8075;
wire n8076;
wire n8077;
wire n8078;
wire n8079;
wire n8080;
wire n8081;
wire n8082;
wire n8083;
wire n8084;
wire n8085;
wire n8086;
wire n8087;
wire n8088;
wire n8089;
wire n8090;
wire n8091;
wire n8092;
wire n8093;
wire n8094;
wire n8095;
wire n8096;
wire n8097;
wire n8098;
wire n8099;
wire n8100;
wire n8101;
wire n8102;
wire n8103;
wire n8104;
wire n8105;
wire n8106;
wire n8107;
wire n8108;
wire n8109;
wire n8110;
wire n8111;
wire n8112;
wire n8113;
wire n8114;
wire n8115;
wire n8116;
wire n8117;
wire n8118;
wire n8119;
wire n8120;
wire n8121;
wire n8122;
wire n8123;
wire n8124;
wire n8125;
wire n8126;
wire n8127;
wire n8128;
wire n8129;
wire n8130;
wire n8131;
wire n8132;
wire n8133;
wire n8134;
wire n8135;
wire n8136;
wire n8137;
wire n8138;
wire n8139;
wire n8140;
wire n8141;
wire n8142;
wire n8143;
wire n8144;
wire n8145;
wire n8146;
wire n8147;
wire n8148;
wire n8149;
wire n8150;
wire n8151;
wire n8152;
wire n8153;
wire n8154;
wire n8155;
wire n8156;
wire n8157;
wire n8158;
wire n8159;
wire n8160;
wire n8161;
wire n8162;
wire n8163;
wire n8164;
wire n8165;
wire n8166;
wire n8167;
wire n8168;
wire n8169;
wire n8170;
wire n8171;
wire n8172;
wire n8173;
wire n8174;
wire n8175;
wire n8176;
wire n8177;
wire n8178;
wire n8179;
wire n8180;
wire n8181;
wire n8182;
wire n8183;
wire n8184;
wire n8185;
wire n8186;
wire n8187;
wire n8188;
wire n8189;
wire n8190;
wire n8191;
wire n8192;
wire n8193;
wire n8194;
wire n8195;
wire n8196;
wire n8197;
wire n8198;
wire n8199;
wire n8200;
wire n8201;
wire n8202;
wire n8203;
wire n8204;
wire n8205;
wire n8206;
wire n8207;
wire n8208;
wire n8209;
wire n8210;
wire n8211;
wire n8212;
wire n8213;
wire n8214;
wire n8215;
wire n8216;
wire n8217;
wire n8218;
wire n8219;
wire n8220;
wire n8221;
wire n8222;
wire n8223;
wire n8224;
wire n8225;
wire n8226;
wire n8227;
wire n8228;
wire n8229;
wire n8230;
wire n8231;
wire n8232;
wire n8233;
wire n8234;
wire n8235;
wire n8236;
wire n8237;
wire n8238;
wire n8239;
wire n8240;
wire n8241;
wire n8242;
wire n8243;
wire n8244;
wire n8245;
wire n8246;
wire n8247;
wire n8248;
wire n8249;
wire n8250;
wire n8251;
wire n8252;
wire n8253;
wire n8254;
wire n8255;
wire n8256;
wire n8257;
wire n8258;
wire n8259;
wire n8260;
wire n8261;
wire n8262;
wire n8263;
wire n8264;
wire n8265;
wire n8266;
wire n8267;
wire n8268;
wire n8269;
wire n8270;
wire n8271;
wire n8272;
wire n8273;
wire n8274;
wire n8275;
wire n8276;
wire n8277;
wire n8278;
wire n8279;
wire n8280;
wire n8281;
wire n8282;
wire n8283;
wire n8284;
wire n8285;
wire n8286;
wire n8287;
wire n8288;
wire n8289;
wire n8290;
wire n8291;
wire n8292;
wire n8293;
wire n8294;
wire n8295;
wire n8296;
wire n8297;
wire n8298;
wire n8299;
wire n8300;
wire n8301;
wire n8302;
wire n8303;
wire n8304;
wire n8305;
wire n8306;
wire n8307;
wire n8308;
wire n8309;
wire n8310;
wire n8311;
wire n8312;
wire n8313;
wire n8314;
wire n8315;
wire n8316;
wire n8317;
wire n8318;
wire n8319;
wire n8320;
wire n8321;
wire n8322;
wire n8323;
wire n8324;
wire n8325;
wire n8326;
wire n8327;
wire n8328;
wire n8329;
wire n8330;
wire n8331;
wire n8332;
wire n8333;
wire n8334;
wire n8335;
wire n8336;
wire n8337;
wire n8338;
wire n8339;
wire n8340;
wire n8341;
wire n8342;
wire n8343;
wire n8344;
wire n8345;
wire n8346;
wire n8347;
wire n8348;
wire n8349;
wire n8350;
wire n8351;
wire n8352;
wire n8353;
wire n8354;
wire n8355;
wire n8356;
wire n8357;
wire n8358;
wire n8359;
wire n8360;
wire n8361;
wire n8362;
wire n8363;
wire n8364;
wire n8365;
wire n8366;
wire n8367;
wire n8368;
wire n8369;
wire n8370;
wire n8371;
wire n8372;
wire n8373;
wire n8374;
wire n8375;
wire n8376;
wire n8377;
wire n8378;
wire n8379;
wire n8380;
wire n8381;
wire n8382;
wire n8383;
wire n8384;
wire n8385;
wire n8386;
wire n8387;
wire n8388;
wire n8389;
wire n8390;
wire n8391;
wire n8392;
wire n8393;
wire n8394;
wire n8395;
wire n8396;
wire n8397;
wire n8398;
wire n8399;
wire n8400;
wire n8401;
wire n8402;
wire n8403;
wire n8404;
wire n8405;
wire n8406;
wire n8407;
wire n8408;
wire n8409;
wire n8410;
wire n8411;
wire n8412;
wire n8413;
wire n8414;
wire n8415;
wire n8416;
wire n8417;
wire n8418;
wire n8419;
wire n8420;
wire n8421;
wire n8422;
wire n8423;
wire n8424;
wire n8425;
wire n8426;
wire n8427;
wire n8428;
wire n8429;
wire n8430;
wire n8431;
wire n8432;
wire n8433;
wire n8434;
wire n8435;
wire n8436;
wire n8437;
wire n8438;
wire n8439;
wire n8440;
wire n8441;
wire n8442;
wire n8443;
wire n8444;
wire n8445;
wire n8446;
wire n8447;
wire n8448;
wire n8449;
wire n8450;
wire n8451;
wire n8452;
wire n8453;
wire n8454;
wire n8455;
wire n8456;
wire n8457;
wire n8458;
wire n8459;
wire n8460;
wire n8461;
wire n8462;
wire n8463;
wire n8464;
wire n8465;
wire n8466;
wire n8467;
wire n8468;
wire n8469;
wire n8470;
wire n8471;
wire n8472;
wire n8473;
wire n8474;
wire n8475;
wire n8476;
wire n8477;
wire n8478;
wire n8479;
wire n8480;
wire n8481;
wire n8482;
wire n8483;
wire n8484;
wire n8485;
wire n8486;
wire n8487;
wire n8488;
wire n8489;
wire n8490;
wire n8491;
wire n8492;
wire n8493;
wire n8494;
wire n8495;
wire n8496;
wire n8497;
wire n8498;
wire n8499;
wire n8500;
wire n8501;
wire n8502;
wire n8503;
wire n8504;
wire n8505;
wire n8506;
wire n8507;
wire n8508;
wire n8509;
wire n8510;
wire n8511;
wire n8512;
wire n8513;
wire n8514;
wire n8515;
wire n8516;
wire n8517;
wire n8518;
wire n8519;
wire n8520;
wire n8521;
wire n8522;
wire n8523;
wire n8524;
wire n8525;
wire n8526;
wire n8527;
wire n8528;
wire n8529;
wire n8530;
wire n8531;
wire n8532;
wire n8533;
wire n8534;
wire n8535;
wire n8536;
wire n8537;
wire n8538;
wire n8539;
wire n8540;
wire n8541;
wire n8542;
wire n8543;
wire n8544;
wire n8545;
wire n8546;
wire n8547;
wire n8548;
wire n8549;
wire n8550;
wire n8551;
wire n8552;
wire n8553;
wire n8554;
wire n8555;
wire n8556;
wire n8557;
wire n8558;
wire n8559;
wire n8560;
wire n8561;
wire n8562;
wire n8563;
wire n8564;
wire n8565;
wire n8566;
wire n8567;
wire n8568;
wire n8569;
wire n8570;
wire n8571;
wire n8572;
wire n8573;
wire n8574;
wire n8575;
wire n8576;
wire n8577;
wire n8578;
wire n8579;
wire n8580;
wire n8581;
wire n8582;
wire n8583;
wire n8584;
wire n8585;
wire n8586;
wire n8587;
wire n8588;
wire n8589;
wire n8590;
wire n8591;
wire n8592;
wire n8593;
wire n8594;
wire n8595;
wire n8596;
wire n8597;
wire n8598;
wire n8599;
wire n8600;
wire n8601;
wire n8602;
wire n8603;
wire n8604;
wire n8605;
wire n8606;
wire n8607;
wire n8608;
wire n8609;
wire n8610;
wire n8611;
wire n8612;
wire n8613;
wire n8614;
wire n8615;
wire n8616;
wire n8617;
wire n8618;
wire n8619;
wire n8620;
wire n8621;
wire n8622;
wire n8623;
wire n8624;
wire n8625;
wire n8626;
wire n8627;
wire n8628;
wire n8629;
wire n8630;
wire n8631;
wire n8632;
wire n8633;
wire n8634;
wire n8635;
wire n8636;
wire n8637;
wire n8638;
wire n8639;
wire n8640;
wire n8641;
wire n8642;
wire n8643;
wire n8644;
wire n8645;
wire n8646;
wire n8647;
wire n8648;
wire n8649;
wire n8650;
wire n8651;
wire n8652;
wire n8653;
wire n8654;
wire n8655;
wire n8656;
wire n8657;
wire n8658;
wire n8659;
wire n8660;
wire n8661;
wire n8662;
wire n8663;
wire n8664;
wire n8665;
wire n8666;
wire n8667;
wire n8668;
wire n8669;
wire n8670;
wire n8671;
wire n8672;
wire n8673;
wire n8674;
wire n8675;
wire n8676;
wire n8677;
wire n8678;
wire n8679;
wire n8680;
wire n8681;
wire n8682;
wire n8683;
wire n8684;
wire n8685;
wire n8686;
wire n8687;
wire n8688;
wire n8689;
wire n8690;
wire n8691;
wire n8692;
wire n8693;
wire n8694;
wire n8695;
wire n8696;
wire n8697;
wire n8698;
wire n8699;
wire n8700;
wire n8701;
wire n8702;
wire n8703;
wire n8704;
wire n8705;
wire n8706;
wire n8707;
wire n8708;
wire n8709;
wire n8710;
wire n8711;
wire n8712;
wire n8713;
wire n8714;
wire n8715;
wire n8716;
wire n8717;
wire n8718;
wire n8719;
wire n8720;
wire n8721;
wire n8722;
wire n8723;
wire n8724;
wire n8725;
wire n8726;
wire n8727;
wire n8728;
wire n8729;
wire n8730;
wire n8731;
wire n8732;
wire n8733;
wire n8734;
wire n8735;
wire n8736;
wire n8737;
wire n8738;
wire n8739;
wire n8740;
wire n8741;
wire n8742;
wire n8743;
wire n8744;
wire n8745;
wire n8746;
wire n8747;
wire n8748;
wire n8749;
wire n8750;
wire n8751;
wire n8752;
wire n8753;
wire n8754;
wire n8755;
wire n8756;
wire n8757;
wire n8758;
wire n8759;
wire n8760;
wire n8761;
wire n8762;
wire n8763;
wire n8764;
wire n8765;
wire n8766;
wire n8767;
wire n8768;
wire n8769;
wire n8770;
wire n8771;
wire n8772;
wire n8773;
wire n8774;
wire n8775;
wire n8776;
wire n8777;
wire n8778;
wire n8779;
wire n8780;
wire n8781;
wire n8782;
wire n8783;
wire n8784;
wire n8785;
wire n8786;
wire n8787;
wire n8788;
wire n8789;
wire n8790;
wire n8791;
wire n8792;
wire n8793;
wire n8794;
wire n8795;
wire n8796;
wire n8797;
wire n8798;
wire n8799;
wire n8800;
wire n8801;
wire n8802;
wire n8803;
wire n8804;
wire n8805;
wire n8806;
wire n8807;
wire n8808;
wire n8809;
wire n8810;
wire n8811;
wire n8812;
wire n8813;
wire n8814;
wire n8815;
wire n8816;
wire n8817;
wire n8818;
wire n8819;
wire n8820;
wire n8821;
wire n8822;
wire n8823;
wire n8824;
wire n8825;
wire n8826;
wire n8827;
wire n8828;
wire n8829;
wire n8830;
wire n8831;
wire n8832;
wire n8833;
wire n8834;
wire n8835;
wire n8836;
wire n8837;
wire n8838;
wire n8839;
wire n8840;
wire n8841;
wire n8842;
wire n8843;
wire n8844;
wire n8845;
wire n8846;
wire n8847;
wire n8848;
wire n8849;
wire n8850;
wire n8851;
wire n8852;
wire n8853;
wire n8854;
wire n8855;
wire n8856;
wire n8857;
wire n8858;
wire n8859;
wire n8860;
wire n8861;
wire n8862;
wire n8863;
wire n8864;
wire n8865;
wire n8866;
wire n8867;
wire n8868;
wire n8869;
wire n8870;
wire n8871;
wire n8872;
wire n8873;
wire n8874;
wire n8875;
wire n8876;
wire n8877;
wire n8878;
wire n8879;
wire n8880;
wire n8881;
wire n8882;
wire n8883;
wire n8884;
wire n8885;
wire n8886;
wire n8887;
wire n8888;
wire n8889;
wire n8890;
wire n8891;
wire n8892;
wire n8893;
wire n8894;
wire n8895;
wire n8896;
wire n8897;
wire n8898;
wire n8899;
wire n8900;
wire n8901;
wire n8902;
wire n8903;
wire n8904;
wire n8905;
wire n8906;
wire n8907;
wire n8908;
wire n8909;
wire n8910;
wire n8911;
wire n8912;
wire n8913;
wire n8914;
wire n8915;
wire n8916;
wire n8917;
wire n8918;
wire n8919;
wire n8920;
wire n8921;
wire n8922;
wire n8923;
wire n8924;
wire n8925;
wire n8926;
wire n8927;
wire n8928;
wire n8929;
wire n8930;
wire n8931;
wire n8932;
wire n8933;
wire n8934;
wire n8935;
wire n8936;
wire n8937;
wire n8938;
wire n8939;
wire n8940;
wire n8941;
wire n8942;
wire n8943;
wire n8944;
wire n8945;
wire n8946;
wire n8947;
wire n8948;
wire n8949;
wire n8950;
wire n8951;
wire n8952;
wire n8953;
wire n8954;
wire n8955;
wire n8956;
wire n8957;
wire n8958;
wire n8959;
wire n8960;
wire n8961;
wire n8962;
wire n8963;
wire n8964;
wire n8965;
wire n8966;
wire n8967;
wire n8968;
wire n8969;
wire n8970;
wire n8971;
wire n8972;
wire n8973;
wire n8974;
wire n8975;
wire n8976;
wire n8977;
wire n8978;
wire n8979;
wire n8980;
wire n8981;
wire n8982;
wire n8983;
wire n8984;
wire n8985;
wire n8986;
wire n8987;
wire n8988;
wire n8989;
wire n8990;
wire n8991;
wire n8992;
wire n8993;
wire n8994;
wire n8995;
wire n8996;
wire n8997;
wire n8998;
wire n8999;
wire n9000;
wire n9001;
wire n9002;
wire n9003;
wire n9004;
wire n9005;
wire n9006;
wire n9007;
wire n9008;
wire n9009;
wire n9010;
wire n9011;
wire n9012;
wire n9013;
wire n9014;
wire n9015;
wire n9016;
wire n9017;
wire n9018;
wire n9019;
wire n9020;
wire n9021;
wire n9022;
wire n9023;
wire n9024;
wire n9025;
wire n9026;
wire n9027;
wire n9028;
wire n9029;
wire n9030;
wire n9031;
wire n9032;
wire n9033;
wire n9034;
wire n9035;
wire n9036;
wire n9037;
wire n9038;
wire n9039;
wire n9040;
wire n9041;
wire n9042;
wire n9043;
wire n9044;
wire n9045;
wire n9046;
wire n9047;
wire n9048;
wire n9049;
wire n9050;
wire n9051;
wire n9052;
wire n9053;
wire n9054;
wire n9055;
wire n9056;
wire n9057;
wire n9058;
wire n9059;
wire n9060;
wire n9061;
wire n9062;
wire n9063;
wire n9064;
wire n9065;
wire n9066;
wire n9067;
wire n9068;
wire n9069;
wire n9070;
wire n9071;
wire n9072;
wire n9073;
wire n9074;
wire n9075;
wire n9076;
wire n9077;
wire n9078;
wire n9079;
wire n9080;
wire n9081;
wire n9082;
wire n9083;
wire n9084;
wire n9085;
wire n9086;
wire n9087;
wire n9088;
wire n9089;
wire n9090;
wire n9091;
wire n9092;
wire n9093;
wire n9094;
wire n9095;
wire n9096;
wire n9097;
wire n9098;
wire n9099;
wire n9100;
wire n9101;
wire n9102;
wire n9103;
wire n9104;
wire n9105;
wire n9106;
wire n9107;
wire n9108;
wire n9109;
wire n9110;
wire n9111;
wire n9112;
wire n9113;
wire n9114;
wire n9115;
wire n9116;
wire n9117;
wire n9118;
wire n9119;
wire n9120;
wire n9121;
wire n9122;
wire n9123;
wire n9124;
wire n9125;
wire n9126;
wire n9127;
wire n9128;
wire n9129;
wire n9130;
wire n9131;
wire n9132;
wire n9133;
wire n9134;
wire n9135;
wire n9136;
wire n9137;
wire n9138;
wire n9139;
wire n9140;
wire n9141;
wire n9142;
wire n9143;
wire n9144;
wire n9145;
wire n9146;
wire n9147;
wire n9148;
wire n9149;
wire n9150;
wire n9151;
wire n9152;
wire n9153;
wire n9154;
wire n9155;
wire n9156;
wire n9157;
wire n9158;
wire n9159;
wire n9160;
wire n9161;
wire n9162;
wire n9163;
wire n9164;
wire n9165;
wire n9166;
wire n9167;
wire n9168;
wire n9169;
wire n9170;
wire n9171;
wire n9172;
wire n9173;
wire n9174;
wire n9175;
wire n9176;
wire n9177;
wire n9178;
wire n9179;
wire n9180;
wire n9181;
wire n9182;
wire n9183;
wire n9184;
wire n9185;
wire n9186;
wire n9187;
wire n9188;
wire n9189;
wire n9190;
wire n9191;
wire n9192;
wire n9193;
wire n9194;
wire n9195;
wire n9196;
wire n9197;
wire n9198;
wire n9199;
wire n9200;
wire n9201;
wire n9202;
wire n9203;
wire n9204;
wire n9205;
wire n9206;
wire n9207;
wire n9208;
wire n9209;
wire n9210;
wire n9211;
wire n9212;
wire n9213;
wire n9214;
wire n9215;
wire n9216;
wire n9217;
wire n9218;
wire n9219;
wire n9220;
wire n9221;
wire n9222;
wire n9223;
wire n9224;
wire n9225;
wire n9226;
wire n9227;
wire n9228;
wire n9229;
wire n9230;
wire n9231;
wire n9232;
wire n9233;
wire n9234;
wire n9235;
wire n9236;
wire n9237;
wire n9238;
wire n9239;
wire n9240;
wire n9241;
wire n9242;
wire n9243;
wire n9244;
wire n9245;
wire n9246;
wire n9247;
wire n9248;
wire n9249;
wire n9250;
wire n9251;
wire n9252;
wire n9253;
wire n9254;
wire n9255;
wire n9256;
wire n9257;
wire n9258;
wire n9259;
wire n9260;
wire n9261;
wire n9262;
wire n9263;
wire n9264;
wire n9265;
wire n9266;
wire n9267;
wire n9268;
wire n9269;
wire n9270;
wire n9271;
wire n9272;
wire n9273;
wire n9274;
wire n9275;
wire n9276;
wire n9277;
wire n9278;
wire n9279;
wire n9280;
wire n9281;
wire n9282;
wire n9283;
wire n9284;
wire n9285;
wire n9286;
wire n9287;
wire n9288;
wire n9289;
wire n9290;
wire n9291;
wire n9292;
wire n9293;
wire n9294;
wire n9295;
wire n9296;
wire n9297;
wire n9298;
wire n9299;
wire n9300;
wire n9301;
wire n9302;
wire n9303;
wire n9304;
wire n9305;
wire n9306;
wire n9307;
wire n9308;
wire n9309;
wire n9310;
wire n9311;
wire n9312;
wire n9313;
wire n9314;
wire n9315;
wire n9316;
wire n9317;
wire n9318;
wire n9319;
wire n9320;
wire n9321;
wire n9322;
wire n9323;
wire n9324;
wire n9325;
wire n9326;
wire n9327;
wire n9328;
wire n9329;
wire n9330;
wire n9331;
wire n9332;
wire n9333;
wire n9334;
wire n9335;
wire n9336;
wire n9337;
wire n9338;
wire n9339;
wire n9340;
wire n9341;
wire n9342;
wire n9343;
wire n9344;
wire n9345;
wire n9346;
wire n9347;
wire n9348;
wire n9349;
wire n9350;
wire n9351;
wire n9352;
wire n9353;
wire n9354;
wire n9355;
wire n9356;
wire n9357;
wire n9358;
wire n9359;
wire n9360;
wire n9361;
wire n9362;
wire n9363;
wire n9364;
wire n9365;
wire n9366;
wire n9367;
wire n9368;
wire n9369;
wire n9370;
wire n9371;
wire n9372;
wire n9373;
wire n9374;
wire n9375;
wire n9376;
wire n9377;
wire n9378;
wire n9379;
wire n9380;
wire n9381;
wire n9382;
wire n9383;
wire n9384;
wire n9385;
wire n9386;
wire n9387;
wire n9388;
wire n9389;
wire n9390;
wire n9391;
wire n9392;
wire n9393;
wire n9394;
wire n9395;
wire n9396;
wire n9397;
wire n9398;
wire n9399;
wire n9400;
wire n9401;
wire n9402;
wire n9403;
wire n9404;
wire n9405;
wire n9406;
wire n9407;
wire n9408;
wire n9409;
wire n9410;
wire n9411;
wire n9412;
wire n9413;
wire n9414;
wire n9415;
wire n9416;
wire n9417;
wire n9418;
wire n9419;
wire n9420;
wire n9421;
wire n9422;
wire n9423;
wire n9424;
wire n9425;
wire n9426;
wire n9427;
wire n9428;
wire n9429;
wire n9430;
wire n9431;
wire n9432;
wire n9433;
wire n9434;
wire n9435;
wire n9436;
wire n9437;
wire n9438;
wire n9439;
wire n9440;
wire n9441;
wire n9442;
wire n9443;
wire n9444;
wire n9445;
wire n9446;
wire n9447;
wire n9448;
wire n9449;
wire n9450;
wire n9451;
wire n9452;
wire n9453;
wire n9454;
wire n9455;
wire n9456;
wire n9457;
wire n9458;
wire n9459;
wire n9460;
wire n9461;
wire n9462;
wire n9463;
wire n9464;
wire n9465;
wire n9466;
wire n9467;
wire n9468;
wire n9469;
wire n9470;
wire n9471;
wire n9472;
wire n9473;
wire n9474;
wire n9475;
wire n9476;
wire n9477;
wire n9478;
wire n9479;
wire n9480;
wire n9481;
wire n9482;
wire n9483;
wire n9484;
wire n9485;
wire n9486;
wire n9487;
wire n9488;
wire n9489;
wire n9490;
wire n9491;
wire n9492;
wire n9493;
wire n9494;
wire n9495;
wire n9496;
wire n9497;
wire n9498;
wire n9499;
wire n9500;
wire n9501;
wire n9502;
wire n9503;
wire n9504;
wire n9505;
wire n9506;
wire n9507;
wire n9508;
wire n9509;
wire n9510;
wire n9511;
wire n9512;
wire n9513;
wire n9514;
xor (out,n0,n8769);
nand (n0,n1,n6828);
not (n1,n2);
or (n2,1'b0,n4,n6815,n6825,n6826,n6827);
and (n4,n5,n904);
wire s0n5,s1n5,notn5;
or (n5,s0n5,s1n5);
not(notn5,n896);
and (s0n5,notn5,1'b0);
and (s1n5,n896,n6);
xor (n6,n7,n6793);
or (n7,n8,n6019,n6792);
and (n8,n9,n3058);
or (n9,1'b0,n10,n893,n907,n2974);
and (n10,n11,n22);
wire s0n11,s1n11,notn11;
or (n11,s0n11,s1n11);
not(notn11,n13);
and (s0n11,notn11,1'b0);
and (s1n11,n13,n12);
and (n13,n14,n21);
nand (n14,n15,n16,n18,n19);
not (n16,n17);
not (n19,n20);
or (n21,n15,n17,n18,n20);
or (n22,n23,n891);
nor (n23,n24,n671,n744,n817);
not (n24,n25);
wire s0n25,s1n25,notn25;
or (n25,s0n25,s1n25);
not(notn25,n594);
and (s0n25,notn25,1'b0);
and (s1n25,n594,n26);
wire s0n26,s1n26,notn26;
or (n26,s0n26,s1n26);
not(notn26,n594);
and (s0n26,notn26,n27);
and (s1n26,n594,n630);
wire s0n27,s1n27,notn27;
or (n27,s0n27,s1n27);
not(notn27,n66);
and (s0n27,notn27,1'b0);
and (s1n27,n66,n28);
wire s0n28,s1n28,notn28;
or (n28,s0n28,s1n28);
not(notn28,n629);
and (s0n28,notn28,n29);
and (s1n28,n629,n620);
or (n29,n30,n596,n607,n618);
and (n30,n31,n53);
wire s0n31,s1n31,notn31;
or (n31,s0n31,s1n31);
not(notn31,n48);
and (s0n31,notn31,n32);
and (s1n31,n48,n33);
or (n33,n34,n39,n43,n46);
and (n34,n35,n36);
nor (n36,n37,n38);
and (n39,n40,n41);
nor (n41,n42,n38);
not (n42,n37);
and (n43,n44,n45);
and (n45,n42,n38);
and (n46,n32,n47);
and (n47,n37,n38);
wire s0n48,s1n48,notn48;
or (n48,s0n48,s1n48);
not(notn48,n594);
and (s0n48,notn48,n49);
and (s1n48,n594,n582);
and (n49,n50,n66);
or (n50,n51,n56,n60,n63);
and (n51,n52,n53);
and (n53,n54,n55);
and (n56,n57,n58);
and (n58,n59,n55);
not (n59,n54);
and (n60,n61,n62);
nor (n62,n59,n55);
and (n63,n64,n65);
nor (n65,n54,n55);
and (n66,n67,n581);
not (n67,n68);
wire s0n68,s1n68,notn68;
or (n68,s0n68,s1n68);
not(notn68,n580);
and (s0n68,notn68,n69);
and (s1n68,n580,1'b0);
wire s0n69,s1n69,notn69;
or (n69,s0n69,s1n69);
not(notn69,n210);
and (s0n69,notn69,n70);
and (s1n69,n210,n71);
wire s0n71,s1n71,notn71;
or (n71,s0n71,s1n71);
not(notn71,n573);
and (s0n71,notn71,n72);
and (s1n71,n573,n547);
or (n72,n73,n515,n546,1'b0,1'b0,1'b0,1'b0,1'b0);
or (n73,n74,n514);
or (n74,n75,n513);
or (n75,n76,n512);
or (n76,n77,n510);
or (n77,n78,n509);
or (n78,n79,n507);
or (n79,n80,n505);
nor (n80,n81,n430,n439,n451,n463,n474,n485,n496);
or (n81,1'b0,n82,n424,n428);
and (n82,n83,n423);
wire s0n83,s1n83,notn83;
or (n83,s0n83,s1n83);
not(notn83,n414);
and (s0n83,notn83,n84);
and (s1n83,n414,n322);
wire s0n84,s1n84,notn84;
or (n84,s0n84,s1n84);
not(notn84,n281);
and (s0n84,notn84,1'b0);
and (s1n84,n281,n85);
or (n85,n86,n262,n266,n270,n273,n276,n278,1'b0);
and (n86,n87,n89);
not (n87,n88);
and (n89,n90,n235,n246,n256);
wire s0n90,s1n90,notn90;
or (n90,s0n90,s1n90);
not(notn90,n124);
and (s0n90,notn90,n91);
and (s1n90,n124,1'b0);
wire s0n91,s1n91,notn91;
or (n91,s0n91,s1n91);
not(notn91,n122);
and (s0n91,notn91,n92);
and (s1n91,n122,n120);
wire s0n92,s1n92,notn92;
or (n92,s0n92,s1n92);
not(notn92,n116);
and (s0n92,notn92,n93);
and (s1n92,n116,n110);
wire s0n93,s1n93,notn93;
or (n93,s0n93,s1n93);
not(notn93,n109);
and (s0n93,notn93,n94);
and (s1n93,n109,1'b0);
wire s0n94,s1n94,notn94;
or (n94,s0n94,s1n94);
not(notn94,n108);
and (s0n94,notn94,n95);
and (s1n94,n108,1'b1);
wire s0n95,s1n95,notn95;
or (n95,s0n95,s1n95);
not(notn95,n107);
and (s0n95,notn95,n96);
and (s1n95,n107,1'b0);
wire s0n96,s1n96,notn96;
or (n96,s0n96,s1n96);
not(notn96,n106);
and (s0n96,notn96,n97);
and (s1n96,n106,1'b1);
wire s0n97,s1n97,notn97;
or (n97,s0n97,s1n97);
not(notn97,n105);
and (s0n97,notn97,n98);
and (s1n97,n105,1'b0);
wire s0n98,s1n98,notn98;
or (n98,s0n98,s1n98);
not(notn98,n104);
and (s0n98,notn98,n99);
and (s1n98,n104,1'b1);
wire s0n99,s1n99,notn99;
or (n99,s0n99,s1n99);
not(notn99,n103);
and (s0n99,notn99,n100);
and (s1n99,n103,1'b0);
wire s0n100,s1n100,notn100;
or (n100,s0n100,s1n100);
not(notn100,n102);
and (s0n100,notn100,n87);
and (s1n100,n102,1'b1);
wire s0n110,s1n110,notn110;
or (n110,s0n110,s1n110);
not(notn110,n115);
and (s0n110,notn110,n111);
and (s1n110,n115,1'b0);
wire s0n111,s1n111,notn111;
or (n111,s0n111,s1n111);
not(notn111,n114);
and (s0n111,notn111,n112);
and (s1n111,n114,1'b1);
not (n112,n113);
or (n116,n117,n119);
or (n117,n118,n113);
or (n118,n115,n114);
not (n120,n121);
or (n122,n121,n123);
not (n124,n125);
or (n125,n126,n233);
or (n126,n127,n231);
or (n127,n128,n225);
or (n128,n129,n224);
or (n129,n130,n220);
or (n130,n131,n219);
or (n131,n132,n214);
or (n132,n133,n213);
or (n133,n134,n212);
or (n134,n135,n210);
or (n135,n136,n204);
or (n136,n137,n203);
or (n137,n138,n202);
or (n138,n139,n201);
or (n139,n140,n200);
or (n140,n141,n199);
or (n141,n142,n198);
or (n142,n143,n197);
or (n143,n144,n194);
or (n144,n145,n188);
or (n145,n146,n187);
or (n146,n147,n186);
or (n147,n148,n185);
or (n148,n149,n184);
or (n149,n150,n183);
or (n150,n151,n181);
or (n151,n152,n179);
or (n152,n153,n173);
or (n153,n154,n172);
or (n154,n155,n171);
or (n155,n156,n170);
or (n156,n157,n169);
or (n157,n158,n167);
or (n158,n159,n165);
nor (n159,n160,n161,n163,n164);
not (n161,n162);
nor (n165,n160,n161,n166,n164);
not (n166,n163);
and (n167,n160,n162,n163,n168);
not (n168,n164);
and (n169,n160,n161,n163,n168);
nor (n170,n160,n162,n166,n164);
and (n171,n160,n161,n163,n164);
and (n172,n160,n162,n163,n164);
nor (n173,n174,n176,n177,n178);
not (n174,n175);
nor (n179,n174,n180,n177,n178);
not (n180,n176);
and (n181,n174,n176,n177,n182);
not (n182,n178);
and (n183,n175,n176,n177,n182);
and (n184,n175,n180,n177,n182);
and (n185,n174,n180,n177,n178);
and (n186,n175,n180,n177,n178);
and (n187,n175,n176,n177,n178);
nor (n188,n189,n191,n192,n193);
not (n189,n190);
and (n194,n190,n191,n195,n196);
not (n195,n192);
not (n196,n193);
and (n197,n189,n191,n195,n196);
and (n198,n190,n191,n192,n196);
nor (n199,n190,n191,n195,n196);
and (n200,n189,n191,n192,n193);
and (n201,n189,n191,n195,n193);
and (n202,n190,n191,n195,n193);
nor (n203,n189,n191,n192,n196);
nor (n204,n205,n207,n208,n209);
not (n205,n206);
nor (n210,n206,n211,n208,n209);
not (n211,n207);
and (n212,n205,n211,n208,n209);
and (n213,n206,n211,n208,n209);
nor (n214,n215,n216,n218);
not (n216,n217);
and (n219,n215,n217,n218);
and (n220,n221,n222);
not (n222,n223);
nor (n224,n221,n222);
nor (n225,n226,n227,n229,n230);
not (n227,n228);
and (n231,n226,n228,n229,n232);
not (n232,n230);
and (n233,n234,n227,n229,n232);
not (n234,n226);
wire s0n235,s1n235,notn235;
or (n235,s0n235,s1n235);
not(notn235,n124);
and (s0n235,notn235,n236);
and (s1n235,n124,1'b0);
wire s0n236,s1n236,notn236;
or (n236,s0n236,s1n236);
not(notn236,n122);
and (s0n236,notn236,n237);
and (s1n236,n122,1'b0);
wire s0n237,s1n237,notn237;
or (n237,s0n237,s1n237);
not(notn237,n116);
and (s0n237,notn237,n238);
and (s1n237,n116,n118);
wire s0n238,s1n238,notn238;
or (n238,s0n238,s1n238);
not(notn238,n109);
and (s0n238,notn238,n239);
and (s1n238,n109,1'b1);
wire s0n239,s1n239,notn239;
or (n239,s0n239,s1n239);
not(notn239,n108);
and (s0n239,notn239,n240);
and (s1n239,n108,1'b1);
wire s0n240,s1n240,notn240;
or (n240,s0n240,s1n240);
not(notn240,n107);
and (s0n240,notn240,n241);
and (s1n240,n107,1'b0);
wire s0n241,s1n241,notn241;
or (n241,s0n241,s1n241);
not(notn241,n106);
and (s0n241,notn241,n242);
and (s1n241,n106,1'b0);
wire s0n242,s1n242,notn242;
or (n242,s0n242,s1n242);
not(notn242,n105);
and (s0n242,notn242,n243);
and (s1n242,n105,1'b1);
wire s0n243,s1n243,notn243;
or (n243,s0n243,s1n243);
not(notn243,n104);
and (s0n243,notn243,n244);
and (s1n243,n104,1'b1);
wire s0n244,s1n244,notn244;
or (n244,s0n244,s1n244);
not(notn244,n103);
and (s0n244,notn244,n245);
and (s1n244,n103,1'b0);
not (n245,n102);
wire s0n246,s1n246,notn246;
or (n246,s0n246,s1n246);
not(notn246,n124);
and (s0n246,notn246,n247);
and (s1n246,n124,1'b0);
wire s0n247,s1n247,notn247;
or (n247,s0n247,s1n247);
not(notn247,n122);
and (s0n247,notn247,n248);
and (s1n247,n122,1'b0);
wire s0n248,s1n248,notn248;
or (n248,s0n248,s1n248);
not(notn248,n116);
and (s0n248,notn248,n249);
and (s1n248,n116,n255);
wire s0n249,s1n249,notn249;
or (n249,s0n249,s1n249);
not(notn249,n109);
and (s0n249,notn249,n250);
and (s1n249,n109,1'b1);
wire s0n250,s1n250,notn250;
or (n250,s0n250,s1n250);
not(notn250,n108);
and (s0n250,notn250,n251);
and (s1n250,n108,1'b1);
wire s0n251,s1n251,notn251;
or (n251,s0n251,s1n251);
not(notn251,n107);
and (s0n251,notn251,n252);
and (s1n251,n107,1'b0);
wire s0n252,s1n252,notn252;
or (n252,s0n252,s1n252);
not(notn252,n106);
and (s0n252,notn252,n253);
and (s1n252,n106,1'b0);
wire s0n253,s1n253,notn253;
or (n253,s0n253,s1n253);
not(notn253,n105);
and (s0n253,notn253,n254);
and (s1n253,n105,1'b0);
not (n254,n104);
not (n255,n118);
not (n256,n257);
wire s0n257,s1n257,notn257;
or (n257,s0n257,s1n257);
not(notn257,n124);
and (s0n257,notn257,n258);
and (s1n257,n124,1'b0);
wire s0n258,s1n258,notn258;
or (n258,s0n258,s1n258);
not(notn258,n122);
and (s0n258,notn258,n259);
and (s1n258,n122,1'b0);
wire s0n259,s1n259,notn259;
or (n259,s0n259,s1n259);
not(notn259,n116);
and (s0n259,notn259,n260);
and (s1n259,n116,1'b0);
wire s0n260,s1n260,notn260;
or (n260,s0n260,s1n260);
not(notn260,n109);
and (s0n260,notn260,n261);
and (s1n260,n109,1'b0);
not (n261,n108);
and (n262,n263,n264);
not (n263,n103);
and (n264,n265,n235,n246,n256);
not (n265,n90);
and (n266,n267,n268);
not (n267,n105);
and (n268,n90,n269,n246,n256);
not (n269,n235);
and (n270,n271,n272);
not (n271,n107);
and (n272,n265,n269,n246,n256);
and (n273,n274,n275);
not (n274,n109);
nor (n275,n265,n269,n246,n257);
and (n276,n112,n277);
nor (n277,n90,n269,n246,n257);
and (n278,n279,n280);
not (n279,n115);
nor (n280,n265,n235,n246,n257);
or (n281,n282,n311);
wire s0n282,s1n282,notn282;
or (n282,s0n282,s1n282);
not(notn282,n309);
and (s0n282,notn282,n283);
and (s1n282,n309,1'b0);
wire s0n283,s1n283,notn283;
or (n283,s0n283,s1n283);
not(notn283,n308);
and (s0n283,notn283,n284);
and (s1n283,n308,n303);
wire s0n284,s1n284,notn284;
or (n284,s0n284,s1n284);
not(notn284,n302);
and (s0n284,notn284,n285);
and (s1n284,n302,n291);
wire s0n285,s1n285,notn285;
or (n285,s0n285,s1n285);
not(notn285,n290);
and (s0n285,notn285,n286);
and (s1n285,n290,n153);
or (n286,n287,n184);
or (n287,n288,n183);
or (n288,n289,n181);
or (n289,n173,n179);
or (n290,n160,n162,n163,n164);
or (n291,1'b0,1'b0,n292,n298,n300);
and (n292,n293,n296);
or (n293,1'b0,1'b0,n294,n214);
and (n294,n295,n217,n218);
not (n295,n215);
and (n296,n205,n211,n208,n297);
not (n297,n209);
and (n298,n221,n299);
and (n299,n206,n211,n208,n297);
or (n300,n301,n212);
or (n301,n204,n210);
or (n302,n206,n207,n208,n209);
or (n303,n304,n203);
or (n304,n305,n201);
or (n305,n306,n198);
or (n306,n307,n197);
or (n307,n188,n194);
or (n308,n190,n191,n192,n193);
not (n309,n310);
wire s0n311,s1n311,notn311;
or (n311,s0n311,s1n311);
not(notn311,n309);
and (s0n311,notn311,n312);
and (s1n311,n309,1'b0);
wire s0n312,s1n312,notn312;
or (n312,s0n312,s1n312);
not(notn312,n308);
and (s0n312,notn312,n313);
and (s1n312,n308,n321);
wire s0n313,s1n313,notn313;
or (n313,s0n313,s1n313);
not(notn313,n302);
and (s0n313,notn313,n314);
and (s1n313,n302,n317);
wire s0n314,s1n314,notn314;
or (n314,s0n314,s1n314);
not(notn314,n290);
and (s0n314,notn314,n315);
and (s1n314,n290,1'b0);
or (n315,n316,n187);
or (n316,n185,n186);
or (n317,1'b0,n213,n318,n320,1'b0);
and (n318,n319,n296);
or (n319,1'b0,n219,n294,1'b0);
and (n320,n223,n299);
or (n321,n200,n202);
not (n322,n323);
nor (n323,n84,n324,n340,n360,n377,n391,n402,n410);
wire s0n324,s1n324,notn324;
or (n324,s0n324,s1n324);
not(notn324,n281);
and (s0n324,notn324,1'b0);
and (s1n324,n281,n325);
or (n325,n326,n328,n330,n332,n334,n336,n338,1'b0);
and (n326,n327,n89);
xnor (n327,n102,n88);
and (n328,n329,n264);
xnor (n329,n104,n103);
and (n330,n331,n268);
xnor (n331,n106,n105);
and (n332,n333,n272);
xnor (n333,n108,n107);
and (n334,n335,n275);
xnor (n335,n119,n109);
and (n336,n337,n277);
xnor (n337,n114,n113);
and (n338,n339,n280);
xnor (n339,n123,n115);
wire s0n340,s1n340,notn340;
or (n340,s0n340,s1n340);
not(notn340,n281);
and (s0n340,notn340,1'b0);
and (s1n340,n281,n341);
or (n341,n342,n345,n348,n351,n354,n357,1'b0,1'b0);
and (n342,n343,n89);
xnor (n343,n103,n344);
or (n344,n102,n88);
and (n345,n346,n264);
xnor (n346,n105,n347);
or (n347,n104,n103);
and (n348,n349,n268);
xnor (n349,n107,n350);
or (n350,n106,n105);
and (n351,n352,n272);
xnor (n352,n109,n353);
or (n353,n108,n107);
and (n354,n355,n275);
xnor (n355,n113,n356);
or (n356,n119,n109);
and (n357,n358,n277);
xnor (n358,n115,n359);
or (n359,n114,n113);
wire s0n360,s1n360,notn360;
or (n360,s0n360,s1n360);
not(notn360,n281);
and (s0n360,notn360,1'b0);
and (s1n360,n281,n361);
or (n361,n362,n365,n368,n371,n374,1'b0,1'b0,1'b0);
and (n362,n363,n89);
xnor (n363,n104,n364);
or (n364,n103,n344);
and (n365,n366,n264);
xnor (n366,n106,n367);
or (n367,n105,n347);
and (n368,n369,n268);
xnor (n369,n108,n370);
or (n370,n107,n350);
and (n371,n372,n272);
xnor (n372,n119,n373);
or (n373,n109,n353);
and (n374,n375,n275);
xnor (n375,n114,n376);
or (n376,n113,n356);
wire s0n377,s1n377,notn377;
or (n377,s0n377,s1n377);
not(notn377,n281);
and (s0n377,notn377,1'b0);
and (s1n377,n281,n378);
or (n378,n379,n382,n385,n388,1'b0,1'b0,1'b0,1'b0);
and (n379,n380,n89);
xnor (n380,n105,n381);
or (n381,n104,n364);
and (n382,n383,n264);
xnor (n383,n107,n384);
or (n384,n106,n367);
and (n385,n386,n268);
xnor (n386,n109,n387);
or (n387,n108,n370);
and (n388,n389,n272);
xnor (n389,n113,n390);
or (n390,n119,n373);
wire s0n391,s1n391,notn391;
or (n391,s0n391,s1n391);
not(notn391,n281);
and (s0n391,notn391,1'b0);
and (s1n391,n281,n392);
or (n392,n393,n396,n399,1'b0,1'b0,1'b0,1'b0,1'b0);
and (n393,n394,n89);
xnor (n394,n106,n395);
or (n395,n105,n381);
and (n396,n397,n264);
xnor (n397,n108,n398);
or (n398,n107,n384);
and (n399,n400,n268);
xnor (n400,n119,n401);
or (n401,n109,n387);
wire s0n402,s1n402,notn402;
or (n402,s0n402,s1n402);
not(notn402,n281);
and (s0n402,notn402,1'b0);
and (s1n402,n281,n403);
or (n403,n404,n407,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0);
and (n404,n405,n89);
xnor (n405,n107,n406);
or (n406,n106,n395);
and (n407,n408,n264);
xnor (n408,n109,n409);
or (n409,n108,n398);
wire s0n410,s1n410,notn410;
or (n410,s0n410,s1n410);
not(notn410,n281);
and (s0n410,notn410,1'b0);
and (s1n410,n281,n411);
and (n411,n412,n89);
xnor (n412,n108,n413);
or (n413,n107,n406);
nor (n414,n415,n417,n420);
not (n415,n416);
not (n417,n418);
xor (n418,n419,n416);
xor (n420,n421,n422);
and (n422,n419,n416);
and (n423,n282,n311);
and (n424,n425,n426);
xor (n425,n324,n84);
nor (n426,n282,n427);
not (n427,n311);
and (n428,n84,n429);
and (n429,n282,n427);
not (n430,n431);
or (n431,1'b0,n432,n434,n438);
and (n432,n433,n423);
wire s0n433,s1n433,notn433;
or (n433,s0n433,s1n433);
not(notn433,n414);
and (s0n433,notn433,n324);
and (s1n433,n414,1'b0);
and (n434,n435,n426);
xor (n435,n436,n437);
not (n436,n340);
not (n437,n324);
and (n438,n324,n429);
or (n439,1'b0,n440,n442,n450);
and (n440,n441,n423);
wire s0n441,s1n441,notn441;
or (n441,s0n441,s1n441);
not(notn441,n414);
and (s0n441,notn441,n340);
and (s1n441,n414,1'b0);
and (n442,n443,n426);
wire s0n443,s1n443,notn443;
or (n443,s0n443,s1n443);
not(notn443,n84);
and (s0n443,notn443,n444);
and (s1n443,n84,n447);
xor (n444,n445,n446);
not (n445,n360);
and (n446,n436,n437);
xor (n447,n360,n448);
and (n448,n340,n449);
and (n449,n324,n84);
and (n450,n340,n429);
not (n451,n452);
or (n452,1'b0,n453,n455,n462);
and (n453,n454,n423);
wire s0n454,s1n454,notn454;
or (n454,s0n454,s1n454);
not(notn454,n414);
and (s0n454,notn454,n360);
and (s1n454,n414,1'b0);
and (n455,n456,n426);
wire s0n456,s1n456,notn456;
or (n456,s0n456,s1n456);
not(notn456,n84);
and (s0n456,notn456,n457);
and (s1n456,n84,n460);
xor (n457,n458,n459);
not (n458,n377);
and (n459,n445,n446);
xor (n460,n377,n461);
and (n461,n360,n448);
and (n462,n360,n429);
or (n463,1'b0,n464,n466,n473);
and (n464,n465,n423);
wire s0n465,s1n465,notn465;
or (n465,s0n465,s1n465);
not(notn465,n414);
and (s0n465,notn465,n377);
and (s1n465,n414,1'b0);
and (n466,n467,n426);
wire s0n467,s1n467,notn467;
or (n467,s0n467,s1n467);
not(notn467,n84);
and (s0n467,notn467,n468);
and (s1n467,n84,n471);
xor (n468,n469,n470);
not (n469,n391);
and (n470,n458,n459);
xor (n471,n391,n472);
and (n472,n377,n461);
and (n473,n377,n429);
or (n474,1'b0,n475,n477,n484);
and (n475,n476,n423);
wire s0n476,s1n476,notn476;
or (n476,s0n476,s1n476);
not(notn476,n414);
and (s0n476,notn476,n391);
and (s1n476,n414,1'b0);
and (n477,n478,n426);
wire s0n478,s1n478,notn478;
or (n478,s0n478,s1n478);
not(notn478,n84);
and (s0n478,notn478,n479);
and (s1n478,n84,n482);
xor (n479,n480,n481);
not (n480,n402);
and (n481,n469,n470);
xor (n482,n402,n483);
and (n483,n391,n472);
and (n484,n391,n429);
or (n485,1'b0,n486,n488,n495);
and (n486,n487,n423);
wire s0n487,s1n487,notn487;
or (n487,s0n487,s1n487);
not(notn487,n414);
and (s0n487,notn487,n402);
and (s1n487,n414,1'b0);
and (n488,n489,n426);
wire s0n489,s1n489,notn489;
or (n489,s0n489,s1n489);
not(notn489,n84);
and (s0n489,notn489,n490);
and (s1n489,n84,n493);
xor (n490,n491,n492);
not (n491,n410);
and (n492,n480,n481);
xor (n493,n410,n494);
and (n494,n402,n483);
and (n495,n402,n429);
or (n496,1'b0,n497,n499,n504);
and (n497,n498,n423);
wire s0n498,s1n498,notn498;
or (n498,s0n498,s1n498);
not(notn498,n414);
and (s0n498,notn498,n410);
and (s1n498,n414,1'b0);
and (n499,n500,n426);
wire s0n500,s1n500,notn500;
or (n500,s0n500,s1n500);
not(notn500,n84);
and (s0n500,notn500,n501);
and (s1n500,n84,n503);
not (n501,n502);
and (n502,n491,n492);
and (n503,n410,n494);
and (n504,n410,n429);
nor (n505,n506,n430,n439,n451,n463,n474,n485,n496);
not (n506,n81);
nor (n507,n81,n431,n508,n451,n463,n474,n485,n496);
not (n508,n439);
nor (n509,n506,n431,n508,n451,n463,n474,n485,n496);
nor (n510,n81,n430,n508,n452,n511,n474,n485,n496);
not (n511,n463);
nor (n512,n506,n430,n508,n452,n511,n474,n485,n496);
nor (n513,n81,n431,n439,n451,n511,n474,n485,n496);
nor (n514,n506,n431,n439,n451,n511,n474,n485,n496);
or (n515,n516,n531);
or (n516,n517,n530);
or (n517,n518,n529);
or (n518,n519,n528);
or (n519,n520,n527);
or (n520,n521,n526);
or (n521,n522,n525);
or (n522,n523,n524);
nor (n523,n81,n430,n508,n452,n463,n474,n485,n496);
nor (n524,n506,n430,n508,n452,n463,n474,n485,n496);
nor (n525,n81,n431,n439,n451,n463,n474,n485,n496);
nor (n526,n506,n431,n439,n451,n463,n474,n485,n496);
nor (n527,n81,n430,n439,n452,n511,n474,n485,n496);
nor (n528,n506,n430,n439,n452,n511,n474,n485,n496);
nor (n529,n81,n431,n508,n452,n511,n474,n485,n496);
nor (n530,n506,n431,n508,n452,n511,n474,n485,n496);
or (n531,n532,n545);
or (n532,n533,n544);
or (n533,n534,n543);
or (n534,n535,n542);
or (n535,n536,n541);
or (n536,n537,n540);
or (n537,n538,n539);
nor (n538,n81,n430,n508,n451,n463,n474,n485,n496);
nor (n539,n506,n430,n508,n451,n463,n474,n485,n496);
nor (n540,n81,n431,n439,n452,n511,n474,n485,n496);
nor (n541,n506,n431,n439,n452,n511,n474,n485,n496);
nor (n542,n81,n430,n439,n451,n511,n474,n485,n496);
nor (n543,n506,n430,n439,n451,n511,n474,n485,n496);
nor (n544,n81,n431,n508,n451,n511,n474,n485,n496);
nor (n545,n506,n431,n508,n451,n511,n474,n485,n496);
nor (n546,n506,n431,n508,n452,n463,n474,n485,n496);
or (n547,1'b0,n548,n555,n562,n323);
or (n548,n549,n513);
or (n549,n550,n512);
or (n550,n551,n510);
or (n551,n552,n530);
or (n552,n553,n507);
or (n553,n554,n505);
or (n554,n526,n80);
or (n555,n556,n529);
or (n556,n557,n528);
or (n557,n558,n527);
or (n558,n559,n541);
or (n559,n560,n525);
or (n560,n561,n524);
or (n561,n546,n523);
or (n562,n563,n540);
or (n563,n564,n539);
or (n564,n565,n538);
or (n565,n566,n509);
or (n566,n567,n572);
or (n567,n568,n571);
or (n568,n569,n570);
nor (n569,n506,n431,n439,n452,n463,n474,n485,n496);
nor (n570,n81,n430,n439,n452,n463,n474,n485,n496);
nor (n571,n506,n430,n439,n452,n463,n474,n485,n496);
nor (n572,n81,n431,n508,n452,n463,n474,n485,n496);
or (n573,n574,n579);
nor (n574,n575,n576,n578);
not (n576,n577);
and (n579,n575,n577,n578);
nor (n580,n205,n211,n208,n209);
or (n582,n583,n587,n590,n592);
and (n583,n52,n584);
and (n584,n585,n586);
and (n587,n57,n588);
and (n588,n589,n586);
not (n589,n585);
and (n590,n61,n591);
nor (n591,n589,n586);
and (n592,n64,n593);
nor (n593,n585,n586);
and (n594,n67,n595);
not (n595,n581);
and (n596,n597,n58);
wire s0n597,s1n597,notn597;
or (n597,s0n597,s1n597);
not(notn597,n48);
and (s0n597,notn597,n598);
and (s1n597,n48,n599);
or (n599,n600,n602,n604,n606);
and (n600,n601,n36);
and (n602,n603,n41);
and (n604,n605,n45);
and (n606,n598,n47);
and (n607,n608,n62);
wire s0n608,s1n608,notn608;
or (n608,s0n608,s1n608);
not(notn608,n48);
and (s0n608,notn608,n609);
and (s1n608,n48,n610);
or (n610,n611,n613,n615,n617);
and (n611,n612,n36);
and (n613,n614,n41);
and (n615,n616,n45);
and (n617,n609,n47);
and (n618,n619,n65);
wire s0n619,s1n619,notn619;
or (n619,s0n619,s1n619);
not(notn619,n48);
and (s0n619,notn619,n620);
and (s1n619,n48,n621);
or (n621,n622,n624,n626,n628);
and (n622,n623,n36);
and (n624,n625,n41);
and (n626,n627,n45);
and (n628,n620,n47);
wire s0n630,s1n630,notn630;
or (n630,s0n630,s1n630);
not(notn630,n629);
and (s0n630,notn630,n631);
and (s1n630,n629,n620);
wire s0n631,s1n631,notn631;
or (n631,s0n631,s1n631);
not(notn631,n48);
and (s0n631,notn631,n632);
and (s1n631,n48,n637);
or (n632,n633,n634,n635,n636);
and (n633,n32,n584);
and (n634,n598,n588);
and (n635,n609,n591);
and (n636,n620,n593);
or (n637,1'b0,n638,n640,n642,n645,n647,n649,n651,n653,n655,n657,n659,n661,n663,n665,n667,n669);
and (n638,n35,n639);
and (n639,n54,n55,n585,n586,n595);
and (n640,n40,n641);
and (n641,n59,n55,n585,n586,n595);
and (n642,n44,n643);
and (n643,n54,n644,n585,n586,n595);
not (n644,n55);
and (n645,n32,n646);
and (n646,n59,n644,n585,n586,n595);
and (n647,n601,n648);
and (n648,n54,n55,n589,n586,n595);
and (n649,n603,n650);
and (n650,n59,n55,n589,n586,n595);
and (n651,n605,n652);
and (n652,n54,n644,n589,n586,n595);
and (n653,n598,n654);
and (n654,n59,n644,n589,n586,n595);
and (n655,n612,n656);
nor (n656,n59,n644,n589,n586,n581);
and (n657,n614,n658);
nor (n658,n54,n644,n589,n586,n581);
and (n659,n616,n660);
nor (n660,n59,n55,n589,n586,n581);
and (n661,n609,n662);
nor (n662,n54,n55,n589,n586,n581);
and (n663,n623,n664);
nor (n664,n59,n644,n585,n586,n581);
and (n665,n625,n666);
nor (n666,n54,n644,n585,n586,n581);
and (n667,n627,n668);
nor (n668,n59,n55,n585,n586,n581);
and (n669,n620,n670);
nor (n670,n54,n55,n585,n586,n581);
wire s0n671,s1n671,notn671;
or (n671,s0n671,s1n671);
not(notn671,n594);
and (s0n671,notn671,1'b0);
and (s1n671,n594,n672);
wire s0n672,s1n672,notn672;
or (n672,s0n672,s1n672);
not(notn672,n594);
and (s0n672,notn672,n673);
and (s1n672,n594,n720);
wire s0n673,s1n673,notn673;
or (n673,s0n673,s1n673);
not(notn673,n66);
and (s0n673,notn673,1'b0);
and (s1n673,n66,n674);
wire s0n674,s1n674,notn674;
or (n674,s0n674,s1n674);
not(notn674,n629);
and (s0n674,notn674,n675);
and (s1n674,n629,n711);
or (n675,n676,n687,n698,n709);
and (n676,n677,n53);
wire s0n677,s1n677,notn677;
or (n677,s0n677,s1n677);
not(notn677,n48);
and (s0n677,notn677,n678);
and (s1n677,n48,n679);
or (n679,n680,n682,n684,n686);
and (n680,n681,n36);
and (n682,n683,n41);
and (n684,n685,n45);
and (n686,n678,n47);
and (n687,n688,n58);
wire s0n688,s1n688,notn688;
or (n688,s0n688,s1n688);
not(notn688,n48);
and (s0n688,notn688,n689);
and (s1n688,n48,n690);
or (n690,n691,n693,n695,n697);
and (n691,n692,n36);
and (n693,n694,n41);
and (n695,n696,n45);
and (n697,n689,n47);
and (n698,n699,n62);
wire s0n699,s1n699,notn699;
or (n699,s0n699,s1n699);
not(notn699,n48);
and (s0n699,notn699,n700);
and (s1n699,n48,n701);
or (n701,n702,n704,n706,n708);
and (n702,n703,n36);
and (n704,n705,n41);
and (n706,n707,n45);
and (n708,n700,n47);
and (n709,n710,n65);
wire s0n710,s1n710,notn710;
or (n710,s0n710,s1n710);
not(notn710,n48);
and (s0n710,notn710,n711);
and (s1n710,n48,n712);
or (n712,n713,n715,n717,n719);
and (n713,n714,n36);
and (n715,n716,n41);
and (n717,n718,n45);
and (n719,n711,n47);
wire s0n720,s1n720,notn720;
or (n720,s0n720,s1n720);
not(notn720,n629);
and (s0n720,notn720,n721);
and (s1n720,n629,n711);
wire s0n721,s1n721,notn721;
or (n721,s0n721,s1n721);
not(notn721,n48);
and (s0n721,notn721,n722);
and (s1n721,n48,n727);
or (n722,n723,n724,n725,n726);
and (n723,n678,n584);
and (n724,n689,n588);
and (n725,n700,n591);
and (n726,n711,n593);
or (n727,1'b0,n728,n729,n730,n731,n732,n733,n734,n735,n736,n737,n738,n739,n740,n741,n742,n743);
and (n728,n681,n639);
and (n729,n683,n641);
and (n730,n685,n643);
and (n731,n678,n646);
and (n732,n692,n648);
and (n733,n694,n650);
and (n734,n696,n652);
and (n735,n689,n654);
and (n736,n703,n656);
and (n737,n705,n658);
and (n738,n707,n660);
and (n739,n700,n662);
and (n740,n714,n664);
and (n741,n716,n666);
and (n742,n718,n668);
and (n743,n711,n670);
wire s0n744,s1n744,notn744;
or (n744,s0n744,s1n744);
not(notn744,n594);
and (s0n744,notn744,1'b0);
and (s1n744,n594,n745);
wire s0n745,s1n745,notn745;
or (n745,s0n745,s1n745);
not(notn745,n594);
and (s0n745,notn745,n746);
and (s1n745,n594,n793);
wire s0n746,s1n746,notn746;
or (n746,s0n746,s1n746);
not(notn746,n66);
and (s0n746,notn746,1'b0);
and (s1n746,n66,n747);
wire s0n747,s1n747,notn747;
or (n747,s0n747,s1n747);
not(notn747,n629);
and (s0n747,notn747,n748);
and (s1n747,n629,n784);
or (n748,n749,n760,n771,n782);
and (n749,n750,n53);
wire s0n750,s1n750,notn750;
or (n750,s0n750,s1n750);
not(notn750,n48);
and (s0n750,notn750,n751);
and (s1n750,n48,n752);
or (n752,n753,n755,n757,n759);
and (n753,n754,n36);
and (n755,n756,n41);
and (n757,n758,n45);
and (n759,n751,n47);
and (n760,n761,n58);
wire s0n761,s1n761,notn761;
or (n761,s0n761,s1n761);
not(notn761,n48);
and (s0n761,notn761,n762);
and (s1n761,n48,n763);
or (n763,n764,n766,n768,n770);
and (n764,n765,n36);
and (n766,n767,n41);
and (n768,n769,n45);
and (n770,n762,n47);
and (n771,n772,n62);
wire s0n772,s1n772,notn772;
or (n772,s0n772,s1n772);
not(notn772,n48);
and (s0n772,notn772,n773);
and (s1n772,n48,n774);
or (n774,n775,n777,n779,n781);
and (n775,n776,n36);
and (n777,n778,n41);
and (n779,n780,n45);
and (n781,n773,n47);
and (n782,n783,n65);
wire s0n783,s1n783,notn783;
or (n783,s0n783,s1n783);
not(notn783,n48);
and (s0n783,notn783,n784);
and (s1n783,n48,n785);
or (n785,n786,n788,n790,n792);
and (n786,n787,n36);
and (n788,n789,n41);
and (n790,n791,n45);
and (n792,n784,n47);
wire s0n793,s1n793,notn793;
or (n793,s0n793,s1n793);
not(notn793,n629);
and (s0n793,notn793,n794);
and (s1n793,n629,n784);
wire s0n794,s1n794,notn794;
or (n794,s0n794,s1n794);
not(notn794,n48);
and (s0n794,notn794,n795);
and (s1n794,n48,n800);
or (n795,n796,n797,n798,n799);
and (n796,n751,n584);
and (n797,n762,n588);
and (n798,n773,n591);
and (n799,n784,n593);
or (n800,1'b0,n801,n802,n803,n804,n805,n806,n807,n808,n809,n810,n811,n812,n813,n814,n815,n816);
and (n801,n754,n639);
and (n802,n756,n641);
and (n803,n758,n643);
and (n804,n751,n646);
and (n805,n765,n648);
and (n806,n767,n650);
and (n807,n769,n652);
and (n808,n762,n654);
and (n809,n776,n656);
and (n810,n778,n658);
and (n811,n780,n660);
and (n812,n773,n662);
and (n813,n787,n664);
and (n814,n789,n666);
and (n815,n791,n668);
and (n816,n784,n670);
not (n817,n818);
wire s0n818,s1n818,notn818;
or (n818,s0n818,s1n818);
not(notn818,n594);
and (s0n818,notn818,1'b0);
and (s1n818,n594,n819);
wire s0n819,s1n819,notn819;
or (n819,s0n819,s1n819);
not(notn819,n594);
and (s0n819,notn819,n820);
and (s1n819,n594,n867);
wire s0n820,s1n820,notn820;
or (n820,s0n820,s1n820);
not(notn820,n66);
and (s0n820,notn820,1'b0);
and (s1n820,n66,n821);
wire s0n821,s1n821,notn821;
or (n821,s0n821,s1n821);
not(notn821,n629);
and (s0n821,notn821,n822);
and (s1n821,n629,n858);
or (n822,n823,n834,n845,n856);
and (n823,n824,n53);
wire s0n824,s1n824,notn824;
or (n824,s0n824,s1n824);
not(notn824,n48);
and (s0n824,notn824,n825);
and (s1n824,n48,n826);
or (n826,n827,n829,n831,n833);
and (n827,n828,n36);
and (n829,n830,n41);
and (n831,n832,n45);
and (n833,n825,n47);
and (n834,n835,n58);
wire s0n835,s1n835,notn835;
or (n835,s0n835,s1n835);
not(notn835,n48);
and (s0n835,notn835,n836);
and (s1n835,n48,n837);
or (n837,n838,n840,n842,n844);
and (n838,n839,n36);
and (n840,n841,n41);
and (n842,n843,n45);
and (n844,n836,n47);
and (n845,n846,n62);
wire s0n846,s1n846,notn846;
or (n846,s0n846,s1n846);
not(notn846,n48);
and (s0n846,notn846,n847);
and (s1n846,n48,n848);
or (n848,n849,n851,n853,n855);
and (n849,n850,n36);
and (n851,n852,n41);
and (n853,n854,n45);
and (n855,n847,n47);
and (n856,n857,n65);
wire s0n857,s1n857,notn857;
or (n857,s0n857,s1n857);
not(notn857,n48);
and (s0n857,notn857,n858);
and (s1n857,n48,n859);
or (n859,n860,n862,n864,n866);
and (n860,n861,n36);
and (n862,n863,n41);
and (n864,n865,n45);
and (n866,n858,n47);
wire s0n867,s1n867,notn867;
or (n867,s0n867,s1n867);
not(notn867,n629);
and (s0n867,notn867,n868);
and (s1n867,n629,n858);
wire s0n868,s1n868,notn868;
or (n868,s0n868,s1n868);
not(notn868,n48);
and (s0n868,notn868,n869);
and (s1n868,n48,n874);
or (n869,n870,n871,n872,n873);
and (n870,n825,n584);
and (n871,n836,n588);
and (n872,n847,n591);
and (n873,n858,n593);
or (n874,1'b0,n875,n876,n877,n878,n879,n880,n881,n882,n883,n884,n885,n886,n887,n888,n889,n890);
and (n875,n828,n639);
and (n876,n830,n641);
and (n877,n832,n643);
and (n878,n825,n646);
and (n879,n839,n648);
and (n880,n841,n650);
and (n881,n843,n652);
and (n882,n836,n654);
and (n883,n850,n656);
and (n884,n852,n658);
and (n885,n854,n660);
and (n886,n847,n662);
and (n887,n861,n664);
and (n888,n863,n666);
and (n889,n865,n668);
and (n890,n858,n670);
and (n891,n25,n671,n892,n818);
not (n892,n744);
and (n893,n894,n904);
wire s0n894,s1n894,notn894;
or (n894,s0n894,s1n894);
not(notn894,n896);
and (s0n894,notn894,1'b0);
and (s1n894,n896,n895);
or (n896,n897,n903);
or (n897,n898,n901);
or (n898,n899,n900);
and (n899,n15,n17,n18,n19);
not (n900,n14);
nor (n901,n902,n16,n18,n20);
not (n902,n15);
nor (n903,n902,n17,n18,n20);
or (n904,n905,n906);
and (n905,n24,n671,n744,n817);
and (n906,n24,n671,n744,n818);
and (n907,n908,n2971);
wire s0n908,s1n908,notn908;
or (n908,s0n908,s1n908);
not(notn908,n2966);
and (s0n908,notn908,n909);
and (s1n908,n2966,1'b0);
wire s0n909,s1n909,notn909;
or (n909,s0n909,s1n909);
not(notn909,n2961);
and (s0n909,notn909,n910);
and (s1n909,n2961,1'b1);
wire s0n910,s1n910,notn910;
or (n910,s0n910,s1n910);
not(notn910,n2948);
and (s0n910,notn910,1'b0);
and (s1n910,n2948,n911);
xor (n911,n912,n2925);
xor (n912,n913,n2872);
xor (n913,n914,n2448);
xor (n914,n915,n2446);
xor (n915,n916,n2416);
not (n916,n917);
or (n917,n918,n1831);
or (n918,n919,n1076,n1830);
and (n919,n920,n1045);
or (n920,1'b0,n921,n984,n1004,n1024);
and (n921,n922,n981);
or (n922,1'b0,n923,n951,n961,n971);
and (n923,n924,n930);
wire s0n924,s1n924,notn924;
or (n924,s0n924,s1n924);
not(notn924,n927);
and (s0n924,notn924,n925);
and (s1n924,n927,n926);
or (n927,n928,n929);
and (n928,n25,n671,n744,n817);
and (n929,n25,n671,n744,n818);
or (n930,n931,n950);
or (n931,n932,n945);
and (n932,n933,n903);
or (n933,n934,n929);
or (n934,n935,n928);
or (n935,n936,n944);
or (n936,n937,n943);
or (n937,n938,n942);
or (n938,n939,n940);
nor (n939,n25,n671,n744,n817);
and (n940,n24,n941,n744,n817);
not (n941,n671);
and (n942,n24,n941,n744,n818);
and (n943,n25,n941,n744,n817);
and (n944,n25,n941,n744,n818);
and (n945,n946,n949);
or (n946,n947,n891);
or (n947,n948,n23);
nor (n948,n25,n941,n744,n817);
nor (n949,n15,n16,n18,n20);
and (n950,n904,n949);
and (n951,n952,n955);
wire s0n952,s1n952,notn952;
or (n952,s0n952,s1n952);
not(notn952,n927);
and (s0n952,notn952,n953);
and (s1n952,n927,n954);
or (n955,n956,n959);
or (n956,n957,n958);
and (n957,n933,n949);
and (n958,n946,n901);
and (n959,n904,n960);
and (n960,n902,n16,n18,n19);
and (n961,n962,n965);
wire s0n962,s1n962,notn962;
or (n962,s0n962,s1n962);
not(notn962,n927);
and (s0n962,notn962,n963);
and (s1n962,n927,n964);
or (n965,n966,n969);
or (n966,n967,n968);
and (n967,n933,n901);
and (n968,n946,n960);
and (n969,n904,n970);
and (n970,n902,n17,n18,n19);
and (n971,n972,n975);
wire s0n972,s1n972,notn972;
or (n972,s0n972,s1n972);
not(notn972,n927);
and (s0n972,notn972,n973);
and (s1n972,n927,n974);
or (n975,n976,n979);
or (n976,n977,n978);
and (n977,n933,n960);
and (n978,n946,n900);
and (n979,n904,n980);
nor (n980,n15,n17,n18,n19);
and (n981,n594,n982);
and (n982,n983,n53);
not (n983,n48);
and (n984,n985,n1002);
or (n985,1'b0,n986,n990,n994,n998);
and (n986,n987,n930);
wire s0n987,s1n987,notn987;
or (n987,s0n987,s1n987);
not(notn987,n927);
and (s0n987,notn987,n988);
and (s1n987,n927,n989);
and (n990,n991,n955);
wire s0n991,s1n991,notn991;
or (n991,s0n991,s1n991);
not(notn991,n927);
and (s0n991,notn991,n992);
and (s1n991,n927,n993);
and (n994,n995,n965);
wire s0n995,s1n995,notn995;
or (n995,s0n995,s1n995);
not(notn995,n927);
and (s0n995,notn995,n996);
and (s1n995,n927,n997);
and (n998,n999,n975);
wire s0n999,s1n999,notn999;
or (n999,s0n999,s1n999);
not(notn999,n927);
and (s0n999,notn999,n1000);
and (s1n999,n927,n1001);
and (n1002,n594,n1003);
and (n1003,n983,n58);
and (n1004,n1005,n1022);
or (n1005,1'b0,n1006,n1010,n1014,n1018);
and (n1006,n1007,n930);
wire s0n1007,s1n1007,notn1007;
or (n1007,s0n1007,s1n1007);
not(notn1007,n927);
and (s0n1007,notn1007,n1008);
and (s1n1007,n927,n1009);
and (n1010,n1011,n955);
wire s0n1011,s1n1011,notn1011;
or (n1011,s0n1011,s1n1011);
not(notn1011,n927);
and (s0n1011,notn1011,n1012);
and (s1n1011,n927,n1013);
and (n1014,n1015,n965);
wire s0n1015,s1n1015,notn1015;
or (n1015,s0n1015,s1n1015);
not(notn1015,n927);
and (s0n1015,notn1015,n1016);
and (s1n1015,n927,n1017);
and (n1018,n1019,n975);
wire s0n1019,s1n1019,notn1019;
or (n1019,s0n1019,s1n1019);
not(notn1019,n927);
and (s0n1019,notn1019,n1020);
and (s1n1019,n927,n1021);
and (n1022,n594,n1023);
and (n1023,n983,n62);
and (n1024,n1025,n1042);
or (n1025,1'b0,n1026,n1030,n1034,n1038);
and (n1026,n1027,n930);
wire s0n1027,s1n1027,notn1027;
or (n1027,s0n1027,s1n1027);
not(notn1027,n927);
and (s0n1027,notn1027,n1028);
and (s1n1027,n927,n1029);
and (n1030,n1031,n955);
wire s0n1031,s1n1031,notn1031;
or (n1031,s0n1031,s1n1031);
not(notn1031,n927);
and (s0n1031,notn1031,n1032);
and (s1n1031,n927,n1033);
and (n1034,n1035,n965);
wire s0n1035,s1n1035,notn1035;
or (n1035,s0n1035,s1n1035);
not(notn1035,n927);
and (s0n1035,notn1035,n1036);
and (s1n1035,n927,n1037);
and (n1038,n1039,n975);
wire s0n1039,s1n1039,notn1039;
or (n1039,s0n1039,s1n1039);
not(notn1039,n927);
and (s0n1039,notn1039,n1040);
and (s1n1039,n927,n1041);
and (n1042,n594,n1043);
or (n1043,n48,n1044);
and (n1044,n983,n65);
or (n1045,1'b0,n1046,n1055,n1061,n1070);
and (n1046,n1047,n981);
or (n1047,1'b0,n1048,n1052,n1053,n1054);
and (n1048,n1049,n930);
wire s0n1049,s1n1049,notn1049;
or (n1049,s0n1049,s1n1049);
not(notn1049,n927);
and (s0n1049,notn1049,n1050);
and (s1n1049,n927,n1051);
and (n1052,n924,n955);
and (n1053,n952,n965);
and (n1054,n962,n975);
and (n1055,n1056,n1002);
or (n1056,1'b0,n1057,n1058,n1059,n1060);
and (n1057,n972,n930);
and (n1058,n987,n955);
and (n1059,n991,n965);
and (n1060,n995,n975);
and (n1061,n1062,n1022);
or (n1062,1'b0,n1063,n1067,n1068,n1069);
and (n1063,n1064,n930);
wire s0n1064,s1n1064,notn1064;
or (n1064,s0n1064,s1n1064);
not(notn1064,n927);
and (s0n1064,notn1064,n1065);
and (s1n1064,n927,n1066);
and (n1067,n1007,n955);
and (n1068,n1011,n965);
and (n1069,n1015,n975);
and (n1070,n1071,n1042);
or (n1071,1'b0,n1072,n1073,n1074,n1075);
and (n1072,n1019,n930);
and (n1073,n1027,n955);
and (n1074,n1031,n965);
and (n1075,n1035,n975);
and (n1076,n1045,n1077);
or (n1077,n1078,n1183,n1829);
and (n1078,n1079,n1152);
or (n1079,1'b0,n1080,n1098,n1116,n1134);
and (n1080,n1081,n981);
or (n1081,1'b0,n1082,n1086,n1090,n1094);
and (n1082,n1083,n930);
wire s0n1083,s1n1083,notn1083;
or (n1083,s0n1083,s1n1083);
not(notn1083,n927);
and (s0n1083,notn1083,n1084);
and (s1n1083,n927,n1085);
and (n1086,n1087,n955);
wire s0n1087,s1n1087,notn1087;
or (n1087,s0n1087,s1n1087);
not(notn1087,n927);
and (s0n1087,notn1087,n1088);
and (s1n1087,n927,n1089);
and (n1090,n1091,n965);
wire s0n1091,s1n1091,notn1091;
or (n1091,s0n1091,s1n1091);
not(notn1091,n927);
and (s0n1091,notn1091,n1092);
and (s1n1091,n927,n1093);
and (n1094,n1095,n975);
wire s0n1095,s1n1095,notn1095;
or (n1095,s0n1095,s1n1095);
not(notn1095,n927);
and (s0n1095,notn1095,n1096);
and (s1n1095,n927,n1097);
and (n1098,n1099,n1002);
or (n1099,1'b0,n1100,n1104,n1108,n1112);
and (n1100,n1101,n930);
wire s0n1101,s1n1101,notn1101;
or (n1101,s0n1101,s1n1101);
not(notn1101,n927);
and (s0n1101,notn1101,n1102);
and (s1n1101,n927,n1103);
and (n1104,n1105,n955);
wire s0n1105,s1n1105,notn1105;
or (n1105,s0n1105,s1n1105);
not(notn1105,n927);
and (s0n1105,notn1105,n1106);
and (s1n1105,n927,n1107);
and (n1108,n1109,n965);
wire s0n1109,s1n1109,notn1109;
or (n1109,s0n1109,s1n1109);
not(notn1109,n927);
and (s0n1109,notn1109,n1110);
and (s1n1109,n927,n1111);
and (n1112,n1113,n975);
wire s0n1113,s1n1113,notn1113;
or (n1113,s0n1113,s1n1113);
not(notn1113,n927);
and (s0n1113,notn1113,n1114);
and (s1n1113,n927,n1115);
and (n1116,n1117,n1022);
or (n1117,1'b0,n1118,n1122,n1126,n1130);
and (n1118,n1119,n930);
wire s0n1119,s1n1119,notn1119;
or (n1119,s0n1119,s1n1119);
not(notn1119,n927);
and (s0n1119,notn1119,n1120);
and (s1n1119,n927,n1121);
and (n1122,n1123,n955);
wire s0n1123,s1n1123,notn1123;
or (n1123,s0n1123,s1n1123);
not(notn1123,n927);
and (s0n1123,notn1123,n1124);
and (s1n1123,n927,n1125);
and (n1126,n1127,n965);
wire s0n1127,s1n1127,notn1127;
or (n1127,s0n1127,s1n1127);
not(notn1127,n927);
and (s0n1127,notn1127,n1128);
and (s1n1127,n927,n1129);
and (n1130,n1131,n975);
wire s0n1131,s1n1131,notn1131;
or (n1131,s0n1131,s1n1131);
not(notn1131,n927);
and (s0n1131,notn1131,n1132);
and (s1n1131,n927,n1133);
and (n1134,n1135,n1042);
or (n1135,1'b0,n1136,n1140,n1144,n1148);
and (n1136,n1137,n930);
wire s0n1137,s1n1137,notn1137;
or (n1137,s0n1137,s1n1137);
not(notn1137,n927);
and (s0n1137,notn1137,n1138);
and (s1n1137,n927,n1139);
and (n1140,n1141,n955);
wire s0n1141,s1n1141,notn1141;
or (n1141,s0n1141,s1n1141);
not(notn1141,n927);
and (s0n1141,notn1141,n1142);
and (s1n1141,n927,n1143);
and (n1144,n1145,n965);
wire s0n1145,s1n1145,notn1145;
or (n1145,s0n1145,s1n1145);
not(notn1145,n927);
and (s0n1145,notn1145,n1146);
and (s1n1145,n927,n1147);
and (n1148,n1149,n975);
wire s0n1149,s1n1149,notn1149;
or (n1149,s0n1149,s1n1149);
not(notn1149,n927);
and (s0n1149,notn1149,n1150);
and (s1n1149,n927,n1151);
or (n1152,1'b0,n1153,n1162,n1168,n1177);
and (n1153,n1154,n981);
or (n1154,1'b0,n1155,n1159,n1160,n1161);
and (n1155,n1156,n930);
wire s0n1156,s1n1156,notn1156;
or (n1156,s0n1156,s1n1156);
not(notn1156,n927);
and (s0n1156,notn1156,n1157);
and (s1n1156,n927,n1158);
and (n1159,n1083,n955);
and (n1160,n1087,n965);
and (n1161,n1091,n975);
and (n1162,n1163,n1002);
or (n1163,1'b0,n1164,n1165,n1166,n1167);
and (n1164,n1095,n930);
and (n1165,n1101,n955);
and (n1166,n1105,n965);
and (n1167,n1109,n975);
and (n1168,n1169,n1022);
or (n1169,1'b0,n1170,n1174,n1175,n1176);
and (n1170,n1171,n930);
wire s0n1171,s1n1171,notn1171;
or (n1171,s0n1171,s1n1171);
not(notn1171,n927);
and (s0n1171,notn1171,n1172);
and (s1n1171,n927,n1173);
and (n1174,n1119,n955);
and (n1175,n1123,n965);
and (n1176,n1127,n975);
and (n1177,n1178,n1042);
or (n1178,1'b0,n1179,n1180,n1181,n1182);
and (n1179,n1131,n930);
and (n1180,n1137,n955);
and (n1181,n1141,n965);
and (n1182,n1145,n975);
and (n1183,n1152,n1184);
or (n1184,n1185,n1290,n1828);
and (n1185,n1186,n1259);
or (n1186,1'b0,n1187,n1205,n1223,n1241);
and (n1187,n1188,n981);
or (n1188,1'b0,n1189,n1193,n1197,n1201);
and (n1189,n1190,n930);
wire s0n1190,s1n1190,notn1190;
or (n1190,s0n1190,s1n1190);
not(notn1190,n927);
and (s0n1190,notn1190,n1191);
and (s1n1190,n927,n1192);
and (n1193,n1194,n955);
wire s0n1194,s1n1194,notn1194;
or (n1194,s0n1194,s1n1194);
not(notn1194,n927);
and (s0n1194,notn1194,n1195);
and (s1n1194,n927,n1196);
and (n1197,n1198,n965);
wire s0n1198,s1n1198,notn1198;
or (n1198,s0n1198,s1n1198);
not(notn1198,n927);
and (s0n1198,notn1198,n1199);
and (s1n1198,n927,n1200);
and (n1201,n1202,n975);
wire s0n1202,s1n1202,notn1202;
or (n1202,s0n1202,s1n1202);
not(notn1202,n927);
and (s0n1202,notn1202,n1203);
and (s1n1202,n927,n1204);
and (n1205,n1206,n1002);
or (n1206,1'b0,n1207,n1211,n1215,n1219);
and (n1207,n1208,n930);
wire s0n1208,s1n1208,notn1208;
or (n1208,s0n1208,s1n1208);
not(notn1208,n927);
and (s0n1208,notn1208,n1209);
and (s1n1208,n927,n1210);
and (n1211,n1212,n955);
wire s0n1212,s1n1212,notn1212;
or (n1212,s0n1212,s1n1212);
not(notn1212,n927);
and (s0n1212,notn1212,n1213);
and (s1n1212,n927,n1214);
and (n1215,n1216,n965);
wire s0n1216,s1n1216,notn1216;
or (n1216,s0n1216,s1n1216);
not(notn1216,n927);
and (s0n1216,notn1216,n1217);
and (s1n1216,n927,n1218);
and (n1219,n1220,n975);
wire s0n1220,s1n1220,notn1220;
or (n1220,s0n1220,s1n1220);
not(notn1220,n927);
and (s0n1220,notn1220,n1221);
and (s1n1220,n927,n1222);
and (n1223,n1224,n1022);
or (n1224,1'b0,n1225,n1229,n1233,n1237);
and (n1225,n1226,n930);
wire s0n1226,s1n1226,notn1226;
or (n1226,s0n1226,s1n1226);
not(notn1226,n927);
and (s0n1226,notn1226,n1227);
and (s1n1226,n927,n1228);
and (n1229,n1230,n955);
wire s0n1230,s1n1230,notn1230;
or (n1230,s0n1230,s1n1230);
not(notn1230,n927);
and (s0n1230,notn1230,n1231);
and (s1n1230,n927,n1232);
and (n1233,n1234,n965);
wire s0n1234,s1n1234,notn1234;
or (n1234,s0n1234,s1n1234);
not(notn1234,n927);
and (s0n1234,notn1234,n1235);
and (s1n1234,n927,n1236);
and (n1237,n1238,n975);
wire s0n1238,s1n1238,notn1238;
or (n1238,s0n1238,s1n1238);
not(notn1238,n927);
and (s0n1238,notn1238,n1239);
and (s1n1238,n927,n1240);
and (n1241,n1242,n1042);
or (n1242,1'b0,n1243,n1247,n1251,n1255);
and (n1243,n1244,n930);
wire s0n1244,s1n1244,notn1244;
or (n1244,s0n1244,s1n1244);
not(notn1244,n927);
and (s0n1244,notn1244,n1245);
and (s1n1244,n927,n1246);
and (n1247,n1248,n955);
wire s0n1248,s1n1248,notn1248;
or (n1248,s0n1248,s1n1248);
not(notn1248,n927);
and (s0n1248,notn1248,n1249);
and (s1n1248,n927,n1250);
and (n1251,n1252,n965);
wire s0n1252,s1n1252,notn1252;
or (n1252,s0n1252,s1n1252);
not(notn1252,n927);
and (s0n1252,notn1252,n1253);
and (s1n1252,n927,n1254);
and (n1255,n1256,n975);
wire s0n1256,s1n1256,notn1256;
or (n1256,s0n1256,s1n1256);
not(notn1256,n927);
and (s0n1256,notn1256,n1257);
and (s1n1256,n927,n1258);
or (n1259,1'b0,n1260,n1269,n1275,n1284);
and (n1260,n1261,n981);
or (n1261,1'b0,n1262,n1266,n1267,n1268);
and (n1262,n1263,n930);
wire s0n1263,s1n1263,notn1263;
or (n1263,s0n1263,s1n1263);
not(notn1263,n927);
and (s0n1263,notn1263,n1264);
and (s1n1263,n927,n1265);
and (n1266,n1190,n955);
and (n1267,n1194,n965);
and (n1268,n1198,n975);
and (n1269,n1270,n1002);
or (n1270,1'b0,n1271,n1272,n1273,n1274);
and (n1271,n1202,n930);
and (n1272,n1208,n955);
and (n1273,n1212,n965);
and (n1274,n1216,n975);
and (n1275,n1276,n1022);
or (n1276,1'b0,n1277,n1281,n1282,n1283);
and (n1277,n1278,n930);
wire s0n1278,s1n1278,notn1278;
or (n1278,s0n1278,s1n1278);
not(notn1278,n927);
and (s0n1278,notn1278,n1279);
and (s1n1278,n927,n1280);
and (n1281,n1226,n955);
and (n1282,n1230,n965);
and (n1283,n1234,n975);
and (n1284,n1285,n1042);
or (n1285,1'b0,n1286,n1287,n1288,n1289);
and (n1286,n1238,n930);
and (n1287,n1244,n955);
and (n1288,n1248,n965);
and (n1289,n1252,n975);
and (n1290,n1259,n1291);
or (n1291,n1292,n1397,n1827);
and (n1292,n1293,n1366);
or (n1293,1'b0,n1294,n1312,n1330,n1348);
and (n1294,n1295,n981);
or (n1295,1'b0,n1296,n1300,n1304,n1308);
and (n1296,n1297,n930);
wire s0n1297,s1n1297,notn1297;
or (n1297,s0n1297,s1n1297);
not(notn1297,n927);
and (s0n1297,notn1297,n1298);
and (s1n1297,n927,n1299);
and (n1300,n1301,n955);
wire s0n1301,s1n1301,notn1301;
or (n1301,s0n1301,s1n1301);
not(notn1301,n927);
and (s0n1301,notn1301,n1302);
and (s1n1301,n927,n1303);
and (n1304,n1305,n965);
wire s0n1305,s1n1305,notn1305;
or (n1305,s0n1305,s1n1305);
not(notn1305,n927);
and (s0n1305,notn1305,n1306);
and (s1n1305,n927,n1307);
and (n1308,n1309,n975);
wire s0n1309,s1n1309,notn1309;
or (n1309,s0n1309,s1n1309);
not(notn1309,n927);
and (s0n1309,notn1309,n1310);
and (s1n1309,n927,n1311);
and (n1312,n1313,n1002);
or (n1313,1'b0,n1314,n1318,n1322,n1326);
and (n1314,n1315,n930);
wire s0n1315,s1n1315,notn1315;
or (n1315,s0n1315,s1n1315);
not(notn1315,n927);
and (s0n1315,notn1315,n1316);
and (s1n1315,n927,n1317);
and (n1318,n1319,n955);
wire s0n1319,s1n1319,notn1319;
or (n1319,s0n1319,s1n1319);
not(notn1319,n927);
and (s0n1319,notn1319,n1320);
and (s1n1319,n927,n1321);
and (n1322,n1323,n965);
wire s0n1323,s1n1323,notn1323;
or (n1323,s0n1323,s1n1323);
not(notn1323,n927);
and (s0n1323,notn1323,n1324);
and (s1n1323,n927,n1325);
and (n1326,n1327,n975);
wire s0n1327,s1n1327,notn1327;
or (n1327,s0n1327,s1n1327);
not(notn1327,n927);
and (s0n1327,notn1327,n1328);
and (s1n1327,n927,n1329);
and (n1330,n1331,n1022);
or (n1331,1'b0,n1332,n1336,n1340,n1344);
and (n1332,n1333,n930);
wire s0n1333,s1n1333,notn1333;
or (n1333,s0n1333,s1n1333);
not(notn1333,n927);
and (s0n1333,notn1333,n1334);
and (s1n1333,n927,n1335);
and (n1336,n1337,n955);
wire s0n1337,s1n1337,notn1337;
or (n1337,s0n1337,s1n1337);
not(notn1337,n927);
and (s0n1337,notn1337,n1338);
and (s1n1337,n927,n1339);
and (n1340,n1341,n965);
wire s0n1341,s1n1341,notn1341;
or (n1341,s0n1341,s1n1341);
not(notn1341,n927);
and (s0n1341,notn1341,n1342);
and (s1n1341,n927,n1343);
and (n1344,n1345,n975);
wire s0n1345,s1n1345,notn1345;
or (n1345,s0n1345,s1n1345);
not(notn1345,n927);
and (s0n1345,notn1345,n1346);
and (s1n1345,n927,n1347);
and (n1348,n1349,n1042);
or (n1349,1'b0,n1350,n1354,n1358,n1362);
and (n1350,n1351,n930);
wire s0n1351,s1n1351,notn1351;
or (n1351,s0n1351,s1n1351);
not(notn1351,n927);
and (s0n1351,notn1351,n1352);
and (s1n1351,n927,n1353);
and (n1354,n1355,n955);
wire s0n1355,s1n1355,notn1355;
or (n1355,s0n1355,s1n1355);
not(notn1355,n927);
and (s0n1355,notn1355,n1356);
and (s1n1355,n927,n1357);
and (n1358,n1359,n965);
wire s0n1359,s1n1359,notn1359;
or (n1359,s0n1359,s1n1359);
not(notn1359,n927);
and (s0n1359,notn1359,n1360);
and (s1n1359,n927,n1361);
and (n1362,n1363,n975);
wire s0n1363,s1n1363,notn1363;
or (n1363,s0n1363,s1n1363);
not(notn1363,n927);
and (s0n1363,notn1363,n1364);
and (s1n1363,n927,n1365);
or (n1366,1'b0,n1367,n1376,n1382,n1391);
and (n1367,n1368,n981);
or (n1368,1'b0,n1369,n1373,n1374,n1375);
and (n1369,n1370,n930);
wire s0n1370,s1n1370,notn1370;
or (n1370,s0n1370,s1n1370);
not(notn1370,n927);
and (s0n1370,notn1370,n1371);
and (s1n1370,n927,n1372);
and (n1373,n1297,n955);
and (n1374,n1301,n965);
and (n1375,n1305,n975);
and (n1376,n1377,n1002);
or (n1377,1'b0,n1378,n1379,n1380,n1381);
and (n1378,n1309,n930);
and (n1379,n1315,n955);
and (n1380,n1319,n965);
and (n1381,n1323,n975);
and (n1382,n1383,n1022);
or (n1383,1'b0,n1384,n1388,n1389,n1390);
and (n1384,n1385,n930);
wire s0n1385,s1n1385,notn1385;
or (n1385,s0n1385,s1n1385);
not(notn1385,n927);
and (s0n1385,notn1385,n1386);
and (s1n1385,n927,n1387);
and (n1388,n1333,n955);
and (n1389,n1337,n965);
and (n1390,n1341,n975);
and (n1391,n1392,n1042);
or (n1392,1'b0,n1393,n1394,n1395,n1396);
and (n1393,n1345,n930);
and (n1394,n1351,n955);
and (n1395,n1355,n965);
and (n1396,n1359,n975);
and (n1397,n1366,n1398);
or (n1398,n1399,n1504,n1826);
and (n1399,n1400,n1473);
or (n1400,1'b0,n1401,n1419,n1437,n1455);
and (n1401,n1402,n981);
or (n1402,1'b0,n1403,n1407,n1411,n1415);
and (n1403,n1404,n930);
wire s0n1404,s1n1404,notn1404;
or (n1404,s0n1404,s1n1404);
not(notn1404,n927);
and (s0n1404,notn1404,n1405);
and (s1n1404,n927,n1406);
and (n1407,n1408,n955);
wire s0n1408,s1n1408,notn1408;
or (n1408,s0n1408,s1n1408);
not(notn1408,n927);
and (s0n1408,notn1408,n1409);
and (s1n1408,n927,n1410);
and (n1411,n1412,n965);
wire s0n1412,s1n1412,notn1412;
or (n1412,s0n1412,s1n1412);
not(notn1412,n927);
and (s0n1412,notn1412,n1413);
and (s1n1412,n927,n1414);
and (n1415,n1416,n975);
wire s0n1416,s1n1416,notn1416;
or (n1416,s0n1416,s1n1416);
not(notn1416,n927);
and (s0n1416,notn1416,n1417);
and (s1n1416,n927,n1418);
and (n1419,n1420,n1002);
or (n1420,1'b0,n1421,n1425,n1429,n1433);
and (n1421,n1422,n930);
wire s0n1422,s1n1422,notn1422;
or (n1422,s0n1422,s1n1422);
not(notn1422,n927);
and (s0n1422,notn1422,n1423);
and (s1n1422,n927,n1424);
and (n1425,n1426,n955);
wire s0n1426,s1n1426,notn1426;
or (n1426,s0n1426,s1n1426);
not(notn1426,n927);
and (s0n1426,notn1426,n1427);
and (s1n1426,n927,n1428);
and (n1429,n1430,n965);
wire s0n1430,s1n1430,notn1430;
or (n1430,s0n1430,s1n1430);
not(notn1430,n927);
and (s0n1430,notn1430,n1431);
and (s1n1430,n927,n1432);
and (n1433,n1434,n975);
wire s0n1434,s1n1434,notn1434;
or (n1434,s0n1434,s1n1434);
not(notn1434,n927);
and (s0n1434,notn1434,n1435);
and (s1n1434,n927,n1436);
and (n1437,n1438,n1022);
or (n1438,1'b0,n1439,n1443,n1447,n1451);
and (n1439,n1440,n930);
wire s0n1440,s1n1440,notn1440;
or (n1440,s0n1440,s1n1440);
not(notn1440,n927);
and (s0n1440,notn1440,n1441);
and (s1n1440,n927,n1442);
and (n1443,n1444,n955);
wire s0n1444,s1n1444,notn1444;
or (n1444,s0n1444,s1n1444);
not(notn1444,n927);
and (s0n1444,notn1444,n1445);
and (s1n1444,n927,n1446);
and (n1447,n1448,n965);
wire s0n1448,s1n1448,notn1448;
or (n1448,s0n1448,s1n1448);
not(notn1448,n927);
and (s0n1448,notn1448,n1449);
and (s1n1448,n927,n1450);
and (n1451,n1452,n975);
wire s0n1452,s1n1452,notn1452;
or (n1452,s0n1452,s1n1452);
not(notn1452,n927);
and (s0n1452,notn1452,n1453);
and (s1n1452,n927,n1454);
and (n1455,n1456,n1042);
or (n1456,1'b0,n1457,n1461,n1465,n1469);
and (n1457,n1458,n930);
wire s0n1458,s1n1458,notn1458;
or (n1458,s0n1458,s1n1458);
not(notn1458,n927);
and (s0n1458,notn1458,n1459);
and (s1n1458,n927,n1460);
and (n1461,n1462,n955);
wire s0n1462,s1n1462,notn1462;
or (n1462,s0n1462,s1n1462);
not(notn1462,n927);
and (s0n1462,notn1462,n1463);
and (s1n1462,n927,n1464);
and (n1465,n1466,n965);
wire s0n1466,s1n1466,notn1466;
or (n1466,s0n1466,s1n1466);
not(notn1466,n927);
and (s0n1466,notn1466,n1467);
and (s1n1466,n927,n1468);
and (n1469,n1470,n975);
wire s0n1470,s1n1470,notn1470;
or (n1470,s0n1470,s1n1470);
not(notn1470,n927);
and (s0n1470,notn1470,n1471);
and (s1n1470,n927,n1472);
or (n1473,1'b0,n1474,n1483,n1489,n1498);
and (n1474,n1475,n981);
or (n1475,1'b0,n1476,n1480,n1481,n1482);
and (n1476,n1477,n930);
wire s0n1477,s1n1477,notn1477;
or (n1477,s0n1477,s1n1477);
not(notn1477,n927);
and (s0n1477,notn1477,n1478);
and (s1n1477,n927,n1479);
and (n1480,n1404,n955);
and (n1481,n1408,n965);
and (n1482,n1412,n975);
and (n1483,n1484,n1002);
or (n1484,1'b0,n1485,n1486,n1487,n1488);
and (n1485,n1416,n930);
and (n1486,n1422,n955);
and (n1487,n1426,n965);
and (n1488,n1430,n975);
and (n1489,n1490,n1022);
or (n1490,1'b0,n1491,n1495,n1496,n1497);
and (n1491,n1492,n930);
wire s0n1492,s1n1492,notn1492;
or (n1492,s0n1492,s1n1492);
not(notn1492,n927);
and (s0n1492,notn1492,n1493);
and (s1n1492,n927,n1494);
and (n1495,n1440,n955);
and (n1496,n1444,n965);
and (n1497,n1448,n975);
and (n1498,n1499,n1042);
or (n1499,1'b0,n1500,n1501,n1502,n1503);
and (n1500,n1452,n930);
and (n1501,n1458,n955);
and (n1502,n1462,n965);
and (n1503,n1466,n975);
and (n1504,n1473,n1505);
or (n1505,n1506,n1611,n1825);
and (n1506,n1507,n1580);
or (n1507,1'b0,n1508,n1526,n1544,n1562);
and (n1508,n1509,n981);
or (n1509,1'b0,n1510,n1514,n1518,n1522);
and (n1510,n1511,n930);
wire s0n1511,s1n1511,notn1511;
or (n1511,s0n1511,s1n1511);
not(notn1511,n927);
and (s0n1511,notn1511,n1512);
and (s1n1511,n927,n1513);
and (n1514,n1515,n955);
wire s0n1515,s1n1515,notn1515;
or (n1515,s0n1515,s1n1515);
not(notn1515,n927);
and (s0n1515,notn1515,n1516);
and (s1n1515,n927,n1517);
and (n1518,n1519,n965);
wire s0n1519,s1n1519,notn1519;
or (n1519,s0n1519,s1n1519);
not(notn1519,n927);
and (s0n1519,notn1519,n1520);
and (s1n1519,n927,n1521);
and (n1522,n1523,n975);
wire s0n1523,s1n1523,notn1523;
or (n1523,s0n1523,s1n1523);
not(notn1523,n927);
and (s0n1523,notn1523,n1524);
and (s1n1523,n927,n1525);
and (n1526,n1527,n1002);
or (n1527,1'b0,n1528,n1532,n1536,n1540);
and (n1528,n1529,n930);
wire s0n1529,s1n1529,notn1529;
or (n1529,s0n1529,s1n1529);
not(notn1529,n927);
and (s0n1529,notn1529,n1530);
and (s1n1529,n927,n1531);
and (n1532,n1533,n955);
wire s0n1533,s1n1533,notn1533;
or (n1533,s0n1533,s1n1533);
not(notn1533,n927);
and (s0n1533,notn1533,n1534);
and (s1n1533,n927,n1535);
and (n1536,n1537,n965);
wire s0n1537,s1n1537,notn1537;
or (n1537,s0n1537,s1n1537);
not(notn1537,n927);
and (s0n1537,notn1537,n1538);
and (s1n1537,n927,n1539);
and (n1540,n1541,n975);
wire s0n1541,s1n1541,notn1541;
or (n1541,s0n1541,s1n1541);
not(notn1541,n927);
and (s0n1541,notn1541,n1542);
and (s1n1541,n927,n1543);
and (n1544,n1545,n1022);
or (n1545,1'b0,n1546,n1550,n1554,n1558);
and (n1546,n1547,n930);
wire s0n1547,s1n1547,notn1547;
or (n1547,s0n1547,s1n1547);
not(notn1547,n927);
and (s0n1547,notn1547,n1548);
and (s1n1547,n927,n1549);
and (n1550,n1551,n955);
wire s0n1551,s1n1551,notn1551;
or (n1551,s0n1551,s1n1551);
not(notn1551,n927);
and (s0n1551,notn1551,n1552);
and (s1n1551,n927,n1553);
and (n1554,n1555,n965);
wire s0n1555,s1n1555,notn1555;
or (n1555,s0n1555,s1n1555);
not(notn1555,n927);
and (s0n1555,notn1555,n1556);
and (s1n1555,n927,n1557);
and (n1558,n1559,n975);
wire s0n1559,s1n1559,notn1559;
or (n1559,s0n1559,s1n1559);
not(notn1559,n927);
and (s0n1559,notn1559,n1560);
and (s1n1559,n927,n1561);
and (n1562,n1563,n1042);
or (n1563,1'b0,n1564,n1568,n1572,n1576);
and (n1564,n1565,n930);
wire s0n1565,s1n1565,notn1565;
or (n1565,s0n1565,s1n1565);
not(notn1565,n927);
and (s0n1565,notn1565,n1566);
and (s1n1565,n927,n1567);
and (n1568,n1569,n955);
wire s0n1569,s1n1569,notn1569;
or (n1569,s0n1569,s1n1569);
not(notn1569,n927);
and (s0n1569,notn1569,n1570);
and (s1n1569,n927,n1571);
and (n1572,n1573,n965);
wire s0n1573,s1n1573,notn1573;
or (n1573,s0n1573,s1n1573);
not(notn1573,n927);
and (s0n1573,notn1573,n1574);
and (s1n1573,n927,n1575);
and (n1576,n1577,n975);
wire s0n1577,s1n1577,notn1577;
or (n1577,s0n1577,s1n1577);
not(notn1577,n927);
and (s0n1577,notn1577,n1578);
and (s1n1577,n927,n1579);
or (n1580,1'b0,n1581,n1590,n1596,n1605);
and (n1581,n1582,n981);
or (n1582,1'b0,n1583,n1587,n1588,n1589);
and (n1583,n1584,n930);
wire s0n1584,s1n1584,notn1584;
or (n1584,s0n1584,s1n1584);
not(notn1584,n927);
and (s0n1584,notn1584,n1585);
and (s1n1584,n927,n1586);
and (n1587,n1511,n955);
and (n1588,n1515,n965);
and (n1589,n1519,n975);
and (n1590,n1591,n1002);
or (n1591,1'b0,n1592,n1593,n1594,n1595);
and (n1592,n1523,n930);
and (n1593,n1529,n955);
and (n1594,n1533,n965);
and (n1595,n1537,n975);
and (n1596,n1597,n1022);
or (n1597,1'b0,n1598,n1602,n1603,n1604);
and (n1598,n1599,n930);
wire s0n1599,s1n1599,notn1599;
or (n1599,s0n1599,s1n1599);
not(notn1599,n927);
and (s0n1599,notn1599,n1600);
and (s1n1599,n927,n1601);
and (n1602,n1547,n955);
and (n1603,n1551,n965);
and (n1604,n1555,n975);
and (n1605,n1606,n1042);
or (n1606,1'b0,n1607,n1608,n1609,n1610);
and (n1607,n1559,n930);
and (n1608,n1565,n955);
and (n1609,n1569,n965);
and (n1610,n1573,n975);
and (n1611,n1580,n1612);
or (n1612,n1613,n1718,n1824);
and (n1613,n1614,n1687);
or (n1614,1'b0,n1615,n1633,n1651,n1669);
and (n1615,n1616,n981);
or (n1616,1'b0,n1617,n1621,n1625,n1629);
and (n1617,n1618,n930);
wire s0n1618,s1n1618,notn1618;
or (n1618,s0n1618,s1n1618);
not(notn1618,n927);
and (s0n1618,notn1618,n1619);
and (s1n1618,n927,n1620);
and (n1621,n1622,n955);
wire s0n1622,s1n1622,notn1622;
or (n1622,s0n1622,s1n1622);
not(notn1622,n927);
and (s0n1622,notn1622,n1623);
and (s1n1622,n927,n1624);
and (n1625,n1626,n965);
wire s0n1626,s1n1626,notn1626;
or (n1626,s0n1626,s1n1626);
not(notn1626,n927);
and (s0n1626,notn1626,n1627);
and (s1n1626,n927,n1628);
and (n1629,n1630,n975);
wire s0n1630,s1n1630,notn1630;
or (n1630,s0n1630,s1n1630);
not(notn1630,n927);
and (s0n1630,notn1630,n1631);
and (s1n1630,n927,n1632);
and (n1633,n1634,n1002);
or (n1634,1'b0,n1635,n1639,n1643,n1647);
and (n1635,n1636,n930);
wire s0n1636,s1n1636,notn1636;
or (n1636,s0n1636,s1n1636);
not(notn1636,n927);
and (s0n1636,notn1636,n1637);
and (s1n1636,n927,n1638);
and (n1639,n1640,n955);
wire s0n1640,s1n1640,notn1640;
or (n1640,s0n1640,s1n1640);
not(notn1640,n927);
and (s0n1640,notn1640,n1641);
and (s1n1640,n927,n1642);
and (n1643,n1644,n965);
wire s0n1644,s1n1644,notn1644;
or (n1644,s0n1644,s1n1644);
not(notn1644,n927);
and (s0n1644,notn1644,n1645);
and (s1n1644,n927,n1646);
and (n1647,n1648,n975);
wire s0n1648,s1n1648,notn1648;
or (n1648,s0n1648,s1n1648);
not(notn1648,n927);
and (s0n1648,notn1648,n1649);
and (s1n1648,n927,n1650);
and (n1651,n1652,n1022);
or (n1652,1'b0,n1653,n1657,n1661,n1665);
and (n1653,n1654,n930);
wire s0n1654,s1n1654,notn1654;
or (n1654,s0n1654,s1n1654);
not(notn1654,n927);
and (s0n1654,notn1654,n1655);
and (s1n1654,n927,n1656);
and (n1657,n1658,n955);
wire s0n1658,s1n1658,notn1658;
or (n1658,s0n1658,s1n1658);
not(notn1658,n927);
and (s0n1658,notn1658,n1659);
and (s1n1658,n927,n1660);
and (n1661,n1662,n965);
wire s0n1662,s1n1662,notn1662;
or (n1662,s0n1662,s1n1662);
not(notn1662,n927);
and (s0n1662,notn1662,n1663);
and (s1n1662,n927,n1664);
and (n1665,n1666,n975);
wire s0n1666,s1n1666,notn1666;
or (n1666,s0n1666,s1n1666);
not(notn1666,n927);
and (s0n1666,notn1666,n1667);
and (s1n1666,n927,n1668);
and (n1669,n1670,n1042);
or (n1670,1'b0,n1671,n1675,n1679,n1683);
and (n1671,n1672,n930);
wire s0n1672,s1n1672,notn1672;
or (n1672,s0n1672,s1n1672);
not(notn1672,n927);
and (s0n1672,notn1672,n1673);
and (s1n1672,n927,n1674);
and (n1675,n1676,n955);
wire s0n1676,s1n1676,notn1676;
or (n1676,s0n1676,s1n1676);
not(notn1676,n927);
and (s0n1676,notn1676,n1677);
and (s1n1676,n927,n1678);
and (n1679,n1680,n965);
wire s0n1680,s1n1680,notn1680;
or (n1680,s0n1680,s1n1680);
not(notn1680,n927);
and (s0n1680,notn1680,n1681);
and (s1n1680,n927,n1682);
and (n1683,n1684,n975);
wire s0n1684,s1n1684,notn1684;
or (n1684,s0n1684,s1n1684);
not(notn1684,n927);
and (s0n1684,notn1684,n1685);
and (s1n1684,n927,n1686);
or (n1687,1'b0,n1688,n1697,n1703,n1712);
and (n1688,n1689,n981);
or (n1689,1'b0,n1690,n1694,n1695,n1696);
and (n1690,n1691,n930);
wire s0n1691,s1n1691,notn1691;
or (n1691,s0n1691,s1n1691);
not(notn1691,n927);
and (s0n1691,notn1691,n1692);
and (s1n1691,n927,n1693);
and (n1694,n1618,n955);
and (n1695,n1622,n965);
and (n1696,n1626,n975);
and (n1697,n1698,n1002);
or (n1698,1'b0,n1699,n1700,n1701,n1702);
and (n1699,n1630,n930);
and (n1700,n1636,n955);
and (n1701,n1640,n965);
and (n1702,n1644,n975);
and (n1703,n1704,n1022);
or (n1704,1'b0,n1705,n1709,n1710,n1711);
and (n1705,n1706,n930);
wire s0n1706,s1n1706,notn1706;
or (n1706,s0n1706,s1n1706);
not(notn1706,n927);
and (s0n1706,notn1706,n1707);
and (s1n1706,n927,n1708);
and (n1709,n1654,n955);
and (n1710,n1658,n965);
and (n1711,n1662,n975);
and (n1712,n1713,n1042);
or (n1713,1'b0,n1714,n1715,n1716,n1717);
and (n1714,n1666,n930);
and (n1715,n1672,n955);
and (n1716,n1676,n965);
and (n1717,n1680,n975);
and (n1718,n1687,n1719);
and (n1719,n1720,n1793);
or (n1720,1'b0,n1721,n1739,n1757,n1775);
and (n1721,n1722,n981);
or (n1722,1'b0,n1723,n1727,n1731,n1735);
and (n1723,n1724,n930);
wire s0n1724,s1n1724,notn1724;
or (n1724,s0n1724,s1n1724);
not(notn1724,n927);
and (s0n1724,notn1724,n1725);
and (s1n1724,n927,n1726);
and (n1727,n1728,n955);
wire s0n1728,s1n1728,notn1728;
or (n1728,s0n1728,s1n1728);
not(notn1728,n927);
and (s0n1728,notn1728,n1729);
and (s1n1728,n927,n1730);
and (n1731,n1732,n965);
wire s0n1732,s1n1732,notn1732;
or (n1732,s0n1732,s1n1732);
not(notn1732,n927);
and (s0n1732,notn1732,n1733);
and (s1n1732,n927,n1734);
and (n1735,n1736,n975);
wire s0n1736,s1n1736,notn1736;
or (n1736,s0n1736,s1n1736);
not(notn1736,n927);
and (s0n1736,notn1736,n1737);
and (s1n1736,n927,n1738);
and (n1739,n1740,n1002);
or (n1740,1'b0,n1741,n1745,n1749,n1753);
and (n1741,n1742,n930);
wire s0n1742,s1n1742,notn1742;
or (n1742,s0n1742,s1n1742);
not(notn1742,n927);
and (s0n1742,notn1742,n1743);
and (s1n1742,n927,n1744);
and (n1745,n1746,n955);
wire s0n1746,s1n1746,notn1746;
or (n1746,s0n1746,s1n1746);
not(notn1746,n927);
and (s0n1746,notn1746,n1747);
and (s1n1746,n927,n1748);
and (n1749,n1750,n965);
wire s0n1750,s1n1750,notn1750;
or (n1750,s0n1750,s1n1750);
not(notn1750,n927);
and (s0n1750,notn1750,n1751);
and (s1n1750,n927,n1752);
and (n1753,n1754,n975);
wire s0n1754,s1n1754,notn1754;
or (n1754,s0n1754,s1n1754);
not(notn1754,n927);
and (s0n1754,notn1754,n1755);
and (s1n1754,n927,n1756);
and (n1757,n1758,n1022);
or (n1758,1'b0,n1759,n1763,n1767,n1771);
and (n1759,n1760,n930);
wire s0n1760,s1n1760,notn1760;
or (n1760,s0n1760,s1n1760);
not(notn1760,n927);
and (s0n1760,notn1760,n1761);
and (s1n1760,n927,n1762);
and (n1763,n1764,n955);
wire s0n1764,s1n1764,notn1764;
or (n1764,s0n1764,s1n1764);
not(notn1764,n927);
and (s0n1764,notn1764,n1765);
and (s1n1764,n927,n1766);
and (n1767,n1768,n965);
wire s0n1768,s1n1768,notn1768;
or (n1768,s0n1768,s1n1768);
not(notn1768,n927);
and (s0n1768,notn1768,n1769);
and (s1n1768,n927,n1770);
and (n1771,n1772,n975);
wire s0n1772,s1n1772,notn1772;
or (n1772,s0n1772,s1n1772);
not(notn1772,n927);
and (s0n1772,notn1772,n1773);
and (s1n1772,n927,n1774);
and (n1775,n1776,n1042);
or (n1776,1'b0,n1777,n1781,n1785,n1789);
and (n1777,n1778,n930);
wire s0n1778,s1n1778,notn1778;
or (n1778,s0n1778,s1n1778);
not(notn1778,n927);
and (s0n1778,notn1778,n1779);
and (s1n1778,n927,n1780);
and (n1781,n1782,n955);
wire s0n1782,s1n1782,notn1782;
or (n1782,s0n1782,s1n1782);
not(notn1782,n927);
and (s0n1782,notn1782,n1783);
and (s1n1782,n927,n1784);
and (n1785,n1786,n965);
wire s0n1786,s1n1786,notn1786;
or (n1786,s0n1786,s1n1786);
not(notn1786,n927);
and (s0n1786,notn1786,n1787);
and (s1n1786,n927,n1788);
and (n1789,n1790,n975);
wire s0n1790,s1n1790,notn1790;
or (n1790,s0n1790,s1n1790);
not(notn1790,n927);
and (s0n1790,notn1790,n1791);
and (s1n1790,n927,n1792);
or (n1793,1'b0,n1794,n1803,n1809,n1818);
and (n1794,n1795,n981);
or (n1795,1'b0,n1796,n1800,n1801,n1802);
and (n1796,n1797,n930);
wire s0n1797,s1n1797,notn1797;
or (n1797,s0n1797,s1n1797);
not(notn1797,n927);
and (s0n1797,notn1797,n1798);
and (s1n1797,n927,n1799);
and (n1800,n1724,n955);
and (n1801,n1728,n965);
and (n1802,n1732,n975);
and (n1803,n1804,n1002);
or (n1804,1'b0,n1805,n1806,n1807,n1808);
and (n1805,n1736,n930);
and (n1806,n1742,n955);
and (n1807,n1746,n965);
and (n1808,n1750,n975);
and (n1809,n1810,n1022);
or (n1810,1'b0,n1811,n1815,n1816,n1817);
and (n1811,n1812,n930);
wire s0n1812,s1n1812,notn1812;
or (n1812,s0n1812,s1n1812);
not(notn1812,n927);
and (s0n1812,notn1812,n1813);
and (s1n1812,n927,n1814);
and (n1815,n1760,n955);
and (n1816,n1764,n965);
and (n1817,n1768,n975);
and (n1818,n1819,n1042);
or (n1819,1'b0,n1820,n1821,n1822,n1823);
and (n1820,n1772,n930);
and (n1821,n1778,n955);
and (n1822,n1782,n965);
and (n1823,n1786,n975);
and (n1824,n1614,n1719);
and (n1825,n1507,n1612);
and (n1826,n1400,n1505);
and (n1827,n1293,n1398);
and (n1828,n1186,n1291);
and (n1829,n1079,n1184);
and (n1830,n920,n1077);
or (n1831,n1832,n1834);
xor (n1832,n1833,n1077);
xor (n1833,n920,n1045);
or (n1834,n1835,n2364,n2415);
and (n1835,n1836,n1838);
xor (n1836,n1837,n1184);
xor (n1837,n1079,n1152);
not (n1838,n1839);
or (n1839,n1840,n1903,n2363);
and (n1840,n1841,n1872);
or (n1841,1'b0,n1842,n1848,n1857,n1863);
and (n1842,n1843,n981);
or (n1843,1'b0,n1844,n1845,n1846,n1847);
and (n1844,n952,n930);
and (n1845,n962,n955);
and (n1846,n972,n965);
and (n1847,n987,n975);
and (n1848,n1849,n1002);
or (n1849,1'b0,n1850,n1851,n1852,n1853);
and (n1850,n991,n930);
and (n1851,n995,n955);
and (n1852,n999,n965);
and (n1853,n1854,n975);
wire s0n1854,s1n1854,notn1854;
or (n1854,s0n1854,s1n1854);
not(notn1854,n927);
and (s0n1854,notn1854,n1855);
and (s1n1854,n927,n1856);
and (n1857,n1858,n1022);
or (n1858,1'b0,n1859,n1860,n1861,n1862);
and (n1859,n1011,n930);
and (n1860,n1015,n955);
and (n1861,n1019,n965);
and (n1862,n1027,n975);
and (n1863,n1864,n1042);
or (n1864,1'b0,n1865,n1866,n1867,n1868);
and (n1865,n1031,n930);
and (n1866,n1035,n955);
and (n1867,n1039,n965);
and (n1868,n1869,n975);
wire s0n1869,s1n1869,notn1869;
or (n1869,s0n1869,s1n1869);
not(notn1869,n927);
and (s0n1869,notn1869,n1870);
and (s1n1869,n927,n1871);
or (n1872,1'b0,n1873,n1882,n1888,n1897);
and (n1873,n1874,n981);
or (n1874,1'b0,n1875,n1879,n1880,n1881);
and (n1875,n1876,n930);
wire s0n1876,s1n1876,notn1876;
or (n1876,s0n1876,s1n1876);
not(notn1876,n927);
and (s0n1876,notn1876,n1877);
and (s1n1876,n927,n1878);
and (n1879,n1049,n955);
and (n1880,n924,n965);
and (n1881,n952,n975);
and (n1882,n1883,n1002);
or (n1883,1'b0,n1884,n1885,n1886,n1887);
and (n1884,n962,n930);
and (n1885,n972,n955);
and (n1886,n987,n965);
and (n1887,n991,n975);
and (n1888,n1889,n1022);
or (n1889,1'b0,n1890,n1894,n1895,n1896);
and (n1890,n1891,n930);
wire s0n1891,s1n1891,notn1891;
or (n1891,s0n1891,s1n1891);
not(notn1891,n927);
and (s0n1891,notn1891,n1892);
and (s1n1891,n927,n1893);
and (n1894,n1064,n955);
and (n1895,n1007,n965);
and (n1896,n1011,n975);
and (n1897,n1898,n1042);
or (n1898,1'b0,n1899,n1900,n1901,n1902);
and (n1899,n1015,n930);
and (n1900,n1019,n955);
and (n1901,n1027,n965);
and (n1902,n1031,n975);
and (n1903,n1872,n1904);
or (n1904,n1905,n1968,n2362);
and (n1905,n1906,n1937);
or (n1906,1'b0,n1907,n1913,n1922,n1928);
and (n1907,n1908,n981);
or (n1908,1'b0,n1909,n1910,n1911,n1912);
and (n1909,n1087,n930);
and (n1910,n1091,n955);
and (n1911,n1095,n965);
and (n1912,n1101,n975);
and (n1913,n1914,n1002);
or (n1914,1'b0,n1915,n1916,n1917,n1918);
and (n1915,n1105,n930);
and (n1916,n1109,n955);
and (n1917,n1113,n965);
and (n1918,n1919,n975);
wire s0n1919,s1n1919,notn1919;
or (n1919,s0n1919,s1n1919);
not(notn1919,n927);
and (s0n1919,notn1919,n1920);
and (s1n1919,n927,n1921);
and (n1922,n1923,n1022);
or (n1923,1'b0,n1924,n1925,n1926,n1927);
and (n1924,n1123,n930);
and (n1925,n1127,n955);
and (n1926,n1131,n965);
and (n1927,n1137,n975);
and (n1928,n1929,n1042);
or (n1929,1'b0,n1930,n1931,n1932,n1933);
and (n1930,n1141,n930);
and (n1931,n1145,n955);
and (n1932,n1149,n965);
and (n1933,n1934,n975);
wire s0n1934,s1n1934,notn1934;
or (n1934,s0n1934,s1n1934);
not(notn1934,n927);
and (s0n1934,notn1934,n1935);
and (s1n1934,n927,n1936);
or (n1937,1'b0,n1938,n1947,n1953,n1962);
and (n1938,n1939,n981);
or (n1939,1'b0,n1940,n1944,n1945,n1946);
and (n1940,n1941,n930);
wire s0n1941,s1n1941,notn1941;
or (n1941,s0n1941,s1n1941);
not(notn1941,n927);
and (s0n1941,notn1941,n1942);
and (s1n1941,n927,n1943);
and (n1944,n1156,n955);
and (n1945,n1083,n965);
and (n1946,n1087,n975);
and (n1947,n1948,n1002);
or (n1948,1'b0,n1949,n1950,n1951,n1952);
and (n1949,n1091,n930);
and (n1950,n1095,n955);
and (n1951,n1101,n965);
and (n1952,n1105,n975);
and (n1953,n1954,n1022);
or (n1954,1'b0,n1955,n1959,n1960,n1961);
and (n1955,n1956,n930);
wire s0n1956,s1n1956,notn1956;
or (n1956,s0n1956,s1n1956);
not(notn1956,n927);
and (s0n1956,notn1956,n1957);
and (s1n1956,n927,n1958);
and (n1959,n1171,n955);
and (n1960,n1119,n965);
and (n1961,n1123,n975);
and (n1962,n1963,n1042);
or (n1963,1'b0,n1964,n1965,n1966,n1967);
and (n1964,n1127,n930);
and (n1965,n1131,n955);
and (n1966,n1137,n965);
and (n1967,n1141,n975);
and (n1968,n1937,n1969);
or (n1969,n1970,n2033,n2361);
and (n1970,n1971,n2002);
or (n1971,1'b0,n1972,n1978,n1987,n1993);
and (n1972,n1973,n981);
or (n1973,1'b0,n1974,n1975,n1976,n1977);
and (n1974,n1194,n930);
and (n1975,n1198,n955);
and (n1976,n1202,n965);
and (n1977,n1208,n975);
and (n1978,n1979,n1002);
or (n1979,1'b0,n1980,n1981,n1982,n1983);
and (n1980,n1212,n930);
and (n1981,n1216,n955);
and (n1982,n1220,n965);
and (n1983,n1984,n975);
wire s0n1984,s1n1984,notn1984;
or (n1984,s0n1984,s1n1984);
not(notn1984,n927);
and (s0n1984,notn1984,n1985);
and (s1n1984,n927,n1986);
and (n1987,n1988,n1022);
or (n1988,1'b0,n1989,n1990,n1991,n1992);
and (n1989,n1230,n930);
and (n1990,n1234,n955);
and (n1991,n1238,n965);
and (n1992,n1244,n975);
and (n1993,n1994,n1042);
or (n1994,1'b0,n1995,n1996,n1997,n1998);
and (n1995,n1248,n930);
and (n1996,n1252,n955);
and (n1997,n1256,n965);
and (n1998,n1999,n975);
wire s0n1999,s1n1999,notn1999;
or (n1999,s0n1999,s1n1999);
not(notn1999,n927);
and (s0n1999,notn1999,n2000);
and (s1n1999,n927,n2001);
or (n2002,1'b0,n2003,n2012,n2018,n2027);
and (n2003,n2004,n981);
or (n2004,1'b0,n2005,n2009,n2010,n2011);
and (n2005,n2006,n930);
wire s0n2006,s1n2006,notn2006;
or (n2006,s0n2006,s1n2006);
not(notn2006,n927);
and (s0n2006,notn2006,n2007);
and (s1n2006,n927,n2008);
and (n2009,n1263,n955);
and (n2010,n1190,n965);
and (n2011,n1194,n975);
and (n2012,n2013,n1002);
or (n2013,1'b0,n2014,n2015,n2016,n2017);
and (n2014,n1198,n930);
and (n2015,n1202,n955);
and (n2016,n1208,n965);
and (n2017,n1212,n975);
and (n2018,n2019,n1022);
or (n2019,1'b0,n2020,n2024,n2025,n2026);
and (n2020,n2021,n930);
wire s0n2021,s1n2021,notn2021;
or (n2021,s0n2021,s1n2021);
not(notn2021,n927);
and (s0n2021,notn2021,n2022);
and (s1n2021,n927,n2023);
and (n2024,n1278,n955);
and (n2025,n1226,n965);
and (n2026,n1230,n975);
and (n2027,n2028,n1042);
or (n2028,1'b0,n2029,n2030,n2031,n2032);
and (n2029,n1234,n930);
and (n2030,n1238,n955);
and (n2031,n1244,n965);
and (n2032,n1248,n975);
and (n2033,n2002,n2034);
or (n2034,n2035,n2098,n2360);
and (n2035,n2036,n2067);
or (n2036,1'b0,n2037,n2043,n2052,n2058);
and (n2037,n2038,n981);
or (n2038,1'b0,n2039,n2040,n2041,n2042);
and (n2039,n1301,n930);
and (n2040,n1305,n955);
and (n2041,n1309,n965);
and (n2042,n1315,n975);
and (n2043,n2044,n1002);
or (n2044,1'b0,n2045,n2046,n2047,n2048);
and (n2045,n1319,n930);
and (n2046,n1323,n955);
and (n2047,n1327,n965);
and (n2048,n2049,n975);
wire s0n2049,s1n2049,notn2049;
or (n2049,s0n2049,s1n2049);
not(notn2049,n927);
and (s0n2049,notn2049,n2050);
and (s1n2049,n927,n2051);
and (n2052,n2053,n1022);
or (n2053,1'b0,n2054,n2055,n2056,n2057);
and (n2054,n1337,n930);
and (n2055,n1341,n955);
and (n2056,n1345,n965);
and (n2057,n1351,n975);
and (n2058,n2059,n1042);
or (n2059,1'b0,n2060,n2061,n2062,n2063);
and (n2060,n1355,n930);
and (n2061,n1359,n955);
and (n2062,n1363,n965);
and (n2063,n2064,n975);
wire s0n2064,s1n2064,notn2064;
or (n2064,s0n2064,s1n2064);
not(notn2064,n927);
and (s0n2064,notn2064,n2065);
and (s1n2064,n927,n2066);
or (n2067,1'b0,n2068,n2077,n2083,n2092);
and (n2068,n2069,n981);
or (n2069,1'b0,n2070,n2074,n2075,n2076);
and (n2070,n2071,n930);
wire s0n2071,s1n2071,notn2071;
or (n2071,s0n2071,s1n2071);
not(notn2071,n927);
and (s0n2071,notn2071,n2072);
and (s1n2071,n927,n2073);
and (n2074,n1370,n955);
and (n2075,n1297,n965);
and (n2076,n1301,n975);
and (n2077,n2078,n1002);
or (n2078,1'b0,n2079,n2080,n2081,n2082);
and (n2079,n1305,n930);
and (n2080,n1309,n955);
and (n2081,n1315,n965);
and (n2082,n1319,n975);
and (n2083,n2084,n1022);
or (n2084,1'b0,n2085,n2089,n2090,n2091);
and (n2085,n2086,n930);
wire s0n2086,s1n2086,notn2086;
or (n2086,s0n2086,s1n2086);
not(notn2086,n927);
and (s0n2086,notn2086,n2087);
and (s1n2086,n927,n2088);
and (n2089,n1385,n955);
and (n2090,n1333,n965);
and (n2091,n1337,n975);
and (n2092,n2093,n1042);
or (n2093,1'b0,n2094,n2095,n2096,n2097);
and (n2094,n1341,n930);
and (n2095,n1345,n955);
and (n2096,n1351,n965);
and (n2097,n1355,n975);
and (n2098,n2067,n2099);
or (n2099,n2100,n2163,n2359);
and (n2100,n2101,n2132);
or (n2101,1'b0,n2102,n2108,n2117,n2123);
and (n2102,n2103,n981);
or (n2103,1'b0,n2104,n2105,n2106,n2107);
and (n2104,n1408,n930);
and (n2105,n1412,n955);
and (n2106,n1416,n965);
and (n2107,n1422,n975);
and (n2108,n2109,n1002);
or (n2109,1'b0,n2110,n2111,n2112,n2113);
and (n2110,n1426,n930);
and (n2111,n1430,n955);
and (n2112,n1434,n965);
and (n2113,n2114,n975);
wire s0n2114,s1n2114,notn2114;
or (n2114,s0n2114,s1n2114);
not(notn2114,n927);
and (s0n2114,notn2114,n2115);
and (s1n2114,n927,n2116);
and (n2117,n2118,n1022);
or (n2118,1'b0,n2119,n2120,n2121,n2122);
and (n2119,n1444,n930);
and (n2120,n1448,n955);
and (n2121,n1452,n965);
and (n2122,n1458,n975);
and (n2123,n2124,n1042);
or (n2124,1'b0,n2125,n2126,n2127,n2128);
and (n2125,n1462,n930);
and (n2126,n1466,n955);
and (n2127,n1470,n965);
and (n2128,n2129,n975);
wire s0n2129,s1n2129,notn2129;
or (n2129,s0n2129,s1n2129);
not(notn2129,n927);
and (s0n2129,notn2129,n2130);
and (s1n2129,n927,n2131);
or (n2132,1'b0,n2133,n2142,n2148,n2157);
and (n2133,n2134,n981);
or (n2134,1'b0,n2135,n2139,n2140,n2141);
and (n2135,n2136,n930);
wire s0n2136,s1n2136,notn2136;
or (n2136,s0n2136,s1n2136);
not(notn2136,n927);
and (s0n2136,notn2136,n2137);
and (s1n2136,n927,n2138);
and (n2139,n1477,n955);
and (n2140,n1404,n965);
and (n2141,n1408,n975);
and (n2142,n2143,n1002);
or (n2143,1'b0,n2144,n2145,n2146,n2147);
and (n2144,n1412,n930);
and (n2145,n1416,n955);
and (n2146,n1422,n965);
and (n2147,n1426,n975);
and (n2148,n2149,n1022);
or (n2149,1'b0,n2150,n2154,n2155,n2156);
and (n2150,n2151,n930);
wire s0n2151,s1n2151,notn2151;
or (n2151,s0n2151,s1n2151);
not(notn2151,n927);
and (s0n2151,notn2151,n2152);
and (s1n2151,n927,n2153);
and (n2154,n1492,n955);
and (n2155,n1440,n965);
and (n2156,n1444,n975);
and (n2157,n2158,n1042);
or (n2158,1'b0,n2159,n2160,n2161,n2162);
and (n2159,n1448,n930);
and (n2160,n1452,n955);
and (n2161,n1458,n965);
and (n2162,n1462,n975);
and (n2163,n2132,n2164);
or (n2164,n2165,n2228,n2358);
and (n2165,n2166,n2197);
or (n2166,1'b0,n2167,n2173,n2182,n2188);
and (n2167,n2168,n981);
or (n2168,1'b0,n2169,n2170,n2171,n2172);
and (n2169,n1515,n930);
and (n2170,n1519,n955);
and (n2171,n1523,n965);
and (n2172,n1529,n975);
and (n2173,n2174,n1002);
or (n2174,1'b0,n2175,n2176,n2177,n2178);
and (n2175,n1533,n930);
and (n2176,n1537,n955);
and (n2177,n1541,n965);
and (n2178,n2179,n975);
wire s0n2179,s1n2179,notn2179;
or (n2179,s0n2179,s1n2179);
not(notn2179,n927);
and (s0n2179,notn2179,n2180);
and (s1n2179,n927,n2181);
and (n2182,n2183,n1022);
or (n2183,1'b0,n2184,n2185,n2186,n2187);
and (n2184,n1551,n930);
and (n2185,n1555,n955);
and (n2186,n1559,n965);
and (n2187,n1565,n975);
and (n2188,n2189,n1042);
or (n2189,1'b0,n2190,n2191,n2192,n2193);
and (n2190,n1569,n930);
and (n2191,n1573,n955);
and (n2192,n1577,n965);
and (n2193,n2194,n975);
wire s0n2194,s1n2194,notn2194;
or (n2194,s0n2194,s1n2194);
not(notn2194,n927);
and (s0n2194,notn2194,n2195);
and (s1n2194,n927,n2196);
or (n2197,1'b0,n2198,n2207,n2213,n2222);
and (n2198,n2199,n981);
or (n2199,1'b0,n2200,n2204,n2205,n2206);
and (n2200,n2201,n930);
wire s0n2201,s1n2201,notn2201;
or (n2201,s0n2201,s1n2201);
not(notn2201,n927);
and (s0n2201,notn2201,n2202);
and (s1n2201,n927,n2203);
and (n2204,n1584,n955);
and (n2205,n1511,n965);
and (n2206,n1515,n975);
and (n2207,n2208,n1002);
or (n2208,1'b0,n2209,n2210,n2211,n2212);
and (n2209,n1519,n930);
and (n2210,n1523,n955);
and (n2211,n1529,n965);
and (n2212,n1533,n975);
and (n2213,n2214,n1022);
or (n2214,1'b0,n2215,n2219,n2220,n2221);
and (n2215,n2216,n930);
wire s0n2216,s1n2216,notn2216;
or (n2216,s0n2216,s1n2216);
not(notn2216,n927);
and (s0n2216,notn2216,n2217);
and (s1n2216,n927,n2218);
and (n2219,n1599,n955);
and (n2220,n1547,n965);
and (n2221,n1551,n975);
and (n2222,n2223,n1042);
or (n2223,1'b0,n2224,n2225,n2226,n2227);
and (n2224,n1555,n930);
and (n2225,n1559,n955);
and (n2226,n1565,n965);
and (n2227,n1569,n975);
and (n2228,n2197,n2229);
or (n2229,n2230,n2293,n2357);
and (n2230,n2231,n2262);
or (n2231,1'b0,n2232,n2238,n2247,n2253);
and (n2232,n2233,n981);
or (n2233,1'b0,n2234,n2235,n2236,n2237);
and (n2234,n1622,n930);
and (n2235,n1626,n955);
and (n2236,n1630,n965);
and (n2237,n1636,n975);
and (n2238,n2239,n1002);
or (n2239,1'b0,n2240,n2241,n2242,n2243);
and (n2240,n1640,n930);
and (n2241,n1644,n955);
and (n2242,n1648,n965);
and (n2243,n2244,n975);
wire s0n2244,s1n2244,notn2244;
or (n2244,s0n2244,s1n2244);
not(notn2244,n927);
and (s0n2244,notn2244,n2245);
and (s1n2244,n927,n2246);
and (n2247,n2248,n1022);
or (n2248,1'b0,n2249,n2250,n2251,n2252);
and (n2249,n1658,n930);
and (n2250,n1662,n955);
and (n2251,n1666,n965);
and (n2252,n1672,n975);
and (n2253,n2254,n1042);
or (n2254,1'b0,n2255,n2256,n2257,n2258);
and (n2255,n1676,n930);
and (n2256,n1680,n955);
and (n2257,n1684,n965);
and (n2258,n2259,n975);
wire s0n2259,s1n2259,notn2259;
or (n2259,s0n2259,s1n2259);
not(notn2259,n927);
and (s0n2259,notn2259,n2260);
and (s1n2259,n927,n2261);
or (n2262,1'b0,n2263,n2272,n2278,n2287);
and (n2263,n2264,n981);
or (n2264,1'b0,n2265,n2269,n2270,n2271);
and (n2265,n2266,n930);
wire s0n2266,s1n2266,notn2266;
or (n2266,s0n2266,s1n2266);
not(notn2266,n927);
and (s0n2266,notn2266,n2267);
and (s1n2266,n927,n2268);
and (n2269,n1691,n955);
and (n2270,n1618,n965);
and (n2271,n1622,n975);
and (n2272,n2273,n1002);
or (n2273,1'b0,n2274,n2275,n2276,n2277);
and (n2274,n1626,n930);
and (n2275,n1630,n955);
and (n2276,n1636,n965);
and (n2277,n1640,n975);
and (n2278,n2279,n1022);
or (n2279,1'b0,n2280,n2284,n2285,n2286);
and (n2280,n2281,n930);
wire s0n2281,s1n2281,notn2281;
or (n2281,s0n2281,s1n2281);
not(notn2281,n927);
and (s0n2281,notn2281,n2282);
and (s1n2281,n927,n2283);
and (n2284,n1706,n955);
and (n2285,n1654,n965);
and (n2286,n1658,n975);
and (n2287,n2288,n1042);
or (n2288,1'b0,n2289,n2290,n2291,n2292);
and (n2289,n1662,n930);
and (n2290,n1666,n955);
and (n2291,n1672,n965);
and (n2292,n1676,n975);
and (n2293,n2262,n2294);
and (n2294,n2295,n2326);
or (n2295,1'b0,n2296,n2302,n2311,n2317);
and (n2296,n2297,n981);
or (n2297,1'b0,n2298,n2299,n2300,n2301);
and (n2298,n1728,n930);
and (n2299,n1732,n955);
and (n2300,n1736,n965);
and (n2301,n1742,n975);
and (n2302,n2303,n1002);
or (n2303,1'b0,n2304,n2305,n2306,n2307);
and (n2304,n1746,n930);
and (n2305,n1750,n955);
and (n2306,n1754,n965);
and (n2307,n2308,n975);
wire s0n2308,s1n2308,notn2308;
or (n2308,s0n2308,s1n2308);
not(notn2308,n927);
and (s0n2308,notn2308,n2309);
and (s1n2308,n927,n2310);
and (n2311,n2312,n1022);
or (n2312,1'b0,n2313,n2314,n2315,n2316);
and (n2313,n1764,n930);
and (n2314,n1768,n955);
and (n2315,n1772,n965);
and (n2316,n1778,n975);
and (n2317,n2318,n1042);
or (n2318,1'b0,n2319,n2320,n2321,n2322);
and (n2319,n1782,n930);
and (n2320,n1786,n955);
and (n2321,n1790,n965);
and (n2322,n2323,n975);
wire s0n2323,s1n2323,notn2323;
or (n2323,s0n2323,s1n2323);
not(notn2323,n927);
and (s0n2323,notn2323,n2324);
and (s1n2323,n927,n2325);
or (n2326,1'b0,n2327,n2336,n2342,n2351);
and (n2327,n2328,n981);
or (n2328,1'b0,n2329,n2333,n2334,n2335);
and (n2329,n2330,n930);
wire s0n2330,s1n2330,notn2330;
or (n2330,s0n2330,s1n2330);
not(notn2330,n927);
and (s0n2330,notn2330,n2331);
and (s1n2330,n927,n2332);
and (n2333,n1797,n955);
and (n2334,n1724,n965);
and (n2335,n1728,n975);
and (n2336,n2337,n1002);
or (n2337,1'b0,n2338,n2339,n2340,n2341);
and (n2338,n1732,n930);
and (n2339,n1736,n955);
and (n2340,n1742,n965);
and (n2341,n1746,n975);
and (n2342,n2343,n1022);
or (n2343,1'b0,n2344,n2348,n2349,n2350);
and (n2344,n2345,n930);
wire s0n2345,s1n2345,notn2345;
or (n2345,s0n2345,s1n2345);
not(notn2345,n927);
and (s0n2345,notn2345,n2346);
and (s1n2345,n927,n2347);
and (n2348,n1812,n955);
and (n2349,n1760,n965);
and (n2350,n1764,n975);
and (n2351,n2352,n1042);
or (n2352,1'b0,n2353,n2354,n2355,n2356);
and (n2353,n1768,n930);
and (n2354,n1772,n955);
and (n2355,n1778,n965);
and (n2356,n1782,n975);
and (n2357,n2231,n2294);
and (n2358,n2166,n2229);
and (n2359,n2101,n2164);
and (n2360,n2036,n2099);
and (n2361,n1971,n2034);
and (n2362,n1906,n1969);
and (n2363,n1841,n1904);
and (n2364,n1838,n2365);
or (n2365,n2366,n2372,n2414);
and (n2366,n2367,n2369);
xor (n2367,n2368,n1291);
xor (n2368,n1186,n1259);
not (n2369,n2370);
xor (n2370,n2371,n1904);
xor (n2371,n1841,n1872);
and (n2372,n2369,n2373);
or (n2373,n2374,n2380,n2413);
and (n2374,n2375,n2377);
xor (n2375,n2376,n1398);
xor (n2376,n1293,n1366);
not (n2377,n2378);
xor (n2378,n2379,n1969);
xor (n2379,n1906,n1937);
and (n2380,n2377,n2381);
or (n2381,n2382,n2388,n2412);
and (n2382,n2383,n2385);
xor (n2383,n2384,n1505);
xor (n2384,n1400,n1473);
not (n2385,n2386);
xor (n2386,n2387,n2034);
xor (n2387,n1971,n2002);
and (n2388,n2385,n2389);
or (n2389,n2390,n2396,n2411);
and (n2390,n2391,n2393);
xor (n2391,n2392,n1612);
xor (n2392,n1507,n1580);
not (n2393,n2394);
xor (n2394,n2395,n2099);
xor (n2395,n2036,n2067);
and (n2396,n2393,n2397);
or (n2397,n2398,n2404,n2410);
and (n2398,n2399,n2401);
xor (n2399,n2400,n1719);
xor (n2400,n1614,n1687);
not (n2401,n2402);
xor (n2402,n2403,n2164);
xor (n2403,n2101,n2132);
and (n2404,n2401,n2405);
and (n2405,n2406,n2407);
xor (n2406,n1720,n1793);
not (n2407,n2408);
xor (n2408,n2409,n2229);
xor (n2409,n2166,n2197);
and (n2410,n2399,n2405);
and (n2411,n2391,n2397);
and (n2412,n2383,n2389);
and (n2413,n2375,n2381);
and (n2414,n2367,n2373);
and (n2415,n1836,n2365);
and (n2416,n2417,n2418);
xnor (n2417,n918,n1831);
and (n2418,n2419,n2420);
xnor (n2419,n1832,n1834);
and (n2420,n2421,n2423);
xor (n2421,n2422,n2365);
xor (n2422,n1836,n1838);
and (n2423,n2424,n2426);
xor (n2424,n2425,n2373);
xor (n2425,n2367,n2369);
and (n2426,n2427,n2429);
xor (n2427,n2428,n2381);
xor (n2428,n2375,n2377);
and (n2429,n2430,n2432);
xor (n2430,n2431,n2389);
xor (n2431,n2383,n2385);
and (n2432,n2433,n2435);
xor (n2433,n2434,n2397);
xor (n2434,n2391,n2393);
and (n2435,n2436,n2438);
xor (n2436,n2437,n2405);
xor (n2437,n2399,n2401);
and (n2438,n2439,n2440);
xor (n2439,n2406,n2407);
and (n2440,n2441,n2444);
not (n2441,n2442);
xor (n2442,n2443,n2294);
xor (n2443,n2231,n2262);
not (n2444,n2445);
xor (n2445,n2295,n2326);
and (n2446,n915,n2447);
and (n2447,n2448,n2449);
xor (n2448,n2417,n2418);
and (n2449,n2450,n2451);
xor (n2450,n2419,n2420);
or (n2451,n2452,n2819,n2871);
and (n2452,n2453,n2818);
or (n2453,n2454,n2497,n2817);
and (n2454,n2455,n2476);
or (n2455,1'b0,n2456,n2457,n2466,n2467);
and (n2456,n1883,n981);
and (n2457,n2458,n1002);
or (n2458,1'b0,n2459,n2460,n2461,n2462);
and (n2459,n995,n930);
and (n2460,n999,n955);
and (n2461,n1854,n965);
and (n2462,n2463,n975);
wire s0n2463,s1n2463,notn2463;
or (n2463,s0n2463,s1n2463);
not(notn2463,n927);
and (s0n2463,notn2463,n2464);
and (s1n2463,n927,n2465);
and (n2466,n1898,n1022);
and (n2467,n2468,n1042);
or (n2468,1'b0,n2469,n2470,n2471,n2472);
and (n2469,n1035,n930);
and (n2470,n1039,n955);
and (n2471,n1869,n965);
and (n2472,n2473,n975);
wire s0n2473,s1n2473,notn2473;
or (n2473,s0n2473,s1n2473);
not(notn2473,n927);
and (s0n2473,notn2473,n2474);
and (s1n2473,n927,n2475);
or (n2476,1'b0,n2477,n2486,n2487,n2496);
and (n2477,n2478,n981);
or (n2478,1'b0,n2479,n2483,n2484,n2485);
and (n2479,n2480,n930);
wire s0n2480,s1n2480,notn2480;
or (n2480,s0n2480,s1n2480);
not(notn2480,n927);
and (s0n2480,notn2480,n2481);
and (s1n2480,n927,n2482);
and (n2483,n1876,n955);
and (n2484,n1049,n965);
and (n2485,n924,n975);
and (n2486,n1843,n1002);
and (n2487,n2488,n1022);
or (n2488,1'b0,n2489,n2493,n2494,n2495);
and (n2489,n2490,n930);
wire s0n2490,s1n2490,notn2490;
or (n2490,s0n2490,s1n2490);
not(notn2490,n927);
and (s0n2490,notn2490,n2491);
and (s1n2490,n927,n2492);
and (n2493,n1891,n955);
and (n2494,n1064,n965);
and (n2495,n1007,n975);
and (n2496,n1858,n1042);
and (n2497,n2476,n2498);
or (n2498,n2499,n2542,n2816);
and (n2499,n2500,n2521);
or (n2500,1'b0,n2501,n2502,n2511,n2512);
and (n2501,n1948,n981);
and (n2502,n2503,n1002);
or (n2503,1'b0,n2504,n2505,n2506,n2507);
and (n2504,n1109,n930);
and (n2505,n1113,n955);
and (n2506,n1919,n965);
and (n2507,n2508,n975);
wire s0n2508,s1n2508,notn2508;
or (n2508,s0n2508,s1n2508);
not(notn2508,n927);
and (s0n2508,notn2508,n2509);
and (s1n2508,n927,n2510);
and (n2511,n1963,n1022);
and (n2512,n2513,n1042);
or (n2513,1'b0,n2514,n2515,n2516,n2517);
and (n2514,n1145,n930);
and (n2515,n1149,n955);
and (n2516,n1934,n965);
and (n2517,n2518,n975);
wire s0n2518,s1n2518,notn2518;
or (n2518,s0n2518,s1n2518);
not(notn2518,n927);
and (s0n2518,notn2518,n2519);
and (s1n2518,n927,n2520);
or (n2521,1'b0,n2522,n2531,n2532,n2541);
and (n2522,n2523,n981);
or (n2523,1'b0,n2524,n2528,n2529,n2530);
and (n2524,n2525,n930);
wire s0n2525,s1n2525,notn2525;
or (n2525,s0n2525,s1n2525);
not(notn2525,n927);
and (s0n2525,notn2525,n2526);
and (s1n2525,n927,n2527);
and (n2528,n1941,n955);
and (n2529,n1156,n965);
and (n2530,n1083,n975);
and (n2531,n1908,n1002);
and (n2532,n2533,n1022);
or (n2533,1'b0,n2534,n2538,n2539,n2540);
and (n2534,n2535,n930);
wire s0n2535,s1n2535,notn2535;
or (n2535,s0n2535,s1n2535);
not(notn2535,n927);
and (s0n2535,notn2535,n2536);
and (s1n2535,n927,n2537);
and (n2538,n1956,n955);
and (n2539,n1171,n965);
and (n2540,n1119,n975);
and (n2541,n1923,n1042);
and (n2542,n2521,n2543);
or (n2543,n2544,n2587,n2815);
and (n2544,n2545,n2566);
or (n2545,1'b0,n2546,n2547,n2556,n2557);
and (n2546,n2013,n981);
and (n2547,n2548,n1002);
or (n2548,1'b0,n2549,n2550,n2551,n2552);
and (n2549,n1216,n930);
and (n2550,n1220,n955);
and (n2551,n1984,n965);
and (n2552,n2553,n975);
wire s0n2553,s1n2553,notn2553;
or (n2553,s0n2553,s1n2553);
not(notn2553,n927);
and (s0n2553,notn2553,n2554);
and (s1n2553,n927,n2555);
and (n2556,n2028,n1022);
and (n2557,n2558,n1042);
or (n2558,1'b0,n2559,n2560,n2561,n2562);
and (n2559,n1252,n930);
and (n2560,n1256,n955);
and (n2561,n1999,n965);
and (n2562,n2563,n975);
wire s0n2563,s1n2563,notn2563;
or (n2563,s0n2563,s1n2563);
not(notn2563,n927);
and (s0n2563,notn2563,n2564);
and (s1n2563,n927,n2565);
or (n2566,1'b0,n2567,n2576,n2577,n2586);
and (n2567,n2568,n981);
or (n2568,1'b0,n2569,n2573,n2574,n2575);
and (n2569,n2570,n930);
wire s0n2570,s1n2570,notn2570;
or (n2570,s0n2570,s1n2570);
not(notn2570,n927);
and (s0n2570,notn2570,n2571);
and (s1n2570,n927,n2572);
and (n2573,n2006,n955);
and (n2574,n1263,n965);
and (n2575,n1190,n975);
and (n2576,n1973,n1002);
and (n2577,n2578,n1022);
or (n2578,1'b0,n2579,n2583,n2584,n2585);
and (n2579,n2580,n930);
wire s0n2580,s1n2580,notn2580;
or (n2580,s0n2580,s1n2580);
not(notn2580,n927);
and (s0n2580,notn2580,n2581);
and (s1n2580,n927,n2582);
and (n2583,n2021,n955);
and (n2584,n1278,n965);
and (n2585,n1226,n975);
and (n2586,n1988,n1042);
and (n2587,n2566,n2588);
or (n2588,n2589,n2632,n2814);
and (n2589,n2590,n2611);
or (n2590,1'b0,n2591,n2592,n2601,n2602);
and (n2591,n2078,n981);
and (n2592,n2593,n1002);
or (n2593,1'b0,n2594,n2595,n2596,n2597);
and (n2594,n1323,n930);
and (n2595,n1327,n955);
and (n2596,n2049,n965);
and (n2597,n2598,n975);
wire s0n2598,s1n2598,notn2598;
or (n2598,s0n2598,s1n2598);
not(notn2598,n927);
and (s0n2598,notn2598,n2599);
and (s1n2598,n927,n2600);
and (n2601,n2093,n1022);
and (n2602,n2603,n1042);
or (n2603,1'b0,n2604,n2605,n2606,n2607);
and (n2604,n1359,n930);
and (n2605,n1363,n955);
and (n2606,n2064,n965);
and (n2607,n2608,n975);
wire s0n2608,s1n2608,notn2608;
or (n2608,s0n2608,s1n2608);
not(notn2608,n927);
and (s0n2608,notn2608,n2609);
and (s1n2608,n927,n2610);
or (n2611,1'b0,n2612,n2621,n2622,n2631);
and (n2612,n2613,n981);
or (n2613,1'b0,n2614,n2618,n2619,n2620);
and (n2614,n2615,n930);
wire s0n2615,s1n2615,notn2615;
or (n2615,s0n2615,s1n2615);
not(notn2615,n927);
and (s0n2615,notn2615,n2616);
and (s1n2615,n927,n2617);
and (n2618,n2071,n955);
and (n2619,n1370,n965);
and (n2620,n1297,n975);
and (n2621,n2038,n1002);
and (n2622,n2623,n1022);
or (n2623,1'b0,n2624,n2628,n2629,n2630);
and (n2624,n2625,n930);
wire s0n2625,s1n2625,notn2625;
or (n2625,s0n2625,s1n2625);
not(notn2625,n927);
and (s0n2625,notn2625,n2626);
and (s1n2625,n927,n2627);
and (n2628,n2086,n955);
and (n2629,n1385,n965);
and (n2630,n1333,n975);
and (n2631,n2053,n1042);
and (n2632,n2611,n2633);
or (n2633,n2634,n2677,n2813);
and (n2634,n2635,n2656);
or (n2635,1'b0,n2636,n2637,n2646,n2647);
and (n2636,n2143,n981);
and (n2637,n2638,n1002);
or (n2638,1'b0,n2639,n2640,n2641,n2642);
and (n2639,n1430,n930);
and (n2640,n1434,n955);
and (n2641,n2114,n965);
and (n2642,n2643,n975);
wire s0n2643,s1n2643,notn2643;
or (n2643,s0n2643,s1n2643);
not(notn2643,n927);
and (s0n2643,notn2643,n2644);
and (s1n2643,n927,n2645);
and (n2646,n2158,n1022);
and (n2647,n2648,n1042);
or (n2648,1'b0,n2649,n2650,n2651,n2652);
and (n2649,n1466,n930);
and (n2650,n1470,n955);
and (n2651,n2129,n965);
and (n2652,n2653,n975);
wire s0n2653,s1n2653,notn2653;
or (n2653,s0n2653,s1n2653);
not(notn2653,n927);
and (s0n2653,notn2653,n2654);
and (s1n2653,n927,n2655);
or (n2656,1'b0,n2657,n2666,n2667,n2676);
and (n2657,n2658,n981);
or (n2658,1'b0,n2659,n2663,n2664,n2665);
and (n2659,n2660,n930);
wire s0n2660,s1n2660,notn2660;
or (n2660,s0n2660,s1n2660);
not(notn2660,n927);
and (s0n2660,notn2660,n2661);
and (s1n2660,n927,n2662);
and (n2663,n2136,n955);
and (n2664,n1477,n965);
and (n2665,n1404,n975);
and (n2666,n2103,n1002);
and (n2667,n2668,n1022);
or (n2668,1'b0,n2669,n2673,n2674,n2675);
and (n2669,n2670,n930);
wire s0n2670,s1n2670,notn2670;
or (n2670,s0n2670,s1n2670);
not(notn2670,n927);
and (s0n2670,notn2670,n2671);
and (s1n2670,n927,n2672);
and (n2673,n2151,n955);
and (n2674,n1492,n965);
and (n2675,n1440,n975);
and (n2676,n2118,n1042);
and (n2677,n2656,n2678);
or (n2678,n2679,n2722,n2812);
and (n2679,n2680,n2701);
or (n2680,1'b0,n2681,n2682,n2691,n2692);
and (n2681,n2208,n981);
and (n2682,n2683,n1002);
or (n2683,1'b0,n2684,n2685,n2686,n2687);
and (n2684,n1537,n930);
and (n2685,n1541,n955);
and (n2686,n2179,n965);
and (n2687,n2688,n975);
wire s0n2688,s1n2688,notn2688;
or (n2688,s0n2688,s1n2688);
not(notn2688,n927);
and (s0n2688,notn2688,n2689);
and (s1n2688,n927,n2690);
and (n2691,n2223,n1022);
and (n2692,n2693,n1042);
or (n2693,1'b0,n2694,n2695,n2696,n2697);
and (n2694,n1573,n930);
and (n2695,n1577,n955);
and (n2696,n2194,n965);
and (n2697,n2698,n975);
wire s0n2698,s1n2698,notn2698;
or (n2698,s0n2698,s1n2698);
not(notn2698,n927);
and (s0n2698,notn2698,n2699);
and (s1n2698,n927,n2700);
or (n2701,1'b0,n2702,n2711,n2712,n2721);
and (n2702,n2703,n981);
or (n2703,1'b0,n2704,n2708,n2709,n2710);
and (n2704,n2705,n930);
wire s0n2705,s1n2705,notn2705;
or (n2705,s0n2705,s1n2705);
not(notn2705,n927);
and (s0n2705,notn2705,n2706);
and (s1n2705,n927,n2707);
and (n2708,n2201,n955);
and (n2709,n1584,n965);
and (n2710,n1511,n975);
and (n2711,n2168,n1002);
and (n2712,n2713,n1022);
or (n2713,1'b0,n2714,n2718,n2719,n2720);
and (n2714,n2715,n930);
wire s0n2715,s1n2715,notn2715;
or (n2715,s0n2715,s1n2715);
not(notn2715,n927);
and (s0n2715,notn2715,n2716);
and (s1n2715,n927,n2717);
and (n2718,n2216,n955);
and (n2719,n1599,n965);
and (n2720,n1547,n975);
and (n2721,n2183,n1042);
and (n2722,n2701,n2723);
or (n2723,n2724,n2767,n2811);
and (n2724,n2725,n2746);
or (n2725,1'b0,n2726,n2727,n2736,n2737);
and (n2726,n2273,n981);
and (n2727,n2728,n1002);
or (n2728,1'b0,n2729,n2730,n2731,n2732);
and (n2729,n1644,n930);
and (n2730,n1648,n955);
and (n2731,n2244,n965);
and (n2732,n2733,n975);
wire s0n2733,s1n2733,notn2733;
or (n2733,s0n2733,s1n2733);
not(notn2733,n927);
and (s0n2733,notn2733,n2734);
and (s1n2733,n927,n2735);
and (n2736,n2288,n1022);
and (n2737,n2738,n1042);
or (n2738,1'b0,n2739,n2740,n2741,n2742);
and (n2739,n1680,n930);
and (n2740,n1684,n955);
and (n2741,n2259,n965);
and (n2742,n2743,n975);
wire s0n2743,s1n2743,notn2743;
or (n2743,s0n2743,s1n2743);
not(notn2743,n927);
and (s0n2743,notn2743,n2744);
and (s1n2743,n927,n2745);
or (n2746,1'b0,n2747,n2756,n2757,n2766);
and (n2747,n2748,n981);
or (n2748,1'b0,n2749,n2753,n2754,n2755);
and (n2749,n2750,n930);
wire s0n2750,s1n2750,notn2750;
or (n2750,s0n2750,s1n2750);
not(notn2750,n927);
and (s0n2750,notn2750,n2751);
and (s1n2750,n927,n2752);
and (n2753,n2266,n955);
and (n2754,n1691,n965);
and (n2755,n1618,n975);
and (n2756,n2233,n1002);
and (n2757,n2758,n1022);
or (n2758,1'b0,n2759,n2763,n2764,n2765);
and (n2759,n2760,n930);
wire s0n2760,s1n2760,notn2760;
or (n2760,s0n2760,s1n2760);
not(notn2760,n927);
and (s0n2760,notn2760,n2761);
and (s1n2760,n927,n2762);
and (n2763,n2281,n955);
and (n2764,n1706,n965);
and (n2765,n1654,n975);
and (n2766,n2248,n1042);
and (n2767,n2746,n2768);
and (n2768,n2769,n2790);
or (n2769,1'b0,n2770,n2771,n2780,n2781);
and (n2770,n2337,n981);
and (n2771,n2772,n1002);
or (n2772,1'b0,n2773,n2774,n2775,n2776);
and (n2773,n1750,n930);
and (n2774,n1754,n955);
and (n2775,n2308,n965);
and (n2776,n2777,n975);
wire s0n2777,s1n2777,notn2777;
or (n2777,s0n2777,s1n2777);
not(notn2777,n927);
and (s0n2777,notn2777,n2778);
and (s1n2777,n927,n2779);
and (n2780,n2352,n1022);
and (n2781,n2782,n1042);
or (n2782,1'b0,n2783,n2784,n2785,n2786);
and (n2783,n1786,n930);
and (n2784,n1790,n955);
and (n2785,n2323,n965);
and (n2786,n2787,n975);
wire s0n2787,s1n2787,notn2787;
or (n2787,s0n2787,s1n2787);
not(notn2787,n927);
and (s0n2787,notn2787,n2788);
and (s1n2787,n927,n2789);
or (n2790,1'b0,n2791,n2800,n2801,n2810);
and (n2791,n2792,n981);
or (n2792,1'b0,n2793,n2797,n2798,n2799);
and (n2793,n2794,n930);
wire s0n2794,s1n2794,notn2794;
or (n2794,s0n2794,s1n2794);
not(notn2794,n927);
and (s0n2794,notn2794,n2795);
and (s1n2794,n927,n2796);
and (n2797,n2330,n955);
and (n2798,n1797,n965);
and (n2799,n1724,n975);
and (n2800,n2297,n1002);
and (n2801,n2802,n1022);
or (n2802,1'b0,n2803,n2807,n2808,n2809);
and (n2803,n2804,n930);
wire s0n2804,s1n2804,notn2804;
or (n2804,s0n2804,s1n2804);
not(notn2804,n927);
and (s0n2804,notn2804,n2805);
and (s1n2804,n927,n2806);
and (n2807,n2345,n955);
and (n2808,n1812,n965);
and (n2809,n1760,n975);
and (n2810,n2312,n1042);
and (n2811,n2725,n2768);
and (n2812,n2680,n2723);
and (n2813,n2635,n2678);
and (n2814,n2590,n2633);
and (n2815,n2545,n2588);
and (n2816,n2500,n2543);
and (n2817,n2455,n2498);
xor (n2818,n2421,n2423);
and (n2819,n2818,n2820);
or (n2820,n2821,n2825,n2870);
and (n2821,n2822,n2824);
xor (n2822,n2823,n2498);
xor (n2823,n2455,n2476);
xor (n2824,n2424,n2426);
and (n2825,n2824,n2826);
or (n2826,n2827,n2831,n2869);
and (n2827,n2828,n2830);
xor (n2828,n2829,n2543);
xor (n2829,n2500,n2521);
xor (n2830,n2427,n2429);
and (n2831,n2830,n2832);
or (n2832,n2833,n2837,n2868);
and (n2833,n2834,n2836);
xor (n2834,n2835,n2588);
xor (n2835,n2545,n2566);
xor (n2836,n2430,n2432);
and (n2837,n2836,n2838);
or (n2838,n2839,n2843,n2867);
and (n2839,n2840,n2842);
xor (n2840,n2841,n2633);
xor (n2841,n2590,n2611);
xor (n2842,n2433,n2435);
and (n2843,n2842,n2844);
or (n2844,n2845,n2849,n2866);
and (n2845,n2846,n2848);
xor (n2846,n2847,n2678);
xor (n2847,n2635,n2656);
xor (n2848,n2436,n2438);
and (n2849,n2848,n2850);
or (n2850,n2851,n2855,n2865);
and (n2851,n2852,n2854);
xor (n2852,n2853,n2723);
xor (n2853,n2680,n2701);
xor (n2854,n2439,n2440);
and (n2855,n2854,n2856);
or (n2856,n2857,n2861,n2864);
and (n2857,n2858,n2860);
xor (n2858,n2859,n2768);
xor (n2859,n2725,n2746);
xor (n2860,n2441,n2444);
and (n2861,n2860,n2862);
and (n2862,n2863,n2445);
xor (n2863,n2769,n2790);
and (n2864,n2858,n2862);
and (n2865,n2852,n2856);
and (n2866,n2846,n2850);
and (n2867,n2840,n2844);
and (n2868,n2834,n2838);
and (n2869,n2828,n2832);
and (n2870,n2822,n2826);
and (n2871,n2453,n2820);
or (n2872,n2873,n2874,n2924);
xor (n2873,n915,n2447);
and (n2874,n2450,n2875);
or (n2875,n2876,n2878,n2923);
and (n2876,n2877,n2818);
xor (n2877,n2448,n2449);
and (n2878,n2818,n2879);
or (n2879,n2880,n2882,n2922);
and (n2880,n2881,n2824);
xor (n2881,n2450,n2451);
and (n2882,n2824,n2883);
or (n2883,n2884,n2887,n2921);
and (n2884,n2885,n2830);
xor (n2885,n2886,n2820);
xor (n2886,n2453,n2818);
and (n2887,n2830,n2888);
or (n2888,n2889,n2892,n2920);
and (n2889,n2890,n2836);
xor (n2890,n2891,n2826);
xor (n2891,n2822,n2824);
and (n2892,n2836,n2893);
or (n2893,n2894,n2897,n2919);
and (n2894,n2895,n2842);
xor (n2895,n2896,n2832);
xor (n2896,n2828,n2830);
and (n2897,n2842,n2898);
or (n2898,n2899,n2902,n2918);
and (n2899,n2900,n2848);
xor (n2900,n2901,n2838);
xor (n2901,n2834,n2836);
and (n2902,n2848,n2903);
or (n2903,n2904,n2907,n2917);
and (n2904,n2905,n2854);
xor (n2905,n2906,n2844);
xor (n2906,n2840,n2842);
and (n2907,n2854,n2908);
or (n2908,n2909,n2912,n2916);
and (n2909,n2910,n2860);
xor (n2910,n2911,n2850);
xor (n2911,n2846,n2848);
and (n2912,n2860,n2913);
and (n2913,n2914,n2445);
xor (n2914,n2915,n2856);
xor (n2915,n2852,n2854);
and (n2916,n2910,n2913);
and (n2917,n2905,n2908);
and (n2918,n2900,n2903);
and (n2919,n2895,n2898);
and (n2920,n2890,n2893);
and (n2921,n2885,n2888);
and (n2922,n2881,n2883);
and (n2923,n2877,n2879);
and (n2924,n2873,n2875);
and (n2925,n2926,n2928);
xor (n2926,n2927,n2875);
xor (n2927,n2873,n2450);
and (n2928,n2929,n2931);
xor (n2929,n2930,n2879);
xor (n2930,n2877,n2818);
and (n2931,n2932,n2934);
xor (n2932,n2933,n2883);
xor (n2933,n2881,n2824);
and (n2934,n2935,n2937);
xor (n2935,n2936,n2888);
xor (n2936,n2885,n2830);
and (n2937,n2938,n2940);
xor (n2938,n2939,n2893);
xor (n2939,n2890,n2836);
and (n2940,n2941,n2943);
xor (n2941,n2942,n2898);
xor (n2942,n2895,n2842);
and (n2943,n2944,n2946);
xor (n2944,n2945,n2903);
xor (n2945,n2900,n2848);
xor (n2946,n2947,n2908);
xor (n2947,n2905,n2854);
and (n2948,n2949,n2960);
and (n2949,n2950,n2959);
and (n2950,n2951,n2958);
and (n2951,n2952,n2957);
and (n2952,n2953,n2956);
and (n2953,n21,n2954);
not (n2954,n2955);
nor (n2955,n25,n671,n744,n818);
not (n2956,n905);
not (n2957,n948);
not (n2958,n906);
or (n2959,n24,n671,n744,n818);
nand (n2960,n25,n671,n892,n817);
wire s0n2961,s1n2961,notn2961;
or (n2961,s0n2961,s1n2961);
not(notn2961,n2948);
and (s0n2961,notn2961,1'b0);
and (s1n2961,n2948,n2962);
xor (n2962,n2963,n2965);
xor (n2963,n2446,n2964);
and (n2964,n2448,n2872);
and (n2965,n912,n2925);
wire s0n2966,s1n2966,notn2966;
or (n2966,s0n2966,s1n2966);
not(notn2966,n2948);
and (s0n2966,notn2966,1'b0);
and (s1n2966,n2948,n2967);
xor (n2967,n2968,n2970);
xor (n2968,n2446,n2969);
and (n2969,n915,n2964);
and (n2970,n2963,n2965);
or (n2971,n2972,n929);
or (n2972,n2973,n928);
or (n2973,n943,n944);
or (n2974,1'b0,n2975,n2998,n3018,n3038);
and (n2975,n2976,n981);
or (n2976,1'b0,n2977,n2984,n2990);
and (n2977,n2978,n2983);
or (n2978,1'b0,n2979,n2980,n2981,n2982);
and (n2979,n926,n903);
and (n2980,n954,n949);
and (n2981,n964,n901);
and (n2982,n974,n960);
not (n2983,n2960);
and (n2984,n2985,n942);
or (n2985,1'b0,n2986,n2987,n2988,n2989);
and (n2986,n1050,n903);
and (n2987,n925,n949);
and (n2988,n953,n901);
and (n2989,n963,n960);
and (n2990,n2991,n2996);
or (n2991,1'b0,n2992,n2993,n2994,n2995);
and (n2992,n925,n903);
and (n2993,n953,n949);
and (n2994,n963,n901);
and (n2995,n973,n960);
or (n2996,n940,n2997);
not (n2997,n2959);
and (n2998,n2999,n1002);
or (n2999,1'b0,n3000,n3006,n3012);
and (n3000,n3001,n2983);
or (n3001,1'b0,n3002,n3003,n3004,n3005);
and (n3002,n989,n903);
and (n3003,n993,n949);
and (n3004,n997,n901);
and (n3005,n1001,n960);
and (n3006,n3007,n942);
or (n3007,1'b0,n3008,n3009,n3010,n3011);
and (n3008,n973,n903);
and (n3009,n988,n949);
and (n3010,n992,n901);
and (n3011,n996,n960);
and (n3012,n3013,n2996);
or (n3013,1'b0,n3014,n3015,n3016,n3017);
and (n3014,n988,n903);
and (n3015,n992,n949);
and (n3016,n996,n901);
and (n3017,n1000,n960);
and (n3018,n3019,n1022);
or (n3019,1'b0,n3020,n3026,n3032);
and (n3020,n3021,n2983);
or (n3021,1'b0,n3022,n3023,n3024,n3025);
and (n3022,n1009,n903);
and (n3023,n1013,n949);
and (n3024,n1017,n901);
and (n3025,n1021,n960);
and (n3026,n3027,n942);
or (n3027,1'b0,n3028,n3029,n3030,n3031);
and (n3028,n1065,n903);
and (n3029,n1008,n949);
and (n3030,n1012,n901);
and (n3031,n1016,n960);
and (n3032,n3033,n2996);
or (n3033,1'b0,n3034,n3035,n3036,n3037);
and (n3034,n1008,n903);
and (n3035,n1012,n949);
and (n3036,n1016,n901);
and (n3037,n1020,n960);
and (n3038,n3039,n1042);
or (n3039,1'b0,n3040,n3046,n3052);
and (n3040,n3041,n2983);
or (n3041,1'b0,n3042,n3043,n3044,n3045);
and (n3042,n1029,n903);
and (n3043,n1033,n949);
and (n3044,n1037,n901);
and (n3045,n1041,n960);
and (n3046,n3047,n942);
or (n3047,1'b0,n3048,n3049,n3050,n3051);
and (n3048,n1020,n903);
and (n3049,n1028,n949);
and (n3050,n1032,n901);
and (n3051,n1036,n960);
and (n3052,n3053,n2996);
or (n3053,1'b0,n3054,n3055,n3056,n3057);
and (n3054,n1028,n903);
and (n3055,n1032,n949);
and (n3056,n1036,n901);
and (n3057,n1040,n960);
or (n3058,1'b0,n3059,n6012,n6014,n6017);
and (n3059,n3060,n22);
wire s0n3060,s1n3060,notn3060;
or (n3060,s0n3060,s1n3060);
not(notn3060,n13);
and (s0n3060,notn3060,1'b0);
and (s1n3060,n13,n3061);
wire s0n3061,s1n3061,notn3061;
or (n3061,s0n3061,s1n3061);
not(notn3061,n6001);
and (s0n3061,notn3061,n3062);
and (s1n3061,n6001,1'b0);
wire s0n3062,s1n3062,notn3062;
or (n3062,s0n3062,s1n3062);
not(notn3062,n5986);
and (s0n3062,notn3062,n3063);
and (s1n3062,n5986,1'b1);
wire s0n3063,s1n3063,notn3063;
or (n3063,s0n3063,s1n3063);
not(notn3063,n3074);
and (s0n3063,notn3063,n3064);
and (s1n3063,n3074,n5775);
wire s0n3064,s1n3064,notn3064;
or (n3064,s0n3064,s1n3064);
not(notn3064,n3074);
and (s0n3064,notn3064,n3065);
and (s1n3064,n3074,n5772);
xor (n3065,n3066,n5749);
xor (n3066,n3067,n5692);
xor (n3067,n3068,n5623);
xor (n3068,n3069,n5613);
xor (n3069,n3070,n4138);
xor (n3070,n3071,n3084);
xor (n3071,n3072,n3082);
wire s0n3072,s1n3072,notn3072;
or (n3072,s0n3072,s1n3072);
not(notn3072,n3074);
and (s0n3072,notn3072,1'b0);
and (s1n3072,n3074,n3073);
or (n3074,n3075,n3081);
or (n3075,n3076,n3080);
and (n3076,n948,n3077);
or (n3077,n3078,n903);
or (n3078,n3079,n949);
or (n3079,n960,n901);
and (n3080,n22,n3077);
and (n3081,n904,n896);
wire s0n3082,s1n3082,notn3082;
or (n3082,s0n3082,s1n3082);
not(notn3082,n3074);
and (s0n3082,notn3082,1'b0);
and (s1n3082,n3074,n3083);
or (n3084,n3085,n3090,n4137);
and (n3085,n3086,n3088);
wire s0n3086,s1n3086,notn3086;
or (n3086,s0n3086,s1n3086);
not(notn3086,n3074);
and (s0n3086,notn3086,1'b0);
and (s1n3086,n3074,n3087);
wire s0n3088,s1n3088,notn3088;
or (n3088,s0n3088,s1n3088);
not(notn3088,n3074);
and (s0n3088,notn3088,1'b0);
and (s1n3088,n3074,n3089);
and (n3090,n3088,n3091);
or (n3091,n3092,n3097,n4136);
and (n3092,n3093,n3095);
wire s0n3093,s1n3093,notn3093;
or (n3093,s0n3093,s1n3093);
not(notn3093,n3074);
and (s0n3093,notn3093,1'b0);
and (s1n3093,n3074,n3094);
wire s0n3095,s1n3095,notn3095;
or (n3095,s0n3095,s1n3095);
not(notn3095,n3074);
and (s0n3095,notn3095,1'b0);
and (s1n3095,n3074,n3096);
and (n3097,n3095,n3098);
or (n3098,n3099,n3104,n4135);
and (n3099,n3100,n3102);
wire s0n3100,s1n3100,notn3100;
or (n3100,s0n3100,s1n3100);
not(notn3100,n3074);
and (s0n3100,notn3100,1'b0);
and (s1n3100,n3074,n3101);
wire s0n3102,s1n3102,notn3102;
or (n3102,s0n3102,s1n3102);
not(notn3102,n3074);
and (s0n3102,notn3102,1'b0);
and (s1n3102,n3074,n3103);
and (n3104,n3102,n3105);
or (n3105,n3106,n3111,n4134);
and (n3106,n3107,n3109);
wire s0n3107,s1n3107,notn3107;
or (n3107,s0n3107,s1n3107);
not(notn3107,n3074);
and (s0n3107,notn3107,1'b0);
and (s1n3107,n3074,n3108);
wire s0n3109,s1n3109,notn3109;
or (n3109,s0n3109,s1n3109);
not(notn3109,n3074);
and (s0n3109,notn3109,1'b0);
and (s1n3109,n3074,n3110);
and (n3111,n3109,n3112);
or (n3112,n3113,n3253,n4133);
and (n3113,n3114,n3192);
wire s0n3114,s1n3114,notn3114;
or (n3114,s0n3114,s1n3114);
not(notn3114,n3074);
and (s0n3114,notn3114,n3115);
and (s1n3114,n3074,n3191);
or (n3115,1'b0,n3116,n3148,n3162,n3177);
and (n3116,n3117,n981);
or (n3117,1'b0,n3118,n3133,n3138,n3143);
and (n3118,n3119,n3124);
wire s0n3119,s1n3119,notn3119;
or (n3119,s0n3119,s1n3119);
not(notn3119,n3122);
and (s0n3119,notn3119,n3120);
and (s1n3119,n3122,n3121);
or (n3122,n3123,n906);
or (n3123,n944,n929);
or (n3124,n3125,n950);
and (n3125,n3126,n903);
or (n3126,n3127,n929);
or (n3127,n3128,n928);
or (n3128,n3129,n944);
or (n3129,n3130,n943);
or (n3130,n3131,n2983);
or (n3131,n3132,n2997);
nor (n3132,n25,n941,n744,n818);
and (n3133,n3134,n3136);
wire s0n3134,s1n3134,notn3134;
or (n3134,s0n3134,s1n3134);
not(notn3134,n3122);
and (s0n3134,notn3134,n3135);
and (s1n3134,n3122,n3120);
or (n3136,n3137,n959);
and (n3137,n3126,n949);
and (n3138,n3139,n3141);
wire s0n3139,s1n3139,notn3139;
or (n3139,s0n3139,s1n3139);
not(notn3139,n3122);
and (s0n3139,notn3139,n3140);
and (s1n3139,n3122,n3135);
or (n3141,n3142,n969);
and (n3142,n3126,n901);
and (n3143,n3144,n3146);
wire s0n3144,s1n3144,notn3144;
or (n3144,s0n3144,s1n3144);
not(notn3144,n3122);
and (s0n3144,notn3144,n3145);
and (s1n3144,n3122,n3140);
or (n3146,n3147,n979);
and (n3147,n3126,n960);
and (n3148,n3149,n1002);
or (n3149,1'b0,n3150,n3153,n3156,n3159);
and (n3150,n3151,n3124);
wire s0n3151,s1n3151,notn3151;
or (n3151,s0n3151,s1n3151);
not(notn3151,n3122);
and (s0n3151,notn3151,n3152);
and (s1n3151,n3122,n3145);
and (n3153,n3154,n3136);
wire s0n3154,s1n3154,notn3154;
or (n3154,s0n3154,s1n3154);
not(notn3154,n3122);
and (s0n3154,notn3154,n3155);
and (s1n3154,n3122,n3152);
and (n3156,n3157,n3141);
wire s0n3157,s1n3157,notn3157;
or (n3157,s0n3157,s1n3157);
not(notn3157,n3122);
and (s0n3157,notn3157,n3158);
and (s1n3157,n3122,n3155);
and (n3159,n3160,n3146);
wire s0n3160,s1n3160,notn3160;
or (n3160,s0n3160,s1n3160);
not(notn3160,n3122);
and (s0n3160,notn3160,n3161);
and (s1n3160,n3122,n3158);
and (n3162,n3163,n1022);
or (n3163,1'b0,n3164,n3168,n3171,n3174);
and (n3164,n3165,n3124);
wire s0n3165,s1n3165,notn3165;
or (n3165,s0n3165,s1n3165);
not(notn3165,n3122);
and (s0n3165,notn3165,n3166);
and (s1n3165,n3122,n3167);
and (n3168,n3169,n3136);
wire s0n3169,s1n3169,notn3169;
or (n3169,s0n3169,s1n3169);
not(notn3169,n3122);
and (s0n3169,notn3169,n3170);
and (s1n3169,n3122,n3166);
and (n3171,n3172,n3141);
wire s0n3172,s1n3172,notn3172;
or (n3172,s0n3172,s1n3172);
not(notn3172,n3122);
and (s0n3172,notn3172,n3173);
and (s1n3172,n3122,n3170);
and (n3174,n3175,n3146);
wire s0n3175,s1n3175,notn3175;
or (n3175,s0n3175,s1n3175);
not(notn3175,n3122);
and (s0n3175,notn3175,n3176);
and (s1n3175,n3122,n3173);
and (n3177,n3178,n1042);
or (n3178,1'b0,n3179,n3182,n3185,n3188);
and (n3179,n3180,n3124);
wire s0n3180,s1n3180,notn3180;
or (n3180,s0n3180,s1n3180);
not(notn3180,n3122);
and (s0n3180,notn3180,n3181);
and (s1n3180,n3122,n3176);
and (n3182,n3183,n3136);
wire s0n3183,s1n3183,notn3183;
or (n3183,s0n3183,s1n3183);
not(notn3183,n3122);
and (s0n3183,notn3183,n3184);
and (s1n3183,n3122,n3181);
and (n3185,n3186,n3141);
wire s0n3186,s1n3186,notn3186;
or (n3186,s0n3186,s1n3186);
not(notn3186,n3122);
and (s0n3186,notn3186,n3187);
and (s1n3186,n3122,n3184);
and (n3188,n3189,n3146);
wire s0n3189,s1n3189,notn3189;
or (n3189,s0n3189,s1n3189);
not(notn3189,n3122);
and (s0n3189,notn3189,n3190);
and (s1n3189,n3122,n3187);
wire s0n3192,s1n3192,notn3192;
or (n3192,s0n3192,s1n3192);
not(notn3192,n3074);
and (s0n3192,notn3192,n3193);
and (s1n3192,n3074,n3252);
or (n3193,1'b0,n3194,n3209,n3223,n3238);
and (n3194,n3195,n981);
or (n3195,1'b0,n3196,n3200,n3203,n3206);
and (n3196,n3197,n3124);
wire s0n3197,s1n3197,notn3197;
or (n3197,s0n3197,s1n3197);
not(notn3197,n3122);
and (s0n3197,notn3197,n3198);
and (s1n3197,n3122,n3199);
and (n3200,n3201,n3136);
wire s0n3201,s1n3201,notn3201;
or (n3201,s0n3201,s1n3201);
not(notn3201,n3122);
and (s0n3201,notn3201,n3202);
and (s1n3201,n3122,n3198);
and (n3203,n3204,n3141);
wire s0n3204,s1n3204,notn3204;
or (n3204,s0n3204,s1n3204);
not(notn3204,n3122);
and (s0n3204,notn3204,n3205);
and (s1n3204,n3122,n3202);
and (n3206,n3207,n3146);
wire s0n3207,s1n3207,notn3207;
or (n3207,s0n3207,s1n3207);
not(notn3207,n3122);
and (s0n3207,notn3207,n3208);
and (s1n3207,n3122,n3205);
and (n3209,n3210,n1002);
or (n3210,1'b0,n3211,n3214,n3217,n3220);
and (n3211,n3212,n3124);
wire s0n3212,s1n3212,notn3212;
or (n3212,s0n3212,s1n3212);
not(notn3212,n3122);
and (s0n3212,notn3212,n3213);
and (s1n3212,n3122,n3208);
and (n3214,n3215,n3136);
wire s0n3215,s1n3215,notn3215;
or (n3215,s0n3215,s1n3215);
not(notn3215,n3122);
and (s0n3215,notn3215,n3216);
and (s1n3215,n3122,n3213);
and (n3217,n3218,n3141);
wire s0n3218,s1n3218,notn3218;
or (n3218,s0n3218,s1n3218);
not(notn3218,n3122);
and (s0n3218,notn3218,n3219);
and (s1n3218,n3122,n3216);
and (n3220,n3221,n3146);
wire s0n3221,s1n3221,notn3221;
or (n3221,s0n3221,s1n3221);
not(notn3221,n3122);
and (s0n3221,notn3221,n3222);
and (s1n3221,n3122,n3219);
and (n3223,n3224,n1022);
or (n3224,1'b0,n3225,n3229,n3232,n3235);
and (n3225,n3226,n3124);
wire s0n3226,s1n3226,notn3226;
or (n3226,s0n3226,s1n3226);
not(notn3226,n3122);
and (s0n3226,notn3226,n3227);
and (s1n3226,n3122,n3228);
and (n3229,n3230,n3136);
wire s0n3230,s1n3230,notn3230;
or (n3230,s0n3230,s1n3230);
not(notn3230,n3122);
and (s0n3230,notn3230,n3231);
and (s1n3230,n3122,n3227);
and (n3232,n3233,n3141);
wire s0n3233,s1n3233,notn3233;
or (n3233,s0n3233,s1n3233);
not(notn3233,n3122);
and (s0n3233,notn3233,n3234);
and (s1n3233,n3122,n3231);
and (n3235,n3236,n3146);
wire s0n3236,s1n3236,notn3236;
or (n3236,s0n3236,s1n3236);
not(notn3236,n3122);
and (s0n3236,notn3236,n3237);
and (s1n3236,n3122,n3234);
and (n3238,n3239,n1042);
or (n3239,1'b0,n3240,n3243,n3246,n3249);
and (n3240,n3241,n3124);
wire s0n3241,s1n3241,notn3241;
or (n3241,s0n3241,s1n3241);
not(notn3241,n3122);
and (s0n3241,notn3241,n3242);
and (s1n3241,n3122,n3237);
and (n3243,n3244,n3136);
wire s0n3244,s1n3244,notn3244;
or (n3244,s0n3244,s1n3244);
not(notn3244,n3122);
and (s0n3244,notn3244,n3245);
and (s1n3244,n3122,n3242);
and (n3246,n3247,n3141);
wire s0n3247,s1n3247,notn3247;
or (n3247,s0n3247,s1n3247);
not(notn3247,n3122);
and (s0n3247,notn3247,n3248);
and (s1n3247,n3122,n3245);
and (n3249,n3250,n3146);
wire s0n3250,s1n3250,notn3250;
or (n3250,s0n3250,s1n3250);
not(notn3250,n3122);
and (s0n3250,notn3250,n3251);
and (s1n3250,n3122,n3248);
and (n3253,n3192,n3254);
or (n3254,n3255,n3378,n4132);
and (n3255,n3256,n3317);
wire s0n3256,s1n3256,notn3256;
or (n3256,s0n3256,s1n3256);
not(notn3256,n3074);
and (s0n3256,notn3256,n3257);
and (s1n3256,n3074,n3316);
or (n3257,1'b0,n3258,n3273,n3287,n3302);
and (n3258,n3259,n981);
or (n3259,1'b0,n3260,n3264,n3267,n3270);
and (n3260,n3261,n3124);
wire s0n3261,s1n3261,notn3261;
or (n3261,s0n3261,s1n3261);
not(notn3261,n3122);
and (s0n3261,notn3261,n3262);
and (s1n3261,n3122,n3263);
and (n3264,n3265,n3136);
wire s0n3265,s1n3265,notn3265;
or (n3265,s0n3265,s1n3265);
not(notn3265,n3122);
and (s0n3265,notn3265,n3266);
and (s1n3265,n3122,n3262);
and (n3267,n3268,n3141);
wire s0n3268,s1n3268,notn3268;
or (n3268,s0n3268,s1n3268);
not(notn3268,n3122);
and (s0n3268,notn3268,n3269);
and (s1n3268,n3122,n3266);
and (n3270,n3271,n3146);
wire s0n3271,s1n3271,notn3271;
or (n3271,s0n3271,s1n3271);
not(notn3271,n3122);
and (s0n3271,notn3271,n3272);
and (s1n3271,n3122,n3269);
and (n3273,n3274,n1002);
or (n3274,1'b0,n3275,n3278,n3281,n3284);
and (n3275,n3276,n3124);
wire s0n3276,s1n3276,notn3276;
or (n3276,s0n3276,s1n3276);
not(notn3276,n3122);
and (s0n3276,notn3276,n3277);
and (s1n3276,n3122,n3272);
and (n3278,n3279,n3136);
wire s0n3279,s1n3279,notn3279;
or (n3279,s0n3279,s1n3279);
not(notn3279,n3122);
and (s0n3279,notn3279,n3280);
and (s1n3279,n3122,n3277);
and (n3281,n3282,n3141);
wire s0n3282,s1n3282,notn3282;
or (n3282,s0n3282,s1n3282);
not(notn3282,n3122);
and (s0n3282,notn3282,n3283);
and (s1n3282,n3122,n3280);
and (n3284,n3285,n3146);
wire s0n3285,s1n3285,notn3285;
or (n3285,s0n3285,s1n3285);
not(notn3285,n3122);
and (s0n3285,notn3285,n3286);
and (s1n3285,n3122,n3283);
and (n3287,n3288,n1022);
or (n3288,1'b0,n3289,n3293,n3296,n3299);
and (n3289,n3290,n3124);
wire s0n3290,s1n3290,notn3290;
or (n3290,s0n3290,s1n3290);
not(notn3290,n3122);
and (s0n3290,notn3290,n3291);
and (s1n3290,n3122,n3292);
and (n3293,n3294,n3136);
wire s0n3294,s1n3294,notn3294;
or (n3294,s0n3294,s1n3294);
not(notn3294,n3122);
and (s0n3294,notn3294,n3295);
and (s1n3294,n3122,n3291);
and (n3296,n3297,n3141);
wire s0n3297,s1n3297,notn3297;
or (n3297,s0n3297,s1n3297);
not(notn3297,n3122);
and (s0n3297,notn3297,n3298);
and (s1n3297,n3122,n3295);
and (n3299,n3300,n3146);
wire s0n3300,s1n3300,notn3300;
or (n3300,s0n3300,s1n3300);
not(notn3300,n3122);
and (s0n3300,notn3300,n3301);
and (s1n3300,n3122,n3298);
and (n3302,n3303,n1042);
or (n3303,1'b0,n3304,n3307,n3310,n3313);
and (n3304,n3305,n3124);
wire s0n3305,s1n3305,notn3305;
or (n3305,s0n3305,s1n3305);
not(notn3305,n3122);
and (s0n3305,notn3305,n3306);
and (s1n3305,n3122,n3301);
and (n3307,n3308,n3136);
wire s0n3308,s1n3308,notn3308;
or (n3308,s0n3308,s1n3308);
not(notn3308,n3122);
and (s0n3308,notn3308,n3309);
and (s1n3308,n3122,n3306);
and (n3310,n3311,n3141);
wire s0n3311,s1n3311,notn3311;
or (n3311,s0n3311,s1n3311);
not(notn3311,n3122);
and (s0n3311,notn3311,n3312);
and (s1n3311,n3122,n3309);
and (n3313,n3314,n3146);
wire s0n3314,s1n3314,notn3314;
or (n3314,s0n3314,s1n3314);
not(notn3314,n3122);
and (s0n3314,notn3314,n3315);
and (s1n3314,n3122,n3312);
wire s0n3317,s1n3317,notn3317;
or (n3317,s0n3317,s1n3317);
not(notn3317,n3074);
and (s0n3317,notn3317,n3318);
and (s1n3317,n3074,n3377);
or (n3318,1'b0,n3319,n3334,n3348,n3363);
and (n3319,n3320,n981);
or (n3320,1'b0,n3321,n3325,n3328,n3331);
and (n3321,n3322,n3124);
wire s0n3322,s1n3322,notn3322;
or (n3322,s0n3322,s1n3322);
not(notn3322,n3122);
and (s0n3322,notn3322,n3323);
and (s1n3322,n3122,n3324);
and (n3325,n3326,n3136);
wire s0n3326,s1n3326,notn3326;
or (n3326,s0n3326,s1n3326);
not(notn3326,n3122);
and (s0n3326,notn3326,n3327);
and (s1n3326,n3122,n3323);
and (n3328,n3329,n3141);
wire s0n3329,s1n3329,notn3329;
or (n3329,s0n3329,s1n3329);
not(notn3329,n3122);
and (s0n3329,notn3329,n3330);
and (s1n3329,n3122,n3327);
and (n3331,n3332,n3146);
wire s0n3332,s1n3332,notn3332;
or (n3332,s0n3332,s1n3332);
not(notn3332,n3122);
and (s0n3332,notn3332,n3333);
and (s1n3332,n3122,n3330);
and (n3334,n3335,n1002);
or (n3335,1'b0,n3336,n3339,n3342,n3345);
and (n3336,n3337,n3124);
wire s0n3337,s1n3337,notn3337;
or (n3337,s0n3337,s1n3337);
not(notn3337,n3122);
and (s0n3337,notn3337,n3338);
and (s1n3337,n3122,n3333);
and (n3339,n3340,n3136);
wire s0n3340,s1n3340,notn3340;
or (n3340,s0n3340,s1n3340);
not(notn3340,n3122);
and (s0n3340,notn3340,n3341);
and (s1n3340,n3122,n3338);
and (n3342,n3343,n3141);
wire s0n3343,s1n3343,notn3343;
or (n3343,s0n3343,s1n3343);
not(notn3343,n3122);
and (s0n3343,notn3343,n3344);
and (s1n3343,n3122,n3341);
and (n3345,n3346,n3146);
wire s0n3346,s1n3346,notn3346;
or (n3346,s0n3346,s1n3346);
not(notn3346,n3122);
and (s0n3346,notn3346,n3347);
and (s1n3346,n3122,n3344);
and (n3348,n3349,n1022);
or (n3349,1'b0,n3350,n3354,n3357,n3360);
and (n3350,n3351,n3124);
wire s0n3351,s1n3351,notn3351;
or (n3351,s0n3351,s1n3351);
not(notn3351,n3122);
and (s0n3351,notn3351,n3352);
and (s1n3351,n3122,n3353);
and (n3354,n3355,n3136);
wire s0n3355,s1n3355,notn3355;
or (n3355,s0n3355,s1n3355);
not(notn3355,n3122);
and (s0n3355,notn3355,n3356);
and (s1n3355,n3122,n3352);
and (n3357,n3358,n3141);
wire s0n3358,s1n3358,notn3358;
or (n3358,s0n3358,s1n3358);
not(notn3358,n3122);
and (s0n3358,notn3358,n3359);
and (s1n3358,n3122,n3356);
and (n3360,n3361,n3146);
wire s0n3361,s1n3361,notn3361;
or (n3361,s0n3361,s1n3361);
not(notn3361,n3122);
and (s0n3361,notn3361,n3362);
and (s1n3361,n3122,n3359);
and (n3363,n3364,n1042);
or (n3364,1'b0,n3365,n3368,n3371,n3374);
and (n3365,n3366,n3124);
wire s0n3366,s1n3366,notn3366;
or (n3366,s0n3366,s1n3366);
not(notn3366,n3122);
and (s0n3366,notn3366,n3367);
and (s1n3366,n3122,n3362);
and (n3368,n3369,n3136);
wire s0n3369,s1n3369,notn3369;
or (n3369,s0n3369,s1n3369);
not(notn3369,n3122);
and (s0n3369,notn3369,n3370);
and (s1n3369,n3122,n3367);
and (n3371,n3372,n3141);
wire s0n3372,s1n3372,notn3372;
or (n3372,s0n3372,s1n3372);
not(notn3372,n3122);
and (s0n3372,notn3372,n3373);
and (s1n3372,n3122,n3370);
and (n3374,n3375,n3146);
wire s0n3375,s1n3375,notn3375;
or (n3375,s0n3375,s1n3375);
not(notn3375,n3122);
and (s0n3375,notn3375,n3376);
and (s1n3375,n3122,n3373);
and (n3378,n3317,n3379);
or (n3379,n3380,n3503,n4131);
and (n3380,n3381,n3442);
wire s0n3381,s1n3381,notn3381;
or (n3381,s0n3381,s1n3381);
not(notn3381,n3074);
and (s0n3381,notn3381,n3382);
and (s1n3381,n3074,n3441);
or (n3382,1'b0,n3383,n3398,n3412,n3427);
and (n3383,n3384,n981);
or (n3384,1'b0,n3385,n3389,n3392,n3395);
and (n3385,n3386,n3124);
wire s0n3386,s1n3386,notn3386;
or (n3386,s0n3386,s1n3386);
not(notn3386,n3122);
and (s0n3386,notn3386,n3387);
and (s1n3386,n3122,n3388);
and (n3389,n3390,n3136);
wire s0n3390,s1n3390,notn3390;
or (n3390,s0n3390,s1n3390);
not(notn3390,n3122);
and (s0n3390,notn3390,n3391);
and (s1n3390,n3122,n3387);
and (n3392,n3393,n3141);
wire s0n3393,s1n3393,notn3393;
or (n3393,s0n3393,s1n3393);
not(notn3393,n3122);
and (s0n3393,notn3393,n3394);
and (s1n3393,n3122,n3391);
and (n3395,n3396,n3146);
wire s0n3396,s1n3396,notn3396;
or (n3396,s0n3396,s1n3396);
not(notn3396,n3122);
and (s0n3396,notn3396,n3397);
and (s1n3396,n3122,n3394);
and (n3398,n3399,n1002);
or (n3399,1'b0,n3400,n3403,n3406,n3409);
and (n3400,n3401,n3124);
wire s0n3401,s1n3401,notn3401;
or (n3401,s0n3401,s1n3401);
not(notn3401,n3122);
and (s0n3401,notn3401,n3402);
and (s1n3401,n3122,n3397);
and (n3403,n3404,n3136);
wire s0n3404,s1n3404,notn3404;
or (n3404,s0n3404,s1n3404);
not(notn3404,n3122);
and (s0n3404,notn3404,n3405);
and (s1n3404,n3122,n3402);
and (n3406,n3407,n3141);
wire s0n3407,s1n3407,notn3407;
or (n3407,s0n3407,s1n3407);
not(notn3407,n3122);
and (s0n3407,notn3407,n3408);
and (s1n3407,n3122,n3405);
and (n3409,n3410,n3146);
wire s0n3410,s1n3410,notn3410;
or (n3410,s0n3410,s1n3410);
not(notn3410,n3122);
and (s0n3410,notn3410,n3411);
and (s1n3410,n3122,n3408);
and (n3412,n3413,n1022);
or (n3413,1'b0,n3414,n3418,n3421,n3424);
and (n3414,n3415,n3124);
wire s0n3415,s1n3415,notn3415;
or (n3415,s0n3415,s1n3415);
not(notn3415,n3122);
and (s0n3415,notn3415,n3416);
and (s1n3415,n3122,n3417);
and (n3418,n3419,n3136);
wire s0n3419,s1n3419,notn3419;
or (n3419,s0n3419,s1n3419);
not(notn3419,n3122);
and (s0n3419,notn3419,n3420);
and (s1n3419,n3122,n3416);
and (n3421,n3422,n3141);
wire s0n3422,s1n3422,notn3422;
or (n3422,s0n3422,s1n3422);
not(notn3422,n3122);
and (s0n3422,notn3422,n3423);
and (s1n3422,n3122,n3420);
and (n3424,n3425,n3146);
wire s0n3425,s1n3425,notn3425;
or (n3425,s0n3425,s1n3425);
not(notn3425,n3122);
and (s0n3425,notn3425,n3426);
and (s1n3425,n3122,n3423);
and (n3427,n3428,n1042);
or (n3428,1'b0,n3429,n3432,n3435,n3438);
and (n3429,n3430,n3124);
wire s0n3430,s1n3430,notn3430;
or (n3430,s0n3430,s1n3430);
not(notn3430,n3122);
and (s0n3430,notn3430,n3431);
and (s1n3430,n3122,n3426);
and (n3432,n3433,n3136);
wire s0n3433,s1n3433,notn3433;
or (n3433,s0n3433,s1n3433);
not(notn3433,n3122);
and (s0n3433,notn3433,n3434);
and (s1n3433,n3122,n3431);
and (n3435,n3436,n3141);
wire s0n3436,s1n3436,notn3436;
or (n3436,s0n3436,s1n3436);
not(notn3436,n3122);
and (s0n3436,notn3436,n3437);
and (s1n3436,n3122,n3434);
and (n3438,n3439,n3146);
wire s0n3439,s1n3439,notn3439;
or (n3439,s0n3439,s1n3439);
not(notn3439,n3122);
and (s0n3439,notn3439,n3440);
and (s1n3439,n3122,n3437);
wire s0n3442,s1n3442,notn3442;
or (n3442,s0n3442,s1n3442);
not(notn3442,n3074);
and (s0n3442,notn3442,n3443);
and (s1n3442,n3074,n3502);
or (n3443,1'b0,n3444,n3459,n3473,n3488);
and (n3444,n3445,n981);
or (n3445,1'b0,n3446,n3450,n3453,n3456);
and (n3446,n3447,n3124);
wire s0n3447,s1n3447,notn3447;
or (n3447,s0n3447,s1n3447);
not(notn3447,n3122);
and (s0n3447,notn3447,n3448);
and (s1n3447,n3122,n3449);
and (n3450,n3451,n3136);
wire s0n3451,s1n3451,notn3451;
or (n3451,s0n3451,s1n3451);
not(notn3451,n3122);
and (s0n3451,notn3451,n3452);
and (s1n3451,n3122,n3448);
and (n3453,n3454,n3141);
wire s0n3454,s1n3454,notn3454;
or (n3454,s0n3454,s1n3454);
not(notn3454,n3122);
and (s0n3454,notn3454,n3455);
and (s1n3454,n3122,n3452);
and (n3456,n3457,n3146);
wire s0n3457,s1n3457,notn3457;
or (n3457,s0n3457,s1n3457);
not(notn3457,n3122);
and (s0n3457,notn3457,n3458);
and (s1n3457,n3122,n3455);
and (n3459,n3460,n1002);
or (n3460,1'b0,n3461,n3464,n3467,n3470);
and (n3461,n3462,n3124);
wire s0n3462,s1n3462,notn3462;
or (n3462,s0n3462,s1n3462);
not(notn3462,n3122);
and (s0n3462,notn3462,n3463);
and (s1n3462,n3122,n3458);
and (n3464,n3465,n3136);
wire s0n3465,s1n3465,notn3465;
or (n3465,s0n3465,s1n3465);
not(notn3465,n3122);
and (s0n3465,notn3465,n3466);
and (s1n3465,n3122,n3463);
and (n3467,n3468,n3141);
wire s0n3468,s1n3468,notn3468;
or (n3468,s0n3468,s1n3468);
not(notn3468,n3122);
and (s0n3468,notn3468,n3469);
and (s1n3468,n3122,n3466);
and (n3470,n3471,n3146);
wire s0n3471,s1n3471,notn3471;
or (n3471,s0n3471,s1n3471);
not(notn3471,n3122);
and (s0n3471,notn3471,n3472);
and (s1n3471,n3122,n3469);
and (n3473,n3474,n1022);
or (n3474,1'b0,n3475,n3479,n3482,n3485);
and (n3475,n3476,n3124);
wire s0n3476,s1n3476,notn3476;
or (n3476,s0n3476,s1n3476);
not(notn3476,n3122);
and (s0n3476,notn3476,n3477);
and (s1n3476,n3122,n3478);
and (n3479,n3480,n3136);
wire s0n3480,s1n3480,notn3480;
or (n3480,s0n3480,s1n3480);
not(notn3480,n3122);
and (s0n3480,notn3480,n3481);
and (s1n3480,n3122,n3477);
and (n3482,n3483,n3141);
wire s0n3483,s1n3483,notn3483;
or (n3483,s0n3483,s1n3483);
not(notn3483,n3122);
and (s0n3483,notn3483,n3484);
and (s1n3483,n3122,n3481);
and (n3485,n3486,n3146);
wire s0n3486,s1n3486,notn3486;
or (n3486,s0n3486,s1n3486);
not(notn3486,n3122);
and (s0n3486,notn3486,n3487);
and (s1n3486,n3122,n3484);
and (n3488,n3489,n1042);
or (n3489,1'b0,n3490,n3493,n3496,n3499);
and (n3490,n3491,n3124);
wire s0n3491,s1n3491,notn3491;
or (n3491,s0n3491,s1n3491);
not(notn3491,n3122);
and (s0n3491,notn3491,n3492);
and (s1n3491,n3122,n3487);
and (n3493,n3494,n3136);
wire s0n3494,s1n3494,notn3494;
or (n3494,s0n3494,s1n3494);
not(notn3494,n3122);
and (s0n3494,notn3494,n3495);
and (s1n3494,n3122,n3492);
and (n3496,n3497,n3141);
wire s0n3497,s1n3497,notn3497;
or (n3497,s0n3497,s1n3497);
not(notn3497,n3122);
and (s0n3497,notn3497,n3498);
and (s1n3497,n3122,n3495);
and (n3499,n3500,n3146);
wire s0n3500,s1n3500,notn3500;
or (n3500,s0n3500,s1n3500);
not(notn3500,n3122);
and (s0n3500,notn3500,n3501);
and (s1n3500,n3122,n3498);
and (n3503,n3442,n3504);
or (n3504,n3505,n3628,n4130);
and (n3505,n3506,n3567);
wire s0n3506,s1n3506,notn3506;
or (n3506,s0n3506,s1n3506);
not(notn3506,n3074);
and (s0n3506,notn3506,n3507);
and (s1n3506,n3074,n3566);
or (n3507,1'b0,n3508,n3523,n3537,n3552);
and (n3508,n3509,n981);
or (n3509,1'b0,n3510,n3514,n3517,n3520);
and (n3510,n3511,n3124);
wire s0n3511,s1n3511,notn3511;
or (n3511,s0n3511,s1n3511);
not(notn3511,n3122);
and (s0n3511,notn3511,n3512);
and (s1n3511,n3122,n3513);
and (n3514,n3515,n3136);
wire s0n3515,s1n3515,notn3515;
or (n3515,s0n3515,s1n3515);
not(notn3515,n3122);
and (s0n3515,notn3515,n3516);
and (s1n3515,n3122,n3512);
and (n3517,n3518,n3141);
wire s0n3518,s1n3518,notn3518;
or (n3518,s0n3518,s1n3518);
not(notn3518,n3122);
and (s0n3518,notn3518,n3519);
and (s1n3518,n3122,n3516);
and (n3520,n3521,n3146);
wire s0n3521,s1n3521,notn3521;
or (n3521,s0n3521,s1n3521);
not(notn3521,n3122);
and (s0n3521,notn3521,n3522);
and (s1n3521,n3122,n3519);
and (n3523,n3524,n1002);
or (n3524,1'b0,n3525,n3528,n3531,n3534);
and (n3525,n3526,n3124);
wire s0n3526,s1n3526,notn3526;
or (n3526,s0n3526,s1n3526);
not(notn3526,n3122);
and (s0n3526,notn3526,n3527);
and (s1n3526,n3122,n3522);
and (n3528,n3529,n3136);
wire s0n3529,s1n3529,notn3529;
or (n3529,s0n3529,s1n3529);
not(notn3529,n3122);
and (s0n3529,notn3529,n3530);
and (s1n3529,n3122,n3527);
and (n3531,n3532,n3141);
wire s0n3532,s1n3532,notn3532;
or (n3532,s0n3532,s1n3532);
not(notn3532,n3122);
and (s0n3532,notn3532,n3533);
and (s1n3532,n3122,n3530);
and (n3534,n3535,n3146);
wire s0n3535,s1n3535,notn3535;
or (n3535,s0n3535,s1n3535);
not(notn3535,n3122);
and (s0n3535,notn3535,n3536);
and (s1n3535,n3122,n3533);
and (n3537,n3538,n1022);
or (n3538,1'b0,n3539,n3543,n3546,n3549);
and (n3539,n3540,n3124);
wire s0n3540,s1n3540,notn3540;
or (n3540,s0n3540,s1n3540);
not(notn3540,n3122);
and (s0n3540,notn3540,n3541);
and (s1n3540,n3122,n3542);
and (n3543,n3544,n3136);
wire s0n3544,s1n3544,notn3544;
or (n3544,s0n3544,s1n3544);
not(notn3544,n3122);
and (s0n3544,notn3544,n3545);
and (s1n3544,n3122,n3541);
and (n3546,n3547,n3141);
wire s0n3547,s1n3547,notn3547;
or (n3547,s0n3547,s1n3547);
not(notn3547,n3122);
and (s0n3547,notn3547,n3548);
and (s1n3547,n3122,n3545);
and (n3549,n3550,n3146);
wire s0n3550,s1n3550,notn3550;
or (n3550,s0n3550,s1n3550);
not(notn3550,n3122);
and (s0n3550,notn3550,n3551);
and (s1n3550,n3122,n3548);
and (n3552,n3553,n1042);
or (n3553,1'b0,n3554,n3557,n3560,n3563);
and (n3554,n3555,n3124);
wire s0n3555,s1n3555,notn3555;
or (n3555,s0n3555,s1n3555);
not(notn3555,n3122);
and (s0n3555,notn3555,n3556);
and (s1n3555,n3122,n3551);
and (n3557,n3558,n3136);
wire s0n3558,s1n3558,notn3558;
or (n3558,s0n3558,s1n3558);
not(notn3558,n3122);
and (s0n3558,notn3558,n3559);
and (s1n3558,n3122,n3556);
and (n3560,n3561,n3141);
wire s0n3561,s1n3561,notn3561;
or (n3561,s0n3561,s1n3561);
not(notn3561,n3122);
and (s0n3561,notn3561,n3562);
and (s1n3561,n3122,n3559);
and (n3563,n3564,n3146);
wire s0n3564,s1n3564,notn3564;
or (n3564,s0n3564,s1n3564);
not(notn3564,n3122);
and (s0n3564,notn3564,n3565);
and (s1n3564,n3122,n3562);
wire s0n3567,s1n3567,notn3567;
or (n3567,s0n3567,s1n3567);
not(notn3567,n3074);
and (s0n3567,notn3567,n3568);
and (s1n3567,n3074,n3627);
or (n3568,1'b0,n3569,n3584,n3598,n3613);
and (n3569,n3570,n981);
or (n3570,1'b0,n3571,n3575,n3578,n3581);
and (n3571,n3572,n3124);
wire s0n3572,s1n3572,notn3572;
or (n3572,s0n3572,s1n3572);
not(notn3572,n3122);
and (s0n3572,notn3572,n3573);
and (s1n3572,n3122,n3574);
and (n3575,n3576,n3136);
wire s0n3576,s1n3576,notn3576;
or (n3576,s0n3576,s1n3576);
not(notn3576,n3122);
and (s0n3576,notn3576,n3577);
and (s1n3576,n3122,n3573);
and (n3578,n3579,n3141);
wire s0n3579,s1n3579,notn3579;
or (n3579,s0n3579,s1n3579);
not(notn3579,n3122);
and (s0n3579,notn3579,n3580);
and (s1n3579,n3122,n3577);
and (n3581,n3582,n3146);
wire s0n3582,s1n3582,notn3582;
or (n3582,s0n3582,s1n3582);
not(notn3582,n3122);
and (s0n3582,notn3582,n3583);
and (s1n3582,n3122,n3580);
and (n3584,n3585,n1002);
or (n3585,1'b0,n3586,n3589,n3592,n3595);
and (n3586,n3587,n3124);
wire s0n3587,s1n3587,notn3587;
or (n3587,s0n3587,s1n3587);
not(notn3587,n3122);
and (s0n3587,notn3587,n3588);
and (s1n3587,n3122,n3583);
and (n3589,n3590,n3136);
wire s0n3590,s1n3590,notn3590;
or (n3590,s0n3590,s1n3590);
not(notn3590,n3122);
and (s0n3590,notn3590,n3591);
and (s1n3590,n3122,n3588);
and (n3592,n3593,n3141);
wire s0n3593,s1n3593,notn3593;
or (n3593,s0n3593,s1n3593);
not(notn3593,n3122);
and (s0n3593,notn3593,n3594);
and (s1n3593,n3122,n3591);
and (n3595,n3596,n3146);
wire s0n3596,s1n3596,notn3596;
or (n3596,s0n3596,s1n3596);
not(notn3596,n3122);
and (s0n3596,notn3596,n3597);
and (s1n3596,n3122,n3594);
and (n3598,n3599,n1022);
or (n3599,1'b0,n3600,n3604,n3607,n3610);
and (n3600,n3601,n3124);
wire s0n3601,s1n3601,notn3601;
or (n3601,s0n3601,s1n3601);
not(notn3601,n3122);
and (s0n3601,notn3601,n3602);
and (s1n3601,n3122,n3603);
and (n3604,n3605,n3136);
wire s0n3605,s1n3605,notn3605;
or (n3605,s0n3605,s1n3605);
not(notn3605,n3122);
and (s0n3605,notn3605,n3606);
and (s1n3605,n3122,n3602);
and (n3607,n3608,n3141);
wire s0n3608,s1n3608,notn3608;
or (n3608,s0n3608,s1n3608);
not(notn3608,n3122);
and (s0n3608,notn3608,n3609);
and (s1n3608,n3122,n3606);
and (n3610,n3611,n3146);
wire s0n3611,s1n3611,notn3611;
or (n3611,s0n3611,s1n3611);
not(notn3611,n3122);
and (s0n3611,notn3611,n3612);
and (s1n3611,n3122,n3609);
and (n3613,n3614,n1042);
or (n3614,1'b0,n3615,n3618,n3621,n3624);
and (n3615,n3616,n3124);
wire s0n3616,s1n3616,notn3616;
or (n3616,s0n3616,s1n3616);
not(notn3616,n3122);
and (s0n3616,notn3616,n3617);
and (s1n3616,n3122,n3612);
and (n3618,n3619,n3136);
wire s0n3619,s1n3619,notn3619;
or (n3619,s0n3619,s1n3619);
not(notn3619,n3122);
and (s0n3619,notn3619,n3620);
and (s1n3619,n3122,n3617);
and (n3621,n3622,n3141);
wire s0n3622,s1n3622,notn3622;
or (n3622,s0n3622,s1n3622);
not(notn3622,n3122);
and (s0n3622,notn3622,n3623);
and (s1n3622,n3122,n3620);
and (n3624,n3625,n3146);
wire s0n3625,s1n3625,notn3625;
or (n3625,s0n3625,s1n3625);
not(notn3625,n3122);
and (s0n3625,notn3625,n3626);
and (s1n3625,n3122,n3623);
and (n3628,n3567,n3629);
or (n3629,n3630,n3753,n4129);
and (n3630,n3631,n3692);
wire s0n3631,s1n3631,notn3631;
or (n3631,s0n3631,s1n3631);
not(notn3631,n3074);
and (s0n3631,notn3631,n3632);
and (s1n3631,n3074,n3691);
or (n3632,1'b0,n3633,n3648,n3662,n3677);
and (n3633,n3634,n981);
or (n3634,1'b0,n3635,n3639,n3642,n3645);
and (n3635,n3636,n3124);
wire s0n3636,s1n3636,notn3636;
or (n3636,s0n3636,s1n3636);
not(notn3636,n3122);
and (s0n3636,notn3636,n3637);
and (s1n3636,n3122,n3638);
and (n3639,n3640,n3136);
wire s0n3640,s1n3640,notn3640;
or (n3640,s0n3640,s1n3640);
not(notn3640,n3122);
and (s0n3640,notn3640,n3641);
and (s1n3640,n3122,n3637);
and (n3642,n3643,n3141);
wire s0n3643,s1n3643,notn3643;
or (n3643,s0n3643,s1n3643);
not(notn3643,n3122);
and (s0n3643,notn3643,n3644);
and (s1n3643,n3122,n3641);
and (n3645,n3646,n3146);
wire s0n3646,s1n3646,notn3646;
or (n3646,s0n3646,s1n3646);
not(notn3646,n3122);
and (s0n3646,notn3646,n3647);
and (s1n3646,n3122,n3644);
and (n3648,n3649,n1002);
or (n3649,1'b0,n3650,n3653,n3656,n3659);
and (n3650,n3651,n3124);
wire s0n3651,s1n3651,notn3651;
or (n3651,s0n3651,s1n3651);
not(notn3651,n3122);
and (s0n3651,notn3651,n3652);
and (s1n3651,n3122,n3647);
and (n3653,n3654,n3136);
wire s0n3654,s1n3654,notn3654;
or (n3654,s0n3654,s1n3654);
not(notn3654,n3122);
and (s0n3654,notn3654,n3655);
and (s1n3654,n3122,n3652);
and (n3656,n3657,n3141);
wire s0n3657,s1n3657,notn3657;
or (n3657,s0n3657,s1n3657);
not(notn3657,n3122);
and (s0n3657,notn3657,n3658);
and (s1n3657,n3122,n3655);
and (n3659,n3660,n3146);
wire s0n3660,s1n3660,notn3660;
or (n3660,s0n3660,s1n3660);
not(notn3660,n3122);
and (s0n3660,notn3660,n3661);
and (s1n3660,n3122,n3658);
and (n3662,n3663,n1022);
or (n3663,1'b0,n3664,n3668,n3671,n3674);
and (n3664,n3665,n3124);
wire s0n3665,s1n3665,notn3665;
or (n3665,s0n3665,s1n3665);
not(notn3665,n3122);
and (s0n3665,notn3665,n3666);
and (s1n3665,n3122,n3667);
and (n3668,n3669,n3136);
wire s0n3669,s1n3669,notn3669;
or (n3669,s0n3669,s1n3669);
not(notn3669,n3122);
and (s0n3669,notn3669,n3670);
and (s1n3669,n3122,n3666);
and (n3671,n3672,n3141);
wire s0n3672,s1n3672,notn3672;
or (n3672,s0n3672,s1n3672);
not(notn3672,n3122);
and (s0n3672,notn3672,n3673);
and (s1n3672,n3122,n3670);
and (n3674,n3675,n3146);
wire s0n3675,s1n3675,notn3675;
or (n3675,s0n3675,s1n3675);
not(notn3675,n3122);
and (s0n3675,notn3675,n3676);
and (s1n3675,n3122,n3673);
and (n3677,n3678,n1042);
or (n3678,1'b0,n3679,n3682,n3685,n3688);
and (n3679,n3680,n3124);
wire s0n3680,s1n3680,notn3680;
or (n3680,s0n3680,s1n3680);
not(notn3680,n3122);
and (s0n3680,notn3680,n3681);
and (s1n3680,n3122,n3676);
and (n3682,n3683,n3136);
wire s0n3683,s1n3683,notn3683;
or (n3683,s0n3683,s1n3683);
not(notn3683,n3122);
and (s0n3683,notn3683,n3684);
and (s1n3683,n3122,n3681);
and (n3685,n3686,n3141);
wire s0n3686,s1n3686,notn3686;
or (n3686,s0n3686,s1n3686);
not(notn3686,n3122);
and (s0n3686,notn3686,n3687);
and (s1n3686,n3122,n3684);
and (n3688,n3689,n3146);
wire s0n3689,s1n3689,notn3689;
or (n3689,s0n3689,s1n3689);
not(notn3689,n3122);
and (s0n3689,notn3689,n3690);
and (s1n3689,n3122,n3687);
wire s0n3692,s1n3692,notn3692;
or (n3692,s0n3692,s1n3692);
not(notn3692,n3074);
and (s0n3692,notn3692,n3693);
and (s1n3692,n3074,n3752);
or (n3693,1'b0,n3694,n3709,n3723,n3738);
and (n3694,n3695,n981);
or (n3695,1'b0,n3696,n3700,n3703,n3706);
and (n3696,n3697,n3124);
wire s0n3697,s1n3697,notn3697;
or (n3697,s0n3697,s1n3697);
not(notn3697,n3122);
and (s0n3697,notn3697,n3698);
and (s1n3697,n3122,n3699);
and (n3700,n3701,n3136);
wire s0n3701,s1n3701,notn3701;
or (n3701,s0n3701,s1n3701);
not(notn3701,n3122);
and (s0n3701,notn3701,n3702);
and (s1n3701,n3122,n3698);
and (n3703,n3704,n3141);
wire s0n3704,s1n3704,notn3704;
or (n3704,s0n3704,s1n3704);
not(notn3704,n3122);
and (s0n3704,notn3704,n3705);
and (s1n3704,n3122,n3702);
and (n3706,n3707,n3146);
wire s0n3707,s1n3707,notn3707;
or (n3707,s0n3707,s1n3707);
not(notn3707,n3122);
and (s0n3707,notn3707,n3708);
and (s1n3707,n3122,n3705);
and (n3709,n3710,n1002);
or (n3710,1'b0,n3711,n3714,n3717,n3720);
and (n3711,n3712,n3124);
wire s0n3712,s1n3712,notn3712;
or (n3712,s0n3712,s1n3712);
not(notn3712,n3122);
and (s0n3712,notn3712,n3713);
and (s1n3712,n3122,n3708);
and (n3714,n3715,n3136);
wire s0n3715,s1n3715,notn3715;
or (n3715,s0n3715,s1n3715);
not(notn3715,n3122);
and (s0n3715,notn3715,n3716);
and (s1n3715,n3122,n3713);
and (n3717,n3718,n3141);
wire s0n3718,s1n3718,notn3718;
or (n3718,s0n3718,s1n3718);
not(notn3718,n3122);
and (s0n3718,notn3718,n3719);
and (s1n3718,n3122,n3716);
and (n3720,n3721,n3146);
wire s0n3721,s1n3721,notn3721;
or (n3721,s0n3721,s1n3721);
not(notn3721,n3122);
and (s0n3721,notn3721,n3722);
and (s1n3721,n3122,n3719);
and (n3723,n3724,n1022);
or (n3724,1'b0,n3725,n3729,n3732,n3735);
and (n3725,n3726,n3124);
wire s0n3726,s1n3726,notn3726;
or (n3726,s0n3726,s1n3726);
not(notn3726,n3122);
and (s0n3726,notn3726,n3727);
and (s1n3726,n3122,n3728);
and (n3729,n3730,n3136);
wire s0n3730,s1n3730,notn3730;
or (n3730,s0n3730,s1n3730);
not(notn3730,n3122);
and (s0n3730,notn3730,n3731);
and (s1n3730,n3122,n3727);
and (n3732,n3733,n3141);
wire s0n3733,s1n3733,notn3733;
or (n3733,s0n3733,s1n3733);
not(notn3733,n3122);
and (s0n3733,notn3733,n3734);
and (s1n3733,n3122,n3731);
and (n3735,n3736,n3146);
wire s0n3736,s1n3736,notn3736;
or (n3736,s0n3736,s1n3736);
not(notn3736,n3122);
and (s0n3736,notn3736,n3737);
and (s1n3736,n3122,n3734);
and (n3738,n3739,n1042);
or (n3739,1'b0,n3740,n3743,n3746,n3749);
and (n3740,n3741,n3124);
wire s0n3741,s1n3741,notn3741;
or (n3741,s0n3741,s1n3741);
not(notn3741,n3122);
and (s0n3741,notn3741,n3742);
and (s1n3741,n3122,n3737);
and (n3743,n3744,n3136);
wire s0n3744,s1n3744,notn3744;
or (n3744,s0n3744,s1n3744);
not(notn3744,n3122);
and (s0n3744,notn3744,n3745);
and (s1n3744,n3122,n3742);
and (n3746,n3747,n3141);
wire s0n3747,s1n3747,notn3747;
or (n3747,s0n3747,s1n3747);
not(notn3747,n3122);
and (s0n3747,notn3747,n3748);
and (s1n3747,n3122,n3745);
and (n3749,n3750,n3146);
wire s0n3750,s1n3750,notn3750;
or (n3750,s0n3750,s1n3750);
not(notn3750,n3122);
and (s0n3750,notn3750,n3751);
and (s1n3750,n3122,n3748);
and (n3753,n3692,n3754);
or (n3754,n3755,n3878,n4128);
and (n3755,n3756,n3817);
wire s0n3756,s1n3756,notn3756;
or (n3756,s0n3756,s1n3756);
not(notn3756,n3074);
and (s0n3756,notn3756,n3757);
and (s1n3756,n3074,n3816);
or (n3757,1'b0,n3758,n3773,n3787,n3802);
and (n3758,n3759,n981);
or (n3759,1'b0,n3760,n3764,n3767,n3770);
and (n3760,n3761,n3124);
wire s0n3761,s1n3761,notn3761;
or (n3761,s0n3761,s1n3761);
not(notn3761,n3122);
and (s0n3761,notn3761,n3762);
and (s1n3761,n3122,n3763);
and (n3764,n3765,n3136);
wire s0n3765,s1n3765,notn3765;
or (n3765,s0n3765,s1n3765);
not(notn3765,n3122);
and (s0n3765,notn3765,n3766);
and (s1n3765,n3122,n3762);
and (n3767,n3768,n3141);
wire s0n3768,s1n3768,notn3768;
or (n3768,s0n3768,s1n3768);
not(notn3768,n3122);
and (s0n3768,notn3768,n3769);
and (s1n3768,n3122,n3766);
and (n3770,n3771,n3146);
wire s0n3771,s1n3771,notn3771;
or (n3771,s0n3771,s1n3771);
not(notn3771,n3122);
and (s0n3771,notn3771,n3772);
and (s1n3771,n3122,n3769);
and (n3773,n3774,n1002);
or (n3774,1'b0,n3775,n3778,n3781,n3784);
and (n3775,n3776,n3124);
wire s0n3776,s1n3776,notn3776;
or (n3776,s0n3776,s1n3776);
not(notn3776,n3122);
and (s0n3776,notn3776,n3777);
and (s1n3776,n3122,n3772);
and (n3778,n3779,n3136);
wire s0n3779,s1n3779,notn3779;
or (n3779,s0n3779,s1n3779);
not(notn3779,n3122);
and (s0n3779,notn3779,n3780);
and (s1n3779,n3122,n3777);
and (n3781,n3782,n3141);
wire s0n3782,s1n3782,notn3782;
or (n3782,s0n3782,s1n3782);
not(notn3782,n3122);
and (s0n3782,notn3782,n3783);
and (s1n3782,n3122,n3780);
and (n3784,n3785,n3146);
wire s0n3785,s1n3785,notn3785;
or (n3785,s0n3785,s1n3785);
not(notn3785,n3122);
and (s0n3785,notn3785,n3786);
and (s1n3785,n3122,n3783);
and (n3787,n3788,n1022);
or (n3788,1'b0,n3789,n3793,n3796,n3799);
and (n3789,n3790,n3124);
wire s0n3790,s1n3790,notn3790;
or (n3790,s0n3790,s1n3790);
not(notn3790,n3122);
and (s0n3790,notn3790,n3791);
and (s1n3790,n3122,n3792);
and (n3793,n3794,n3136);
wire s0n3794,s1n3794,notn3794;
or (n3794,s0n3794,s1n3794);
not(notn3794,n3122);
and (s0n3794,notn3794,n3795);
and (s1n3794,n3122,n3791);
and (n3796,n3797,n3141);
wire s0n3797,s1n3797,notn3797;
or (n3797,s0n3797,s1n3797);
not(notn3797,n3122);
and (s0n3797,notn3797,n3798);
and (s1n3797,n3122,n3795);
and (n3799,n3800,n3146);
wire s0n3800,s1n3800,notn3800;
or (n3800,s0n3800,s1n3800);
not(notn3800,n3122);
and (s0n3800,notn3800,n3801);
and (s1n3800,n3122,n3798);
and (n3802,n3803,n1042);
or (n3803,1'b0,n3804,n3807,n3810,n3813);
and (n3804,n3805,n3124);
wire s0n3805,s1n3805,notn3805;
or (n3805,s0n3805,s1n3805);
not(notn3805,n3122);
and (s0n3805,notn3805,n3806);
and (s1n3805,n3122,n3801);
and (n3807,n3808,n3136);
wire s0n3808,s1n3808,notn3808;
or (n3808,s0n3808,s1n3808);
not(notn3808,n3122);
and (s0n3808,notn3808,n3809);
and (s1n3808,n3122,n3806);
and (n3810,n3811,n3141);
wire s0n3811,s1n3811,notn3811;
or (n3811,s0n3811,s1n3811);
not(notn3811,n3122);
and (s0n3811,notn3811,n3812);
and (s1n3811,n3122,n3809);
and (n3813,n3814,n3146);
wire s0n3814,s1n3814,notn3814;
or (n3814,s0n3814,s1n3814);
not(notn3814,n3122);
and (s0n3814,notn3814,n3815);
and (s1n3814,n3122,n3812);
wire s0n3817,s1n3817,notn3817;
or (n3817,s0n3817,s1n3817);
not(notn3817,n3074);
and (s0n3817,notn3817,n3818);
and (s1n3817,n3074,n3877);
or (n3818,1'b0,n3819,n3834,n3848,n3863);
and (n3819,n3820,n981);
or (n3820,1'b0,n3821,n3825,n3828,n3831);
and (n3821,n3822,n3124);
wire s0n3822,s1n3822,notn3822;
or (n3822,s0n3822,s1n3822);
not(notn3822,n3122);
and (s0n3822,notn3822,n3823);
and (s1n3822,n3122,n3824);
and (n3825,n3826,n3136);
wire s0n3826,s1n3826,notn3826;
or (n3826,s0n3826,s1n3826);
not(notn3826,n3122);
and (s0n3826,notn3826,n3827);
and (s1n3826,n3122,n3823);
and (n3828,n3829,n3141);
wire s0n3829,s1n3829,notn3829;
or (n3829,s0n3829,s1n3829);
not(notn3829,n3122);
and (s0n3829,notn3829,n3830);
and (s1n3829,n3122,n3827);
and (n3831,n3832,n3146);
wire s0n3832,s1n3832,notn3832;
or (n3832,s0n3832,s1n3832);
not(notn3832,n3122);
and (s0n3832,notn3832,n3833);
and (s1n3832,n3122,n3830);
and (n3834,n3835,n1002);
or (n3835,1'b0,n3836,n3839,n3842,n3845);
and (n3836,n3837,n3124);
wire s0n3837,s1n3837,notn3837;
or (n3837,s0n3837,s1n3837);
not(notn3837,n3122);
and (s0n3837,notn3837,n3838);
and (s1n3837,n3122,n3833);
and (n3839,n3840,n3136);
wire s0n3840,s1n3840,notn3840;
or (n3840,s0n3840,s1n3840);
not(notn3840,n3122);
and (s0n3840,notn3840,n3841);
and (s1n3840,n3122,n3838);
and (n3842,n3843,n3141);
wire s0n3843,s1n3843,notn3843;
or (n3843,s0n3843,s1n3843);
not(notn3843,n3122);
and (s0n3843,notn3843,n3844);
and (s1n3843,n3122,n3841);
and (n3845,n3846,n3146);
wire s0n3846,s1n3846,notn3846;
or (n3846,s0n3846,s1n3846);
not(notn3846,n3122);
and (s0n3846,notn3846,n3847);
and (s1n3846,n3122,n3844);
and (n3848,n3849,n1022);
or (n3849,1'b0,n3850,n3854,n3857,n3860);
and (n3850,n3851,n3124);
wire s0n3851,s1n3851,notn3851;
or (n3851,s0n3851,s1n3851);
not(notn3851,n3122);
and (s0n3851,notn3851,n3852);
and (s1n3851,n3122,n3853);
and (n3854,n3855,n3136);
wire s0n3855,s1n3855,notn3855;
or (n3855,s0n3855,s1n3855);
not(notn3855,n3122);
and (s0n3855,notn3855,n3856);
and (s1n3855,n3122,n3852);
and (n3857,n3858,n3141);
wire s0n3858,s1n3858,notn3858;
or (n3858,s0n3858,s1n3858);
not(notn3858,n3122);
and (s0n3858,notn3858,n3859);
and (s1n3858,n3122,n3856);
and (n3860,n3861,n3146);
wire s0n3861,s1n3861,notn3861;
or (n3861,s0n3861,s1n3861);
not(notn3861,n3122);
and (s0n3861,notn3861,n3862);
and (s1n3861,n3122,n3859);
and (n3863,n3864,n1042);
or (n3864,1'b0,n3865,n3868,n3871,n3874);
and (n3865,n3866,n3124);
wire s0n3866,s1n3866,notn3866;
or (n3866,s0n3866,s1n3866);
not(notn3866,n3122);
and (s0n3866,notn3866,n3867);
and (s1n3866,n3122,n3862);
and (n3868,n3869,n3136);
wire s0n3869,s1n3869,notn3869;
or (n3869,s0n3869,s1n3869);
not(notn3869,n3122);
and (s0n3869,notn3869,n3870);
and (s1n3869,n3122,n3867);
and (n3871,n3872,n3141);
wire s0n3872,s1n3872,notn3872;
or (n3872,s0n3872,s1n3872);
not(notn3872,n3122);
and (s0n3872,notn3872,n3873);
and (s1n3872,n3122,n3870);
and (n3874,n3875,n3146);
wire s0n3875,s1n3875,notn3875;
or (n3875,s0n3875,s1n3875);
not(notn3875,n3122);
and (s0n3875,notn3875,n3876);
and (s1n3875,n3122,n3873);
and (n3878,n3817,n3879);
or (n3879,n3880,n4003,n4127);
and (n3880,n3881,n3942);
wire s0n3881,s1n3881,notn3881;
or (n3881,s0n3881,s1n3881);
not(notn3881,n3074);
and (s0n3881,notn3881,n3882);
and (s1n3881,n3074,n3941);
or (n3882,1'b0,n3883,n3898,n3912,n3927);
and (n3883,n3884,n981);
or (n3884,1'b0,n3885,n3889,n3892,n3895);
and (n3885,n3886,n3124);
wire s0n3886,s1n3886,notn3886;
or (n3886,s0n3886,s1n3886);
not(notn3886,n3122);
and (s0n3886,notn3886,n3887);
and (s1n3886,n3122,n3888);
and (n3889,n3890,n3136);
wire s0n3890,s1n3890,notn3890;
or (n3890,s0n3890,s1n3890);
not(notn3890,n3122);
and (s0n3890,notn3890,n3891);
and (s1n3890,n3122,n3887);
and (n3892,n3893,n3141);
wire s0n3893,s1n3893,notn3893;
or (n3893,s0n3893,s1n3893);
not(notn3893,n3122);
and (s0n3893,notn3893,n3894);
and (s1n3893,n3122,n3891);
and (n3895,n3896,n3146);
wire s0n3896,s1n3896,notn3896;
or (n3896,s0n3896,s1n3896);
not(notn3896,n3122);
and (s0n3896,notn3896,n3897);
and (s1n3896,n3122,n3894);
and (n3898,n3899,n1002);
or (n3899,1'b0,n3900,n3903,n3906,n3909);
and (n3900,n3901,n3124);
wire s0n3901,s1n3901,notn3901;
or (n3901,s0n3901,s1n3901);
not(notn3901,n3122);
and (s0n3901,notn3901,n3902);
and (s1n3901,n3122,n3897);
and (n3903,n3904,n3136);
wire s0n3904,s1n3904,notn3904;
or (n3904,s0n3904,s1n3904);
not(notn3904,n3122);
and (s0n3904,notn3904,n3905);
and (s1n3904,n3122,n3902);
and (n3906,n3907,n3141);
wire s0n3907,s1n3907,notn3907;
or (n3907,s0n3907,s1n3907);
not(notn3907,n3122);
and (s0n3907,notn3907,n3908);
and (s1n3907,n3122,n3905);
and (n3909,n3910,n3146);
wire s0n3910,s1n3910,notn3910;
or (n3910,s0n3910,s1n3910);
not(notn3910,n3122);
and (s0n3910,notn3910,n3911);
and (s1n3910,n3122,n3908);
and (n3912,n3913,n1022);
or (n3913,1'b0,n3914,n3918,n3921,n3924);
and (n3914,n3915,n3124);
wire s0n3915,s1n3915,notn3915;
or (n3915,s0n3915,s1n3915);
not(notn3915,n3122);
and (s0n3915,notn3915,n3916);
and (s1n3915,n3122,n3917);
and (n3918,n3919,n3136);
wire s0n3919,s1n3919,notn3919;
or (n3919,s0n3919,s1n3919);
not(notn3919,n3122);
and (s0n3919,notn3919,n3920);
and (s1n3919,n3122,n3916);
and (n3921,n3922,n3141);
wire s0n3922,s1n3922,notn3922;
or (n3922,s0n3922,s1n3922);
not(notn3922,n3122);
and (s0n3922,notn3922,n3923);
and (s1n3922,n3122,n3920);
and (n3924,n3925,n3146);
wire s0n3925,s1n3925,notn3925;
or (n3925,s0n3925,s1n3925);
not(notn3925,n3122);
and (s0n3925,notn3925,n3926);
and (s1n3925,n3122,n3923);
and (n3927,n3928,n1042);
or (n3928,1'b0,n3929,n3932,n3935,n3938);
and (n3929,n3930,n3124);
wire s0n3930,s1n3930,notn3930;
or (n3930,s0n3930,s1n3930);
not(notn3930,n3122);
and (s0n3930,notn3930,n3931);
and (s1n3930,n3122,n3926);
and (n3932,n3933,n3136);
wire s0n3933,s1n3933,notn3933;
or (n3933,s0n3933,s1n3933);
not(notn3933,n3122);
and (s0n3933,notn3933,n3934);
and (s1n3933,n3122,n3931);
and (n3935,n3936,n3141);
wire s0n3936,s1n3936,notn3936;
or (n3936,s0n3936,s1n3936);
not(notn3936,n3122);
and (s0n3936,notn3936,n3937);
and (s1n3936,n3122,n3934);
and (n3938,n3939,n3146);
wire s0n3939,s1n3939,notn3939;
or (n3939,s0n3939,s1n3939);
not(notn3939,n3122);
and (s0n3939,notn3939,n3940);
and (s1n3939,n3122,n3937);
wire s0n3942,s1n3942,notn3942;
or (n3942,s0n3942,s1n3942);
not(notn3942,n3074);
and (s0n3942,notn3942,n3943);
and (s1n3942,n3074,n4002);
or (n3943,1'b0,n3944,n3959,n3973,n3988);
and (n3944,n3945,n981);
or (n3945,1'b0,n3946,n3950,n3953,n3956);
and (n3946,n3947,n3124);
wire s0n3947,s1n3947,notn3947;
or (n3947,s0n3947,s1n3947);
not(notn3947,n3122);
and (s0n3947,notn3947,n3948);
and (s1n3947,n3122,n3949);
and (n3950,n3951,n3136);
wire s0n3951,s1n3951,notn3951;
or (n3951,s0n3951,s1n3951);
not(notn3951,n3122);
and (s0n3951,notn3951,n3952);
and (s1n3951,n3122,n3948);
and (n3953,n3954,n3141);
wire s0n3954,s1n3954,notn3954;
or (n3954,s0n3954,s1n3954);
not(notn3954,n3122);
and (s0n3954,notn3954,n3955);
and (s1n3954,n3122,n3952);
and (n3956,n3957,n3146);
wire s0n3957,s1n3957,notn3957;
or (n3957,s0n3957,s1n3957);
not(notn3957,n3122);
and (s0n3957,notn3957,n3958);
and (s1n3957,n3122,n3955);
and (n3959,n3960,n1002);
or (n3960,1'b0,n3961,n3964,n3967,n3970);
and (n3961,n3962,n3124);
wire s0n3962,s1n3962,notn3962;
or (n3962,s0n3962,s1n3962);
not(notn3962,n3122);
and (s0n3962,notn3962,n3963);
and (s1n3962,n3122,n3958);
and (n3964,n3965,n3136);
wire s0n3965,s1n3965,notn3965;
or (n3965,s0n3965,s1n3965);
not(notn3965,n3122);
and (s0n3965,notn3965,n3966);
and (s1n3965,n3122,n3963);
and (n3967,n3968,n3141);
wire s0n3968,s1n3968,notn3968;
or (n3968,s0n3968,s1n3968);
not(notn3968,n3122);
and (s0n3968,notn3968,n3969);
and (s1n3968,n3122,n3966);
and (n3970,n3971,n3146);
wire s0n3971,s1n3971,notn3971;
or (n3971,s0n3971,s1n3971);
not(notn3971,n3122);
and (s0n3971,notn3971,n3972);
and (s1n3971,n3122,n3969);
and (n3973,n3974,n1022);
or (n3974,1'b0,n3975,n3979,n3982,n3985);
and (n3975,n3976,n3124);
wire s0n3976,s1n3976,notn3976;
or (n3976,s0n3976,s1n3976);
not(notn3976,n3122);
and (s0n3976,notn3976,n3977);
and (s1n3976,n3122,n3978);
and (n3979,n3980,n3136);
wire s0n3980,s1n3980,notn3980;
or (n3980,s0n3980,s1n3980);
not(notn3980,n3122);
and (s0n3980,notn3980,n3981);
and (s1n3980,n3122,n3977);
and (n3982,n3983,n3141);
wire s0n3983,s1n3983,notn3983;
or (n3983,s0n3983,s1n3983);
not(notn3983,n3122);
and (s0n3983,notn3983,n3984);
and (s1n3983,n3122,n3981);
and (n3985,n3986,n3146);
wire s0n3986,s1n3986,notn3986;
or (n3986,s0n3986,s1n3986);
not(notn3986,n3122);
and (s0n3986,notn3986,n3987);
and (s1n3986,n3122,n3984);
and (n3988,n3989,n1042);
or (n3989,1'b0,n3990,n3993,n3996,n3999);
and (n3990,n3991,n3124);
wire s0n3991,s1n3991,notn3991;
or (n3991,s0n3991,s1n3991);
not(notn3991,n3122);
and (s0n3991,notn3991,n3992);
and (s1n3991,n3122,n3987);
and (n3993,n3994,n3136);
wire s0n3994,s1n3994,notn3994;
or (n3994,s0n3994,s1n3994);
not(notn3994,n3122);
and (s0n3994,notn3994,n3995);
and (s1n3994,n3122,n3992);
and (n3996,n3997,n3141);
wire s0n3997,s1n3997,notn3997;
or (n3997,s0n3997,s1n3997);
not(notn3997,n3122);
and (s0n3997,notn3997,n3998);
and (s1n3997,n3122,n3995);
and (n3999,n4000,n3146);
wire s0n4000,s1n4000,notn4000;
or (n4000,s0n4000,s1n4000);
not(notn4000,n3122);
and (s0n4000,notn4000,n4001);
and (s1n4000,n3122,n3998);
and (n4003,n3942,n4004);
and (n4004,n4005,n4066);
wire s0n4005,s1n4005,notn4005;
or (n4005,s0n4005,s1n4005);
not(notn4005,n3074);
and (s0n4005,notn4005,n4006);
and (s1n4005,n3074,n4065);
or (n4006,1'b0,n4007,n4022,n4036,n4051);
and (n4007,n4008,n981);
or (n4008,1'b0,n4009,n4013,n4016,n4019);
and (n4009,n4010,n3124);
wire s0n4010,s1n4010,notn4010;
or (n4010,s0n4010,s1n4010);
not(notn4010,n3122);
and (s0n4010,notn4010,n4011);
and (s1n4010,n3122,n4012);
and (n4013,n4014,n3136);
wire s0n4014,s1n4014,notn4014;
or (n4014,s0n4014,s1n4014);
not(notn4014,n3122);
and (s0n4014,notn4014,n4015);
and (s1n4014,n3122,n4011);
and (n4016,n4017,n3141);
wire s0n4017,s1n4017,notn4017;
or (n4017,s0n4017,s1n4017);
not(notn4017,n3122);
and (s0n4017,notn4017,n4018);
and (s1n4017,n3122,n4015);
and (n4019,n4020,n3146);
wire s0n4020,s1n4020,notn4020;
or (n4020,s0n4020,s1n4020);
not(notn4020,n3122);
and (s0n4020,notn4020,n4021);
and (s1n4020,n3122,n4018);
and (n4022,n4023,n1002);
or (n4023,1'b0,n4024,n4027,n4030,n4033);
and (n4024,n4025,n3124);
wire s0n4025,s1n4025,notn4025;
or (n4025,s0n4025,s1n4025);
not(notn4025,n3122);
and (s0n4025,notn4025,n4026);
and (s1n4025,n3122,n4021);
and (n4027,n4028,n3136);
wire s0n4028,s1n4028,notn4028;
or (n4028,s0n4028,s1n4028);
not(notn4028,n3122);
and (s0n4028,notn4028,n4029);
and (s1n4028,n3122,n4026);
and (n4030,n4031,n3141);
wire s0n4031,s1n4031,notn4031;
or (n4031,s0n4031,s1n4031);
not(notn4031,n3122);
and (s0n4031,notn4031,n4032);
and (s1n4031,n3122,n4029);
and (n4033,n4034,n3146);
wire s0n4034,s1n4034,notn4034;
or (n4034,s0n4034,s1n4034);
not(notn4034,n3122);
and (s0n4034,notn4034,n4035);
and (s1n4034,n3122,n4032);
and (n4036,n4037,n1022);
or (n4037,1'b0,n4038,n4042,n4045,n4048);
and (n4038,n4039,n3124);
wire s0n4039,s1n4039,notn4039;
or (n4039,s0n4039,s1n4039);
not(notn4039,n3122);
and (s0n4039,notn4039,n4040);
and (s1n4039,n3122,n4041);
and (n4042,n4043,n3136);
wire s0n4043,s1n4043,notn4043;
or (n4043,s0n4043,s1n4043);
not(notn4043,n3122);
and (s0n4043,notn4043,n4044);
and (s1n4043,n3122,n4040);
and (n4045,n4046,n3141);
wire s0n4046,s1n4046,notn4046;
or (n4046,s0n4046,s1n4046);
not(notn4046,n3122);
and (s0n4046,notn4046,n4047);
and (s1n4046,n3122,n4044);
and (n4048,n4049,n3146);
wire s0n4049,s1n4049,notn4049;
or (n4049,s0n4049,s1n4049);
not(notn4049,n3122);
and (s0n4049,notn4049,n4050);
and (s1n4049,n3122,n4047);
and (n4051,n4052,n1042);
or (n4052,1'b0,n4053,n4056,n4059,n4062);
and (n4053,n4054,n3124);
wire s0n4054,s1n4054,notn4054;
or (n4054,s0n4054,s1n4054);
not(notn4054,n3122);
and (s0n4054,notn4054,n4055);
and (s1n4054,n3122,n4050);
and (n4056,n4057,n3136);
wire s0n4057,s1n4057,notn4057;
or (n4057,s0n4057,s1n4057);
not(notn4057,n3122);
and (s0n4057,notn4057,n4058);
and (s1n4057,n3122,n4055);
and (n4059,n4060,n3141);
wire s0n4060,s1n4060,notn4060;
or (n4060,s0n4060,s1n4060);
not(notn4060,n3122);
and (s0n4060,notn4060,n4061);
and (s1n4060,n3122,n4058);
and (n4062,n4063,n3146);
wire s0n4063,s1n4063,notn4063;
or (n4063,s0n4063,s1n4063);
not(notn4063,n3122);
and (s0n4063,notn4063,n4064);
and (s1n4063,n3122,n4061);
wire s0n4066,s1n4066,notn4066;
or (n4066,s0n4066,s1n4066);
not(notn4066,n3074);
and (s0n4066,notn4066,n4067);
and (s1n4066,n3074,n4126);
or (n4067,1'b0,n4068,n4083,n4097,n4112);
and (n4068,n4069,n981);
or (n4069,1'b0,n4070,n4074,n4077,n4080);
and (n4070,n4071,n3124);
wire s0n4071,s1n4071,notn4071;
or (n4071,s0n4071,s1n4071);
not(notn4071,n3122);
and (s0n4071,notn4071,n4072);
and (s1n4071,n3122,n4073);
and (n4074,n4075,n3136);
wire s0n4075,s1n4075,notn4075;
or (n4075,s0n4075,s1n4075);
not(notn4075,n3122);
and (s0n4075,notn4075,n4076);
and (s1n4075,n3122,n4072);
and (n4077,n4078,n3141);
wire s0n4078,s1n4078,notn4078;
or (n4078,s0n4078,s1n4078);
not(notn4078,n3122);
and (s0n4078,notn4078,n4079);
and (s1n4078,n3122,n4076);
and (n4080,n4081,n3146);
wire s0n4081,s1n4081,notn4081;
or (n4081,s0n4081,s1n4081);
not(notn4081,n3122);
and (s0n4081,notn4081,n4082);
and (s1n4081,n3122,n4079);
and (n4083,n4084,n1002);
or (n4084,1'b0,n4085,n4088,n4091,n4094);
and (n4085,n4086,n3124);
wire s0n4086,s1n4086,notn4086;
or (n4086,s0n4086,s1n4086);
not(notn4086,n3122);
and (s0n4086,notn4086,n4087);
and (s1n4086,n3122,n4082);
and (n4088,n4089,n3136);
wire s0n4089,s1n4089,notn4089;
or (n4089,s0n4089,s1n4089);
not(notn4089,n3122);
and (s0n4089,notn4089,n4090);
and (s1n4089,n3122,n4087);
and (n4091,n4092,n3141);
wire s0n4092,s1n4092,notn4092;
or (n4092,s0n4092,s1n4092);
not(notn4092,n3122);
and (s0n4092,notn4092,n4093);
and (s1n4092,n3122,n4090);
and (n4094,n4095,n3146);
wire s0n4095,s1n4095,notn4095;
or (n4095,s0n4095,s1n4095);
not(notn4095,n3122);
and (s0n4095,notn4095,n4096);
and (s1n4095,n3122,n4093);
and (n4097,n4098,n1022);
or (n4098,1'b0,n4099,n4103,n4106,n4109);
and (n4099,n4100,n3124);
wire s0n4100,s1n4100,notn4100;
or (n4100,s0n4100,s1n4100);
not(notn4100,n3122);
and (s0n4100,notn4100,n4101);
and (s1n4100,n3122,n4102);
and (n4103,n4104,n3136);
wire s0n4104,s1n4104,notn4104;
or (n4104,s0n4104,s1n4104);
not(notn4104,n3122);
and (s0n4104,notn4104,n4105);
and (s1n4104,n3122,n4101);
and (n4106,n4107,n3141);
wire s0n4107,s1n4107,notn4107;
or (n4107,s0n4107,s1n4107);
not(notn4107,n3122);
and (s0n4107,notn4107,n4108);
and (s1n4107,n3122,n4105);
and (n4109,n4110,n3146);
wire s0n4110,s1n4110,notn4110;
or (n4110,s0n4110,s1n4110);
not(notn4110,n3122);
and (s0n4110,notn4110,n4111);
and (s1n4110,n3122,n4108);
and (n4112,n4113,n1042);
or (n4113,1'b0,n4114,n4117,n4120,n4123);
and (n4114,n4115,n3124);
wire s0n4115,s1n4115,notn4115;
or (n4115,s0n4115,s1n4115);
not(notn4115,n3122);
and (s0n4115,notn4115,n4116);
and (s1n4115,n3122,n4111);
and (n4117,n4118,n3136);
wire s0n4118,s1n4118,notn4118;
or (n4118,s0n4118,s1n4118);
not(notn4118,n3122);
and (s0n4118,notn4118,n4119);
and (s1n4118,n3122,n4116);
and (n4120,n4121,n3141);
wire s0n4121,s1n4121,notn4121;
or (n4121,s0n4121,s1n4121);
not(notn4121,n3122);
and (s0n4121,notn4121,n4122);
and (s1n4121,n3122,n4119);
and (n4123,n4124,n3146);
wire s0n4124,s1n4124,notn4124;
or (n4124,s0n4124,s1n4124);
not(notn4124,n3122);
and (s0n4124,notn4124,n4125);
and (s1n4124,n3122,n4122);
and (n4127,n3881,n4004);
and (n4128,n3756,n3879);
and (n4129,n3631,n3754);
and (n4130,n3506,n3629);
and (n4131,n3381,n3504);
and (n4132,n3256,n3379);
and (n4133,n3114,n3254);
and (n4134,n3107,n3112);
and (n4135,n3100,n3105);
and (n4136,n3093,n3098);
and (n4137,n3086,n3091);
xor (n4138,n4139,n5578);
xor (n4139,n4140,n5492);
xor (n4140,n4141,n4880);
xor (n4141,n4142,n4147);
xor (n4142,n4143,n4145);
wire s0n4143,s1n4143,notn4143;
or (n4143,s0n4143,s1n4143);
not(notn4143,n3074);
and (s0n4143,notn4143,1'b0);
and (s1n4143,n3074,n4144);
wire s0n4145,s1n4145,notn4145;
or (n4145,s0n4145,s1n4145);
not(notn4145,n3074);
and (s0n4145,notn4145,1'b0);
and (s1n4145,n3074,n4146);
or (n4147,n4148,n4153,n4879);
and (n4148,n4149,n4151);
wire s0n4149,s1n4149,notn4149;
or (n4149,s0n4149,s1n4149);
not(notn4149,n3074);
and (s0n4149,notn4149,1'b0);
and (s1n4149,n3074,n4150);
wire s0n4151,s1n4151,notn4151;
or (n4151,s0n4151,s1n4151);
not(notn4151,n3074);
and (s0n4151,notn4151,1'b0);
and (s1n4151,n3074,n4152);
and (n4153,n4151,n4154);
or (n4154,n4155,n4160,n4878);
and (n4155,n4156,n4158);
wire s0n4156,s1n4156,notn4156;
or (n4156,s0n4156,s1n4156);
not(notn4156,n3074);
and (s0n4156,notn4156,1'b0);
and (s1n4156,n3074,n4157);
wire s0n4158,s1n4158,notn4158;
or (n4158,s0n4158,s1n4158);
not(notn4158,n3074);
and (s0n4158,notn4158,1'b0);
and (s1n4158,n3074,n4159);
and (n4160,n4158,n4161);
or (n4161,n4162,n4249,n4877);
and (n4162,n4163,n4206);
wire s0n4163,s1n4163,notn4163;
or (n4163,s0n4163,s1n4163);
not(notn4163,n3074);
and (s0n4163,notn4163,n4164);
and (s1n4163,n3074,n4205);
or (n4164,1'b0,n4165,n4175,n4185,n4195);
and (n4165,n4166,n981);
or (n4166,1'b0,n4167,n4169,n4171,n4173);
and (n4167,n4168,n3124);
wire s0n4168,s1n4168,notn4168;
or (n4168,s0n4168,s1n4168);
not(notn4168,n3122);
and (s0n4168,notn4168,n925);
and (s1n4168,n3122,n1050);
and (n4169,n4170,n3136);
wire s0n4170,s1n4170,notn4170;
or (n4170,s0n4170,s1n4170);
not(notn4170,n3122);
and (s0n4170,notn4170,n953);
and (s1n4170,n3122,n925);
and (n4171,n4172,n3141);
wire s0n4172,s1n4172,notn4172;
or (n4172,s0n4172,s1n4172);
not(notn4172,n3122);
and (s0n4172,notn4172,n963);
and (s1n4172,n3122,n953);
and (n4173,n4174,n3146);
wire s0n4174,s1n4174,notn4174;
or (n4174,s0n4174,s1n4174);
not(notn4174,n3122);
and (s0n4174,notn4174,n973);
and (s1n4174,n3122,n963);
and (n4175,n4176,n1002);
or (n4176,1'b0,n4177,n4179,n4181,n4183);
and (n4177,n4178,n3124);
wire s0n4178,s1n4178,notn4178;
or (n4178,s0n4178,s1n4178);
not(notn4178,n3122);
and (s0n4178,notn4178,n988);
and (s1n4178,n3122,n973);
and (n4179,n4180,n3136);
wire s0n4180,s1n4180,notn4180;
or (n4180,s0n4180,s1n4180);
not(notn4180,n3122);
and (s0n4180,notn4180,n992);
and (s1n4180,n3122,n988);
and (n4181,n4182,n3141);
wire s0n4182,s1n4182,notn4182;
or (n4182,s0n4182,s1n4182);
not(notn4182,n3122);
and (s0n4182,notn4182,n996);
and (s1n4182,n3122,n992);
and (n4183,n4184,n3146);
wire s0n4184,s1n4184,notn4184;
or (n4184,s0n4184,s1n4184);
not(notn4184,n3122);
and (s0n4184,notn4184,n1000);
and (s1n4184,n3122,n996);
and (n4185,n4186,n1022);
or (n4186,1'b0,n4187,n4189,n4191,n4193);
and (n4187,n4188,n3124);
wire s0n4188,s1n4188,notn4188;
or (n4188,s0n4188,s1n4188);
not(notn4188,n3122);
and (s0n4188,notn4188,n1008);
and (s1n4188,n3122,n1065);
and (n4189,n4190,n3136);
wire s0n4190,s1n4190,notn4190;
or (n4190,s0n4190,s1n4190);
not(notn4190,n3122);
and (s0n4190,notn4190,n1012);
and (s1n4190,n3122,n1008);
and (n4191,n4192,n3141);
wire s0n4192,s1n4192,notn4192;
or (n4192,s0n4192,s1n4192);
not(notn4192,n3122);
and (s0n4192,notn4192,n1016);
and (s1n4192,n3122,n1012);
and (n4193,n4194,n3146);
wire s0n4194,s1n4194,notn4194;
or (n4194,s0n4194,s1n4194);
not(notn4194,n3122);
and (s0n4194,notn4194,n1020);
and (s1n4194,n3122,n1016);
and (n4195,n4196,n1042);
or (n4196,1'b0,n4197,n4199,n4201,n4203);
and (n4197,n4198,n3124);
wire s0n4198,s1n4198,notn4198;
or (n4198,s0n4198,s1n4198);
not(notn4198,n3122);
and (s0n4198,notn4198,n1028);
and (s1n4198,n3122,n1020);
and (n4199,n4200,n3136);
wire s0n4200,s1n4200,notn4200;
or (n4200,s0n4200,s1n4200);
not(notn4200,n3122);
and (s0n4200,notn4200,n1032);
and (s1n4200,n3122,n1028);
and (n4201,n4202,n3141);
wire s0n4202,s1n4202,notn4202;
or (n4202,s0n4202,s1n4202);
not(notn4202,n3122);
and (s0n4202,notn4202,n1036);
and (s1n4202,n3122,n1032);
and (n4203,n4204,n3146);
wire s0n4204,s1n4204,notn4204;
or (n4204,s0n4204,s1n4204);
not(notn4204,n3122);
and (s0n4204,notn4204,n1040);
and (s1n4204,n3122,n1036);
wire s0n4206,s1n4206,notn4206;
or (n4206,s0n4206,s1n4206);
not(notn4206,n3074);
and (s0n4206,notn4206,n4207);
and (s1n4206,n3074,n4248);
or (n4207,1'b0,n4208,n4218,n4228,n4238);
and (n4208,n4209,n981);
or (n4209,1'b0,n4210,n4212,n4214,n4216);
and (n4210,n4211,n3124);
wire s0n4211,s1n4211,notn4211;
or (n4211,s0n4211,s1n4211);
not(notn4211,n3122);
and (s0n4211,notn4211,n926);
and (s1n4211,n3122,n1051);
and (n4212,n4213,n3136);
wire s0n4213,s1n4213,notn4213;
or (n4213,s0n4213,s1n4213);
not(notn4213,n3122);
and (s0n4213,notn4213,n954);
and (s1n4213,n3122,n926);
and (n4214,n4215,n3141);
wire s0n4215,s1n4215,notn4215;
or (n4215,s0n4215,s1n4215);
not(notn4215,n3122);
and (s0n4215,notn4215,n964);
and (s1n4215,n3122,n954);
and (n4216,n4217,n3146);
wire s0n4217,s1n4217,notn4217;
or (n4217,s0n4217,s1n4217);
not(notn4217,n3122);
and (s0n4217,notn4217,n974);
and (s1n4217,n3122,n964);
and (n4218,n4219,n1002);
or (n4219,1'b0,n4220,n4222,n4224,n4226);
and (n4220,n4221,n3124);
wire s0n4221,s1n4221,notn4221;
or (n4221,s0n4221,s1n4221);
not(notn4221,n3122);
and (s0n4221,notn4221,n989);
and (s1n4221,n3122,n974);
and (n4222,n4223,n3136);
wire s0n4223,s1n4223,notn4223;
or (n4223,s0n4223,s1n4223);
not(notn4223,n3122);
and (s0n4223,notn4223,n993);
and (s1n4223,n3122,n989);
and (n4224,n4225,n3141);
wire s0n4225,s1n4225,notn4225;
or (n4225,s0n4225,s1n4225);
not(notn4225,n3122);
and (s0n4225,notn4225,n997);
and (s1n4225,n3122,n993);
and (n4226,n4227,n3146);
wire s0n4227,s1n4227,notn4227;
or (n4227,s0n4227,s1n4227);
not(notn4227,n3122);
and (s0n4227,notn4227,n1001);
and (s1n4227,n3122,n997);
and (n4228,n4229,n1022);
or (n4229,1'b0,n4230,n4232,n4234,n4236);
and (n4230,n4231,n3124);
wire s0n4231,s1n4231,notn4231;
or (n4231,s0n4231,s1n4231);
not(notn4231,n3122);
and (s0n4231,notn4231,n1009);
and (s1n4231,n3122,n1066);
and (n4232,n4233,n3136);
wire s0n4233,s1n4233,notn4233;
or (n4233,s0n4233,s1n4233);
not(notn4233,n3122);
and (s0n4233,notn4233,n1013);
and (s1n4233,n3122,n1009);
and (n4234,n4235,n3141);
wire s0n4235,s1n4235,notn4235;
or (n4235,s0n4235,s1n4235);
not(notn4235,n3122);
and (s0n4235,notn4235,n1017);
and (s1n4235,n3122,n1013);
and (n4236,n4237,n3146);
wire s0n4237,s1n4237,notn4237;
or (n4237,s0n4237,s1n4237);
not(notn4237,n3122);
and (s0n4237,notn4237,n1021);
and (s1n4237,n3122,n1017);
and (n4238,n4239,n1042);
or (n4239,1'b0,n4240,n4242,n4244,n4246);
and (n4240,n4241,n3124);
wire s0n4241,s1n4241,notn4241;
or (n4241,s0n4241,s1n4241);
not(notn4241,n3122);
and (s0n4241,notn4241,n1029);
and (s1n4241,n3122,n1021);
and (n4242,n4243,n3136);
wire s0n4243,s1n4243,notn4243;
or (n4243,s0n4243,s1n4243);
not(notn4243,n3122);
and (s0n4243,notn4243,n1033);
and (s1n4243,n3122,n1029);
and (n4244,n4245,n3141);
wire s0n4245,s1n4245,notn4245;
or (n4245,s0n4245,s1n4245);
not(notn4245,n3122);
and (s0n4245,notn4245,n1037);
and (s1n4245,n3122,n1033);
and (n4246,n4247,n3146);
wire s0n4247,s1n4247,notn4247;
or (n4247,s0n4247,s1n4247);
not(notn4247,n3122);
and (s0n4247,notn4247,n1041);
and (s1n4247,n3122,n1037);
and (n4249,n4206,n4250);
or (n4250,n4251,n4338,n4876);
and (n4251,n4252,n4295);
wire s0n4252,s1n4252,notn4252;
or (n4252,s0n4252,s1n4252);
not(notn4252,n3074);
and (s0n4252,notn4252,n4253);
and (s1n4252,n3074,n4294);
or (n4253,1'b0,n4254,n4264,n4274,n4284);
and (n4254,n4255,n981);
or (n4255,1'b0,n4256,n4258,n4260,n4262);
and (n4256,n4257,n3124);
wire s0n4257,s1n4257,notn4257;
or (n4257,s0n4257,s1n4257);
not(notn4257,n3122);
and (s0n4257,notn4257,n1084);
and (s1n4257,n3122,n1157);
and (n4258,n4259,n3136);
wire s0n4259,s1n4259,notn4259;
or (n4259,s0n4259,s1n4259);
not(notn4259,n3122);
and (s0n4259,notn4259,n1088);
and (s1n4259,n3122,n1084);
and (n4260,n4261,n3141);
wire s0n4261,s1n4261,notn4261;
or (n4261,s0n4261,s1n4261);
not(notn4261,n3122);
and (s0n4261,notn4261,n1092);
and (s1n4261,n3122,n1088);
and (n4262,n4263,n3146);
wire s0n4263,s1n4263,notn4263;
or (n4263,s0n4263,s1n4263);
not(notn4263,n3122);
and (s0n4263,notn4263,n1096);
and (s1n4263,n3122,n1092);
and (n4264,n4265,n1002);
or (n4265,1'b0,n4266,n4268,n4270,n4272);
and (n4266,n4267,n3124);
wire s0n4267,s1n4267,notn4267;
or (n4267,s0n4267,s1n4267);
not(notn4267,n3122);
and (s0n4267,notn4267,n1102);
and (s1n4267,n3122,n1096);
and (n4268,n4269,n3136);
wire s0n4269,s1n4269,notn4269;
or (n4269,s0n4269,s1n4269);
not(notn4269,n3122);
and (s0n4269,notn4269,n1106);
and (s1n4269,n3122,n1102);
and (n4270,n4271,n3141);
wire s0n4271,s1n4271,notn4271;
or (n4271,s0n4271,s1n4271);
not(notn4271,n3122);
and (s0n4271,notn4271,n1110);
and (s1n4271,n3122,n1106);
and (n4272,n4273,n3146);
wire s0n4273,s1n4273,notn4273;
or (n4273,s0n4273,s1n4273);
not(notn4273,n3122);
and (s0n4273,notn4273,n1114);
and (s1n4273,n3122,n1110);
and (n4274,n4275,n1022);
or (n4275,1'b0,n4276,n4278,n4280,n4282);
and (n4276,n4277,n3124);
wire s0n4277,s1n4277,notn4277;
or (n4277,s0n4277,s1n4277);
not(notn4277,n3122);
and (s0n4277,notn4277,n1120);
and (s1n4277,n3122,n1172);
and (n4278,n4279,n3136);
wire s0n4279,s1n4279,notn4279;
or (n4279,s0n4279,s1n4279);
not(notn4279,n3122);
and (s0n4279,notn4279,n1124);
and (s1n4279,n3122,n1120);
and (n4280,n4281,n3141);
wire s0n4281,s1n4281,notn4281;
or (n4281,s0n4281,s1n4281);
not(notn4281,n3122);
and (s0n4281,notn4281,n1128);
and (s1n4281,n3122,n1124);
and (n4282,n4283,n3146);
wire s0n4283,s1n4283,notn4283;
or (n4283,s0n4283,s1n4283);
not(notn4283,n3122);
and (s0n4283,notn4283,n1132);
and (s1n4283,n3122,n1128);
and (n4284,n4285,n1042);
or (n4285,1'b0,n4286,n4288,n4290,n4292);
and (n4286,n4287,n3124);
wire s0n4287,s1n4287,notn4287;
or (n4287,s0n4287,s1n4287);
not(notn4287,n3122);
and (s0n4287,notn4287,n1138);
and (s1n4287,n3122,n1132);
and (n4288,n4289,n3136);
wire s0n4289,s1n4289,notn4289;
or (n4289,s0n4289,s1n4289);
not(notn4289,n3122);
and (s0n4289,notn4289,n1142);
and (s1n4289,n3122,n1138);
and (n4290,n4291,n3141);
wire s0n4291,s1n4291,notn4291;
or (n4291,s0n4291,s1n4291);
not(notn4291,n3122);
and (s0n4291,notn4291,n1146);
and (s1n4291,n3122,n1142);
and (n4292,n4293,n3146);
wire s0n4293,s1n4293,notn4293;
or (n4293,s0n4293,s1n4293);
not(notn4293,n3122);
and (s0n4293,notn4293,n1150);
and (s1n4293,n3122,n1146);
wire s0n4295,s1n4295,notn4295;
or (n4295,s0n4295,s1n4295);
not(notn4295,n3074);
and (s0n4295,notn4295,n4296);
and (s1n4295,n3074,n4337);
or (n4296,1'b0,n4297,n4307,n4317,n4327);
and (n4297,n4298,n981);
or (n4298,1'b0,n4299,n4301,n4303,n4305);
and (n4299,n4300,n3124);
wire s0n4300,s1n4300,notn4300;
or (n4300,s0n4300,s1n4300);
not(notn4300,n3122);
and (s0n4300,notn4300,n1085);
and (s1n4300,n3122,n1158);
and (n4301,n4302,n3136);
wire s0n4302,s1n4302,notn4302;
or (n4302,s0n4302,s1n4302);
not(notn4302,n3122);
and (s0n4302,notn4302,n1089);
and (s1n4302,n3122,n1085);
and (n4303,n4304,n3141);
wire s0n4304,s1n4304,notn4304;
or (n4304,s0n4304,s1n4304);
not(notn4304,n3122);
and (s0n4304,notn4304,n1093);
and (s1n4304,n3122,n1089);
and (n4305,n4306,n3146);
wire s0n4306,s1n4306,notn4306;
or (n4306,s0n4306,s1n4306);
not(notn4306,n3122);
and (s0n4306,notn4306,n1097);
and (s1n4306,n3122,n1093);
and (n4307,n4308,n1002);
or (n4308,1'b0,n4309,n4311,n4313,n4315);
and (n4309,n4310,n3124);
wire s0n4310,s1n4310,notn4310;
or (n4310,s0n4310,s1n4310);
not(notn4310,n3122);
and (s0n4310,notn4310,n1103);
and (s1n4310,n3122,n1097);
and (n4311,n4312,n3136);
wire s0n4312,s1n4312,notn4312;
or (n4312,s0n4312,s1n4312);
not(notn4312,n3122);
and (s0n4312,notn4312,n1107);
and (s1n4312,n3122,n1103);
and (n4313,n4314,n3141);
wire s0n4314,s1n4314,notn4314;
or (n4314,s0n4314,s1n4314);
not(notn4314,n3122);
and (s0n4314,notn4314,n1111);
and (s1n4314,n3122,n1107);
and (n4315,n4316,n3146);
wire s0n4316,s1n4316,notn4316;
or (n4316,s0n4316,s1n4316);
not(notn4316,n3122);
and (s0n4316,notn4316,n1115);
and (s1n4316,n3122,n1111);
and (n4317,n4318,n1022);
or (n4318,1'b0,n4319,n4321,n4323,n4325);
and (n4319,n4320,n3124);
wire s0n4320,s1n4320,notn4320;
or (n4320,s0n4320,s1n4320);
not(notn4320,n3122);
and (s0n4320,notn4320,n1121);
and (s1n4320,n3122,n1173);
and (n4321,n4322,n3136);
wire s0n4322,s1n4322,notn4322;
or (n4322,s0n4322,s1n4322);
not(notn4322,n3122);
and (s0n4322,notn4322,n1125);
and (s1n4322,n3122,n1121);
and (n4323,n4324,n3141);
wire s0n4324,s1n4324,notn4324;
or (n4324,s0n4324,s1n4324);
not(notn4324,n3122);
and (s0n4324,notn4324,n1129);
and (s1n4324,n3122,n1125);
and (n4325,n4326,n3146);
wire s0n4326,s1n4326,notn4326;
or (n4326,s0n4326,s1n4326);
not(notn4326,n3122);
and (s0n4326,notn4326,n1133);
and (s1n4326,n3122,n1129);
and (n4327,n4328,n1042);
or (n4328,1'b0,n4329,n4331,n4333,n4335);
and (n4329,n4330,n3124);
wire s0n4330,s1n4330,notn4330;
or (n4330,s0n4330,s1n4330);
not(notn4330,n3122);
and (s0n4330,notn4330,n1139);
and (s1n4330,n3122,n1133);
and (n4331,n4332,n3136);
wire s0n4332,s1n4332,notn4332;
or (n4332,s0n4332,s1n4332);
not(notn4332,n3122);
and (s0n4332,notn4332,n1143);
and (s1n4332,n3122,n1139);
and (n4333,n4334,n3141);
wire s0n4334,s1n4334,notn4334;
or (n4334,s0n4334,s1n4334);
not(notn4334,n3122);
and (s0n4334,notn4334,n1147);
and (s1n4334,n3122,n1143);
and (n4335,n4336,n3146);
wire s0n4336,s1n4336,notn4336;
or (n4336,s0n4336,s1n4336);
not(notn4336,n3122);
and (s0n4336,notn4336,n1151);
and (s1n4336,n3122,n1147);
and (n4338,n4295,n4339);
or (n4339,n4340,n4427,n4875);
and (n4340,n4341,n4384);
wire s0n4341,s1n4341,notn4341;
or (n4341,s0n4341,s1n4341);
not(notn4341,n3074);
and (s0n4341,notn4341,n4342);
and (s1n4341,n3074,n4383);
or (n4342,1'b0,n4343,n4353,n4363,n4373);
and (n4343,n4344,n981);
or (n4344,1'b0,n4345,n4347,n4349,n4351);
and (n4345,n4346,n3124);
wire s0n4346,s1n4346,notn4346;
or (n4346,s0n4346,s1n4346);
not(notn4346,n3122);
and (s0n4346,notn4346,n1191);
and (s1n4346,n3122,n1264);
and (n4347,n4348,n3136);
wire s0n4348,s1n4348,notn4348;
or (n4348,s0n4348,s1n4348);
not(notn4348,n3122);
and (s0n4348,notn4348,n1195);
and (s1n4348,n3122,n1191);
and (n4349,n4350,n3141);
wire s0n4350,s1n4350,notn4350;
or (n4350,s0n4350,s1n4350);
not(notn4350,n3122);
and (s0n4350,notn4350,n1199);
and (s1n4350,n3122,n1195);
and (n4351,n4352,n3146);
wire s0n4352,s1n4352,notn4352;
or (n4352,s0n4352,s1n4352);
not(notn4352,n3122);
and (s0n4352,notn4352,n1203);
and (s1n4352,n3122,n1199);
and (n4353,n4354,n1002);
or (n4354,1'b0,n4355,n4357,n4359,n4361);
and (n4355,n4356,n3124);
wire s0n4356,s1n4356,notn4356;
or (n4356,s0n4356,s1n4356);
not(notn4356,n3122);
and (s0n4356,notn4356,n1209);
and (s1n4356,n3122,n1203);
and (n4357,n4358,n3136);
wire s0n4358,s1n4358,notn4358;
or (n4358,s0n4358,s1n4358);
not(notn4358,n3122);
and (s0n4358,notn4358,n1213);
and (s1n4358,n3122,n1209);
and (n4359,n4360,n3141);
wire s0n4360,s1n4360,notn4360;
or (n4360,s0n4360,s1n4360);
not(notn4360,n3122);
and (s0n4360,notn4360,n1217);
and (s1n4360,n3122,n1213);
and (n4361,n4362,n3146);
wire s0n4362,s1n4362,notn4362;
or (n4362,s0n4362,s1n4362);
not(notn4362,n3122);
and (s0n4362,notn4362,n1221);
and (s1n4362,n3122,n1217);
and (n4363,n4364,n1022);
or (n4364,1'b0,n4365,n4367,n4369,n4371);
and (n4365,n4366,n3124);
wire s0n4366,s1n4366,notn4366;
or (n4366,s0n4366,s1n4366);
not(notn4366,n3122);
and (s0n4366,notn4366,n1227);
and (s1n4366,n3122,n1279);
and (n4367,n4368,n3136);
wire s0n4368,s1n4368,notn4368;
or (n4368,s0n4368,s1n4368);
not(notn4368,n3122);
and (s0n4368,notn4368,n1231);
and (s1n4368,n3122,n1227);
and (n4369,n4370,n3141);
wire s0n4370,s1n4370,notn4370;
or (n4370,s0n4370,s1n4370);
not(notn4370,n3122);
and (s0n4370,notn4370,n1235);
and (s1n4370,n3122,n1231);
and (n4371,n4372,n3146);
wire s0n4372,s1n4372,notn4372;
or (n4372,s0n4372,s1n4372);
not(notn4372,n3122);
and (s0n4372,notn4372,n1239);
and (s1n4372,n3122,n1235);
and (n4373,n4374,n1042);
or (n4374,1'b0,n4375,n4377,n4379,n4381);
and (n4375,n4376,n3124);
wire s0n4376,s1n4376,notn4376;
or (n4376,s0n4376,s1n4376);
not(notn4376,n3122);
and (s0n4376,notn4376,n1245);
and (s1n4376,n3122,n1239);
and (n4377,n4378,n3136);
wire s0n4378,s1n4378,notn4378;
or (n4378,s0n4378,s1n4378);
not(notn4378,n3122);
and (s0n4378,notn4378,n1249);
and (s1n4378,n3122,n1245);
and (n4379,n4380,n3141);
wire s0n4380,s1n4380,notn4380;
or (n4380,s0n4380,s1n4380);
not(notn4380,n3122);
and (s0n4380,notn4380,n1253);
and (s1n4380,n3122,n1249);
and (n4381,n4382,n3146);
wire s0n4382,s1n4382,notn4382;
or (n4382,s0n4382,s1n4382);
not(notn4382,n3122);
and (s0n4382,notn4382,n1257);
and (s1n4382,n3122,n1253);
wire s0n4384,s1n4384,notn4384;
or (n4384,s0n4384,s1n4384);
not(notn4384,n3074);
and (s0n4384,notn4384,n4385);
and (s1n4384,n3074,n4426);
or (n4385,1'b0,n4386,n4396,n4406,n4416);
and (n4386,n4387,n981);
or (n4387,1'b0,n4388,n4390,n4392,n4394);
and (n4388,n4389,n3124);
wire s0n4389,s1n4389,notn4389;
or (n4389,s0n4389,s1n4389);
not(notn4389,n3122);
and (s0n4389,notn4389,n1192);
and (s1n4389,n3122,n1265);
and (n4390,n4391,n3136);
wire s0n4391,s1n4391,notn4391;
or (n4391,s0n4391,s1n4391);
not(notn4391,n3122);
and (s0n4391,notn4391,n1196);
and (s1n4391,n3122,n1192);
and (n4392,n4393,n3141);
wire s0n4393,s1n4393,notn4393;
or (n4393,s0n4393,s1n4393);
not(notn4393,n3122);
and (s0n4393,notn4393,n1200);
and (s1n4393,n3122,n1196);
and (n4394,n4395,n3146);
wire s0n4395,s1n4395,notn4395;
or (n4395,s0n4395,s1n4395);
not(notn4395,n3122);
and (s0n4395,notn4395,n1204);
and (s1n4395,n3122,n1200);
and (n4396,n4397,n1002);
or (n4397,1'b0,n4398,n4400,n4402,n4404);
and (n4398,n4399,n3124);
wire s0n4399,s1n4399,notn4399;
or (n4399,s0n4399,s1n4399);
not(notn4399,n3122);
and (s0n4399,notn4399,n1210);
and (s1n4399,n3122,n1204);
and (n4400,n4401,n3136);
wire s0n4401,s1n4401,notn4401;
or (n4401,s0n4401,s1n4401);
not(notn4401,n3122);
and (s0n4401,notn4401,n1214);
and (s1n4401,n3122,n1210);
and (n4402,n4403,n3141);
wire s0n4403,s1n4403,notn4403;
or (n4403,s0n4403,s1n4403);
not(notn4403,n3122);
and (s0n4403,notn4403,n1218);
and (s1n4403,n3122,n1214);
and (n4404,n4405,n3146);
wire s0n4405,s1n4405,notn4405;
or (n4405,s0n4405,s1n4405);
not(notn4405,n3122);
and (s0n4405,notn4405,n1222);
and (s1n4405,n3122,n1218);
and (n4406,n4407,n1022);
or (n4407,1'b0,n4408,n4410,n4412,n4414);
and (n4408,n4409,n3124);
wire s0n4409,s1n4409,notn4409;
or (n4409,s0n4409,s1n4409);
not(notn4409,n3122);
and (s0n4409,notn4409,n1228);
and (s1n4409,n3122,n1280);
and (n4410,n4411,n3136);
wire s0n4411,s1n4411,notn4411;
or (n4411,s0n4411,s1n4411);
not(notn4411,n3122);
and (s0n4411,notn4411,n1232);
and (s1n4411,n3122,n1228);
and (n4412,n4413,n3141);
wire s0n4413,s1n4413,notn4413;
or (n4413,s0n4413,s1n4413);
not(notn4413,n3122);
and (s0n4413,notn4413,n1236);
and (s1n4413,n3122,n1232);
and (n4414,n4415,n3146);
wire s0n4415,s1n4415,notn4415;
or (n4415,s0n4415,s1n4415);
not(notn4415,n3122);
and (s0n4415,notn4415,n1240);
and (s1n4415,n3122,n1236);
and (n4416,n4417,n1042);
or (n4417,1'b0,n4418,n4420,n4422,n4424);
and (n4418,n4419,n3124);
wire s0n4419,s1n4419,notn4419;
or (n4419,s0n4419,s1n4419);
not(notn4419,n3122);
and (s0n4419,notn4419,n1246);
and (s1n4419,n3122,n1240);
and (n4420,n4421,n3136);
wire s0n4421,s1n4421,notn4421;
or (n4421,s0n4421,s1n4421);
not(notn4421,n3122);
and (s0n4421,notn4421,n1250);
and (s1n4421,n3122,n1246);
and (n4422,n4423,n3141);
wire s0n4423,s1n4423,notn4423;
or (n4423,s0n4423,s1n4423);
not(notn4423,n3122);
and (s0n4423,notn4423,n1254);
and (s1n4423,n3122,n1250);
and (n4424,n4425,n3146);
wire s0n4425,s1n4425,notn4425;
or (n4425,s0n4425,s1n4425);
not(notn4425,n3122);
and (s0n4425,notn4425,n1258);
and (s1n4425,n3122,n1254);
and (n4427,n4384,n4428);
or (n4428,n4429,n4516,n4874);
and (n4429,n4430,n4473);
wire s0n4430,s1n4430,notn4430;
or (n4430,s0n4430,s1n4430);
not(notn4430,n3074);
and (s0n4430,notn4430,n4431);
and (s1n4430,n3074,n4472);
or (n4431,1'b0,n4432,n4442,n4452,n4462);
and (n4432,n4433,n981);
or (n4433,1'b0,n4434,n4436,n4438,n4440);
and (n4434,n4435,n3124);
wire s0n4435,s1n4435,notn4435;
or (n4435,s0n4435,s1n4435);
not(notn4435,n3122);
and (s0n4435,notn4435,n1298);
and (s1n4435,n3122,n1371);
and (n4436,n4437,n3136);
wire s0n4437,s1n4437,notn4437;
or (n4437,s0n4437,s1n4437);
not(notn4437,n3122);
and (s0n4437,notn4437,n1302);
and (s1n4437,n3122,n1298);
and (n4438,n4439,n3141);
wire s0n4439,s1n4439,notn4439;
or (n4439,s0n4439,s1n4439);
not(notn4439,n3122);
and (s0n4439,notn4439,n1306);
and (s1n4439,n3122,n1302);
and (n4440,n4441,n3146);
wire s0n4441,s1n4441,notn4441;
or (n4441,s0n4441,s1n4441);
not(notn4441,n3122);
and (s0n4441,notn4441,n1310);
and (s1n4441,n3122,n1306);
and (n4442,n4443,n1002);
or (n4443,1'b0,n4444,n4446,n4448,n4450);
and (n4444,n4445,n3124);
wire s0n4445,s1n4445,notn4445;
or (n4445,s0n4445,s1n4445);
not(notn4445,n3122);
and (s0n4445,notn4445,n1316);
and (s1n4445,n3122,n1310);
and (n4446,n4447,n3136);
wire s0n4447,s1n4447,notn4447;
or (n4447,s0n4447,s1n4447);
not(notn4447,n3122);
and (s0n4447,notn4447,n1320);
and (s1n4447,n3122,n1316);
and (n4448,n4449,n3141);
wire s0n4449,s1n4449,notn4449;
or (n4449,s0n4449,s1n4449);
not(notn4449,n3122);
and (s0n4449,notn4449,n1324);
and (s1n4449,n3122,n1320);
and (n4450,n4451,n3146);
wire s0n4451,s1n4451,notn4451;
or (n4451,s0n4451,s1n4451);
not(notn4451,n3122);
and (s0n4451,notn4451,n1328);
and (s1n4451,n3122,n1324);
and (n4452,n4453,n1022);
or (n4453,1'b0,n4454,n4456,n4458,n4460);
and (n4454,n4455,n3124);
wire s0n4455,s1n4455,notn4455;
or (n4455,s0n4455,s1n4455);
not(notn4455,n3122);
and (s0n4455,notn4455,n1334);
and (s1n4455,n3122,n1386);
and (n4456,n4457,n3136);
wire s0n4457,s1n4457,notn4457;
or (n4457,s0n4457,s1n4457);
not(notn4457,n3122);
and (s0n4457,notn4457,n1338);
and (s1n4457,n3122,n1334);
and (n4458,n4459,n3141);
wire s0n4459,s1n4459,notn4459;
or (n4459,s0n4459,s1n4459);
not(notn4459,n3122);
and (s0n4459,notn4459,n1342);
and (s1n4459,n3122,n1338);
and (n4460,n4461,n3146);
wire s0n4461,s1n4461,notn4461;
or (n4461,s0n4461,s1n4461);
not(notn4461,n3122);
and (s0n4461,notn4461,n1346);
and (s1n4461,n3122,n1342);
and (n4462,n4463,n1042);
or (n4463,1'b0,n4464,n4466,n4468,n4470);
and (n4464,n4465,n3124);
wire s0n4465,s1n4465,notn4465;
or (n4465,s0n4465,s1n4465);
not(notn4465,n3122);
and (s0n4465,notn4465,n1352);
and (s1n4465,n3122,n1346);
and (n4466,n4467,n3136);
wire s0n4467,s1n4467,notn4467;
or (n4467,s0n4467,s1n4467);
not(notn4467,n3122);
and (s0n4467,notn4467,n1356);
and (s1n4467,n3122,n1352);
and (n4468,n4469,n3141);
wire s0n4469,s1n4469,notn4469;
or (n4469,s0n4469,s1n4469);
not(notn4469,n3122);
and (s0n4469,notn4469,n1360);
and (s1n4469,n3122,n1356);
and (n4470,n4471,n3146);
wire s0n4471,s1n4471,notn4471;
or (n4471,s0n4471,s1n4471);
not(notn4471,n3122);
and (s0n4471,notn4471,n1364);
and (s1n4471,n3122,n1360);
wire s0n4473,s1n4473,notn4473;
or (n4473,s0n4473,s1n4473);
not(notn4473,n3074);
and (s0n4473,notn4473,n4474);
and (s1n4473,n3074,n4515);
or (n4474,1'b0,n4475,n4485,n4495,n4505);
and (n4475,n4476,n981);
or (n4476,1'b0,n4477,n4479,n4481,n4483);
and (n4477,n4478,n3124);
wire s0n4478,s1n4478,notn4478;
or (n4478,s0n4478,s1n4478);
not(notn4478,n3122);
and (s0n4478,notn4478,n1299);
and (s1n4478,n3122,n1372);
and (n4479,n4480,n3136);
wire s0n4480,s1n4480,notn4480;
or (n4480,s0n4480,s1n4480);
not(notn4480,n3122);
and (s0n4480,notn4480,n1303);
and (s1n4480,n3122,n1299);
and (n4481,n4482,n3141);
wire s0n4482,s1n4482,notn4482;
or (n4482,s0n4482,s1n4482);
not(notn4482,n3122);
and (s0n4482,notn4482,n1307);
and (s1n4482,n3122,n1303);
and (n4483,n4484,n3146);
wire s0n4484,s1n4484,notn4484;
or (n4484,s0n4484,s1n4484);
not(notn4484,n3122);
and (s0n4484,notn4484,n1311);
and (s1n4484,n3122,n1307);
and (n4485,n4486,n1002);
or (n4486,1'b0,n4487,n4489,n4491,n4493);
and (n4487,n4488,n3124);
wire s0n4488,s1n4488,notn4488;
or (n4488,s0n4488,s1n4488);
not(notn4488,n3122);
and (s0n4488,notn4488,n1317);
and (s1n4488,n3122,n1311);
and (n4489,n4490,n3136);
wire s0n4490,s1n4490,notn4490;
or (n4490,s0n4490,s1n4490);
not(notn4490,n3122);
and (s0n4490,notn4490,n1321);
and (s1n4490,n3122,n1317);
and (n4491,n4492,n3141);
wire s0n4492,s1n4492,notn4492;
or (n4492,s0n4492,s1n4492);
not(notn4492,n3122);
and (s0n4492,notn4492,n1325);
and (s1n4492,n3122,n1321);
and (n4493,n4494,n3146);
wire s0n4494,s1n4494,notn4494;
or (n4494,s0n4494,s1n4494);
not(notn4494,n3122);
and (s0n4494,notn4494,n1329);
and (s1n4494,n3122,n1325);
and (n4495,n4496,n1022);
or (n4496,1'b0,n4497,n4499,n4501,n4503);
and (n4497,n4498,n3124);
wire s0n4498,s1n4498,notn4498;
or (n4498,s0n4498,s1n4498);
not(notn4498,n3122);
and (s0n4498,notn4498,n1335);
and (s1n4498,n3122,n1387);
and (n4499,n4500,n3136);
wire s0n4500,s1n4500,notn4500;
or (n4500,s0n4500,s1n4500);
not(notn4500,n3122);
and (s0n4500,notn4500,n1339);
and (s1n4500,n3122,n1335);
and (n4501,n4502,n3141);
wire s0n4502,s1n4502,notn4502;
or (n4502,s0n4502,s1n4502);
not(notn4502,n3122);
and (s0n4502,notn4502,n1343);
and (s1n4502,n3122,n1339);
and (n4503,n4504,n3146);
wire s0n4504,s1n4504,notn4504;
or (n4504,s0n4504,s1n4504);
not(notn4504,n3122);
and (s0n4504,notn4504,n1347);
and (s1n4504,n3122,n1343);
and (n4505,n4506,n1042);
or (n4506,1'b0,n4507,n4509,n4511,n4513);
and (n4507,n4508,n3124);
wire s0n4508,s1n4508,notn4508;
or (n4508,s0n4508,s1n4508);
not(notn4508,n3122);
and (s0n4508,notn4508,n1353);
and (s1n4508,n3122,n1347);
and (n4509,n4510,n3136);
wire s0n4510,s1n4510,notn4510;
or (n4510,s0n4510,s1n4510);
not(notn4510,n3122);
and (s0n4510,notn4510,n1357);
and (s1n4510,n3122,n1353);
and (n4511,n4512,n3141);
wire s0n4512,s1n4512,notn4512;
or (n4512,s0n4512,s1n4512);
not(notn4512,n3122);
and (s0n4512,notn4512,n1361);
and (s1n4512,n3122,n1357);
and (n4513,n4514,n3146);
wire s0n4514,s1n4514,notn4514;
or (n4514,s0n4514,s1n4514);
not(notn4514,n3122);
and (s0n4514,notn4514,n1365);
and (s1n4514,n3122,n1361);
and (n4516,n4473,n4517);
or (n4517,n4518,n4605,n4873);
and (n4518,n4519,n4562);
wire s0n4519,s1n4519,notn4519;
or (n4519,s0n4519,s1n4519);
not(notn4519,n3074);
and (s0n4519,notn4519,n4520);
and (s1n4519,n3074,n4561);
or (n4520,1'b0,n4521,n4531,n4541,n4551);
and (n4521,n4522,n981);
or (n4522,1'b0,n4523,n4525,n4527,n4529);
and (n4523,n4524,n3124);
wire s0n4524,s1n4524,notn4524;
or (n4524,s0n4524,s1n4524);
not(notn4524,n3122);
and (s0n4524,notn4524,n1405);
and (s1n4524,n3122,n1478);
and (n4525,n4526,n3136);
wire s0n4526,s1n4526,notn4526;
or (n4526,s0n4526,s1n4526);
not(notn4526,n3122);
and (s0n4526,notn4526,n1409);
and (s1n4526,n3122,n1405);
and (n4527,n4528,n3141);
wire s0n4528,s1n4528,notn4528;
or (n4528,s0n4528,s1n4528);
not(notn4528,n3122);
and (s0n4528,notn4528,n1413);
and (s1n4528,n3122,n1409);
and (n4529,n4530,n3146);
wire s0n4530,s1n4530,notn4530;
or (n4530,s0n4530,s1n4530);
not(notn4530,n3122);
and (s0n4530,notn4530,n1417);
and (s1n4530,n3122,n1413);
and (n4531,n4532,n1002);
or (n4532,1'b0,n4533,n4535,n4537,n4539);
and (n4533,n4534,n3124);
wire s0n4534,s1n4534,notn4534;
or (n4534,s0n4534,s1n4534);
not(notn4534,n3122);
and (s0n4534,notn4534,n1423);
and (s1n4534,n3122,n1417);
and (n4535,n4536,n3136);
wire s0n4536,s1n4536,notn4536;
or (n4536,s0n4536,s1n4536);
not(notn4536,n3122);
and (s0n4536,notn4536,n1427);
and (s1n4536,n3122,n1423);
and (n4537,n4538,n3141);
wire s0n4538,s1n4538,notn4538;
or (n4538,s0n4538,s1n4538);
not(notn4538,n3122);
and (s0n4538,notn4538,n1431);
and (s1n4538,n3122,n1427);
and (n4539,n4540,n3146);
wire s0n4540,s1n4540,notn4540;
or (n4540,s0n4540,s1n4540);
not(notn4540,n3122);
and (s0n4540,notn4540,n1435);
and (s1n4540,n3122,n1431);
and (n4541,n4542,n1022);
or (n4542,1'b0,n4543,n4545,n4547,n4549);
and (n4543,n4544,n3124);
wire s0n4544,s1n4544,notn4544;
or (n4544,s0n4544,s1n4544);
not(notn4544,n3122);
and (s0n4544,notn4544,n1441);
and (s1n4544,n3122,n1493);
and (n4545,n4546,n3136);
wire s0n4546,s1n4546,notn4546;
or (n4546,s0n4546,s1n4546);
not(notn4546,n3122);
and (s0n4546,notn4546,n1445);
and (s1n4546,n3122,n1441);
and (n4547,n4548,n3141);
wire s0n4548,s1n4548,notn4548;
or (n4548,s0n4548,s1n4548);
not(notn4548,n3122);
and (s0n4548,notn4548,n1449);
and (s1n4548,n3122,n1445);
and (n4549,n4550,n3146);
wire s0n4550,s1n4550,notn4550;
or (n4550,s0n4550,s1n4550);
not(notn4550,n3122);
and (s0n4550,notn4550,n1453);
and (s1n4550,n3122,n1449);
and (n4551,n4552,n1042);
or (n4552,1'b0,n4553,n4555,n4557,n4559);
and (n4553,n4554,n3124);
wire s0n4554,s1n4554,notn4554;
or (n4554,s0n4554,s1n4554);
not(notn4554,n3122);
and (s0n4554,notn4554,n1459);
and (s1n4554,n3122,n1453);
and (n4555,n4556,n3136);
wire s0n4556,s1n4556,notn4556;
or (n4556,s0n4556,s1n4556);
not(notn4556,n3122);
and (s0n4556,notn4556,n1463);
and (s1n4556,n3122,n1459);
and (n4557,n4558,n3141);
wire s0n4558,s1n4558,notn4558;
or (n4558,s0n4558,s1n4558);
not(notn4558,n3122);
and (s0n4558,notn4558,n1467);
and (s1n4558,n3122,n1463);
and (n4559,n4560,n3146);
wire s0n4560,s1n4560,notn4560;
or (n4560,s0n4560,s1n4560);
not(notn4560,n3122);
and (s0n4560,notn4560,n1471);
and (s1n4560,n3122,n1467);
wire s0n4562,s1n4562,notn4562;
or (n4562,s0n4562,s1n4562);
not(notn4562,n3074);
and (s0n4562,notn4562,n4563);
and (s1n4562,n3074,n4604);
or (n4563,1'b0,n4564,n4574,n4584,n4594);
and (n4564,n4565,n981);
or (n4565,1'b0,n4566,n4568,n4570,n4572);
and (n4566,n4567,n3124);
wire s0n4567,s1n4567,notn4567;
or (n4567,s0n4567,s1n4567);
not(notn4567,n3122);
and (s0n4567,notn4567,n1406);
and (s1n4567,n3122,n1479);
and (n4568,n4569,n3136);
wire s0n4569,s1n4569,notn4569;
or (n4569,s0n4569,s1n4569);
not(notn4569,n3122);
and (s0n4569,notn4569,n1410);
and (s1n4569,n3122,n1406);
and (n4570,n4571,n3141);
wire s0n4571,s1n4571,notn4571;
or (n4571,s0n4571,s1n4571);
not(notn4571,n3122);
and (s0n4571,notn4571,n1414);
and (s1n4571,n3122,n1410);
and (n4572,n4573,n3146);
wire s0n4573,s1n4573,notn4573;
or (n4573,s0n4573,s1n4573);
not(notn4573,n3122);
and (s0n4573,notn4573,n1418);
and (s1n4573,n3122,n1414);
and (n4574,n4575,n1002);
or (n4575,1'b0,n4576,n4578,n4580,n4582);
and (n4576,n4577,n3124);
wire s0n4577,s1n4577,notn4577;
or (n4577,s0n4577,s1n4577);
not(notn4577,n3122);
and (s0n4577,notn4577,n1424);
and (s1n4577,n3122,n1418);
and (n4578,n4579,n3136);
wire s0n4579,s1n4579,notn4579;
or (n4579,s0n4579,s1n4579);
not(notn4579,n3122);
and (s0n4579,notn4579,n1428);
and (s1n4579,n3122,n1424);
and (n4580,n4581,n3141);
wire s0n4581,s1n4581,notn4581;
or (n4581,s0n4581,s1n4581);
not(notn4581,n3122);
and (s0n4581,notn4581,n1432);
and (s1n4581,n3122,n1428);
and (n4582,n4583,n3146);
wire s0n4583,s1n4583,notn4583;
or (n4583,s0n4583,s1n4583);
not(notn4583,n3122);
and (s0n4583,notn4583,n1436);
and (s1n4583,n3122,n1432);
and (n4584,n4585,n1022);
or (n4585,1'b0,n4586,n4588,n4590,n4592);
and (n4586,n4587,n3124);
wire s0n4587,s1n4587,notn4587;
or (n4587,s0n4587,s1n4587);
not(notn4587,n3122);
and (s0n4587,notn4587,n1442);
and (s1n4587,n3122,n1494);
and (n4588,n4589,n3136);
wire s0n4589,s1n4589,notn4589;
or (n4589,s0n4589,s1n4589);
not(notn4589,n3122);
and (s0n4589,notn4589,n1446);
and (s1n4589,n3122,n1442);
and (n4590,n4591,n3141);
wire s0n4591,s1n4591,notn4591;
or (n4591,s0n4591,s1n4591);
not(notn4591,n3122);
and (s0n4591,notn4591,n1450);
and (s1n4591,n3122,n1446);
and (n4592,n4593,n3146);
wire s0n4593,s1n4593,notn4593;
or (n4593,s0n4593,s1n4593);
not(notn4593,n3122);
and (s0n4593,notn4593,n1454);
and (s1n4593,n3122,n1450);
and (n4594,n4595,n1042);
or (n4595,1'b0,n4596,n4598,n4600,n4602);
and (n4596,n4597,n3124);
wire s0n4597,s1n4597,notn4597;
or (n4597,s0n4597,s1n4597);
not(notn4597,n3122);
and (s0n4597,notn4597,n1460);
and (s1n4597,n3122,n1454);
and (n4598,n4599,n3136);
wire s0n4599,s1n4599,notn4599;
or (n4599,s0n4599,s1n4599);
not(notn4599,n3122);
and (s0n4599,notn4599,n1464);
and (s1n4599,n3122,n1460);
and (n4600,n4601,n3141);
wire s0n4601,s1n4601,notn4601;
or (n4601,s0n4601,s1n4601);
not(notn4601,n3122);
and (s0n4601,notn4601,n1468);
and (s1n4601,n3122,n1464);
and (n4602,n4603,n3146);
wire s0n4603,s1n4603,notn4603;
or (n4603,s0n4603,s1n4603);
not(notn4603,n3122);
and (s0n4603,notn4603,n1472);
and (s1n4603,n3122,n1468);
and (n4605,n4562,n4606);
or (n4606,n4607,n4694,n4872);
and (n4607,n4608,n4651);
wire s0n4608,s1n4608,notn4608;
or (n4608,s0n4608,s1n4608);
not(notn4608,n3074);
and (s0n4608,notn4608,n4609);
and (s1n4608,n3074,n4650);
or (n4609,1'b0,n4610,n4620,n4630,n4640);
and (n4610,n4611,n981);
or (n4611,1'b0,n4612,n4614,n4616,n4618);
and (n4612,n4613,n3124);
wire s0n4613,s1n4613,notn4613;
or (n4613,s0n4613,s1n4613);
not(notn4613,n3122);
and (s0n4613,notn4613,n1512);
and (s1n4613,n3122,n1585);
and (n4614,n4615,n3136);
wire s0n4615,s1n4615,notn4615;
or (n4615,s0n4615,s1n4615);
not(notn4615,n3122);
and (s0n4615,notn4615,n1516);
and (s1n4615,n3122,n1512);
and (n4616,n4617,n3141);
wire s0n4617,s1n4617,notn4617;
or (n4617,s0n4617,s1n4617);
not(notn4617,n3122);
and (s0n4617,notn4617,n1520);
and (s1n4617,n3122,n1516);
and (n4618,n4619,n3146);
wire s0n4619,s1n4619,notn4619;
or (n4619,s0n4619,s1n4619);
not(notn4619,n3122);
and (s0n4619,notn4619,n1524);
and (s1n4619,n3122,n1520);
and (n4620,n4621,n1002);
or (n4621,1'b0,n4622,n4624,n4626,n4628);
and (n4622,n4623,n3124);
wire s0n4623,s1n4623,notn4623;
or (n4623,s0n4623,s1n4623);
not(notn4623,n3122);
and (s0n4623,notn4623,n1530);
and (s1n4623,n3122,n1524);
and (n4624,n4625,n3136);
wire s0n4625,s1n4625,notn4625;
or (n4625,s0n4625,s1n4625);
not(notn4625,n3122);
and (s0n4625,notn4625,n1534);
and (s1n4625,n3122,n1530);
and (n4626,n4627,n3141);
wire s0n4627,s1n4627,notn4627;
or (n4627,s0n4627,s1n4627);
not(notn4627,n3122);
and (s0n4627,notn4627,n1538);
and (s1n4627,n3122,n1534);
and (n4628,n4629,n3146);
wire s0n4629,s1n4629,notn4629;
or (n4629,s0n4629,s1n4629);
not(notn4629,n3122);
and (s0n4629,notn4629,n1542);
and (s1n4629,n3122,n1538);
and (n4630,n4631,n1022);
or (n4631,1'b0,n4632,n4634,n4636,n4638);
and (n4632,n4633,n3124);
wire s0n4633,s1n4633,notn4633;
or (n4633,s0n4633,s1n4633);
not(notn4633,n3122);
and (s0n4633,notn4633,n1548);
and (s1n4633,n3122,n1600);
and (n4634,n4635,n3136);
wire s0n4635,s1n4635,notn4635;
or (n4635,s0n4635,s1n4635);
not(notn4635,n3122);
and (s0n4635,notn4635,n1552);
and (s1n4635,n3122,n1548);
and (n4636,n4637,n3141);
wire s0n4637,s1n4637,notn4637;
or (n4637,s0n4637,s1n4637);
not(notn4637,n3122);
and (s0n4637,notn4637,n1556);
and (s1n4637,n3122,n1552);
and (n4638,n4639,n3146);
wire s0n4639,s1n4639,notn4639;
or (n4639,s0n4639,s1n4639);
not(notn4639,n3122);
and (s0n4639,notn4639,n1560);
and (s1n4639,n3122,n1556);
and (n4640,n4641,n1042);
or (n4641,1'b0,n4642,n4644,n4646,n4648);
and (n4642,n4643,n3124);
wire s0n4643,s1n4643,notn4643;
or (n4643,s0n4643,s1n4643);
not(notn4643,n3122);
and (s0n4643,notn4643,n1566);
and (s1n4643,n3122,n1560);
and (n4644,n4645,n3136);
wire s0n4645,s1n4645,notn4645;
or (n4645,s0n4645,s1n4645);
not(notn4645,n3122);
and (s0n4645,notn4645,n1570);
and (s1n4645,n3122,n1566);
and (n4646,n4647,n3141);
wire s0n4647,s1n4647,notn4647;
or (n4647,s0n4647,s1n4647);
not(notn4647,n3122);
and (s0n4647,notn4647,n1574);
and (s1n4647,n3122,n1570);
and (n4648,n4649,n3146);
wire s0n4649,s1n4649,notn4649;
or (n4649,s0n4649,s1n4649);
not(notn4649,n3122);
and (s0n4649,notn4649,n1578);
and (s1n4649,n3122,n1574);
wire s0n4651,s1n4651,notn4651;
or (n4651,s0n4651,s1n4651);
not(notn4651,n3074);
and (s0n4651,notn4651,n4652);
and (s1n4651,n3074,n4693);
or (n4652,1'b0,n4653,n4663,n4673,n4683);
and (n4653,n4654,n981);
or (n4654,1'b0,n4655,n4657,n4659,n4661);
and (n4655,n4656,n3124);
wire s0n4656,s1n4656,notn4656;
or (n4656,s0n4656,s1n4656);
not(notn4656,n3122);
and (s0n4656,notn4656,n1513);
and (s1n4656,n3122,n1586);
and (n4657,n4658,n3136);
wire s0n4658,s1n4658,notn4658;
or (n4658,s0n4658,s1n4658);
not(notn4658,n3122);
and (s0n4658,notn4658,n1517);
and (s1n4658,n3122,n1513);
and (n4659,n4660,n3141);
wire s0n4660,s1n4660,notn4660;
or (n4660,s0n4660,s1n4660);
not(notn4660,n3122);
and (s0n4660,notn4660,n1521);
and (s1n4660,n3122,n1517);
and (n4661,n4662,n3146);
wire s0n4662,s1n4662,notn4662;
or (n4662,s0n4662,s1n4662);
not(notn4662,n3122);
and (s0n4662,notn4662,n1525);
and (s1n4662,n3122,n1521);
and (n4663,n4664,n1002);
or (n4664,1'b0,n4665,n4667,n4669,n4671);
and (n4665,n4666,n3124);
wire s0n4666,s1n4666,notn4666;
or (n4666,s0n4666,s1n4666);
not(notn4666,n3122);
and (s0n4666,notn4666,n1531);
and (s1n4666,n3122,n1525);
and (n4667,n4668,n3136);
wire s0n4668,s1n4668,notn4668;
or (n4668,s0n4668,s1n4668);
not(notn4668,n3122);
and (s0n4668,notn4668,n1535);
and (s1n4668,n3122,n1531);
and (n4669,n4670,n3141);
wire s0n4670,s1n4670,notn4670;
or (n4670,s0n4670,s1n4670);
not(notn4670,n3122);
and (s0n4670,notn4670,n1539);
and (s1n4670,n3122,n1535);
and (n4671,n4672,n3146);
wire s0n4672,s1n4672,notn4672;
or (n4672,s0n4672,s1n4672);
not(notn4672,n3122);
and (s0n4672,notn4672,n1543);
and (s1n4672,n3122,n1539);
and (n4673,n4674,n1022);
or (n4674,1'b0,n4675,n4677,n4679,n4681);
and (n4675,n4676,n3124);
wire s0n4676,s1n4676,notn4676;
or (n4676,s0n4676,s1n4676);
not(notn4676,n3122);
and (s0n4676,notn4676,n1549);
and (s1n4676,n3122,n1601);
and (n4677,n4678,n3136);
wire s0n4678,s1n4678,notn4678;
or (n4678,s0n4678,s1n4678);
not(notn4678,n3122);
and (s0n4678,notn4678,n1553);
and (s1n4678,n3122,n1549);
and (n4679,n4680,n3141);
wire s0n4680,s1n4680,notn4680;
or (n4680,s0n4680,s1n4680);
not(notn4680,n3122);
and (s0n4680,notn4680,n1557);
and (s1n4680,n3122,n1553);
and (n4681,n4682,n3146);
wire s0n4682,s1n4682,notn4682;
or (n4682,s0n4682,s1n4682);
not(notn4682,n3122);
and (s0n4682,notn4682,n1561);
and (s1n4682,n3122,n1557);
and (n4683,n4684,n1042);
or (n4684,1'b0,n4685,n4687,n4689,n4691);
and (n4685,n4686,n3124);
wire s0n4686,s1n4686,notn4686;
or (n4686,s0n4686,s1n4686);
not(notn4686,n3122);
and (s0n4686,notn4686,n1567);
and (s1n4686,n3122,n1561);
and (n4687,n4688,n3136);
wire s0n4688,s1n4688,notn4688;
or (n4688,s0n4688,s1n4688);
not(notn4688,n3122);
and (s0n4688,notn4688,n1571);
and (s1n4688,n3122,n1567);
and (n4689,n4690,n3141);
wire s0n4690,s1n4690,notn4690;
or (n4690,s0n4690,s1n4690);
not(notn4690,n3122);
and (s0n4690,notn4690,n1575);
and (s1n4690,n3122,n1571);
and (n4691,n4692,n3146);
wire s0n4692,s1n4692,notn4692;
or (n4692,s0n4692,s1n4692);
not(notn4692,n3122);
and (s0n4692,notn4692,n1579);
and (s1n4692,n3122,n1575);
and (n4694,n4651,n4695);
or (n4695,n4696,n4783,n4871);
and (n4696,n4697,n4740);
wire s0n4697,s1n4697,notn4697;
or (n4697,s0n4697,s1n4697);
not(notn4697,n3074);
and (s0n4697,notn4697,n4698);
and (s1n4697,n3074,n4739);
or (n4698,1'b0,n4699,n4709,n4719,n4729);
and (n4699,n4700,n981);
or (n4700,1'b0,n4701,n4703,n4705,n4707);
and (n4701,n4702,n3124);
wire s0n4702,s1n4702,notn4702;
or (n4702,s0n4702,s1n4702);
not(notn4702,n3122);
and (s0n4702,notn4702,n1619);
and (s1n4702,n3122,n1692);
and (n4703,n4704,n3136);
wire s0n4704,s1n4704,notn4704;
or (n4704,s0n4704,s1n4704);
not(notn4704,n3122);
and (s0n4704,notn4704,n1623);
and (s1n4704,n3122,n1619);
and (n4705,n4706,n3141);
wire s0n4706,s1n4706,notn4706;
or (n4706,s0n4706,s1n4706);
not(notn4706,n3122);
and (s0n4706,notn4706,n1627);
and (s1n4706,n3122,n1623);
and (n4707,n4708,n3146);
wire s0n4708,s1n4708,notn4708;
or (n4708,s0n4708,s1n4708);
not(notn4708,n3122);
and (s0n4708,notn4708,n1631);
and (s1n4708,n3122,n1627);
and (n4709,n4710,n1002);
or (n4710,1'b0,n4711,n4713,n4715,n4717);
and (n4711,n4712,n3124);
wire s0n4712,s1n4712,notn4712;
or (n4712,s0n4712,s1n4712);
not(notn4712,n3122);
and (s0n4712,notn4712,n1637);
and (s1n4712,n3122,n1631);
and (n4713,n4714,n3136);
wire s0n4714,s1n4714,notn4714;
or (n4714,s0n4714,s1n4714);
not(notn4714,n3122);
and (s0n4714,notn4714,n1641);
and (s1n4714,n3122,n1637);
and (n4715,n4716,n3141);
wire s0n4716,s1n4716,notn4716;
or (n4716,s0n4716,s1n4716);
not(notn4716,n3122);
and (s0n4716,notn4716,n1645);
and (s1n4716,n3122,n1641);
and (n4717,n4718,n3146);
wire s0n4718,s1n4718,notn4718;
or (n4718,s0n4718,s1n4718);
not(notn4718,n3122);
and (s0n4718,notn4718,n1649);
and (s1n4718,n3122,n1645);
and (n4719,n4720,n1022);
or (n4720,1'b0,n4721,n4723,n4725,n4727);
and (n4721,n4722,n3124);
wire s0n4722,s1n4722,notn4722;
or (n4722,s0n4722,s1n4722);
not(notn4722,n3122);
and (s0n4722,notn4722,n1655);
and (s1n4722,n3122,n1707);
and (n4723,n4724,n3136);
wire s0n4724,s1n4724,notn4724;
or (n4724,s0n4724,s1n4724);
not(notn4724,n3122);
and (s0n4724,notn4724,n1659);
and (s1n4724,n3122,n1655);
and (n4725,n4726,n3141);
wire s0n4726,s1n4726,notn4726;
or (n4726,s0n4726,s1n4726);
not(notn4726,n3122);
and (s0n4726,notn4726,n1663);
and (s1n4726,n3122,n1659);
and (n4727,n4728,n3146);
wire s0n4728,s1n4728,notn4728;
or (n4728,s0n4728,s1n4728);
not(notn4728,n3122);
and (s0n4728,notn4728,n1667);
and (s1n4728,n3122,n1663);
and (n4729,n4730,n1042);
or (n4730,1'b0,n4731,n4733,n4735,n4737);
and (n4731,n4732,n3124);
wire s0n4732,s1n4732,notn4732;
or (n4732,s0n4732,s1n4732);
not(notn4732,n3122);
and (s0n4732,notn4732,n1673);
and (s1n4732,n3122,n1667);
and (n4733,n4734,n3136);
wire s0n4734,s1n4734,notn4734;
or (n4734,s0n4734,s1n4734);
not(notn4734,n3122);
and (s0n4734,notn4734,n1677);
and (s1n4734,n3122,n1673);
and (n4735,n4736,n3141);
wire s0n4736,s1n4736,notn4736;
or (n4736,s0n4736,s1n4736);
not(notn4736,n3122);
and (s0n4736,notn4736,n1681);
and (s1n4736,n3122,n1677);
and (n4737,n4738,n3146);
wire s0n4738,s1n4738,notn4738;
or (n4738,s0n4738,s1n4738);
not(notn4738,n3122);
and (s0n4738,notn4738,n1685);
and (s1n4738,n3122,n1681);
wire s0n4740,s1n4740,notn4740;
or (n4740,s0n4740,s1n4740);
not(notn4740,n3074);
and (s0n4740,notn4740,n4741);
and (s1n4740,n3074,n4782);
or (n4741,1'b0,n4742,n4752,n4762,n4772);
and (n4742,n4743,n981);
or (n4743,1'b0,n4744,n4746,n4748,n4750);
and (n4744,n4745,n3124);
wire s0n4745,s1n4745,notn4745;
or (n4745,s0n4745,s1n4745);
not(notn4745,n3122);
and (s0n4745,notn4745,n1620);
and (s1n4745,n3122,n1693);
and (n4746,n4747,n3136);
wire s0n4747,s1n4747,notn4747;
or (n4747,s0n4747,s1n4747);
not(notn4747,n3122);
and (s0n4747,notn4747,n1624);
and (s1n4747,n3122,n1620);
and (n4748,n4749,n3141);
wire s0n4749,s1n4749,notn4749;
or (n4749,s0n4749,s1n4749);
not(notn4749,n3122);
and (s0n4749,notn4749,n1628);
and (s1n4749,n3122,n1624);
and (n4750,n4751,n3146);
wire s0n4751,s1n4751,notn4751;
or (n4751,s0n4751,s1n4751);
not(notn4751,n3122);
and (s0n4751,notn4751,n1632);
and (s1n4751,n3122,n1628);
and (n4752,n4753,n1002);
or (n4753,1'b0,n4754,n4756,n4758,n4760);
and (n4754,n4755,n3124);
wire s0n4755,s1n4755,notn4755;
or (n4755,s0n4755,s1n4755);
not(notn4755,n3122);
and (s0n4755,notn4755,n1638);
and (s1n4755,n3122,n1632);
and (n4756,n4757,n3136);
wire s0n4757,s1n4757,notn4757;
or (n4757,s0n4757,s1n4757);
not(notn4757,n3122);
and (s0n4757,notn4757,n1642);
and (s1n4757,n3122,n1638);
and (n4758,n4759,n3141);
wire s0n4759,s1n4759,notn4759;
or (n4759,s0n4759,s1n4759);
not(notn4759,n3122);
and (s0n4759,notn4759,n1646);
and (s1n4759,n3122,n1642);
and (n4760,n4761,n3146);
wire s0n4761,s1n4761,notn4761;
or (n4761,s0n4761,s1n4761);
not(notn4761,n3122);
and (s0n4761,notn4761,n1650);
and (s1n4761,n3122,n1646);
and (n4762,n4763,n1022);
or (n4763,1'b0,n4764,n4766,n4768,n4770);
and (n4764,n4765,n3124);
wire s0n4765,s1n4765,notn4765;
or (n4765,s0n4765,s1n4765);
not(notn4765,n3122);
and (s0n4765,notn4765,n1656);
and (s1n4765,n3122,n1708);
and (n4766,n4767,n3136);
wire s0n4767,s1n4767,notn4767;
or (n4767,s0n4767,s1n4767);
not(notn4767,n3122);
and (s0n4767,notn4767,n1660);
and (s1n4767,n3122,n1656);
and (n4768,n4769,n3141);
wire s0n4769,s1n4769,notn4769;
or (n4769,s0n4769,s1n4769);
not(notn4769,n3122);
and (s0n4769,notn4769,n1664);
and (s1n4769,n3122,n1660);
and (n4770,n4771,n3146);
wire s0n4771,s1n4771,notn4771;
or (n4771,s0n4771,s1n4771);
not(notn4771,n3122);
and (s0n4771,notn4771,n1668);
and (s1n4771,n3122,n1664);
and (n4772,n4773,n1042);
or (n4773,1'b0,n4774,n4776,n4778,n4780);
and (n4774,n4775,n3124);
wire s0n4775,s1n4775,notn4775;
or (n4775,s0n4775,s1n4775);
not(notn4775,n3122);
and (s0n4775,notn4775,n1674);
and (s1n4775,n3122,n1668);
and (n4776,n4777,n3136);
wire s0n4777,s1n4777,notn4777;
or (n4777,s0n4777,s1n4777);
not(notn4777,n3122);
and (s0n4777,notn4777,n1678);
and (s1n4777,n3122,n1674);
and (n4778,n4779,n3141);
wire s0n4779,s1n4779,notn4779;
or (n4779,s0n4779,s1n4779);
not(notn4779,n3122);
and (s0n4779,notn4779,n1682);
and (s1n4779,n3122,n1678);
and (n4780,n4781,n3146);
wire s0n4781,s1n4781,notn4781;
or (n4781,s0n4781,s1n4781);
not(notn4781,n3122);
and (s0n4781,notn4781,n1686);
and (s1n4781,n3122,n1682);
and (n4783,n4740,n4784);
and (n4784,n4785,n4828);
wire s0n4785,s1n4785,notn4785;
or (n4785,s0n4785,s1n4785);
not(notn4785,n3074);
and (s0n4785,notn4785,n4786);
and (s1n4785,n3074,n4827);
or (n4786,1'b0,n4787,n4797,n4807,n4817);
and (n4787,n4788,n981);
or (n4788,1'b0,n4789,n4791,n4793,n4795);
and (n4789,n4790,n3124);
wire s0n4790,s1n4790,notn4790;
or (n4790,s0n4790,s1n4790);
not(notn4790,n3122);
and (s0n4790,notn4790,n1725);
and (s1n4790,n3122,n1798);
and (n4791,n4792,n3136);
wire s0n4792,s1n4792,notn4792;
or (n4792,s0n4792,s1n4792);
not(notn4792,n3122);
and (s0n4792,notn4792,n1729);
and (s1n4792,n3122,n1725);
and (n4793,n4794,n3141);
wire s0n4794,s1n4794,notn4794;
or (n4794,s0n4794,s1n4794);
not(notn4794,n3122);
and (s0n4794,notn4794,n1733);
and (s1n4794,n3122,n1729);
and (n4795,n4796,n3146);
wire s0n4796,s1n4796,notn4796;
or (n4796,s0n4796,s1n4796);
not(notn4796,n3122);
and (s0n4796,notn4796,n1737);
and (s1n4796,n3122,n1733);
and (n4797,n4798,n1002);
or (n4798,1'b0,n4799,n4801,n4803,n4805);
and (n4799,n4800,n3124);
wire s0n4800,s1n4800,notn4800;
or (n4800,s0n4800,s1n4800);
not(notn4800,n3122);
and (s0n4800,notn4800,n1743);
and (s1n4800,n3122,n1737);
and (n4801,n4802,n3136);
wire s0n4802,s1n4802,notn4802;
or (n4802,s0n4802,s1n4802);
not(notn4802,n3122);
and (s0n4802,notn4802,n1747);
and (s1n4802,n3122,n1743);
and (n4803,n4804,n3141);
wire s0n4804,s1n4804,notn4804;
or (n4804,s0n4804,s1n4804);
not(notn4804,n3122);
and (s0n4804,notn4804,n1751);
and (s1n4804,n3122,n1747);
and (n4805,n4806,n3146);
wire s0n4806,s1n4806,notn4806;
or (n4806,s0n4806,s1n4806);
not(notn4806,n3122);
and (s0n4806,notn4806,n1755);
and (s1n4806,n3122,n1751);
and (n4807,n4808,n1022);
or (n4808,1'b0,n4809,n4811,n4813,n4815);
and (n4809,n4810,n3124);
wire s0n4810,s1n4810,notn4810;
or (n4810,s0n4810,s1n4810);
not(notn4810,n3122);
and (s0n4810,notn4810,n1761);
and (s1n4810,n3122,n1813);
and (n4811,n4812,n3136);
wire s0n4812,s1n4812,notn4812;
or (n4812,s0n4812,s1n4812);
not(notn4812,n3122);
and (s0n4812,notn4812,n1765);
and (s1n4812,n3122,n1761);
and (n4813,n4814,n3141);
wire s0n4814,s1n4814,notn4814;
or (n4814,s0n4814,s1n4814);
not(notn4814,n3122);
and (s0n4814,notn4814,n1769);
and (s1n4814,n3122,n1765);
and (n4815,n4816,n3146);
wire s0n4816,s1n4816,notn4816;
or (n4816,s0n4816,s1n4816);
not(notn4816,n3122);
and (s0n4816,notn4816,n1773);
and (s1n4816,n3122,n1769);
and (n4817,n4818,n1042);
or (n4818,1'b0,n4819,n4821,n4823,n4825);
and (n4819,n4820,n3124);
wire s0n4820,s1n4820,notn4820;
or (n4820,s0n4820,s1n4820);
not(notn4820,n3122);
and (s0n4820,notn4820,n1779);
and (s1n4820,n3122,n1773);
and (n4821,n4822,n3136);
wire s0n4822,s1n4822,notn4822;
or (n4822,s0n4822,s1n4822);
not(notn4822,n3122);
and (s0n4822,notn4822,n1783);
and (s1n4822,n3122,n1779);
and (n4823,n4824,n3141);
wire s0n4824,s1n4824,notn4824;
or (n4824,s0n4824,s1n4824);
not(notn4824,n3122);
and (s0n4824,notn4824,n1787);
and (s1n4824,n3122,n1783);
and (n4825,n4826,n3146);
wire s0n4826,s1n4826,notn4826;
or (n4826,s0n4826,s1n4826);
not(notn4826,n3122);
and (s0n4826,notn4826,n1791);
and (s1n4826,n3122,n1787);
wire s0n4828,s1n4828,notn4828;
or (n4828,s0n4828,s1n4828);
not(notn4828,n3074);
and (s0n4828,notn4828,n4829);
and (s1n4828,n3074,n4870);
or (n4829,1'b0,n4830,n4840,n4850,n4860);
and (n4830,n4831,n981);
or (n4831,1'b0,n4832,n4834,n4836,n4838);
and (n4832,n4833,n3124);
wire s0n4833,s1n4833,notn4833;
or (n4833,s0n4833,s1n4833);
not(notn4833,n3122);
and (s0n4833,notn4833,n1726);
and (s1n4833,n3122,n1799);
and (n4834,n4835,n3136);
wire s0n4835,s1n4835,notn4835;
or (n4835,s0n4835,s1n4835);
not(notn4835,n3122);
and (s0n4835,notn4835,n1730);
and (s1n4835,n3122,n1726);
and (n4836,n4837,n3141);
wire s0n4837,s1n4837,notn4837;
or (n4837,s0n4837,s1n4837);
not(notn4837,n3122);
and (s0n4837,notn4837,n1734);
and (s1n4837,n3122,n1730);
and (n4838,n4839,n3146);
wire s0n4839,s1n4839,notn4839;
or (n4839,s0n4839,s1n4839);
not(notn4839,n3122);
and (s0n4839,notn4839,n1738);
and (s1n4839,n3122,n1734);
and (n4840,n4841,n1002);
or (n4841,1'b0,n4842,n4844,n4846,n4848);
and (n4842,n4843,n3124);
wire s0n4843,s1n4843,notn4843;
or (n4843,s0n4843,s1n4843);
not(notn4843,n3122);
and (s0n4843,notn4843,n1744);
and (s1n4843,n3122,n1738);
and (n4844,n4845,n3136);
wire s0n4845,s1n4845,notn4845;
or (n4845,s0n4845,s1n4845);
not(notn4845,n3122);
and (s0n4845,notn4845,n1748);
and (s1n4845,n3122,n1744);
and (n4846,n4847,n3141);
wire s0n4847,s1n4847,notn4847;
or (n4847,s0n4847,s1n4847);
not(notn4847,n3122);
and (s0n4847,notn4847,n1752);
and (s1n4847,n3122,n1748);
and (n4848,n4849,n3146);
wire s0n4849,s1n4849,notn4849;
or (n4849,s0n4849,s1n4849);
not(notn4849,n3122);
and (s0n4849,notn4849,n1756);
and (s1n4849,n3122,n1752);
and (n4850,n4851,n1022);
or (n4851,1'b0,n4852,n4854,n4856,n4858);
and (n4852,n4853,n3124);
wire s0n4853,s1n4853,notn4853;
or (n4853,s0n4853,s1n4853);
not(notn4853,n3122);
and (s0n4853,notn4853,n1762);
and (s1n4853,n3122,n1814);
and (n4854,n4855,n3136);
wire s0n4855,s1n4855,notn4855;
or (n4855,s0n4855,s1n4855);
not(notn4855,n3122);
and (s0n4855,notn4855,n1766);
and (s1n4855,n3122,n1762);
and (n4856,n4857,n3141);
wire s0n4857,s1n4857,notn4857;
or (n4857,s0n4857,s1n4857);
not(notn4857,n3122);
and (s0n4857,notn4857,n1770);
and (s1n4857,n3122,n1766);
and (n4858,n4859,n3146);
wire s0n4859,s1n4859,notn4859;
or (n4859,s0n4859,s1n4859);
not(notn4859,n3122);
and (s0n4859,notn4859,n1774);
and (s1n4859,n3122,n1770);
and (n4860,n4861,n1042);
or (n4861,1'b0,n4862,n4864,n4866,n4868);
and (n4862,n4863,n3124);
wire s0n4863,s1n4863,notn4863;
or (n4863,s0n4863,s1n4863);
not(notn4863,n3122);
and (s0n4863,notn4863,n1780);
and (s1n4863,n3122,n1774);
and (n4864,n4865,n3136);
wire s0n4865,s1n4865,notn4865;
or (n4865,s0n4865,s1n4865);
not(notn4865,n3122);
and (s0n4865,notn4865,n1784);
and (s1n4865,n3122,n1780);
and (n4866,n4867,n3141);
wire s0n4867,s1n4867,notn4867;
or (n4867,s0n4867,s1n4867);
not(notn4867,n3122);
and (s0n4867,notn4867,n1788);
and (s1n4867,n3122,n1784);
and (n4868,n4869,n3146);
wire s0n4869,s1n4869,notn4869;
or (n4869,s0n4869,s1n4869);
not(notn4869,n3122);
and (s0n4869,notn4869,n1792);
and (s1n4869,n3122,n1788);
and (n4871,n4697,n4784);
and (n4872,n4608,n4695);
and (n4873,n4519,n4606);
and (n4874,n4430,n4517);
and (n4875,n4341,n4428);
and (n4876,n4252,n4339);
and (n4877,n4163,n4250);
and (n4878,n4156,n4161);
and (n4879,n4149,n4154);
not (n4880,n4881);
xor (n4881,n4882,n4887);
xor (n4882,n4883,n4885);
wire s0n4883,s1n4883,notn4883;
or (n4883,s0n4883,s1n4883);
not(notn4883,n3074);
and (s0n4883,notn4883,1'b0);
and (s1n4883,n3074,n4884);
wire s0n4885,s1n4885,notn4885;
or (n4885,s0n4885,s1n4885);
not(notn4885,n3074);
and (s0n4885,notn4885,1'b0);
and (s1n4885,n3074,n4886);
or (n4887,n4888,n4893,n5491);
and (n4888,n4889,n4891);
wire s0n4889,s1n4889,notn4889;
or (n4889,s0n4889,s1n4889);
not(notn4889,n3074);
and (s0n4889,notn4889,1'b0);
and (s1n4889,n3074,n4890);
wire s0n4891,s1n4891,notn4891;
or (n4891,s0n4891,s1n4891);
not(notn4891,n3074);
and (s0n4891,notn4891,1'b0);
and (s1n4891,n3074,n4892);
and (n4893,n4891,n4894);
or (n4894,n4895,n4900,n5490);
and (n4895,n4896,n4898);
wire s0n4896,s1n4896,notn4896;
or (n4896,s0n4896,s1n4896);
not(notn4896,n3074);
and (s0n4896,notn4896,1'b0);
and (s1n4896,n3074,n4897);
wire s0n4898,s1n4898,notn4898;
or (n4898,s0n4898,s1n4898);
not(notn4898,n3074);
and (s0n4898,notn4898,1'b0);
and (s1n4898,n3074,n4899);
and (n4900,n4898,n4901);
or (n4901,n4902,n4907,n5489);
and (n4902,n4903,n4905);
wire s0n4903,s1n4903,notn4903;
or (n4903,s0n4903,s1n4903);
not(notn4903,n3074);
and (s0n4903,notn4903,1'b0);
and (s1n4903,n3074,n4904);
wire s0n4905,s1n4905,notn4905;
or (n4905,s0n4905,s1n4905);
not(notn4905,n3074);
and (s0n4905,notn4905,1'b0);
and (s1n4905,n3074,n4906);
and (n4907,n4905,n4908);
or (n4908,n4909,n4914,n5488);
and (n4909,n4910,n4912);
wire s0n4910,s1n4910,notn4910;
or (n4910,s0n4910,s1n4910);
not(notn4910,n3074);
and (s0n4910,notn4910,1'b0);
and (s1n4910,n3074,n4911);
wire s0n4912,s1n4912,notn4912;
or (n4912,s0n4912,s1n4912);
not(notn4912,n3074);
and (s0n4912,notn4912,1'b0);
and (s1n4912,n3074,n4913);
and (n4914,n4912,n4915);
or (n4915,n4916,n4985,n5487);
and (n4916,n4917,n4951);
wire s0n4917,s1n4917,notn4917;
or (n4917,s0n4917,s1n4917);
not(notn4917,n3074);
and (s0n4917,notn4917,n4918);
and (s1n4917,n3074,n4950);
or (n4918,1'b0,n4919,n4920,n4921,n4936);
and (n4919,n3224,n981);
and (n4920,n3239,n1002);
and (n4921,n4922,n1022);
or (n4922,1'b0,n4923,n4927,n4930,n4933);
and (n4923,n4924,n3124);
wire s0n4924,s1n4924,notn4924;
or (n4924,s0n4924,s1n4924);
not(notn4924,n3122);
and (s0n4924,notn4924,n4925);
and (s1n4924,n3122,n4926);
and (n4927,n4928,n3136);
wire s0n4928,s1n4928,notn4928;
or (n4928,s0n4928,s1n4928);
not(notn4928,n3122);
and (s0n4928,notn4928,n4929);
and (s1n4928,n3122,n4925);
and (n4930,n4931,n3141);
wire s0n4931,s1n4931,notn4931;
or (n4931,s0n4931,s1n4931);
not(notn4931,n3122);
and (s0n4931,notn4931,n4932);
and (s1n4931,n3122,n4929);
and (n4933,n4934,n3146);
wire s0n4934,s1n4934,notn4934;
or (n4934,s0n4934,s1n4934);
not(notn4934,n3122);
and (s0n4934,notn4934,n4935);
and (s1n4934,n3122,n4932);
and (n4936,n4937,n1042);
or (n4937,1'b0,n4938,n4941,n4944,n4947);
and (n4938,n4939,n3124);
wire s0n4939,s1n4939,notn4939;
or (n4939,s0n4939,s1n4939);
not(notn4939,n3122);
and (s0n4939,notn4939,n4940);
and (s1n4939,n3122,n4935);
and (n4941,n4942,n3136);
wire s0n4942,s1n4942,notn4942;
or (n4942,s0n4942,s1n4942);
not(notn4942,n3122);
and (s0n4942,notn4942,n4943);
and (s1n4942,n3122,n4940);
and (n4944,n4945,n3141);
wire s0n4945,s1n4945,notn4945;
or (n4945,s0n4945,s1n4945);
not(notn4945,n3122);
and (s0n4945,notn4945,n4946);
and (s1n4945,n3122,n4943);
and (n4947,n4948,n3146);
wire s0n4948,s1n4948,notn4948;
or (n4948,s0n4948,s1n4948);
not(notn4948,n3122);
and (s0n4948,notn4948,n4949);
and (s1n4948,n3122,n4946);
wire s0n4951,s1n4951,notn4951;
or (n4951,s0n4951,s1n4951);
not(notn4951,n3074);
and (s0n4951,notn4951,n4952);
and (s1n4951,n3074,n4984);
or (n4952,1'b0,n4953,n4968,n4982,n4983);
and (n4953,n4954,n981);
or (n4954,1'b0,n4955,n4959,n4962,n4965);
and (n4955,n4956,n3124);
wire s0n4956,s1n4956,notn4956;
or (n4956,s0n4956,s1n4956);
not(notn4956,n3122);
and (s0n4956,notn4956,n4957);
and (s1n4956,n3122,n4958);
and (n4959,n4960,n3136);
wire s0n4960,s1n4960,notn4960;
or (n4960,s0n4960,s1n4960);
not(notn4960,n3122);
and (s0n4960,notn4960,n4961);
and (s1n4960,n3122,n4957);
and (n4962,n4963,n3141);
wire s0n4963,s1n4963,notn4963;
or (n4963,s0n4963,s1n4963);
not(notn4963,n3122);
and (s0n4963,notn4963,n4964);
and (s1n4963,n3122,n4961);
and (n4965,n4966,n3146);
wire s0n4966,s1n4966,notn4966;
or (n4966,s0n4966,s1n4966);
not(notn4966,n3122);
and (s0n4966,notn4966,n4967);
and (s1n4966,n3122,n4964);
and (n4968,n4969,n1002);
or (n4969,1'b0,n4970,n4973,n4976,n4979);
and (n4970,n4971,n3124);
wire s0n4971,s1n4971,notn4971;
or (n4971,s0n4971,s1n4971);
not(notn4971,n3122);
and (s0n4971,notn4971,n4972);
and (s1n4971,n3122,n4967);
and (n4973,n4974,n3136);
wire s0n4974,s1n4974,notn4974;
or (n4974,s0n4974,s1n4974);
not(notn4974,n3122);
and (s0n4974,notn4974,n4975);
and (s1n4974,n3122,n4972);
and (n4976,n4977,n3141);
wire s0n4977,s1n4977,notn4977;
or (n4977,s0n4977,s1n4977);
not(notn4977,n3122);
and (s0n4977,notn4977,n4978);
and (s1n4977,n3122,n4975);
and (n4979,n4980,n3146);
wire s0n4980,s1n4980,notn4980;
or (n4980,s0n4980,s1n4980);
not(notn4980,n3122);
and (s0n4980,notn4980,n4981);
and (s1n4980,n3122,n4978);
and (n4982,n3117,n1022);
and (n4983,n3149,n1042);
and (n4985,n4951,n4986);
or (n4986,n4987,n5056,n5486);
and (n4987,n4988,n5022);
wire s0n4988,s1n4988,notn4988;
or (n4988,s0n4988,s1n4988);
not(notn4988,n3074);
and (s0n4988,notn4988,n4989);
and (s1n4988,n3074,n5021);
or (n4989,1'b0,n4990,n4991,n4992,n5007);
and (n4990,n3349,n981);
and (n4991,n3364,n1002);
and (n4992,n4993,n1022);
or (n4993,1'b0,n4994,n4998,n5001,n5004);
and (n4994,n4995,n3124);
wire s0n4995,s1n4995,notn4995;
or (n4995,s0n4995,s1n4995);
not(notn4995,n3122);
and (s0n4995,notn4995,n4996);
and (s1n4995,n3122,n4997);
and (n4998,n4999,n3136);
wire s0n4999,s1n4999,notn4999;
or (n4999,s0n4999,s1n4999);
not(notn4999,n3122);
and (s0n4999,notn4999,n5000);
and (s1n4999,n3122,n4996);
and (n5001,n5002,n3141);
wire s0n5002,s1n5002,notn5002;
or (n5002,s0n5002,s1n5002);
not(notn5002,n3122);
and (s0n5002,notn5002,n5003);
and (s1n5002,n3122,n5000);
and (n5004,n5005,n3146);
wire s0n5005,s1n5005,notn5005;
or (n5005,s0n5005,s1n5005);
not(notn5005,n3122);
and (s0n5005,notn5005,n5006);
and (s1n5005,n3122,n5003);
and (n5007,n5008,n1042);
or (n5008,1'b0,n5009,n5012,n5015,n5018);
and (n5009,n5010,n3124);
wire s0n5010,s1n5010,notn5010;
or (n5010,s0n5010,s1n5010);
not(notn5010,n3122);
and (s0n5010,notn5010,n5011);
and (s1n5010,n3122,n5006);
and (n5012,n5013,n3136);
wire s0n5013,s1n5013,notn5013;
or (n5013,s0n5013,s1n5013);
not(notn5013,n3122);
and (s0n5013,notn5013,n5014);
and (s1n5013,n3122,n5011);
and (n5015,n5016,n3141);
wire s0n5016,s1n5016,notn5016;
or (n5016,s0n5016,s1n5016);
not(notn5016,n3122);
and (s0n5016,notn5016,n5017);
and (s1n5016,n3122,n5014);
and (n5018,n5019,n3146);
wire s0n5019,s1n5019,notn5019;
or (n5019,s0n5019,s1n5019);
not(notn5019,n3122);
and (s0n5019,notn5019,n5020);
and (s1n5019,n3122,n5017);
wire s0n5022,s1n5022,notn5022;
or (n5022,s0n5022,s1n5022);
not(notn5022,n3074);
and (s0n5022,notn5022,n5023);
and (s1n5022,n3074,n5055);
or (n5023,1'b0,n5024,n5039,n5053,n5054);
and (n5024,n5025,n981);
or (n5025,1'b0,n5026,n5030,n5033,n5036);
and (n5026,n5027,n3124);
wire s0n5027,s1n5027,notn5027;
or (n5027,s0n5027,s1n5027);
not(notn5027,n3122);
and (s0n5027,notn5027,n5028);
and (s1n5027,n3122,n5029);
and (n5030,n5031,n3136);
wire s0n5031,s1n5031,notn5031;
or (n5031,s0n5031,s1n5031);
not(notn5031,n3122);
and (s0n5031,notn5031,n5032);
and (s1n5031,n3122,n5028);
and (n5033,n5034,n3141);
wire s0n5034,s1n5034,notn5034;
or (n5034,s0n5034,s1n5034);
not(notn5034,n3122);
and (s0n5034,notn5034,n5035);
and (s1n5034,n3122,n5032);
and (n5036,n5037,n3146);
wire s0n5037,s1n5037,notn5037;
or (n5037,s0n5037,s1n5037);
not(notn5037,n3122);
and (s0n5037,notn5037,n5038);
and (s1n5037,n3122,n5035);
and (n5039,n5040,n1002);
or (n5040,1'b0,n5041,n5044,n5047,n5050);
and (n5041,n5042,n3124);
wire s0n5042,s1n5042,notn5042;
or (n5042,s0n5042,s1n5042);
not(notn5042,n3122);
and (s0n5042,notn5042,n5043);
and (s1n5042,n3122,n5038);
and (n5044,n5045,n3136);
wire s0n5045,s1n5045,notn5045;
or (n5045,s0n5045,s1n5045);
not(notn5045,n3122);
and (s0n5045,notn5045,n5046);
and (s1n5045,n3122,n5043);
and (n5047,n5048,n3141);
wire s0n5048,s1n5048,notn5048;
or (n5048,s0n5048,s1n5048);
not(notn5048,n3122);
and (s0n5048,notn5048,n5049);
and (s1n5048,n3122,n5046);
and (n5050,n5051,n3146);
wire s0n5051,s1n5051,notn5051;
or (n5051,s0n5051,s1n5051);
not(notn5051,n3122);
and (s0n5051,notn5051,n5052);
and (s1n5051,n3122,n5049);
and (n5053,n3259,n1022);
and (n5054,n3274,n1042);
and (n5056,n5022,n5057);
or (n5057,n5058,n5127,n5485);
and (n5058,n5059,n5093);
wire s0n5059,s1n5059,notn5059;
or (n5059,s0n5059,s1n5059);
not(notn5059,n3074);
and (s0n5059,notn5059,n5060);
and (s1n5059,n3074,n5092);
or (n5060,1'b0,n5061,n5062,n5063,n5078);
and (n5061,n3474,n981);
and (n5062,n3489,n1002);
and (n5063,n5064,n1022);
or (n5064,1'b0,n5065,n5069,n5072,n5075);
and (n5065,n5066,n3124);
wire s0n5066,s1n5066,notn5066;
or (n5066,s0n5066,s1n5066);
not(notn5066,n3122);
and (s0n5066,notn5066,n5067);
and (s1n5066,n3122,n5068);
and (n5069,n5070,n3136);
wire s0n5070,s1n5070,notn5070;
or (n5070,s0n5070,s1n5070);
not(notn5070,n3122);
and (s0n5070,notn5070,n5071);
and (s1n5070,n3122,n5067);
and (n5072,n5073,n3141);
wire s0n5073,s1n5073,notn5073;
or (n5073,s0n5073,s1n5073);
not(notn5073,n3122);
and (s0n5073,notn5073,n5074);
and (s1n5073,n3122,n5071);
and (n5075,n5076,n3146);
wire s0n5076,s1n5076,notn5076;
or (n5076,s0n5076,s1n5076);
not(notn5076,n3122);
and (s0n5076,notn5076,n5077);
and (s1n5076,n3122,n5074);
and (n5078,n5079,n1042);
or (n5079,1'b0,n5080,n5083,n5086,n5089);
and (n5080,n5081,n3124);
wire s0n5081,s1n5081,notn5081;
or (n5081,s0n5081,s1n5081);
not(notn5081,n3122);
and (s0n5081,notn5081,n5082);
and (s1n5081,n3122,n5077);
and (n5083,n5084,n3136);
wire s0n5084,s1n5084,notn5084;
or (n5084,s0n5084,s1n5084);
not(notn5084,n3122);
and (s0n5084,notn5084,n5085);
and (s1n5084,n3122,n5082);
and (n5086,n5087,n3141);
wire s0n5087,s1n5087,notn5087;
or (n5087,s0n5087,s1n5087);
not(notn5087,n3122);
and (s0n5087,notn5087,n5088);
and (s1n5087,n3122,n5085);
and (n5089,n5090,n3146);
wire s0n5090,s1n5090,notn5090;
or (n5090,s0n5090,s1n5090);
not(notn5090,n3122);
and (s0n5090,notn5090,n5091);
and (s1n5090,n3122,n5088);
wire s0n5093,s1n5093,notn5093;
or (n5093,s0n5093,s1n5093);
not(notn5093,n3074);
and (s0n5093,notn5093,n5094);
and (s1n5093,n3074,n5126);
or (n5094,1'b0,n5095,n5110,n5124,n5125);
and (n5095,n5096,n981);
or (n5096,1'b0,n5097,n5101,n5104,n5107);
and (n5097,n5098,n3124);
wire s0n5098,s1n5098,notn5098;
or (n5098,s0n5098,s1n5098);
not(notn5098,n3122);
and (s0n5098,notn5098,n5099);
and (s1n5098,n3122,n5100);
and (n5101,n5102,n3136);
wire s0n5102,s1n5102,notn5102;
or (n5102,s0n5102,s1n5102);
not(notn5102,n3122);
and (s0n5102,notn5102,n5103);
and (s1n5102,n3122,n5099);
and (n5104,n5105,n3141);
wire s0n5105,s1n5105,notn5105;
or (n5105,s0n5105,s1n5105);
not(notn5105,n3122);
and (s0n5105,notn5105,n5106);
and (s1n5105,n3122,n5103);
and (n5107,n5108,n3146);
wire s0n5108,s1n5108,notn5108;
or (n5108,s0n5108,s1n5108);
not(notn5108,n3122);
and (s0n5108,notn5108,n5109);
and (s1n5108,n3122,n5106);
and (n5110,n5111,n1002);
or (n5111,1'b0,n5112,n5115,n5118,n5121);
and (n5112,n5113,n3124);
wire s0n5113,s1n5113,notn5113;
or (n5113,s0n5113,s1n5113);
not(notn5113,n3122);
and (s0n5113,notn5113,n5114);
and (s1n5113,n3122,n5109);
and (n5115,n5116,n3136);
wire s0n5116,s1n5116,notn5116;
or (n5116,s0n5116,s1n5116);
not(notn5116,n3122);
and (s0n5116,notn5116,n5117);
and (s1n5116,n3122,n5114);
and (n5118,n5119,n3141);
wire s0n5119,s1n5119,notn5119;
or (n5119,s0n5119,s1n5119);
not(notn5119,n3122);
and (s0n5119,notn5119,n5120);
and (s1n5119,n3122,n5117);
and (n5121,n5122,n3146);
wire s0n5122,s1n5122,notn5122;
or (n5122,s0n5122,s1n5122);
not(notn5122,n3122);
and (s0n5122,notn5122,n5123);
and (s1n5122,n3122,n5120);
and (n5124,n3384,n1022);
and (n5125,n3399,n1042);
and (n5127,n5093,n5128);
or (n5128,n5129,n5198,n5484);
and (n5129,n5130,n5164);
wire s0n5130,s1n5130,notn5130;
or (n5130,s0n5130,s1n5130);
not(notn5130,n3074);
and (s0n5130,notn5130,n5131);
and (s1n5130,n3074,n5163);
or (n5131,1'b0,n5132,n5133,n5134,n5149);
and (n5132,n3599,n981);
and (n5133,n3614,n1002);
and (n5134,n5135,n1022);
or (n5135,1'b0,n5136,n5140,n5143,n5146);
and (n5136,n5137,n3124);
wire s0n5137,s1n5137,notn5137;
or (n5137,s0n5137,s1n5137);
not(notn5137,n3122);
and (s0n5137,notn5137,n5138);
and (s1n5137,n3122,n5139);
and (n5140,n5141,n3136);
wire s0n5141,s1n5141,notn5141;
or (n5141,s0n5141,s1n5141);
not(notn5141,n3122);
and (s0n5141,notn5141,n5142);
and (s1n5141,n3122,n5138);
and (n5143,n5144,n3141);
wire s0n5144,s1n5144,notn5144;
or (n5144,s0n5144,s1n5144);
not(notn5144,n3122);
and (s0n5144,notn5144,n5145);
and (s1n5144,n3122,n5142);
and (n5146,n5147,n3146);
wire s0n5147,s1n5147,notn5147;
or (n5147,s0n5147,s1n5147);
not(notn5147,n3122);
and (s0n5147,notn5147,n5148);
and (s1n5147,n3122,n5145);
and (n5149,n5150,n1042);
or (n5150,1'b0,n5151,n5154,n5157,n5160);
and (n5151,n5152,n3124);
wire s0n5152,s1n5152,notn5152;
or (n5152,s0n5152,s1n5152);
not(notn5152,n3122);
and (s0n5152,notn5152,n5153);
and (s1n5152,n3122,n5148);
and (n5154,n5155,n3136);
wire s0n5155,s1n5155,notn5155;
or (n5155,s0n5155,s1n5155);
not(notn5155,n3122);
and (s0n5155,notn5155,n5156);
and (s1n5155,n3122,n5153);
and (n5157,n5158,n3141);
wire s0n5158,s1n5158,notn5158;
or (n5158,s0n5158,s1n5158);
not(notn5158,n3122);
and (s0n5158,notn5158,n5159);
and (s1n5158,n3122,n5156);
and (n5160,n5161,n3146);
wire s0n5161,s1n5161,notn5161;
or (n5161,s0n5161,s1n5161);
not(notn5161,n3122);
and (s0n5161,notn5161,n5162);
and (s1n5161,n3122,n5159);
wire s0n5164,s1n5164,notn5164;
or (n5164,s0n5164,s1n5164);
not(notn5164,n3074);
and (s0n5164,notn5164,n5165);
and (s1n5164,n3074,n5197);
or (n5165,1'b0,n5166,n5181,n5195,n5196);
and (n5166,n5167,n981);
or (n5167,1'b0,n5168,n5172,n5175,n5178);
and (n5168,n5169,n3124);
wire s0n5169,s1n5169,notn5169;
or (n5169,s0n5169,s1n5169);
not(notn5169,n3122);
and (s0n5169,notn5169,n5170);
and (s1n5169,n3122,n5171);
and (n5172,n5173,n3136);
wire s0n5173,s1n5173,notn5173;
or (n5173,s0n5173,s1n5173);
not(notn5173,n3122);
and (s0n5173,notn5173,n5174);
and (s1n5173,n3122,n5170);
and (n5175,n5176,n3141);
wire s0n5176,s1n5176,notn5176;
or (n5176,s0n5176,s1n5176);
not(notn5176,n3122);
and (s0n5176,notn5176,n5177);
and (s1n5176,n3122,n5174);
and (n5178,n5179,n3146);
wire s0n5179,s1n5179,notn5179;
or (n5179,s0n5179,s1n5179);
not(notn5179,n3122);
and (s0n5179,notn5179,n5180);
and (s1n5179,n3122,n5177);
and (n5181,n5182,n1002);
or (n5182,1'b0,n5183,n5186,n5189,n5192);
and (n5183,n5184,n3124);
wire s0n5184,s1n5184,notn5184;
or (n5184,s0n5184,s1n5184);
not(notn5184,n3122);
and (s0n5184,notn5184,n5185);
and (s1n5184,n3122,n5180);
and (n5186,n5187,n3136);
wire s0n5187,s1n5187,notn5187;
or (n5187,s0n5187,s1n5187);
not(notn5187,n3122);
and (s0n5187,notn5187,n5188);
and (s1n5187,n3122,n5185);
and (n5189,n5190,n3141);
wire s0n5190,s1n5190,notn5190;
or (n5190,s0n5190,s1n5190);
not(notn5190,n3122);
and (s0n5190,notn5190,n5191);
and (s1n5190,n3122,n5188);
and (n5192,n5193,n3146);
wire s0n5193,s1n5193,notn5193;
or (n5193,s0n5193,s1n5193);
not(notn5193,n3122);
and (s0n5193,notn5193,n5194);
and (s1n5193,n3122,n5191);
and (n5195,n3509,n1022);
and (n5196,n3524,n1042);
and (n5198,n5164,n5199);
or (n5199,n5200,n5269,n5483);
and (n5200,n5201,n5235);
wire s0n5201,s1n5201,notn5201;
or (n5201,s0n5201,s1n5201);
not(notn5201,n3074);
and (s0n5201,notn5201,n5202);
and (s1n5201,n3074,n5234);
or (n5202,1'b0,n5203,n5204,n5205,n5220);
and (n5203,n3724,n981);
and (n5204,n3739,n1002);
and (n5205,n5206,n1022);
or (n5206,1'b0,n5207,n5211,n5214,n5217);
and (n5207,n5208,n3124);
wire s0n5208,s1n5208,notn5208;
or (n5208,s0n5208,s1n5208);
not(notn5208,n3122);
and (s0n5208,notn5208,n5209);
and (s1n5208,n3122,n5210);
and (n5211,n5212,n3136);
wire s0n5212,s1n5212,notn5212;
or (n5212,s0n5212,s1n5212);
not(notn5212,n3122);
and (s0n5212,notn5212,n5213);
and (s1n5212,n3122,n5209);
and (n5214,n5215,n3141);
wire s0n5215,s1n5215,notn5215;
or (n5215,s0n5215,s1n5215);
not(notn5215,n3122);
and (s0n5215,notn5215,n5216);
and (s1n5215,n3122,n5213);
and (n5217,n5218,n3146);
wire s0n5218,s1n5218,notn5218;
or (n5218,s0n5218,s1n5218);
not(notn5218,n3122);
and (s0n5218,notn5218,n5219);
and (s1n5218,n3122,n5216);
and (n5220,n5221,n1042);
or (n5221,1'b0,n5222,n5225,n5228,n5231);
and (n5222,n5223,n3124);
wire s0n5223,s1n5223,notn5223;
or (n5223,s0n5223,s1n5223);
not(notn5223,n3122);
and (s0n5223,notn5223,n5224);
and (s1n5223,n3122,n5219);
and (n5225,n5226,n3136);
wire s0n5226,s1n5226,notn5226;
or (n5226,s0n5226,s1n5226);
not(notn5226,n3122);
and (s0n5226,notn5226,n5227);
and (s1n5226,n3122,n5224);
and (n5228,n5229,n3141);
wire s0n5229,s1n5229,notn5229;
or (n5229,s0n5229,s1n5229);
not(notn5229,n3122);
and (s0n5229,notn5229,n5230);
and (s1n5229,n3122,n5227);
and (n5231,n5232,n3146);
wire s0n5232,s1n5232,notn5232;
or (n5232,s0n5232,s1n5232);
not(notn5232,n3122);
and (s0n5232,notn5232,n5233);
and (s1n5232,n3122,n5230);
wire s0n5235,s1n5235,notn5235;
or (n5235,s0n5235,s1n5235);
not(notn5235,n3074);
and (s0n5235,notn5235,n5236);
and (s1n5235,n3074,n5268);
or (n5236,1'b0,n5237,n5252,n5266,n5267);
and (n5237,n5238,n981);
or (n5238,1'b0,n5239,n5243,n5246,n5249);
and (n5239,n5240,n3124);
wire s0n5240,s1n5240,notn5240;
or (n5240,s0n5240,s1n5240);
not(notn5240,n3122);
and (s0n5240,notn5240,n5241);
and (s1n5240,n3122,n5242);
and (n5243,n5244,n3136);
wire s0n5244,s1n5244,notn5244;
or (n5244,s0n5244,s1n5244);
not(notn5244,n3122);
and (s0n5244,notn5244,n5245);
and (s1n5244,n3122,n5241);
and (n5246,n5247,n3141);
wire s0n5247,s1n5247,notn5247;
or (n5247,s0n5247,s1n5247);
not(notn5247,n3122);
and (s0n5247,notn5247,n5248);
and (s1n5247,n3122,n5245);
and (n5249,n5250,n3146);
wire s0n5250,s1n5250,notn5250;
or (n5250,s0n5250,s1n5250);
not(notn5250,n3122);
and (s0n5250,notn5250,n5251);
and (s1n5250,n3122,n5248);
and (n5252,n5253,n1002);
or (n5253,1'b0,n5254,n5257,n5260,n5263);
and (n5254,n5255,n3124);
wire s0n5255,s1n5255,notn5255;
or (n5255,s0n5255,s1n5255);
not(notn5255,n3122);
and (s0n5255,notn5255,n5256);
and (s1n5255,n3122,n5251);
and (n5257,n5258,n3136);
wire s0n5258,s1n5258,notn5258;
or (n5258,s0n5258,s1n5258);
not(notn5258,n3122);
and (s0n5258,notn5258,n5259);
and (s1n5258,n3122,n5256);
and (n5260,n5261,n3141);
wire s0n5261,s1n5261,notn5261;
or (n5261,s0n5261,s1n5261);
not(notn5261,n3122);
and (s0n5261,notn5261,n5262);
and (s1n5261,n3122,n5259);
and (n5263,n5264,n3146);
wire s0n5264,s1n5264,notn5264;
or (n5264,s0n5264,s1n5264);
not(notn5264,n3122);
and (s0n5264,notn5264,n5265);
and (s1n5264,n3122,n5262);
and (n5266,n3634,n1022);
and (n5267,n3649,n1042);
and (n5269,n5235,n5270);
or (n5270,n5271,n5340,n5482);
and (n5271,n5272,n5306);
wire s0n5272,s1n5272,notn5272;
or (n5272,s0n5272,s1n5272);
not(notn5272,n3074);
and (s0n5272,notn5272,n5273);
and (s1n5272,n3074,n5305);
or (n5273,1'b0,n5274,n5275,n5276,n5291);
and (n5274,n3849,n981);
and (n5275,n3864,n1002);
and (n5276,n5277,n1022);
or (n5277,1'b0,n5278,n5282,n5285,n5288);
and (n5278,n5279,n3124);
wire s0n5279,s1n5279,notn5279;
or (n5279,s0n5279,s1n5279);
not(notn5279,n3122);
and (s0n5279,notn5279,n5280);
and (s1n5279,n3122,n5281);
and (n5282,n5283,n3136);
wire s0n5283,s1n5283,notn5283;
or (n5283,s0n5283,s1n5283);
not(notn5283,n3122);
and (s0n5283,notn5283,n5284);
and (s1n5283,n3122,n5280);
and (n5285,n5286,n3141);
wire s0n5286,s1n5286,notn5286;
or (n5286,s0n5286,s1n5286);
not(notn5286,n3122);
and (s0n5286,notn5286,n5287);
and (s1n5286,n3122,n5284);
and (n5288,n5289,n3146);
wire s0n5289,s1n5289,notn5289;
or (n5289,s0n5289,s1n5289);
not(notn5289,n3122);
and (s0n5289,notn5289,n5290);
and (s1n5289,n3122,n5287);
and (n5291,n5292,n1042);
or (n5292,1'b0,n5293,n5296,n5299,n5302);
and (n5293,n5294,n3124);
wire s0n5294,s1n5294,notn5294;
or (n5294,s0n5294,s1n5294);
not(notn5294,n3122);
and (s0n5294,notn5294,n5295);
and (s1n5294,n3122,n5290);
and (n5296,n5297,n3136);
wire s0n5297,s1n5297,notn5297;
or (n5297,s0n5297,s1n5297);
not(notn5297,n3122);
and (s0n5297,notn5297,n5298);
and (s1n5297,n3122,n5295);
and (n5299,n5300,n3141);
wire s0n5300,s1n5300,notn5300;
or (n5300,s0n5300,s1n5300);
not(notn5300,n3122);
and (s0n5300,notn5300,n5301);
and (s1n5300,n3122,n5298);
and (n5302,n5303,n3146);
wire s0n5303,s1n5303,notn5303;
or (n5303,s0n5303,s1n5303);
not(notn5303,n3122);
and (s0n5303,notn5303,n5304);
and (s1n5303,n3122,n5301);
wire s0n5306,s1n5306,notn5306;
or (n5306,s0n5306,s1n5306);
not(notn5306,n3074);
and (s0n5306,notn5306,n5307);
and (s1n5306,n3074,n5339);
or (n5307,1'b0,n5308,n5323,n5337,n5338);
and (n5308,n5309,n981);
or (n5309,1'b0,n5310,n5314,n5317,n5320);
and (n5310,n5311,n3124);
wire s0n5311,s1n5311,notn5311;
or (n5311,s0n5311,s1n5311);
not(notn5311,n3122);
and (s0n5311,notn5311,n5312);
and (s1n5311,n3122,n5313);
and (n5314,n5315,n3136);
wire s0n5315,s1n5315,notn5315;
or (n5315,s0n5315,s1n5315);
not(notn5315,n3122);
and (s0n5315,notn5315,n5316);
and (s1n5315,n3122,n5312);
and (n5317,n5318,n3141);
wire s0n5318,s1n5318,notn5318;
or (n5318,s0n5318,s1n5318);
not(notn5318,n3122);
and (s0n5318,notn5318,n5319);
and (s1n5318,n3122,n5316);
and (n5320,n5321,n3146);
wire s0n5321,s1n5321,notn5321;
or (n5321,s0n5321,s1n5321);
not(notn5321,n3122);
and (s0n5321,notn5321,n5322);
and (s1n5321,n3122,n5319);
and (n5323,n5324,n1002);
or (n5324,1'b0,n5325,n5328,n5331,n5334);
and (n5325,n5326,n3124);
wire s0n5326,s1n5326,notn5326;
or (n5326,s0n5326,s1n5326);
not(notn5326,n3122);
and (s0n5326,notn5326,n5327);
and (s1n5326,n3122,n5322);
and (n5328,n5329,n3136);
wire s0n5329,s1n5329,notn5329;
or (n5329,s0n5329,s1n5329);
not(notn5329,n3122);
and (s0n5329,notn5329,n5330);
and (s1n5329,n3122,n5327);
and (n5331,n5332,n3141);
wire s0n5332,s1n5332,notn5332;
or (n5332,s0n5332,s1n5332);
not(notn5332,n3122);
and (s0n5332,notn5332,n5333);
and (s1n5332,n3122,n5330);
and (n5334,n5335,n3146);
wire s0n5335,s1n5335,notn5335;
or (n5335,s0n5335,s1n5335);
not(notn5335,n3122);
and (s0n5335,notn5335,n5336);
and (s1n5335,n3122,n5333);
and (n5337,n3759,n1022);
and (n5338,n3774,n1042);
and (n5340,n5306,n5341);
or (n5341,n5342,n5411,n5481);
and (n5342,n5343,n5377);
wire s0n5343,s1n5343,notn5343;
or (n5343,s0n5343,s1n5343);
not(notn5343,n3074);
and (s0n5343,notn5343,n5344);
and (s1n5343,n3074,n5376);
or (n5344,1'b0,n5345,n5346,n5347,n5362);
and (n5345,n3974,n981);
and (n5346,n3989,n1002);
and (n5347,n5348,n1022);
or (n5348,1'b0,n5349,n5353,n5356,n5359);
and (n5349,n5350,n3124);
wire s0n5350,s1n5350,notn5350;
or (n5350,s0n5350,s1n5350);
not(notn5350,n3122);
and (s0n5350,notn5350,n5351);
and (s1n5350,n3122,n5352);
and (n5353,n5354,n3136);
wire s0n5354,s1n5354,notn5354;
or (n5354,s0n5354,s1n5354);
not(notn5354,n3122);
and (s0n5354,notn5354,n5355);
and (s1n5354,n3122,n5351);
and (n5356,n5357,n3141);
wire s0n5357,s1n5357,notn5357;
or (n5357,s0n5357,s1n5357);
not(notn5357,n3122);
and (s0n5357,notn5357,n5358);
and (s1n5357,n3122,n5355);
and (n5359,n5360,n3146);
wire s0n5360,s1n5360,notn5360;
or (n5360,s0n5360,s1n5360);
not(notn5360,n3122);
and (s0n5360,notn5360,n5361);
and (s1n5360,n3122,n5358);
and (n5362,n5363,n1042);
or (n5363,1'b0,n5364,n5367,n5370,n5373);
and (n5364,n5365,n3124);
wire s0n5365,s1n5365,notn5365;
or (n5365,s0n5365,s1n5365);
not(notn5365,n3122);
and (s0n5365,notn5365,n5366);
and (s1n5365,n3122,n5361);
and (n5367,n5368,n3136);
wire s0n5368,s1n5368,notn5368;
or (n5368,s0n5368,s1n5368);
not(notn5368,n3122);
and (s0n5368,notn5368,n5369);
and (s1n5368,n3122,n5366);
and (n5370,n5371,n3141);
wire s0n5371,s1n5371,notn5371;
or (n5371,s0n5371,s1n5371);
not(notn5371,n3122);
and (s0n5371,notn5371,n5372);
and (s1n5371,n3122,n5369);
and (n5373,n5374,n3146);
wire s0n5374,s1n5374,notn5374;
or (n5374,s0n5374,s1n5374);
not(notn5374,n3122);
and (s0n5374,notn5374,n5375);
and (s1n5374,n3122,n5372);
wire s0n5377,s1n5377,notn5377;
or (n5377,s0n5377,s1n5377);
not(notn5377,n3074);
and (s0n5377,notn5377,n5378);
and (s1n5377,n3074,n5410);
or (n5378,1'b0,n5379,n5394,n5408,n5409);
and (n5379,n5380,n981);
or (n5380,1'b0,n5381,n5385,n5388,n5391);
and (n5381,n5382,n3124);
wire s0n5382,s1n5382,notn5382;
or (n5382,s0n5382,s1n5382);
not(notn5382,n3122);
and (s0n5382,notn5382,n5383);
and (s1n5382,n3122,n5384);
and (n5385,n5386,n3136);
wire s0n5386,s1n5386,notn5386;
or (n5386,s0n5386,s1n5386);
not(notn5386,n3122);
and (s0n5386,notn5386,n5387);
and (s1n5386,n3122,n5383);
and (n5388,n5389,n3141);
wire s0n5389,s1n5389,notn5389;
or (n5389,s0n5389,s1n5389);
not(notn5389,n3122);
and (s0n5389,notn5389,n5390);
and (s1n5389,n3122,n5387);
and (n5391,n5392,n3146);
wire s0n5392,s1n5392,notn5392;
or (n5392,s0n5392,s1n5392);
not(notn5392,n3122);
and (s0n5392,notn5392,n5393);
and (s1n5392,n3122,n5390);
and (n5394,n5395,n1002);
or (n5395,1'b0,n5396,n5399,n5402,n5405);
and (n5396,n5397,n3124);
wire s0n5397,s1n5397,notn5397;
or (n5397,s0n5397,s1n5397);
not(notn5397,n3122);
and (s0n5397,notn5397,n5398);
and (s1n5397,n3122,n5393);
and (n5399,n5400,n3136);
wire s0n5400,s1n5400,notn5400;
or (n5400,s0n5400,s1n5400);
not(notn5400,n3122);
and (s0n5400,notn5400,n5401);
and (s1n5400,n3122,n5398);
and (n5402,n5403,n3141);
wire s0n5403,s1n5403,notn5403;
or (n5403,s0n5403,s1n5403);
not(notn5403,n3122);
and (s0n5403,notn5403,n5404);
and (s1n5403,n3122,n5401);
and (n5405,n5406,n3146);
wire s0n5406,s1n5406,notn5406;
or (n5406,s0n5406,s1n5406);
not(notn5406,n3122);
and (s0n5406,notn5406,n5407);
and (s1n5406,n3122,n5404);
and (n5408,n3884,n1022);
and (n5409,n3899,n1042);
and (n5411,n5377,n5412);
and (n5412,n5413,n5447);
wire s0n5413,s1n5413,notn5413;
or (n5413,s0n5413,s1n5413);
not(notn5413,n3074);
and (s0n5413,notn5413,n5414);
and (s1n5413,n3074,n5446);
or (n5414,1'b0,n5415,n5416,n5417,n5432);
and (n5415,n4098,n981);
and (n5416,n4113,n1002);
and (n5417,n5418,n1022);
or (n5418,1'b0,n5419,n5423,n5426,n5429);
and (n5419,n5420,n3124);
wire s0n5420,s1n5420,notn5420;
or (n5420,s0n5420,s1n5420);
not(notn5420,n3122);
and (s0n5420,notn5420,n5421);
and (s1n5420,n3122,n5422);
and (n5423,n5424,n3136);
wire s0n5424,s1n5424,notn5424;
or (n5424,s0n5424,s1n5424);
not(notn5424,n3122);
and (s0n5424,notn5424,n5425);
and (s1n5424,n3122,n5421);
and (n5426,n5427,n3141);
wire s0n5427,s1n5427,notn5427;
or (n5427,s0n5427,s1n5427);
not(notn5427,n3122);
and (s0n5427,notn5427,n5428);
and (s1n5427,n3122,n5425);
and (n5429,n5430,n3146);
wire s0n5430,s1n5430,notn5430;
or (n5430,s0n5430,s1n5430);
not(notn5430,n3122);
and (s0n5430,notn5430,n5431);
and (s1n5430,n3122,n5428);
and (n5432,n5433,n1042);
or (n5433,1'b0,n5434,n5437,n5440,n5443);
and (n5434,n5435,n3124);
wire s0n5435,s1n5435,notn5435;
or (n5435,s0n5435,s1n5435);
not(notn5435,n3122);
and (s0n5435,notn5435,n5436);
and (s1n5435,n3122,n5431);
and (n5437,n5438,n3136);
wire s0n5438,s1n5438,notn5438;
or (n5438,s0n5438,s1n5438);
not(notn5438,n3122);
and (s0n5438,notn5438,n5439);
and (s1n5438,n3122,n5436);
and (n5440,n5441,n3141);
wire s0n5441,s1n5441,notn5441;
or (n5441,s0n5441,s1n5441);
not(notn5441,n3122);
and (s0n5441,notn5441,n5442);
and (s1n5441,n3122,n5439);
and (n5443,n5444,n3146);
wire s0n5444,s1n5444,notn5444;
or (n5444,s0n5444,s1n5444);
not(notn5444,n3122);
and (s0n5444,notn5444,n5445);
and (s1n5444,n3122,n5442);
wire s0n5447,s1n5447,notn5447;
or (n5447,s0n5447,s1n5447);
not(notn5447,n3074);
and (s0n5447,notn5447,n5448);
and (s1n5447,n3074,n5480);
or (n5448,1'b0,n5449,n5464,n5478,n5479);
and (n5449,n5450,n981);
or (n5450,1'b0,n5451,n5455,n5458,n5461);
and (n5451,n5452,n3124);
wire s0n5452,s1n5452,notn5452;
or (n5452,s0n5452,s1n5452);
not(notn5452,n3122);
and (s0n5452,notn5452,n5453);
and (s1n5452,n3122,n5454);
and (n5455,n5456,n3136);
wire s0n5456,s1n5456,notn5456;
or (n5456,s0n5456,s1n5456);
not(notn5456,n3122);
and (s0n5456,notn5456,n5457);
and (s1n5456,n3122,n5453);
and (n5458,n5459,n3141);
wire s0n5459,s1n5459,notn5459;
or (n5459,s0n5459,s1n5459);
not(notn5459,n3122);
and (s0n5459,notn5459,n5460);
and (s1n5459,n3122,n5457);
and (n5461,n5462,n3146);
wire s0n5462,s1n5462,notn5462;
or (n5462,s0n5462,s1n5462);
not(notn5462,n3122);
and (s0n5462,notn5462,n5463);
and (s1n5462,n3122,n5460);
and (n5464,n5465,n1002);
or (n5465,1'b0,n5466,n5469,n5472,n5475);
and (n5466,n5467,n3124);
wire s0n5467,s1n5467,notn5467;
or (n5467,s0n5467,s1n5467);
not(notn5467,n3122);
and (s0n5467,notn5467,n5468);
and (s1n5467,n3122,n5463);
and (n5469,n5470,n3136);
wire s0n5470,s1n5470,notn5470;
or (n5470,s0n5470,s1n5470);
not(notn5470,n3122);
and (s0n5470,notn5470,n5471);
and (s1n5470,n3122,n5468);
and (n5472,n5473,n3141);
wire s0n5473,s1n5473,notn5473;
or (n5473,s0n5473,s1n5473);
not(notn5473,n3122);
and (s0n5473,notn5473,n5474);
and (s1n5473,n3122,n5471);
and (n5475,n5476,n3146);
wire s0n5476,s1n5476,notn5476;
or (n5476,s0n5476,s1n5476);
not(notn5476,n3122);
and (s0n5476,notn5476,n5477);
and (s1n5476,n3122,n5474);
and (n5478,n4008,n1022);
and (n5479,n4023,n1042);
and (n5481,n5343,n5412);
and (n5482,n5272,n5341);
and (n5483,n5201,n5270);
and (n5484,n5130,n5199);
and (n5485,n5059,n5128);
and (n5486,n4988,n5057);
and (n5487,n4917,n4986);
and (n5488,n4910,n4915);
and (n5489,n4903,n4908);
and (n5490,n4896,n4901);
and (n5491,n4889,n4894);
or (n5492,n5493,n5499,n5577);
and (n5493,n5494,n5496);
xor (n5494,n5495,n4154);
xor (n5495,n4149,n4151);
not (n5496,n5497);
xor (n5497,n5498,n4894);
xor (n5498,n4889,n4891);
and (n5499,n5496,n5500);
or (n5500,n5501,n5507,n5576);
and (n5501,n5502,n5504);
xor (n5502,n5503,n4161);
xor (n5503,n4156,n4158);
not (n5504,n5505);
xor (n5505,n5506,n4901);
xor (n5506,n4896,n4898);
and (n5507,n5504,n5508);
or (n5508,n5509,n5515,n5575);
and (n5509,n5510,n5512);
xor (n5510,n5511,n4250);
xor (n5511,n4163,n4206);
not (n5512,n5513);
xor (n5513,n5514,n4908);
xor (n5514,n4903,n4905);
and (n5515,n5512,n5516);
or (n5516,n5517,n5523,n5574);
and (n5517,n5518,n5520);
xor (n5518,n5519,n4339);
xor (n5519,n4252,n4295);
not (n5520,n5521);
xor (n5521,n5522,n4915);
xor (n5522,n4910,n4912);
and (n5523,n5520,n5524);
or (n5524,n5525,n5531,n5573);
and (n5525,n5526,n5528);
xor (n5526,n5527,n4428);
xor (n5527,n4341,n4384);
not (n5528,n5529);
xor (n5529,n5530,n4986);
xor (n5530,n4917,n4951);
and (n5531,n5528,n5532);
or (n5532,n5533,n5539,n5572);
and (n5533,n5534,n5536);
xor (n5534,n5535,n4517);
xor (n5535,n4430,n4473);
not (n5536,n5537);
xor (n5537,n5538,n5057);
xor (n5538,n4988,n5022);
and (n5539,n5536,n5540);
or (n5540,n5541,n5547,n5571);
and (n5541,n5542,n5544);
xor (n5542,n5543,n4606);
xor (n5543,n4519,n4562);
not (n5544,n5545);
xor (n5545,n5546,n5128);
xor (n5546,n5059,n5093);
and (n5547,n5544,n5548);
or (n5548,n5549,n5555,n5570);
and (n5549,n5550,n5552);
xor (n5550,n5551,n4695);
xor (n5551,n4608,n4651);
not (n5552,n5553);
xor (n5553,n5554,n5199);
xor (n5554,n5130,n5164);
and (n5555,n5552,n5556);
or (n5556,n5557,n5563,n5569);
and (n5557,n5558,n5560);
xor (n5558,n5559,n4784);
xor (n5559,n4697,n4740);
not (n5560,n5561);
xor (n5561,n5562,n5270);
xor (n5562,n5201,n5235);
and (n5563,n5560,n5564);
and (n5564,n5565,n5566);
xor (n5565,n4785,n4828);
not (n5566,n5567);
xor (n5567,n5568,n5341);
xor (n5568,n5272,n5306);
and (n5569,n5558,n5564);
and (n5570,n5550,n5556);
and (n5571,n5542,n5548);
and (n5572,n5534,n5540);
and (n5573,n5526,n5532);
and (n5574,n5518,n5524);
and (n5575,n5510,n5516);
and (n5576,n5502,n5508);
and (n5577,n5494,n5500);
and (n5578,n5579,n5581);
xor (n5579,n5580,n5500);
xor (n5580,n5494,n5496);
and (n5581,n5582,n5584);
xor (n5582,n5583,n5508);
xor (n5583,n5502,n5504);
and (n5584,n5585,n5587);
xor (n5585,n5586,n5516);
xor (n5586,n5510,n5512);
and (n5587,n5588,n5590);
xor (n5588,n5589,n5524);
xor (n5589,n5518,n5520);
and (n5590,n5591,n5593);
xor (n5591,n5592,n5532);
xor (n5592,n5526,n5528);
and (n5593,n5594,n5596);
xor (n5594,n5595,n5540);
xor (n5595,n5534,n5536);
and (n5596,n5597,n5599);
xor (n5597,n5598,n5548);
xor (n5598,n5542,n5544);
and (n5599,n5600,n5602);
xor (n5600,n5601,n5556);
xor (n5601,n5550,n5552);
and (n5602,n5603,n5605);
xor (n5603,n5604,n5564);
xor (n5604,n5558,n5560);
and (n5605,n5606,n5607);
xor (n5606,n5565,n5566);
and (n5607,n5608,n5611);
not (n5608,n5609);
xor (n5609,n5610,n5412);
xor (n5610,n5343,n5377);
not (n5611,n5612);
xor (n5612,n5413,n5447);
or (n5613,n5614,n5618,n5691);
and (n5614,n5615,n5617);
xor (n5615,n5616,n3091);
xor (n5616,n3086,n3088);
xor (n5617,n5579,n5581);
and (n5618,n5617,n5619);
or (n5619,n5620,n5624,n5690);
and (n5620,n5621,n5623);
xor (n5621,n5622,n3098);
xor (n5622,n3093,n3095);
xor (n5623,n5582,n5584);
and (n5624,n5623,n5625);
or (n5625,n5626,n5630,n5689);
and (n5626,n5627,n5629);
xor (n5627,n5628,n3105);
xor (n5628,n3100,n3102);
xor (n5629,n5585,n5587);
and (n5630,n5629,n5631);
or (n5631,n5632,n5636,n5688);
and (n5632,n5633,n5635);
xor (n5633,n5634,n3112);
xor (n5634,n3107,n3109);
xor (n5635,n5588,n5590);
and (n5636,n5635,n5637);
or (n5637,n5638,n5642,n5687);
and (n5638,n5639,n5641);
xor (n5639,n5640,n3254);
xor (n5640,n3114,n3192);
xor (n5641,n5591,n5593);
and (n5642,n5641,n5643);
or (n5643,n5644,n5648,n5686);
and (n5644,n5645,n5647);
xor (n5645,n5646,n3379);
xor (n5646,n3256,n3317);
xor (n5647,n5594,n5596);
and (n5648,n5647,n5649);
or (n5649,n5650,n5654,n5685);
and (n5650,n5651,n5653);
xor (n5651,n5652,n3504);
xor (n5652,n3381,n3442);
xor (n5653,n5597,n5599);
and (n5654,n5653,n5655);
or (n5655,n5656,n5660,n5684);
and (n5656,n5657,n5659);
xor (n5657,n5658,n3629);
xor (n5658,n3506,n3567);
xor (n5659,n5600,n5602);
and (n5660,n5659,n5661);
or (n5661,n5662,n5666,n5683);
and (n5662,n5663,n5665);
xor (n5663,n5664,n3754);
xor (n5664,n3631,n3692);
xor (n5665,n5603,n5605);
and (n5666,n5665,n5667);
or (n5667,n5668,n5672,n5682);
and (n5668,n5669,n5671);
xor (n5669,n5670,n3879);
xor (n5670,n3756,n3817);
xor (n5671,n5606,n5607);
and (n5672,n5671,n5673);
or (n5673,n5674,n5678,n5681);
and (n5674,n5675,n5677);
xor (n5675,n5676,n4004);
xor (n5676,n3881,n3942);
xor (n5677,n5608,n5611);
and (n5678,n5677,n5679);
and (n5679,n5680,n5612);
xor (n5680,n4005,n4066);
and (n5681,n5675,n5679);
and (n5682,n5669,n5673);
and (n5683,n5663,n5667);
and (n5684,n5657,n5661);
and (n5685,n5651,n5655);
and (n5686,n5645,n5649);
and (n5687,n5639,n5643);
and (n5688,n5633,n5637);
and (n5689,n5627,n5631);
and (n5690,n5621,n5625);
and (n5691,n5615,n5619);
or (n5692,n5693,n5696,n5748);
and (n5693,n5694,n5629);
xor (n5694,n5695,n5619);
xor (n5695,n5615,n5617);
and (n5696,n5629,n5697);
or (n5697,n5698,n5701,n5747);
and (n5698,n5699,n5635);
xor (n5699,n5700,n5625);
xor (n5700,n5621,n5623);
and (n5701,n5635,n5702);
or (n5702,n5703,n5706,n5746);
and (n5703,n5704,n5641);
xor (n5704,n5705,n5631);
xor (n5705,n5627,n5629);
and (n5706,n5641,n5707);
or (n5707,n5708,n5711,n5745);
and (n5708,n5709,n5647);
xor (n5709,n5710,n5637);
xor (n5710,n5633,n5635);
and (n5711,n5647,n5712);
or (n5712,n5713,n5716,n5744);
and (n5713,n5714,n5653);
xor (n5714,n5715,n5643);
xor (n5715,n5639,n5641);
and (n5716,n5653,n5717);
or (n5717,n5718,n5721,n5743);
and (n5718,n5719,n5659);
xor (n5719,n5720,n5649);
xor (n5720,n5645,n5647);
and (n5721,n5659,n5722);
or (n5722,n5723,n5726,n5742);
and (n5723,n5724,n5665);
xor (n5724,n5725,n5655);
xor (n5725,n5651,n5653);
and (n5726,n5665,n5727);
or (n5727,n5728,n5731,n5741);
and (n5728,n5729,n5671);
xor (n5729,n5730,n5661);
xor (n5730,n5657,n5659);
and (n5731,n5671,n5732);
or (n5732,n5733,n5736,n5740);
and (n5733,n5734,n5677);
xor (n5734,n5735,n5667);
xor (n5735,n5663,n5665);
and (n5736,n5677,n5737);
and (n5737,n5738,n5612);
xor (n5738,n5739,n5673);
xor (n5739,n5669,n5671);
and (n5740,n5734,n5737);
and (n5741,n5729,n5732);
and (n5742,n5724,n5727);
and (n5743,n5719,n5722);
and (n5744,n5714,n5717);
and (n5745,n5709,n5712);
and (n5746,n5704,n5707);
and (n5747,n5699,n5702);
and (n5748,n5694,n5697);
and (n5749,n5750,n5752);
xor (n5750,n5751,n5697);
xor (n5751,n5694,n5629);
and (n5752,n5753,n5755);
xor (n5753,n5754,n5702);
xor (n5754,n5699,n5635);
and (n5755,n5756,n5758);
xor (n5756,n5757,n5707);
xor (n5757,n5704,n5641);
and (n5758,n5759,n5761);
xor (n5759,n5760,n5712);
xor (n5760,n5709,n5647);
and (n5761,n5762,n5764);
xor (n5762,n5763,n5717);
xor (n5763,n5714,n5653);
and (n5764,n5765,n5767);
xor (n5765,n5766,n5722);
xor (n5766,n5719,n5659);
and (n5767,n5768,n5770);
xor (n5768,n5769,n5727);
xor (n5769,n5724,n5665);
xor (n5770,n5771,n5732);
xor (n5771,n5729,n5671);
xor (n5772,n3066,n5773);
and (n5773,n5750,n5774);
and (n5774,n5753,n5756);
wire s0n5775,s1n5775,notn5775;
or (n5775,s0n5775,s1n5775);
not(notn5775,n3074);
and (s0n5775,notn5775,n5776);
and (s1n5775,n3074,n5980);
xor (n5776,n5777,n5967);
xor (n5777,n5778,n5939);
xor (n5778,n5779,n5918);
xor (n5779,n5780,n5912);
xor (n5780,n5781,n5803);
xor (n5781,n5782,n5787);
xor (n5782,n5783,n5785);
wire s0n5783,s1n5783,notn5783;
or (n5783,s0n5783,s1n5783);
not(notn5783,n3074);
and (s0n5783,notn5783,1'b0);
and (s1n5783,n3074,n5784);
wire s0n5785,s1n5785,notn5785;
or (n5785,s0n5785,s1n5785);
not(notn5785,n3074);
and (s0n5785,notn5785,1'b0);
and (s1n5785,n3074,n5786);
or (n5787,n5788,n5789,n5802);
and (n5788,n5783,n5785);
and (n5789,n5785,n5790);
or (n5790,n5791,n5796,n5801);
and (n5791,n5792,n5794);
wire s0n5792,s1n5792,notn5792;
or (n5792,s0n5792,s1n5792);
not(notn5792,n3074);
and (s0n5792,notn5792,1'b0);
and (s1n5792,n3074,n5793);
wire s0n5794,s1n5794,notn5794;
or (n5794,s0n5794,s1n5794);
not(notn5794,n3074);
and (s0n5794,notn5794,1'b0);
and (s1n5794,n3074,n5795);
and (n5796,n5794,n5797);
or (n5797,n5798,n5799,n5800);
and (n5798,n3072,n3082);
and (n5799,n3082,n3084);
and (n5800,n3072,n3084);
and (n5801,n5792,n5797);
and (n5802,n5783,n5790);
xor (n5803,n5804,n5899);
xor (n5804,n5805,n5867);
xor (n5805,n5806,n5844);
xor (n5806,n5807,n5812);
xor (n5807,n5808,n5810);
wire s0n5808,s1n5808,notn5808;
or (n5808,s0n5808,s1n5808);
not(notn5808,n3074);
and (s0n5808,notn5808,1'b0);
and (s1n5808,n3074,n5809);
wire s0n5810,s1n5810,notn5810;
or (n5810,s0n5810,s1n5810);
not(notn5810,n3074);
and (s0n5810,notn5810,1'b0);
and (s1n5810,n3074,n5811);
or (n5812,n5813,n5814,n5843);
and (n5813,n5808,n5810);
and (n5814,n5810,n5815);
or (n5815,n5816,n5821,n5842);
and (n5816,n5817,n5819);
wire s0n5817,s1n5817,notn5817;
or (n5817,s0n5817,s1n5817);
not(notn5817,n3074);
and (s0n5817,notn5817,1'b0);
and (s1n5817,n3074,n5818);
wire s0n5819,s1n5819,notn5819;
or (n5819,s0n5819,s1n5819);
not(notn5819,n3074);
and (s0n5819,notn5819,1'b0);
and (s1n5819,n3074,n5820);
and (n5821,n5819,n5822);
or (n5822,n5823,n5828,n5841);
and (n5823,n5824,n5826);
wire s0n5824,s1n5824,notn5824;
or (n5824,s0n5824,s1n5824);
not(notn5824,n3074);
and (s0n5824,notn5824,1'b0);
and (s1n5824,n3074,n5825);
wire s0n5826,s1n5826,notn5826;
or (n5826,s0n5826,s1n5826);
not(notn5826,n3074);
and (s0n5826,notn5826,1'b0);
and (s1n5826,n3074,n5827);
and (n5828,n5826,n5829);
or (n5829,n5830,n5835,n5840);
and (n5830,n5831,n5833);
wire s0n5831,s1n5831,notn5831;
or (n5831,s0n5831,s1n5831);
not(notn5831,n3074);
and (s0n5831,notn5831,1'b0);
and (s1n5831,n3074,n5832);
wire s0n5833,s1n5833,notn5833;
or (n5833,s0n5833,s1n5833);
not(notn5833,n3074);
and (s0n5833,notn5833,1'b0);
and (s1n5833,n3074,n5834);
and (n5835,n5833,n5836);
or (n5836,n5837,n5838,n5839);
and (n5837,n4143,n4145);
and (n5838,n4145,n4147);
and (n5839,n4143,n4147);
and (n5840,n5831,n5836);
and (n5841,n5824,n5829);
and (n5842,n5817,n5822);
and (n5843,n5808,n5815);
not (n5844,n5845);
xor (n5845,n5846,n5851);
xor (n5846,n5847,n5849);
wire s0n5847,s1n5847,notn5847;
or (n5847,s0n5847,s1n5847);
not(notn5847,n3074);
and (s0n5847,notn5847,1'b0);
and (s1n5847,n3074,n5848);
wire s0n5849,s1n5849,notn5849;
or (n5849,s0n5849,s1n5849);
not(notn5849,n3074);
and (s0n5849,notn5849,1'b0);
and (s1n5849,n3074,n5850);
or (n5851,n5852,n5853,n5866);
and (n5852,n5847,n5849);
and (n5853,n5849,n5854);
or (n5854,n5855,n5860,n5865);
and (n5855,n5856,n5858);
wire s0n5856,s1n5856,notn5856;
or (n5856,s0n5856,s1n5856);
not(notn5856,n3074);
and (s0n5856,notn5856,1'b0);
and (s1n5856,n3074,n5857);
wire s0n5858,s1n5858,notn5858;
or (n5858,s0n5858,s1n5858);
not(notn5858,n3074);
and (s0n5858,notn5858,1'b0);
and (s1n5858,n3074,n5859);
and (n5860,n5858,n5861);
or (n5861,n5862,n5863,n5864);
and (n5862,n4883,n4885);
and (n5863,n4885,n4887);
and (n5864,n4883,n4887);
and (n5865,n5856,n5861);
and (n5866,n5847,n5854);
or (n5867,n5868,n5870,n5898);
and (n5868,n5869,n5844);
xor (n5869,n5807,n5815);
and (n5870,n5844,n5871);
or (n5871,n5872,n5875,n5897);
and (n5872,n5873,n5844);
xor (n5873,n5874,n5822);
xor (n5874,n5817,n5819);
and (n5875,n5844,n5876);
or (n5876,n5877,n5882,n5896);
and (n5877,n5878,n5880);
xor (n5878,n5879,n5829);
xor (n5879,n5824,n5826);
not (n5880,n5881);
xor (n5881,n5846,n5854);
and (n5882,n5880,n5883);
or (n5883,n5884,n5890,n5895);
and (n5884,n5885,n5887);
xor (n5885,n5886,n5836);
xor (n5886,n5831,n5833);
not (n5887,n5888);
xor (n5888,n5889,n5861);
xor (n5889,n5856,n5858);
and (n5890,n5887,n5891);
or (n5891,n5892,n5893,n5894);
and (n5892,n4141,n4880);
and (n5893,n4880,n5492);
and (n5894,n4141,n5492);
and (n5895,n5885,n5891);
and (n5896,n5878,n5883);
and (n5897,n5873,n5876);
and (n5898,n5869,n5871);
and (n5899,n5900,n5902);
xor (n5900,n5901,n5871);
xor (n5901,n5869,n5844);
and (n5902,n5903,n5905);
xor (n5903,n5904,n5876);
xor (n5904,n5873,n5844);
and (n5905,n5906,n5908);
xor (n5906,n5907,n5883);
xor (n5907,n5878,n5880);
and (n5908,n5909,n5911);
xor (n5909,n5910,n5891);
xor (n5910,n5885,n5887);
and (n5911,n4139,n5578);
or (n5912,n5913,n5915,n5938);
and (n5913,n5781,n5914);
xor (n5914,n5900,n5902);
and (n5915,n5914,n5916);
or (n5916,n5917,n5919,n5937);
and (n5917,n5781,n5918);
xor (n5918,n5903,n5905);
and (n5919,n5918,n5920);
or (n5920,n5921,n5924,n5936);
and (n5921,n5922,n5923);
xor (n5922,n5782,n5790);
xor (n5923,n5906,n5908);
and (n5924,n5923,n5925);
or (n5925,n5926,n5930,n5935);
and (n5926,n5927,n5929);
xor (n5927,n5928,n5797);
xor (n5928,n5792,n5794);
xor (n5929,n5909,n5911);
and (n5930,n5929,n5931);
or (n5931,n5932,n5933,n5934);
and (n5932,n3070,n4138);
and (n5933,n4138,n5613);
and (n5934,n3070,n5613);
and (n5935,n5927,n5931);
and (n5936,n5922,n5925);
and (n5937,n5781,n5920);
and (n5938,n5781,n5916);
or (n5939,n5940,n5943,n5966);
and (n5940,n5941,n5923);
xor (n5941,n5942,n5916);
xor (n5942,n5781,n5914);
and (n5943,n5923,n5944);
or (n5944,n5945,n5948,n5965);
and (n5945,n5946,n5929);
xor (n5946,n5947,n5920);
xor (n5947,n5781,n5918);
and (n5948,n5929,n5949);
or (n5949,n5950,n5953,n5964);
and (n5950,n5951,n4138);
xor (n5951,n5952,n5925);
xor (n5952,n5922,n5923);
and (n5953,n4138,n5954);
or (n5954,n5955,n5958,n5963);
and (n5955,n5956,n5617);
xor (n5956,n5957,n5931);
xor (n5957,n5927,n5929);
and (n5958,n5617,n5959);
or (n5959,n5960,n5961,n5962);
and (n5960,n3068,n5623);
and (n5961,n5623,n5692);
and (n5962,n3068,n5692);
and (n5963,n5956,n5959);
and (n5964,n5951,n5954);
and (n5965,n5946,n5949);
and (n5966,n5941,n5944);
and (n5967,n5968,n5970);
xor (n5968,n5969,n5944);
xor (n5969,n5941,n5923);
and (n5970,n5971,n5973);
xor (n5971,n5972,n5949);
xor (n5972,n5946,n5929);
and (n5973,n5974,n5976);
xor (n5974,n5975,n5954);
xor (n5975,n5951,n4138);
and (n5976,n5977,n5979);
xor (n5977,n5978,n5959);
xor (n5978,n5956,n5617);
and (n5979,n3066,n5749);
xor (n5980,n5777,n5981);
and (n5981,n5968,n5982);
and (n5982,n5971,n5983);
and (n5983,n5974,n5984);
and (n5984,n5977,n5985);
and (n5985,n3066,n5773);
wire s0n5986,s1n5986,notn5986;
or (n5986,s0n5986,s1n5986);
not(notn5986,n3074);
and (s0n5986,notn5986,n5987);
and (s1n5986,n3074,n5990);
wire s0n5987,s1n5987,notn5987;
or (n5987,s0n5987,s1n5987);
not(notn5987,n3074);
and (s0n5987,notn5987,n5988);
and (s1n5987,n3074,n5989);
xor (n5988,n5977,n5979);
xor (n5989,n5977,n5985);
wire s0n5990,s1n5990,notn5990;
or (n5990,s0n5990,s1n5990);
not(notn5990,n3074);
and (s0n5990,notn5990,n5991);
and (s1n5990,n3074,n5999);
xor (n5991,n5992,n5998);
xor (n5992,n5993,n5994);
xor (n5993,n5779,n5914);
or (n5994,n5995,n5996,n5997);
and (n5995,n5779,n5918);
and (n5996,n5918,n5939);
and (n5997,n5779,n5939);
and (n5998,n5777,n5967);
xor (n5999,n5992,n6000);
and (n6000,n5777,n5981);
wire s0n6001,s1n6001,notn6001;
or (n6001,s0n6001,s1n6001);
not(notn6001,n3074);
and (s0n6001,notn6001,n6002);
and (s1n6001,n3074,n6010);
xor (n6002,n6003,n6009);
xor (n6003,n6004,n6005);
xor (n6004,n5779,n5803);
or (n6005,n6006,n6007,n6008);
and (n6006,n5779,n5914);
and (n6007,n5914,n5994);
and (n6008,n5779,n5994);
and (n6009,n5992,n5998);
xor (n6010,n6003,n6011);
and (n6011,n5992,n6000);
and (n6012,n6013,n904);
wire s0n6013,s1n6013,notn6013;
or (n6013,s0n6013,s1n6013);
not(notn6013,n896);
and (s0n6013,notn6013,1'b0);
and (s1n6013,n896,n3061);
and (n6014,n3061,n6015);
or (n6015,n6016,n2971);
or (n6016,n2997,n2983);
and (n6017,n908,n6018);
or (n6018,n940,n942);
and (n6019,n3058,n6020);
or (n6020,n6021,n6131,n6791);
and (n6021,n6022,n6115);
or (n6022,1'b0,n6023,n6026,n6029,n6034);
and (n6023,n6024,n22);
wire s0n6024,s1n6024,notn6024;
or (n6024,s0n6024,s1n6024);
not(notn6024,n13);
and (s0n6024,notn6024,1'b0);
and (s1n6024,n13,n6025);
and (n6026,n6027,n904);
wire s0n6027,s1n6027,notn6027;
or (n6027,s0n6027,s1n6027);
not(notn6027,n896);
and (s0n6027,notn6027,1'b0);
and (s1n6027,n896,n6028);
and (n6029,n6030,n2971);
wire s0n6030,s1n6030,notn6030;
or (n6030,s0n6030,s1n6030);
not(notn6030,n2966);
and (s0n6030,notn6030,n6031);
and (s1n6030,n2966,1'b0);
wire s0n6031,s1n6031,notn6031;
or (n6031,s0n6031,s1n6031);
not(notn6031,n2961);
and (s0n6031,notn6031,n6032);
and (s1n6031,n2961,1'b1);
wire s0n6032,s1n6032,notn6032;
or (n6032,s0n6032,s1n6032);
not(notn6032,n2948);
and (s0n6032,notn6032,1'b0);
and (s1n6032,n2948,n6033);
xor (n6033,n2926,n2928);
or (n6034,1'b0,n6035,n6055,n6075,n6095);
and (n6035,n6036,n981);
or (n6036,1'b0,n6037,n6043,n6049);
and (n6037,n6038,n2983);
or (n6038,1'b0,n6039,n6040,n6041,n6042);
and (n6039,n1085,n903);
and (n6040,n1089,n949);
and (n6041,n1093,n901);
and (n6042,n1097,n960);
and (n6043,n6044,n942);
or (n6044,1'b0,n6045,n6046,n6047,n6048);
and (n6045,n1157,n903);
and (n6046,n1084,n949);
and (n6047,n1088,n901);
and (n6048,n1092,n960);
and (n6049,n6050,n2996);
or (n6050,1'b0,n6051,n6052,n6053,n6054);
and (n6051,n1084,n903);
and (n6052,n1088,n949);
and (n6053,n1092,n901);
and (n6054,n1096,n960);
and (n6055,n6056,n1002);
or (n6056,1'b0,n6057,n6063,n6069);
and (n6057,n6058,n2983);
or (n6058,1'b0,n6059,n6060,n6061,n6062);
and (n6059,n1103,n903);
and (n6060,n1107,n949);
and (n6061,n1111,n901);
and (n6062,n1115,n960);
and (n6063,n6064,n942);
or (n6064,1'b0,n6065,n6066,n6067,n6068);
and (n6065,n1096,n903);
and (n6066,n1102,n949);
and (n6067,n1106,n901);
and (n6068,n1110,n960);
and (n6069,n6070,n2996);
or (n6070,1'b0,n6071,n6072,n6073,n6074);
and (n6071,n1102,n903);
and (n6072,n1106,n949);
and (n6073,n1110,n901);
and (n6074,n1114,n960);
and (n6075,n6076,n1022);
or (n6076,1'b0,n6077,n6083,n6089);
and (n6077,n6078,n2983);
or (n6078,1'b0,n6079,n6080,n6081,n6082);
and (n6079,n1121,n903);
and (n6080,n1125,n949);
and (n6081,n1129,n901);
and (n6082,n1133,n960);
and (n6083,n6084,n942);
or (n6084,1'b0,n6085,n6086,n6087,n6088);
and (n6085,n1172,n903);
and (n6086,n1120,n949);
and (n6087,n1124,n901);
and (n6088,n1128,n960);
and (n6089,n6090,n2996);
or (n6090,1'b0,n6091,n6092,n6093,n6094);
and (n6091,n1120,n903);
and (n6092,n1124,n949);
and (n6093,n1128,n901);
and (n6094,n1132,n960);
and (n6095,n6096,n1042);
or (n6096,1'b0,n6097,n6103,n6109);
and (n6097,n6098,n2983);
or (n6098,1'b0,n6099,n6100,n6101,n6102);
and (n6099,n1139,n903);
and (n6100,n1143,n949);
and (n6101,n1147,n901);
and (n6102,n1151,n960);
and (n6103,n6104,n942);
or (n6104,1'b0,n6105,n6106,n6107,n6108);
and (n6105,n1132,n903);
and (n6106,n1138,n949);
and (n6107,n1142,n901);
and (n6108,n1146,n960);
and (n6109,n6110,n2996);
or (n6110,1'b0,n6111,n6112,n6113,n6114);
and (n6111,n1138,n903);
and (n6112,n1142,n949);
and (n6113,n1146,n901);
and (n6114,n1150,n960);
or (n6115,1'b0,n6116,n6127,n6129,n6130);
and (n6116,n6117,n22);
wire s0n6117,s1n6117,notn6117;
or (n6117,s0n6117,s1n6117);
not(notn6117,n13);
and (s0n6117,notn6117,1'b0);
and (s1n6117,n13,n6118);
wire s0n6118,s1n6118,notn6118;
or (n6118,s0n6118,s1n6118);
not(notn6118,n6001);
and (s0n6118,notn6118,n6119);
and (s1n6118,n6001,1'b0);
wire s0n6119,s1n6119,notn6119;
or (n6119,s0n6119,s1n6119);
not(notn6119,n5986);
and (s0n6119,notn6119,n6120);
and (s1n6119,n5986,1'b1);
wire s0n6120,s1n6120,notn6120;
or (n6120,s0n6120,s1n6120);
not(notn6120,n3074);
and (s0n6120,notn6120,n6121);
and (s1n6120,n3074,n6124);
wire s0n6121,s1n6121,notn6121;
or (n6121,s0n6121,s1n6121);
not(notn6121,n3074);
and (s0n6121,notn6121,n6122);
and (s1n6121,n3074,n6123);
xor (n6122,n5750,n5752);
xor (n6123,n5750,n5774);
wire s0n6124,s1n6124,notn6124;
or (n6124,s0n6124,s1n6124);
not(notn6124,n3074);
and (s0n6124,notn6124,n6125);
and (s1n6124,n3074,n6126);
xor (n6125,n5968,n5970);
xor (n6126,n5968,n5982);
and (n6127,n6128,n904);
wire s0n6128,s1n6128,notn6128;
or (n6128,s0n6128,s1n6128);
not(notn6128,n896);
and (s0n6128,notn6128,1'b0);
and (s1n6128,n896,n6118);
and (n6129,n6118,n6015);
and (n6130,n6030,n6018);
and (n6131,n6115,n6132);
or (n6132,n6133,n6243,n6790);
and (n6133,n6134,n6227);
or (n6134,1'b0,n6135,n6138,n6141,n6146);
and (n6135,n6136,n22);
wire s0n6136,s1n6136,notn6136;
or (n6136,s0n6136,s1n6136);
not(notn6136,n13);
and (s0n6136,notn6136,1'b0);
and (s1n6136,n13,n6137);
and (n6138,n6139,n904);
wire s0n6139,s1n6139,notn6139;
or (n6139,s0n6139,s1n6139);
not(notn6139,n896);
and (s0n6139,notn6139,1'b0);
and (s1n6139,n896,n6140);
and (n6141,n6142,n2971);
wire s0n6142,s1n6142,notn6142;
or (n6142,s0n6142,s1n6142);
not(notn6142,n2966);
and (s0n6142,notn6142,n6143);
and (s1n6142,n2966,1'b0);
wire s0n6143,s1n6143,notn6143;
or (n6143,s0n6143,s1n6143);
not(notn6143,n2961);
and (s0n6143,notn6143,n6144);
and (s1n6143,n2961,1'b1);
wire s0n6144,s1n6144,notn6144;
or (n6144,s0n6144,s1n6144);
not(notn6144,n2948);
and (s0n6144,notn6144,1'b0);
and (s1n6144,n2948,n6145);
xor (n6145,n2929,n2931);
or (n6146,1'b0,n6147,n6167,n6187,n6207);
and (n6147,n6148,n981);
or (n6148,1'b0,n6149,n6155,n6161);
and (n6149,n6150,n2983);
or (n6150,1'b0,n6151,n6152,n6153,n6154);
and (n6151,n1192,n903);
and (n6152,n1196,n949);
and (n6153,n1200,n901);
and (n6154,n1204,n960);
and (n6155,n6156,n942);
or (n6156,1'b0,n6157,n6158,n6159,n6160);
and (n6157,n1264,n903);
and (n6158,n1191,n949);
and (n6159,n1195,n901);
and (n6160,n1199,n960);
and (n6161,n6162,n2996);
or (n6162,1'b0,n6163,n6164,n6165,n6166);
and (n6163,n1191,n903);
and (n6164,n1195,n949);
and (n6165,n1199,n901);
and (n6166,n1203,n960);
and (n6167,n6168,n1002);
or (n6168,1'b0,n6169,n6175,n6181);
and (n6169,n6170,n2983);
or (n6170,1'b0,n6171,n6172,n6173,n6174);
and (n6171,n1210,n903);
and (n6172,n1214,n949);
and (n6173,n1218,n901);
and (n6174,n1222,n960);
and (n6175,n6176,n942);
or (n6176,1'b0,n6177,n6178,n6179,n6180);
and (n6177,n1203,n903);
and (n6178,n1209,n949);
and (n6179,n1213,n901);
and (n6180,n1217,n960);
and (n6181,n6182,n2996);
or (n6182,1'b0,n6183,n6184,n6185,n6186);
and (n6183,n1209,n903);
and (n6184,n1213,n949);
and (n6185,n1217,n901);
and (n6186,n1221,n960);
and (n6187,n6188,n1022);
or (n6188,1'b0,n6189,n6195,n6201);
and (n6189,n6190,n2983);
or (n6190,1'b0,n6191,n6192,n6193,n6194);
and (n6191,n1228,n903);
and (n6192,n1232,n949);
and (n6193,n1236,n901);
and (n6194,n1240,n960);
and (n6195,n6196,n942);
or (n6196,1'b0,n6197,n6198,n6199,n6200);
and (n6197,n1279,n903);
and (n6198,n1227,n949);
and (n6199,n1231,n901);
and (n6200,n1235,n960);
and (n6201,n6202,n2996);
or (n6202,1'b0,n6203,n6204,n6205,n6206);
and (n6203,n1227,n903);
and (n6204,n1231,n949);
and (n6205,n1235,n901);
and (n6206,n1239,n960);
and (n6207,n6208,n1042);
or (n6208,1'b0,n6209,n6215,n6221);
and (n6209,n6210,n2983);
or (n6210,1'b0,n6211,n6212,n6213,n6214);
and (n6211,n1246,n903);
and (n6212,n1250,n949);
and (n6213,n1254,n901);
and (n6214,n1258,n960);
and (n6215,n6216,n942);
or (n6216,1'b0,n6217,n6218,n6219,n6220);
and (n6217,n1239,n903);
and (n6218,n1245,n949);
and (n6219,n1249,n901);
and (n6220,n1253,n960);
and (n6221,n6222,n2996);
or (n6222,1'b0,n6223,n6224,n6225,n6226);
and (n6223,n1245,n903);
and (n6224,n1249,n949);
and (n6225,n1253,n901);
and (n6226,n1257,n960);
or (n6227,1'b0,n6228,n6239,n6241,n6242);
and (n6228,n6229,n22);
wire s0n6229,s1n6229,notn6229;
or (n6229,s0n6229,s1n6229);
not(notn6229,n13);
and (s0n6229,notn6229,1'b0);
and (s1n6229,n13,n6230);
wire s0n6230,s1n6230,notn6230;
or (n6230,s0n6230,s1n6230);
not(notn6230,n6001);
and (s0n6230,notn6230,n6231);
and (s1n6230,n6001,1'b0);
wire s0n6231,s1n6231,notn6231;
or (n6231,s0n6231,s1n6231);
not(notn6231,n5986);
and (s0n6231,notn6231,n6232);
and (s1n6231,n5986,1'b1);
wire s0n6232,s1n6232,notn6232;
or (n6232,s0n6232,s1n6232);
not(notn6232,n3074);
and (s0n6232,notn6232,n6233);
and (s1n6232,n3074,n6236);
wire s0n6233,s1n6233,notn6233;
or (n6233,s0n6233,s1n6233);
not(notn6233,n3074);
and (s0n6233,notn6233,n6234);
and (s1n6233,n3074,n6235);
xor (n6234,n5753,n5755);
xor (n6235,n5753,n5756);
wire s0n6236,s1n6236,notn6236;
or (n6236,s0n6236,s1n6236);
not(notn6236,n3074);
and (s0n6236,notn6236,n6237);
and (s1n6236,n3074,n6238);
xor (n6237,n5971,n5973);
xor (n6238,n5971,n5983);
and (n6239,n6240,n904);
wire s0n6240,s1n6240,notn6240;
or (n6240,s0n6240,s1n6240);
not(notn6240,n896);
and (s0n6240,notn6240,1'b0);
and (s1n6240,n896,n6230);
and (n6241,n6230,n6015);
and (n6242,n6142,n6018);
and (n6243,n6227,n6244);
or (n6244,n6245,n6355,n6789);
and (n6245,n6246,n6339);
or (n6246,1'b0,n6247,n6250,n6253,n6258);
and (n6247,n6248,n22);
wire s0n6248,s1n6248,notn6248;
or (n6248,s0n6248,s1n6248);
not(notn6248,n13);
and (s0n6248,notn6248,1'b0);
and (s1n6248,n13,n6249);
and (n6250,n6251,n904);
wire s0n6251,s1n6251,notn6251;
or (n6251,s0n6251,s1n6251);
not(notn6251,n896);
and (s0n6251,notn6251,1'b0);
and (s1n6251,n896,n6252);
and (n6253,n6254,n2971);
wire s0n6254,s1n6254,notn6254;
or (n6254,s0n6254,s1n6254);
not(notn6254,n2966);
and (s0n6254,notn6254,n6255);
and (s1n6254,n2966,1'b0);
wire s0n6255,s1n6255,notn6255;
or (n6255,s0n6255,s1n6255);
not(notn6255,n2961);
and (s0n6255,notn6255,n6256);
and (s1n6255,n2961,1'b1);
wire s0n6256,s1n6256,notn6256;
or (n6256,s0n6256,s1n6256);
not(notn6256,n2948);
and (s0n6256,notn6256,1'b0);
and (s1n6256,n2948,n6257);
xor (n6257,n2932,n2934);
or (n6258,1'b0,n6259,n6279,n6299,n6319);
and (n6259,n6260,n981);
or (n6260,1'b0,n6261,n6267,n6273);
and (n6261,n6262,n2983);
or (n6262,1'b0,n6263,n6264,n6265,n6266);
and (n6263,n1299,n903);
and (n6264,n1303,n949);
and (n6265,n1307,n901);
and (n6266,n1311,n960);
and (n6267,n6268,n942);
or (n6268,1'b0,n6269,n6270,n6271,n6272);
and (n6269,n1371,n903);
and (n6270,n1298,n949);
and (n6271,n1302,n901);
and (n6272,n1306,n960);
and (n6273,n6274,n2996);
or (n6274,1'b0,n6275,n6276,n6277,n6278);
and (n6275,n1298,n903);
and (n6276,n1302,n949);
and (n6277,n1306,n901);
and (n6278,n1310,n960);
and (n6279,n6280,n1002);
or (n6280,1'b0,n6281,n6287,n6293);
and (n6281,n6282,n2983);
or (n6282,1'b0,n6283,n6284,n6285,n6286);
and (n6283,n1317,n903);
and (n6284,n1321,n949);
and (n6285,n1325,n901);
and (n6286,n1329,n960);
and (n6287,n6288,n942);
or (n6288,1'b0,n6289,n6290,n6291,n6292);
and (n6289,n1310,n903);
and (n6290,n1316,n949);
and (n6291,n1320,n901);
and (n6292,n1324,n960);
and (n6293,n6294,n2996);
or (n6294,1'b0,n6295,n6296,n6297,n6298);
and (n6295,n1316,n903);
and (n6296,n1320,n949);
and (n6297,n1324,n901);
and (n6298,n1328,n960);
and (n6299,n6300,n1022);
or (n6300,1'b0,n6301,n6307,n6313);
and (n6301,n6302,n2983);
or (n6302,1'b0,n6303,n6304,n6305,n6306);
and (n6303,n1335,n903);
and (n6304,n1339,n949);
and (n6305,n1343,n901);
and (n6306,n1347,n960);
and (n6307,n6308,n942);
or (n6308,1'b0,n6309,n6310,n6311,n6312);
and (n6309,n1386,n903);
and (n6310,n1334,n949);
and (n6311,n1338,n901);
and (n6312,n1342,n960);
and (n6313,n6314,n2996);
or (n6314,1'b0,n6315,n6316,n6317,n6318);
and (n6315,n1334,n903);
and (n6316,n1338,n949);
and (n6317,n1342,n901);
and (n6318,n1346,n960);
and (n6319,n6320,n1042);
or (n6320,1'b0,n6321,n6327,n6333);
and (n6321,n6322,n2983);
or (n6322,1'b0,n6323,n6324,n6325,n6326);
and (n6323,n1353,n903);
and (n6324,n1357,n949);
and (n6325,n1361,n901);
and (n6326,n1365,n960);
and (n6327,n6328,n942);
or (n6328,1'b0,n6329,n6330,n6331,n6332);
and (n6329,n1346,n903);
and (n6330,n1352,n949);
and (n6331,n1356,n901);
and (n6332,n1360,n960);
and (n6333,n6334,n2996);
or (n6334,1'b0,n6335,n6336,n6337,n6338);
and (n6335,n1352,n903);
and (n6336,n1356,n949);
and (n6337,n1360,n901);
and (n6338,n1364,n960);
or (n6339,1'b0,n6340,n6351,n6353,n6354);
and (n6340,n6341,n22);
wire s0n6341,s1n6341,notn6341;
or (n6341,s0n6341,s1n6341);
not(notn6341,n13);
and (s0n6341,notn6341,1'b0);
and (s1n6341,n13,n6342);
wire s0n6342,s1n6342,notn6342;
or (n6342,s0n6342,s1n6342);
not(notn6342,n6001);
and (s0n6342,notn6342,n6343);
and (s1n6342,n6001,1'b0);
wire s0n6343,s1n6343,notn6343;
or (n6343,s0n6343,s1n6343);
not(notn6343,n5986);
and (s0n6343,notn6343,n6344);
and (s1n6343,n5986,1'b1);
wire s0n6344,s1n6344,notn6344;
or (n6344,s0n6344,s1n6344);
not(notn6344,n3074);
and (s0n6344,notn6344,n6345);
and (s1n6344,n3074,n6348);
wire s0n6345,s1n6345,notn6345;
or (n6345,s0n6345,s1n6345);
not(notn6345,n3074);
and (s0n6345,notn6345,n6346);
and (s1n6345,n3074,n6347);
xor (n6346,n5756,n5758);
not (n6347,n5756);
wire s0n6348,s1n6348,notn6348;
or (n6348,s0n6348,s1n6348);
not(notn6348,n3074);
and (s0n6348,notn6348,n6349);
and (s1n6348,n3074,n6350);
xor (n6349,n5974,n5976);
xor (n6350,n5974,n5984);
and (n6351,n6352,n904);
wire s0n6352,s1n6352,notn6352;
or (n6352,s0n6352,s1n6352);
not(notn6352,n896);
and (s0n6352,notn6352,1'b0);
and (s1n6352,n896,n6342);
and (n6353,n6342,n6015);
and (n6354,n6254,n6018);
and (n6355,n6339,n6356);
or (n6356,n6357,n6463,n6788);
and (n6357,n6358,n6451);
or (n6358,1'b0,n6359,n6362,n6365,n6370);
and (n6359,n6360,n22);
wire s0n6360,s1n6360,notn6360;
or (n6360,s0n6360,s1n6360);
not(notn6360,n13);
and (s0n6360,notn6360,1'b0);
and (s1n6360,n13,n6361);
and (n6362,n6363,n904);
wire s0n6363,s1n6363,notn6363;
or (n6363,s0n6363,s1n6363);
not(notn6363,n896);
and (s0n6363,notn6363,1'b0);
and (s1n6363,n896,n6364);
and (n6365,n6366,n2971);
wire s0n6366,s1n6366,notn6366;
or (n6366,s0n6366,s1n6366);
not(notn6366,n2966);
and (s0n6366,notn6366,n6367);
and (s1n6366,n2966,1'b0);
wire s0n6367,s1n6367,notn6367;
or (n6367,s0n6367,s1n6367);
not(notn6367,n2961);
and (s0n6367,notn6367,n6368);
and (s1n6367,n2961,1'b1);
wire s0n6368,s1n6368,notn6368;
or (n6368,s0n6368,s1n6368);
not(notn6368,n2948);
and (s0n6368,notn6368,1'b0);
and (s1n6368,n2948,n6369);
xor (n6369,n2935,n2937);
or (n6370,1'b0,n6371,n6391,n6411,n6431);
and (n6371,n6372,n981);
or (n6372,1'b0,n6373,n6379,n6385);
and (n6373,n6374,n2983);
or (n6374,1'b0,n6375,n6376,n6377,n6378);
and (n6375,n1406,n903);
and (n6376,n1410,n949);
and (n6377,n1414,n901);
and (n6378,n1418,n960);
and (n6379,n6380,n942);
or (n6380,1'b0,n6381,n6382,n6383,n6384);
and (n6381,n1478,n903);
and (n6382,n1405,n949);
and (n6383,n1409,n901);
and (n6384,n1413,n960);
and (n6385,n6386,n2996);
or (n6386,1'b0,n6387,n6388,n6389,n6390);
and (n6387,n1405,n903);
and (n6388,n1409,n949);
and (n6389,n1413,n901);
and (n6390,n1417,n960);
and (n6391,n6392,n1002);
or (n6392,1'b0,n6393,n6399,n6405);
and (n6393,n6394,n2983);
or (n6394,1'b0,n6395,n6396,n6397,n6398);
and (n6395,n1424,n903);
and (n6396,n1428,n949);
and (n6397,n1432,n901);
and (n6398,n1436,n960);
and (n6399,n6400,n942);
or (n6400,1'b0,n6401,n6402,n6403,n6404);
and (n6401,n1417,n903);
and (n6402,n1423,n949);
and (n6403,n1427,n901);
and (n6404,n1431,n960);
and (n6405,n6406,n2996);
or (n6406,1'b0,n6407,n6408,n6409,n6410);
and (n6407,n1423,n903);
and (n6408,n1427,n949);
and (n6409,n1431,n901);
and (n6410,n1435,n960);
and (n6411,n6412,n1022);
or (n6412,1'b0,n6413,n6419,n6425);
and (n6413,n6414,n2983);
or (n6414,1'b0,n6415,n6416,n6417,n6418);
and (n6415,n1442,n903);
and (n6416,n1446,n949);
and (n6417,n1450,n901);
and (n6418,n1454,n960);
and (n6419,n6420,n942);
or (n6420,1'b0,n6421,n6422,n6423,n6424);
and (n6421,n1493,n903);
and (n6422,n1441,n949);
and (n6423,n1445,n901);
and (n6424,n1449,n960);
and (n6425,n6426,n2996);
or (n6426,1'b0,n6427,n6428,n6429,n6430);
and (n6427,n1441,n903);
and (n6428,n1445,n949);
and (n6429,n1449,n901);
and (n6430,n1453,n960);
and (n6431,n6432,n1042);
or (n6432,1'b0,n6433,n6439,n6445);
and (n6433,n6434,n2983);
or (n6434,1'b0,n6435,n6436,n6437,n6438);
and (n6435,n1460,n903);
and (n6436,n1464,n949);
and (n6437,n1468,n901);
and (n6438,n1472,n960);
and (n6439,n6440,n942);
or (n6440,1'b0,n6441,n6442,n6443,n6444);
and (n6441,n1453,n903);
and (n6442,n1459,n949);
and (n6443,n1463,n901);
and (n6444,n1467,n960);
and (n6445,n6446,n2996);
or (n6446,1'b0,n6447,n6448,n6449,n6450);
and (n6447,n1459,n903);
and (n6448,n1463,n949);
and (n6449,n1467,n901);
and (n6450,n1471,n960);
or (n6451,1'b0,n6452,n6459,n6461,n6462);
and (n6452,n6453,n22);
wire s0n6453,s1n6453,notn6453;
or (n6453,s0n6453,s1n6453);
not(notn6453,n13);
and (s0n6453,notn6453,1'b0);
and (s1n6453,n13,n6454);
wire s0n6454,s1n6454,notn6454;
or (n6454,s0n6454,s1n6454);
not(notn6454,n6001);
and (s0n6454,notn6454,n6455);
and (s1n6454,n6001,1'b0);
wire s0n6455,s1n6455,notn6455;
or (n6455,s0n6455,s1n6455);
not(notn6455,n5986);
and (s0n6455,notn6455,n6456);
and (s1n6455,n5986,1'b1);
wire s0n6456,s1n6456,notn6456;
or (n6456,s0n6456,s1n6456);
not(notn6456,n3074);
and (s0n6456,notn6456,n6457);
and (s1n6456,n3074,n5987);
wire s0n6457,s1n6457,notn6457;
or (n6457,s0n6457,s1n6457);
not(notn6457,n3074);
and (s0n6457,notn6457,n6458);
and (s1n6457,n3074,n5759);
xor (n6458,n5759,n5761);
and (n6459,n6460,n904);
wire s0n6460,s1n6460,notn6460;
or (n6460,s0n6460,s1n6460);
not(notn6460,n896);
and (s0n6460,notn6460,1'b0);
and (s1n6460,n896,n6454);
and (n6461,n6454,n6015);
and (n6462,n6366,n6018);
and (n6463,n6451,n6464);
or (n6464,n6465,n6571,n6787);
and (n6465,n6466,n6559);
or (n6466,1'b0,n6467,n6470,n6473,n6478);
and (n6467,n6468,n22);
wire s0n6468,s1n6468,notn6468;
or (n6468,s0n6468,s1n6468);
not(notn6468,n13);
and (s0n6468,notn6468,1'b0);
and (s1n6468,n13,n6469);
and (n6470,n6471,n904);
wire s0n6471,s1n6471,notn6471;
or (n6471,s0n6471,s1n6471);
not(notn6471,n896);
and (s0n6471,notn6471,1'b0);
and (s1n6471,n896,n6472);
and (n6473,n6474,n2971);
wire s0n6474,s1n6474,notn6474;
or (n6474,s0n6474,s1n6474);
not(notn6474,n2966);
and (s0n6474,notn6474,n6475);
and (s1n6474,n2966,1'b0);
wire s0n6475,s1n6475,notn6475;
or (n6475,s0n6475,s1n6475);
not(notn6475,n2961);
and (s0n6475,notn6475,n6476);
and (s1n6475,n2961,1'b1);
wire s0n6476,s1n6476,notn6476;
or (n6476,s0n6476,s1n6476);
not(notn6476,n2948);
and (s0n6476,notn6476,1'b0);
and (s1n6476,n2948,n6477);
xor (n6477,n2938,n2940);
or (n6478,1'b0,n6479,n6499,n6519,n6539);
and (n6479,n6480,n981);
or (n6480,1'b0,n6481,n6487,n6493);
and (n6481,n6482,n2983);
or (n6482,1'b0,n6483,n6484,n6485,n6486);
and (n6483,n1513,n903);
and (n6484,n1517,n949);
and (n6485,n1521,n901);
and (n6486,n1525,n960);
and (n6487,n6488,n942);
or (n6488,1'b0,n6489,n6490,n6491,n6492);
and (n6489,n1585,n903);
and (n6490,n1512,n949);
and (n6491,n1516,n901);
and (n6492,n1520,n960);
and (n6493,n6494,n2996);
or (n6494,1'b0,n6495,n6496,n6497,n6498);
and (n6495,n1512,n903);
and (n6496,n1516,n949);
and (n6497,n1520,n901);
and (n6498,n1524,n960);
and (n6499,n6500,n1002);
or (n6500,1'b0,n6501,n6507,n6513);
and (n6501,n6502,n2983);
or (n6502,1'b0,n6503,n6504,n6505,n6506);
and (n6503,n1531,n903);
and (n6504,n1535,n949);
and (n6505,n1539,n901);
and (n6506,n1543,n960);
and (n6507,n6508,n942);
or (n6508,1'b0,n6509,n6510,n6511,n6512);
and (n6509,n1524,n903);
and (n6510,n1530,n949);
and (n6511,n1534,n901);
and (n6512,n1538,n960);
and (n6513,n6514,n2996);
or (n6514,1'b0,n6515,n6516,n6517,n6518);
and (n6515,n1530,n903);
and (n6516,n1534,n949);
and (n6517,n1538,n901);
and (n6518,n1542,n960);
and (n6519,n6520,n1022);
or (n6520,1'b0,n6521,n6527,n6533);
and (n6521,n6522,n2983);
or (n6522,1'b0,n6523,n6524,n6525,n6526);
and (n6523,n1549,n903);
and (n6524,n1553,n949);
and (n6525,n1557,n901);
and (n6526,n1561,n960);
and (n6527,n6528,n942);
or (n6528,1'b0,n6529,n6530,n6531,n6532);
and (n6529,n1600,n903);
and (n6530,n1548,n949);
and (n6531,n1552,n901);
and (n6532,n1556,n960);
and (n6533,n6534,n2996);
or (n6534,1'b0,n6535,n6536,n6537,n6538);
and (n6535,n1548,n903);
and (n6536,n1552,n949);
and (n6537,n1556,n901);
and (n6538,n1560,n960);
and (n6539,n6540,n1042);
or (n6540,1'b0,n6541,n6547,n6553);
and (n6541,n6542,n2983);
or (n6542,1'b0,n6543,n6544,n6545,n6546);
and (n6543,n1567,n903);
and (n6544,n1571,n949);
and (n6545,n1575,n901);
and (n6546,n1579,n960);
and (n6547,n6548,n942);
or (n6548,1'b0,n6549,n6550,n6551,n6552);
and (n6549,n1560,n903);
and (n6550,n1566,n949);
and (n6551,n1570,n901);
and (n6552,n1574,n960);
and (n6553,n6554,n2996);
or (n6554,1'b0,n6555,n6556,n6557,n6558);
and (n6555,n1566,n903);
and (n6556,n1570,n949);
and (n6557,n1574,n901);
and (n6558,n1578,n960);
or (n6559,1'b0,n6560,n6567,n6569,n6570);
and (n6560,n6561,n22);
wire s0n6561,s1n6561,notn6561;
or (n6561,s0n6561,s1n6561);
not(notn6561,n13);
and (s0n6561,notn6561,1'b0);
and (s1n6561,n13,n6562);
wire s0n6562,s1n6562,notn6562;
or (n6562,s0n6562,s1n6562);
not(notn6562,n6001);
and (s0n6562,notn6562,n6563);
and (s1n6562,n6001,1'b0);
wire s0n6563,s1n6563,notn6563;
or (n6563,s0n6563,s1n6563);
not(notn6563,n5986);
and (s0n6563,notn6563,n6564);
and (s1n6563,n5986,1'b1);
wire s0n6564,s1n6564,notn6564;
or (n6564,s0n6564,s1n6564);
not(notn6564,n3074);
and (s0n6564,notn6564,n6565);
and (s1n6564,n3074,n3064);
wire s0n6565,s1n6565,notn6565;
or (n6565,s0n6565,s1n6565);
not(notn6565,n3074);
and (s0n6565,notn6565,n6566);
and (s1n6565,n3074,n5762);
xor (n6566,n5762,n5764);
and (n6567,n6568,n904);
wire s0n6568,s1n6568,notn6568;
or (n6568,s0n6568,s1n6568);
not(notn6568,n896);
and (s0n6568,notn6568,1'b0);
and (s1n6568,n896,n6562);
and (n6569,n6562,n6015);
and (n6570,n6474,n6018);
and (n6571,n6559,n6572);
or (n6572,n6573,n6679,n6786);
and (n6573,n6574,n6667);
or (n6574,1'b0,n6575,n6578,n6581,n6586);
and (n6575,n6576,n22);
wire s0n6576,s1n6576,notn6576;
or (n6576,s0n6576,s1n6576);
not(notn6576,n13);
and (s0n6576,notn6576,1'b0);
and (s1n6576,n13,n6577);
and (n6578,n6579,n904);
wire s0n6579,s1n6579,notn6579;
or (n6579,s0n6579,s1n6579);
not(notn6579,n896);
and (s0n6579,notn6579,1'b0);
and (s1n6579,n896,n6580);
and (n6581,n6582,n2971);
wire s0n6582,s1n6582,notn6582;
or (n6582,s0n6582,s1n6582);
not(notn6582,n2966);
and (s0n6582,notn6582,n6583);
and (s1n6582,n2966,1'b0);
wire s0n6583,s1n6583,notn6583;
or (n6583,s0n6583,s1n6583);
not(notn6583,n2961);
and (s0n6583,notn6583,n6584);
and (s1n6583,n2961,1'b1);
wire s0n6584,s1n6584,notn6584;
or (n6584,s0n6584,s1n6584);
not(notn6584,n2948);
and (s0n6584,notn6584,1'b0);
and (s1n6584,n2948,n6585);
xor (n6585,n2941,n2943);
or (n6586,1'b0,n6587,n6607,n6627,n6647);
and (n6587,n6588,n981);
or (n6588,1'b0,n6589,n6595,n6601);
and (n6589,n6590,n2983);
or (n6590,1'b0,n6591,n6592,n6593,n6594);
and (n6591,n1620,n903);
and (n6592,n1624,n949);
and (n6593,n1628,n901);
and (n6594,n1632,n960);
and (n6595,n6596,n942);
or (n6596,1'b0,n6597,n6598,n6599,n6600);
and (n6597,n1692,n903);
and (n6598,n1619,n949);
and (n6599,n1623,n901);
and (n6600,n1627,n960);
and (n6601,n6602,n2996);
or (n6602,1'b0,n6603,n6604,n6605,n6606);
and (n6603,n1619,n903);
and (n6604,n1623,n949);
and (n6605,n1627,n901);
and (n6606,n1631,n960);
and (n6607,n6608,n1002);
or (n6608,1'b0,n6609,n6615,n6621);
and (n6609,n6610,n2983);
or (n6610,1'b0,n6611,n6612,n6613,n6614);
and (n6611,n1638,n903);
and (n6612,n1642,n949);
and (n6613,n1646,n901);
and (n6614,n1650,n960);
and (n6615,n6616,n942);
or (n6616,1'b0,n6617,n6618,n6619,n6620);
and (n6617,n1631,n903);
and (n6618,n1637,n949);
and (n6619,n1641,n901);
and (n6620,n1645,n960);
and (n6621,n6622,n2996);
or (n6622,1'b0,n6623,n6624,n6625,n6626);
and (n6623,n1637,n903);
and (n6624,n1641,n949);
and (n6625,n1645,n901);
and (n6626,n1649,n960);
and (n6627,n6628,n1022);
or (n6628,1'b0,n6629,n6635,n6641);
and (n6629,n6630,n2983);
or (n6630,1'b0,n6631,n6632,n6633,n6634);
and (n6631,n1656,n903);
and (n6632,n1660,n949);
and (n6633,n1664,n901);
and (n6634,n1668,n960);
and (n6635,n6636,n942);
or (n6636,1'b0,n6637,n6638,n6639,n6640);
and (n6637,n1707,n903);
and (n6638,n1655,n949);
and (n6639,n1659,n901);
and (n6640,n1663,n960);
and (n6641,n6642,n2996);
or (n6642,1'b0,n6643,n6644,n6645,n6646);
and (n6643,n1655,n903);
and (n6644,n1659,n949);
and (n6645,n1663,n901);
and (n6646,n1667,n960);
and (n6647,n6648,n1042);
or (n6648,1'b0,n6649,n6655,n6661);
and (n6649,n6650,n2983);
or (n6650,1'b0,n6651,n6652,n6653,n6654);
and (n6651,n1674,n903);
and (n6652,n1678,n949);
and (n6653,n1682,n901);
and (n6654,n1686,n960);
and (n6655,n6656,n942);
or (n6656,1'b0,n6657,n6658,n6659,n6660);
and (n6657,n1667,n903);
and (n6658,n1673,n949);
and (n6659,n1677,n901);
and (n6660,n1681,n960);
and (n6661,n6662,n2996);
or (n6662,1'b0,n6663,n6664,n6665,n6666);
and (n6663,n1673,n903);
and (n6664,n1677,n949);
and (n6665,n1681,n901);
and (n6666,n1685,n960);
or (n6667,1'b0,n6668,n6675,n6677,n6678);
and (n6668,n6669,n22);
wire s0n6669,s1n6669,notn6669;
or (n6669,s0n6669,s1n6669);
not(notn6669,n13);
and (s0n6669,notn6669,1'b0);
and (s1n6669,n13,n6670);
wire s0n6670,s1n6670,notn6670;
or (n6670,s0n6670,s1n6670);
not(notn6670,n6001);
and (s0n6670,notn6670,n6671);
and (s1n6670,n6001,1'b0);
wire s0n6671,s1n6671,notn6671;
or (n6671,s0n6671,s1n6671);
not(notn6671,n5986);
and (s0n6671,notn6671,n6672);
and (s1n6671,n5986,1'b1);
wire s0n6672,s1n6672,notn6672;
or (n6672,s0n6672,s1n6672);
not(notn6672,n3074);
and (s0n6672,notn6672,n6673);
and (s1n6672,n3074,n6121);
wire s0n6673,s1n6673,notn6673;
or (n6673,s0n6673,s1n6673);
not(notn6673,n3074);
and (s0n6673,notn6673,n6674);
and (s1n6673,n3074,n5765);
xor (n6674,n5765,n5767);
and (n6675,n6676,n904);
wire s0n6676,s1n6676,notn6676;
or (n6676,s0n6676,s1n6676);
not(notn6676,n896);
and (s0n6676,notn6676,1'b0);
and (s1n6676,n896,n6670);
and (n6677,n6670,n6015);
and (n6678,n6582,n6018);
and (n6679,n6667,n6680);
and (n6680,n6681,n6774);
or (n6681,1'b0,n6682,n6685,n6688,n6693);
and (n6682,n6683,n22);
wire s0n6683,s1n6683,notn6683;
or (n6683,s0n6683,s1n6683);
not(notn6683,n13);
and (s0n6683,notn6683,1'b0);
and (s1n6683,n13,n6684);
and (n6685,n6686,n904);
wire s0n6686,s1n6686,notn6686;
or (n6686,s0n6686,s1n6686);
not(notn6686,n896);
and (s0n6686,notn6686,1'b0);
and (s1n6686,n896,n6687);
and (n6688,n6689,n2971);
wire s0n6689,s1n6689,notn6689;
or (n6689,s0n6689,s1n6689);
not(notn6689,n2966);
and (s0n6689,notn6689,n6690);
and (s1n6689,n2966,1'b0);
wire s0n6690,s1n6690,notn6690;
or (n6690,s0n6690,s1n6690);
not(notn6690,n2961);
and (s0n6690,notn6690,n6691);
and (s1n6690,n2961,1'b1);
wire s0n6691,s1n6691,notn6691;
or (n6691,s0n6691,s1n6691);
not(notn6691,n2948);
and (s0n6691,notn6691,1'b0);
and (s1n6691,n2948,n6692);
xor (n6692,n2944,n2946);
or (n6693,1'b0,n6694,n6714,n6734,n6754);
and (n6694,n6695,n981);
or (n6695,1'b0,n6696,n6702,n6708);
and (n6696,n6697,n2983);
or (n6697,1'b0,n6698,n6699,n6700,n6701);
and (n6698,n1726,n903);
and (n6699,n1730,n949);
and (n6700,n1734,n901);
and (n6701,n1738,n960);
and (n6702,n6703,n942);
or (n6703,1'b0,n6704,n6705,n6706,n6707);
and (n6704,n1798,n903);
and (n6705,n1725,n949);
and (n6706,n1729,n901);
and (n6707,n1733,n960);
and (n6708,n6709,n2996);
or (n6709,1'b0,n6710,n6711,n6712,n6713);
and (n6710,n1725,n903);
and (n6711,n1729,n949);
and (n6712,n1733,n901);
and (n6713,n1737,n960);
and (n6714,n6715,n1002);
or (n6715,1'b0,n6716,n6722,n6728);
and (n6716,n6717,n2983);
or (n6717,1'b0,n6718,n6719,n6720,n6721);
and (n6718,n1744,n903);
and (n6719,n1748,n949);
and (n6720,n1752,n901);
and (n6721,n1756,n960);
and (n6722,n6723,n942);
or (n6723,1'b0,n6724,n6725,n6726,n6727);
and (n6724,n1737,n903);
and (n6725,n1743,n949);
and (n6726,n1747,n901);
and (n6727,n1751,n960);
and (n6728,n6729,n2996);
or (n6729,1'b0,n6730,n6731,n6732,n6733);
and (n6730,n1743,n903);
and (n6731,n1747,n949);
and (n6732,n1751,n901);
and (n6733,n1755,n960);
and (n6734,n6735,n1022);
or (n6735,1'b0,n6736,n6742,n6748);
and (n6736,n6737,n2983);
or (n6737,1'b0,n6738,n6739,n6740,n6741);
and (n6738,n1762,n903);
and (n6739,n1766,n949);
and (n6740,n1770,n901);
and (n6741,n1774,n960);
and (n6742,n6743,n942);
or (n6743,1'b0,n6744,n6745,n6746,n6747);
and (n6744,n1813,n903);
and (n6745,n1761,n949);
and (n6746,n1765,n901);
and (n6747,n1769,n960);
and (n6748,n6749,n2996);
or (n6749,1'b0,n6750,n6751,n6752,n6753);
and (n6750,n1761,n903);
and (n6751,n1765,n949);
and (n6752,n1769,n901);
and (n6753,n1773,n960);
and (n6754,n6755,n1042);
or (n6755,1'b0,n6756,n6762,n6768);
and (n6756,n6757,n2983);
or (n6757,1'b0,n6758,n6759,n6760,n6761);
and (n6758,n1780,n903);
and (n6759,n1784,n949);
and (n6760,n1788,n901);
and (n6761,n1792,n960);
and (n6762,n6763,n942);
or (n6763,1'b0,n6764,n6765,n6766,n6767);
and (n6764,n1773,n903);
and (n6765,n1779,n949);
and (n6766,n1783,n901);
and (n6767,n1787,n960);
and (n6768,n6769,n2996);
or (n6769,1'b0,n6770,n6771,n6772,n6773);
and (n6770,n1779,n903);
and (n6771,n1783,n949);
and (n6772,n1787,n901);
and (n6773,n1791,n960);
or (n6774,1'b0,n6775,n6782,n6784,n6785);
and (n6775,n6776,n22);
wire s0n6776,s1n6776,notn6776;
or (n6776,s0n6776,s1n6776);
not(notn6776,n13);
and (s0n6776,notn6776,1'b0);
and (s1n6776,n13,n6777);
wire s0n6777,s1n6777,notn6777;
or (n6777,s0n6777,s1n6777);
not(notn6777,n6001);
and (s0n6777,notn6777,n6778);
and (s1n6777,n6001,1'b0);
wire s0n6778,s1n6778,notn6778;
or (n6778,s0n6778,s1n6778);
not(notn6778,n5986);
and (s0n6778,notn6778,n6779);
and (s1n6778,n5986,1'b1);
wire s0n6779,s1n6779,notn6779;
or (n6779,s0n6779,s1n6779);
not(notn6779,n3074);
and (s0n6779,notn6779,n6780);
and (s1n6779,n3074,n6233);
wire s0n6780,s1n6780,notn6780;
or (n6780,s0n6780,s1n6780);
not(notn6780,n3074);
and (s0n6780,notn6780,n6781);
and (s1n6780,n3074,n5768);
xor (n6781,n5768,n5770);
and (n6782,n6783,n904);
wire s0n6783,s1n6783,notn6783;
or (n6783,s0n6783,s1n6783);
not(notn6783,n896);
and (s0n6783,notn6783,1'b0);
and (s1n6783,n896,n6777);
and (n6784,n6777,n6015);
and (n6785,n6689,n6018);
and (n6786,n6574,n6680);
and (n6787,n6466,n6572);
and (n6788,n6358,n6464);
and (n6789,n6246,n6356);
and (n6790,n6134,n6244);
and (n6791,n6022,n6132);
and (n6792,n9,n6020);
and (n6793,n6794,n6796);
xor (n6794,n6795,n6020);
xor (n6795,n9,n3058);
and (n6796,n6797,n6799);
xor (n6797,n6798,n6132);
xor (n6798,n6022,n6115);
and (n6799,n6800,n6802);
xor (n6800,n6801,n6244);
xor (n6801,n6134,n6227);
and (n6802,n6803,n6805);
xor (n6803,n6804,n6356);
xor (n6804,n6246,n6339);
and (n6805,n6806,n6808);
xor (n6806,n6807,n6464);
xor (n6807,n6358,n6451);
and (n6808,n6809,n6811);
xor (n6809,n6810,n6572);
xor (n6810,n6466,n6559);
and (n6811,n6812,n6814);
xor (n6812,n6813,n6680);
xor (n6813,n6574,n6667);
xor (n6814,n6681,n6774);
and (n6815,n6816,n6817);
wire s0n6816,s1n6816,notn6816;
or (n6816,s0n6816,s1n6816);
not(notn6816,n3077);
and (s0n6816,notn6816,1'b0);
and (s1n6816,n3077,n6);
or (n6817,n6818,n891);
or (n6818,n6819,n23);
or (n6819,n6820,n929);
or (n6820,n6821,n928);
or (n6821,n6822,n2983);
or (n6822,n6823,n944);
or (n6823,n6824,n943);
or (n6824,n6018,n2997);
and (n6825,n3060,n948);
and (n6826,n3061,n3132);
and (n6827,n908,n939);
nor (n6828,n6829,n6951);
wire s0n6829,s1n6829,notn6829;
or (n6829,s0n6829,s1n6829);
not(notn6829,n6950);
and (s0n6829,notn6829,n6830);
and (s1n6829,n6950,n6945);
wire s0n6830,s1n6830,notn6830;
or (n6830,s0n6830,s1n6830);
not(notn6830,n6839);
and (s0n6830,notn6830,1'b0);
and (s1n6830,n6839,n6831);
wire s0n6831,s1n6831,notn6831;
or (n6831,s0n6831,s1n6831);
not(notn6831,n48);
and (s0n6831,notn6831,n6832);
and (s1n6831,n48,n6838);
or (n6832,1'b0,n6833,n6834,n6835,n6836);
and (n6833,n1040,n903);
and (n6834,n2474,n949);
and (n6835,n3190,n901);
and (n6836,n6837,n960);
wire s0n6838,s1n6838,notn6838;
or (n6838,s0n6838,s1n6838);
not(notn6838,n21);
and (s0n6838,notn6838,1'b0);
and (s1n6838,n21,n6837);
and (n6839,n6840,n6893);
and (n6840,n66,n6841);
and (n6841,n6842,n6890);
not (n6842,n6843);
wire s0n6843,s1n6843,notn6843;
or (n6843,s0n6843,s1n6843);
not(notn6843,n66);
and (s0n6843,notn6843,1'b0);
and (s1n6843,n66,n6844);
wire s0n6844,s1n6844,notn6844;
or (n6844,s0n6844,s1n6844);
not(notn6844,n629);
and (s0n6844,notn6844,n6845);
and (s1n6844,n629,n6881);
or (n6845,n6846,n6857,n6868,n6879);
and (n6846,n6847,n53);
wire s0n6847,s1n6847,notn6847;
or (n6847,s0n6847,s1n6847);
not(notn6847,n48);
and (s0n6847,notn6847,n6848);
and (s1n6847,n48,n6849);
or (n6849,n6850,n6852,n6854,n6856);
and (n6850,n6851,n36);
and (n6852,n6853,n41);
and (n6854,n6855,n45);
and (n6856,n6848,n47);
and (n6857,n6858,n58);
wire s0n6858,s1n6858,notn6858;
or (n6858,s0n6858,s1n6858);
not(notn6858,n48);
and (s0n6858,notn6858,n6859);
and (s1n6858,n48,n6860);
or (n6860,n6861,n6863,n6865,n6867);
and (n6861,n6862,n36);
and (n6863,n6864,n41);
and (n6865,n6866,n45);
and (n6867,n6859,n47);
and (n6868,n6869,n62);
wire s0n6869,s1n6869,notn6869;
or (n6869,s0n6869,s1n6869);
not(notn6869,n48);
and (s0n6869,notn6869,n6870);
and (s1n6869,n48,n6871);
or (n6871,n6872,n6874,n6876,n6878);
and (n6872,n6873,n36);
and (n6874,n6875,n41);
and (n6876,n6877,n45);
and (n6878,n6870,n47);
and (n6879,n6880,n65);
wire s0n6880,s1n6880,notn6880;
or (n6880,s0n6880,s1n6880);
not(notn6880,n48);
and (s0n6880,notn6880,n6881);
and (s1n6880,n48,n6882);
or (n6882,n6883,n6885,n6887,n6889);
and (n6883,n6884,n36);
and (n6885,n6886,n41);
and (n6887,n6888,n45);
and (n6889,n6881,n47);
and (n6890,n6891,n6892);
not (n6891,n820);
not (n6892,n746);
and (n6893,n6894,n6942);
not (n6894,n6895);
wire s0n6895,s1n6895,notn6895;
or (n6895,s0n6895,s1n6895);
not(notn6895,n66);
and (s0n6895,notn6895,1'b0);
and (s1n6895,n66,n6896);
wire s0n6896,s1n6896,notn6896;
or (n6896,s0n6896,s1n6896);
not(notn6896,n629);
and (s0n6896,notn6896,n6897);
and (s1n6896,n629,n6933);
or (n6897,n6898,n6909,n6920,n6931);
and (n6898,n6899,n53);
wire s0n6899,s1n6899,notn6899;
or (n6899,s0n6899,s1n6899);
not(notn6899,n48);
and (s0n6899,notn6899,n6900);
and (s1n6899,n48,n6901);
or (n6901,n6902,n6904,n6906,n6908);
and (n6902,n6903,n36);
and (n6904,n6905,n41);
and (n6906,n6907,n45);
and (n6908,n6900,n47);
and (n6909,n6910,n58);
wire s0n6910,s1n6910,notn6910;
or (n6910,s0n6910,s1n6910);
not(notn6910,n48);
and (s0n6910,notn6910,n6911);
and (s1n6910,n48,n6912);
or (n6912,n6913,n6915,n6917,n6919);
and (n6913,n6914,n36);
and (n6915,n6916,n41);
and (n6917,n6918,n45);
and (n6919,n6911,n47);
and (n6920,n6921,n62);
wire s0n6921,s1n6921,notn6921;
or (n6921,s0n6921,s1n6921);
not(notn6921,n48);
and (s0n6921,notn6921,n6922);
and (s1n6921,n48,n6923);
or (n6923,n6924,n6926,n6928,n6930);
and (n6924,n6925,n36);
and (n6926,n6927,n41);
and (n6928,n6929,n45);
and (n6930,n6922,n47);
and (n6931,n6932,n65);
wire s0n6932,s1n6932,notn6932;
or (n6932,s0n6932,s1n6932);
not(notn6932,n48);
and (s0n6932,notn6932,n6933);
and (s1n6932,n48,n6934);
or (n6934,n6935,n6937,n6939,n6941);
and (n6935,n6936,n36);
and (n6937,n6938,n41);
and (n6939,n6940,n45);
and (n6941,n6933,n47);
and (n6942,n6943,n6944);
not (n6943,n673);
not (n6944,n27);
or (n6945,1'b0,n6946,n6947,n6948,n6949);
and (n6946,n2991,n981);
and (n6947,n3013,n1002);
and (n6948,n3033,n1022);
and (n6949,n3053,n1042);
and (n6950,n594,n2955);
and (n6951,n6952,n8766);
nand (n6952,n6953,n8737);
not (n6953,n6954);
or (n6954,n6955,n8736);
and (n6955,n6956,n8272);
xor (n6956,n6957,n8199);
xor (n6957,n6958,n8136);
xor (n6958,n6959,n8105);
or (n6959,n6960,n8104);
and (n6960,n6961,n7932);
xor (n6961,n6962,n7889);
xor (n6962,n6963,n7756);
xor (n6963,n6964,n7313);
xor (n6964,n6965,n7309);
xor (n6965,n6966,n7135);
wire s0n6966,s1n6966,notn6966;
or (n6966,s0n6966,s1n6966);
not(notn6966,n7134);
and (s0n6966,notn6966,1'b0);
and (s1n6966,n7134,n6967);
xor (n6967,n6968,n6973);
wire s0n6968,s1n6968,notn6968;
or (n6968,s0n6968,s1n6968);
not(notn6968,n6841);
and (s0n6968,notn6968,1'b0);
and (s1n6968,n6841,n6969);
wire s0n6969,s1n6969,notn6969;
or (n6969,s0n6969,s1n6969);
not(notn6969,n6972);
and (s0n6969,notn6969,n6970);
and (s1n6969,n6972,n6832);
wire s0n6970,s1n6970,notn6970;
or (n6970,s0n6970,s1n6970);
not(notn6970,n6971);
and (s0n6970,notn6970,1'b0);
and (s1n6970,n6971,n6837);
and (n6971,n49,n903);
and (n6972,n66,n983);
or (n6973,n6974,n7075,n7133);
and (n6974,n6975,n6987);
xor (n6975,n6976,n6985);
wire s0n6976,s1n6976,notn6976;
or (n6976,s0n6976,s1n6976);
not(notn6976,n6841);
and (s0n6976,notn6976,1'b0);
and (s1n6976,n6841,n6977);
wire s0n6977,s1n6977,notn6977;
or (n6977,s0n6977,s1n6977);
not(notn6977,n6972);
and (s0n6977,notn6977,n6978);
and (s1n6977,n6972,n6980);
wire s0n6978,s1n6978,notn6978;
or (n6978,s0n6978,s1n6978);
not(notn6978,n6971);
and (s0n6978,notn6978,1'b0);
and (s1n6978,n6971,n6979);
or (n6980,1'b0,n6981,n6982,n6983,n6984);
and (n6981,n1150,n903);
and (n6982,n2519,n949);
and (n6983,n3315,n901);
and (n6984,n6979,n960);
wire s0n6985,s1n6985,notn6985;
or (n6985,s0n6985,s1n6985);
not(notn6985,n6986);
and (s0n6985,notn6985,1'b0);
and (s1n6985,n6986,n6969);
xor (n6986,n6842,n6890);
and (n6987,n6988,n6990);
wire s0n6988,s1n6988,notn6988;
or (n6988,s0n6988,s1n6988);
not(notn6988,n6989);
and (s0n6988,notn6988,1'b0);
and (s1n6988,n6989,n6969);
xor (n6989,n6891,n6892);
or (n6990,n6991,n6994,n7074);
and (n6991,n6992,n6993);
wire s0n6992,s1n6992,notn6992;
or (n6992,s0n6992,s1n6992);
not(notn6992,n6989);
and (s0n6992,notn6992,1'b0);
and (s1n6992,n6989,n6977);
wire s0n6993,s1n6993,notn6993;
or (n6993,s0n6993,s1n6993);
not(notn6993,n746);
and (s0n6993,notn6993,1'b0);
and (s1n6993,n746,n6969);
and (n6994,n6993,n6995);
or (n6995,n6996,n7007,n7073);
and (n6996,n6997,n7006);
wire s0n6997,s1n6997,notn6997;
or (n6997,s0n6997,s1n6997);
not(notn6997,n6989);
and (s0n6997,notn6997,1'b0);
and (s1n6997,n6989,n6998);
wire s0n6998,s1n6998,notn6998;
or (n6998,s0n6998,s1n6998);
not(notn6998,n6972);
and (s0n6998,notn6998,n6999);
and (s1n6998,n6972,n7001);
wire s0n6999,s1n6999,notn6999;
or (n6999,s0n6999,s1n6999);
not(notn6999,n6971);
and (s0n6999,notn6999,1'b0);
and (s1n6999,n6971,n7000);
or (n7001,1'b0,n7002,n7003,n7004,n7005);
and (n7002,n1257,n903);
and (n7003,n2564,n949);
and (n7004,n3440,n901);
and (n7005,n7000,n960);
wire s0n7006,s1n7006,notn7006;
or (n7006,s0n7006,s1n7006);
not(notn7006,n746);
and (s0n7006,notn7006,1'b0);
and (s1n7006,n746,n6977);
and (n7007,n7006,n7008);
or (n7008,n7009,n7020,n7072);
and (n7009,n7010,n7019);
wire s0n7010,s1n7010,notn7010;
or (n7010,s0n7010,s1n7010);
not(notn7010,n6989);
and (s0n7010,notn7010,1'b0);
and (s1n7010,n6989,n7011);
wire s0n7011,s1n7011,notn7011;
or (n7011,s0n7011,s1n7011);
not(notn7011,n6972);
and (s0n7011,notn7011,n7012);
and (s1n7011,n6972,n7014);
wire s0n7012,s1n7012,notn7012;
or (n7012,s0n7012,s1n7012);
not(notn7012,n6971);
and (s0n7012,notn7012,1'b0);
and (s1n7012,n6971,n7013);
or (n7014,1'b0,n7015,n7016,n7017,n7018);
and (n7015,n1364,n903);
and (n7016,n2609,n949);
and (n7017,n3565,n901);
and (n7018,n7013,n960);
wire s0n7019,s1n7019,notn7019;
or (n7019,s0n7019,s1n7019);
not(notn7019,n746);
and (s0n7019,notn7019,1'b0);
and (s1n7019,n746,n6998);
and (n7020,n7019,n7021);
or (n7021,n7022,n7033,n7071);
and (n7022,n7023,n7032);
wire s0n7023,s1n7023,notn7023;
or (n7023,s0n7023,s1n7023);
not(notn7023,n6989);
and (s0n7023,notn7023,1'b0);
and (s1n7023,n6989,n7024);
wire s0n7024,s1n7024,notn7024;
or (n7024,s0n7024,s1n7024);
not(notn7024,n6972);
and (s0n7024,notn7024,n7025);
and (s1n7024,n6972,n7027);
wire s0n7025,s1n7025,notn7025;
or (n7025,s0n7025,s1n7025);
not(notn7025,n6971);
and (s0n7025,notn7025,1'b0);
and (s1n7025,n6971,n7026);
or (n7027,1'b0,n7028,n7029,n7030,n7031);
and (n7028,n1471,n903);
and (n7029,n2654,n949);
and (n7030,n3690,n901);
and (n7031,n7026,n960);
wire s0n7032,s1n7032,notn7032;
or (n7032,s0n7032,s1n7032);
not(notn7032,n746);
and (s0n7032,notn7032,1'b0);
and (s1n7032,n746,n7011);
and (n7033,n7032,n7034);
or (n7034,n7035,n7046,n7048);
and (n7035,n7036,n7045);
wire s0n7036,s1n7036,notn7036;
or (n7036,s0n7036,s1n7036);
not(notn7036,n6989);
and (s0n7036,notn7036,1'b0);
and (s1n7036,n6989,n7037);
wire s0n7037,s1n7037,notn7037;
or (n7037,s0n7037,s1n7037);
not(notn7037,n6972);
and (s0n7037,notn7037,n7038);
and (s1n7037,n6972,n7040);
wire s0n7038,s1n7038,notn7038;
or (n7038,s0n7038,s1n7038);
not(notn7038,n6971);
and (s0n7038,notn7038,1'b0);
and (s1n7038,n6971,n7039);
or (n7040,1'b0,n7041,n7042,n7043,n7044);
and (n7041,n1578,n903);
and (n7042,n2699,n949);
and (n7043,n3815,n901);
and (n7044,n7039,n960);
wire s0n7045,s1n7045,notn7045;
or (n7045,s0n7045,s1n7045);
not(notn7045,n746);
and (s0n7045,notn7045,1'b0);
and (s1n7045,n746,n7024);
and (n7046,n7045,n7047);
or (n7047,n7048,n7059,n7060);
and (n7048,n7049,n7058);
wire s0n7049,s1n7049,notn7049;
or (n7049,s0n7049,s1n7049);
not(notn7049,n6989);
and (s0n7049,notn7049,1'b0);
and (s1n7049,n6989,n7050);
wire s0n7050,s1n7050,notn7050;
or (n7050,s0n7050,s1n7050);
not(notn7050,n6972);
and (s0n7050,notn7050,n7051);
and (s1n7050,n6972,n7053);
wire s0n7051,s1n7051,notn7051;
or (n7051,s0n7051,s1n7051);
not(notn7051,n6971);
and (s0n7051,notn7051,1'b0);
and (s1n7051,n6971,n7052);
or (n7053,1'b0,n7054,n7055,n7056,n7057);
and (n7054,n1685,n903);
and (n7055,n2744,n949);
and (n7056,n3940,n901);
and (n7057,n7052,n960);
wire s0n7058,s1n7058,notn7058;
or (n7058,s0n7058,s1n7058);
not(notn7058,n746);
and (s0n7058,notn7058,1'b0);
and (s1n7058,n746,n7037);
and (n7059,n7058,n7060);
and (n7060,n7061,n7070);
wire s0n7061,s1n7061,notn7061;
or (n7061,s0n7061,s1n7061);
not(notn7061,n6989);
and (s0n7061,notn7061,1'b0);
and (s1n7061,n6989,n7062);
wire s0n7062,s1n7062,notn7062;
or (n7062,s0n7062,s1n7062);
not(notn7062,n6972);
and (s0n7062,notn7062,n7063);
and (s1n7062,n6972,n7065);
wire s0n7063,s1n7063,notn7063;
or (n7063,s0n7063,s1n7063);
not(notn7063,n6971);
and (s0n7063,notn7063,1'b0);
and (s1n7063,n6971,n7064);
or (n7065,1'b0,n7066,n7067,n7068,n7069);
and (n7066,n1791,n903);
and (n7067,n2788,n949);
and (n7068,n4064,n901);
and (n7069,n7064,n960);
wire s0n7070,s1n7070,notn7070;
or (n7070,s0n7070,s1n7070);
not(notn7070,n746);
and (s0n7070,notn7070,1'b0);
and (s1n7070,n746,n7050);
and (n7071,n7023,n7034);
and (n7072,n7010,n7021);
and (n7073,n6997,n7008);
and (n7074,n6992,n6995);
and (n7075,n6987,n7076);
or (n7076,n7077,n7082,n7132);
and (n7077,n7078,n7081);
xor (n7078,n7079,n7080);
wire s0n7079,s1n7079,notn7079;
or (n7079,s0n7079,s1n7079);
not(notn7079,n6841);
and (s0n7079,notn7079,1'b0);
and (s1n7079,n6841,n6998);
wire s0n7080,s1n7080,notn7080;
or (n7080,s0n7080,s1n7080);
not(notn7080,n6986);
and (s0n7080,notn7080,1'b0);
and (s1n7080,n6986,n6977);
xor (n7081,n6988,n6990);
and (n7082,n7081,n7083);
or (n7083,n7084,n7090,n7131);
and (n7084,n7085,n7088);
xor (n7085,n7086,n7087);
wire s0n7086,s1n7086,notn7086;
or (n7086,s0n7086,s1n7086);
not(notn7086,n6841);
and (s0n7086,notn7086,1'b0);
and (s1n7086,n6841,n7011);
wire s0n7087,s1n7087,notn7087;
or (n7087,s0n7087,s1n7087);
not(notn7087,n6986);
and (s0n7087,notn7087,1'b0);
and (s1n7087,n6986,n6998);
xor (n7088,n7089,n6995);
xor (n7089,n6992,n6993);
and (n7090,n7088,n7091);
or (n7091,n7092,n7098,n7130);
and (n7092,n7093,n7096);
xor (n7093,n7094,n7095);
wire s0n7094,s1n7094,notn7094;
or (n7094,s0n7094,s1n7094);
not(notn7094,n6841);
and (s0n7094,notn7094,1'b0);
and (s1n7094,n6841,n7024);
wire s0n7095,s1n7095,notn7095;
or (n7095,s0n7095,s1n7095);
not(notn7095,n6986);
and (s0n7095,notn7095,1'b0);
and (s1n7095,n6986,n7011);
xor (n7096,n7097,n7008);
xor (n7097,n6997,n7006);
and (n7098,n7096,n7099);
or (n7099,n7100,n7106,n7129);
and (n7100,n7101,n7104);
xor (n7101,n7102,n7103);
wire s0n7102,s1n7102,notn7102;
or (n7102,s0n7102,s1n7102);
not(notn7102,n6841);
and (s0n7102,notn7102,1'b0);
and (s1n7102,n6841,n7037);
wire s0n7103,s1n7103,notn7103;
or (n7103,s0n7103,s1n7103);
not(notn7103,n6986);
and (s0n7103,notn7103,1'b0);
and (s1n7103,n6986,n7024);
xor (n7104,n7105,n7021);
xor (n7105,n7010,n7019);
and (n7106,n7104,n7107);
or (n7107,n7108,n7114,n7128);
and (n7108,n7109,n7112);
xor (n7109,n7110,n7111);
wire s0n7110,s1n7110,notn7110;
or (n7110,s0n7110,s1n7110);
not(notn7110,n6841);
and (s0n7110,notn7110,1'b0);
and (s1n7110,n6841,n7050);
wire s0n7111,s1n7111,notn7111;
or (n7111,s0n7111,s1n7111);
not(notn7111,n6986);
and (s0n7111,notn7111,1'b0);
and (s1n7111,n6986,n7037);
xor (n7112,n7113,n7034);
xor (n7113,n7023,n7032);
and (n7114,n7112,n7115);
or (n7115,n7116,n7122,n7127);
and (n7116,n7117,n7120);
xor (n7117,n7118,n7119);
wire s0n7118,s1n7118,notn7118;
or (n7118,s0n7118,s1n7118);
not(notn7118,n6841);
and (s0n7118,notn7118,1'b0);
and (s1n7118,n6841,n7062);
wire s0n7119,s1n7119,notn7119;
or (n7119,s0n7119,s1n7119);
not(notn7119,n6986);
and (s0n7119,notn7119,1'b0);
and (s1n7119,n6986,n7050);
xor (n7120,n7121,n7047);
xor (n7121,n7036,n7045);
and (n7122,n7120,n7123);
and (n7123,n7124,n7125);
wire s0n7124,s1n7124,notn7124;
or (n7124,s0n7124,s1n7124);
not(notn7124,n6986);
and (s0n7124,notn7124,1'b0);
and (s1n7124,n6986,n7062);
xor (n7125,n7126,n7060);
xor (n7126,n7049,n7058);
and (n7127,n7117,n7123);
and (n7128,n7109,n7115);
and (n7129,n7101,n7107);
and (n7130,n7093,n7099);
and (n7131,n7085,n7091);
and (n7132,n7078,n7083);
and (n7133,n6975,n7076);
xor (n7134,n6943,n6944);
wire s0n7135,s1n7135,notn7135;
or (n7135,s0n7135,s1n7135);
not(notn7135,n6895);
and (s0n7135,notn7135,1'b0);
and (s1n7135,n6895,n7136);
xor (n7136,n7137,n7176);
xor (n7137,n7138,n7157);
xor (n7138,n7139,n7148);
wire s0n7139,s1n7139,notn7139;
or (n7139,s0n7139,s1n7139);
not(notn7139,n6841);
and (s0n7139,notn7139,1'b0);
and (s1n7139,n6841,n7140);
wire s0n7140,s1n7140,notn7140;
or (n7140,s0n7140,s1n7140);
not(notn7140,n6972);
and (s0n7140,notn7140,n7141);
and (s1n7140,n6972,n7143);
wire s0n7141,s1n7141,notn7141;
or (n7141,s0n7141,s1n7141);
not(notn7141,n6971);
and (s0n7141,notn7141,1'b0);
and (s1n7141,n6971,n7142);
or (n7143,1'b0,n7144,n7145,n7146,n7147);
and (n7144,n1151,n903);
and (n7145,n2520,n949);
and (n7146,n5020,n901);
and (n7147,n7142,n960);
wire s0n7148,s1n7148,notn7148;
or (n7148,s0n7148,s1n7148);
not(notn7148,n6986);
and (s0n7148,notn7148,1'b0);
and (s1n7148,n6986,n7149);
wire s0n7149,s1n7149,notn7149;
or (n7149,s0n7149,s1n7149);
not(notn7149,n6972);
and (s0n7149,notn7149,n7150);
and (s1n7149,n6972,n7152);
wire s0n7150,s1n7150,notn7150;
or (n7150,s0n7150,s1n7150);
not(notn7150,n6971);
and (s0n7150,notn7150,1'b0);
and (s1n7150,n6971,n7151);
or (n7152,1'b0,n7153,n7154,n7155,n7156);
and (n7153,n1041,n903);
and (n7154,n2475,n949);
and (n7155,n4949,n901);
and (n7156,n7151,n960);
or (n7157,n7158,n7175);
and (n7158,n7159,n7172);
xor (n7159,n7160,n7161);
wire s0n7160,s1n7160,notn7160;
or (n7160,s0n7160,s1n7160);
not(notn7160,n6986);
and (s0n7160,notn7160,1'b0);
and (s1n7160,n6986,n7140);
xor (n7161,n7162,n7163);
wire s0n7162,s1n7162,notn7162;
or (n7162,s0n7162,s1n7162);
not(notn7162,n6989);
and (s0n7162,notn7162,1'b0);
and (s1n7162,n6989,n7149);
wire s0n7163,s1n7163,notn7163;
or (n7163,s0n7163,s1n7163);
not(notn7163,n6841);
and (s0n7163,notn7163,1'b0);
and (s1n7163,n6841,n7164);
wire s0n7164,s1n7164,notn7164;
or (n7164,s0n7164,s1n7164);
not(notn7164,n6972);
and (s0n7164,notn7164,n7165);
and (s1n7164,n6972,n7167);
wire s0n7165,s1n7165,notn7165;
or (n7165,s0n7165,s1n7165);
not(notn7165,n6971);
and (s0n7165,notn7165,1'b0);
and (s1n7165,n6971,n7166);
or (n7167,1'b0,n7168,n7169,n7170,n7171);
and (n7168,n1258,n903);
and (n7169,n2565,n949);
and (n7170,n5091,n901);
and (n7171,n7166,n960);
and (n7172,n7173,n7174);
wire s0n7173,s1n7173,notn7173;
or (n7173,s0n7173,s1n7173);
not(notn7173,n6989);
and (s0n7173,notn7173,1'b0);
and (s1n7173,n6989,n7140);
wire s0n7174,s1n7174,notn7174;
or (n7174,s0n7174,s1n7174);
not(notn7174,n746);
and (s0n7174,notn7174,1'b0);
and (s1n7174,n746,n7149);
and (n7175,n7160,n7161);
nand (n7176,n7177,n7308);
or (n7177,n7178,n7303);
nor (n7178,n7179,n7302);
and (n7179,n7180,n7291);
nand (n7180,n7181,n7290);
or (n7181,n7182,n7230);
not (n7182,n7183);
or (n7183,n7184,n7211);
xor (n7184,n7185,n7208);
xor (n7185,n7186,n7195);
wire s0n7186,s1n7186,notn7186;
or (n7186,s0n7186,s1n7186);
not(notn7186,n6986);
and (s0n7186,notn7186,1'b0);
and (s1n7186,n6986,n7187);
wire s0n7187,s1n7187,notn7187;
or (n7187,s0n7187,s1n7187);
not(notn7187,n6972);
and (s0n7187,notn7187,n7188);
and (s1n7187,n6972,n7190);
wire s0n7188,s1n7188,notn7188;
or (n7188,s0n7188,s1n7188);
not(notn7188,n6971);
and (s0n7188,notn7188,1'b0);
and (s1n7188,n6971,n7189);
or (n7190,1'b0,n7191,n7192,n7193,n7194);
and (n7191,n1365,n903);
and (n7192,n2610,n949);
and (n7193,n5162,n901);
and (n7194,n7189,n960);
xor (n7195,n7196,n7199);
xor (n7196,n7197,n7198);
wire s0n7197,s1n7197,notn7197;
or (n7197,s0n7197,s1n7197);
not(notn7197,n6989);
and (s0n7197,notn7197,1'b0);
and (s1n7197,n6989,n7164);
wire s0n7198,s1n7198,notn7198;
or (n7198,s0n7198,s1n7198);
not(notn7198,n746);
and (s0n7198,notn7198,1'b0);
and (s1n7198,n746,n7140);
wire s0n7199,s1n7199,notn7199;
or (n7199,s0n7199,s1n7199);
not(notn7199,n6841);
and (s0n7199,notn7199,1'b0);
and (s1n7199,n6841,n7200);
wire s0n7200,s1n7200,notn7200;
or (n7200,s0n7200,s1n7200);
not(notn7200,n6972);
and (s0n7200,notn7200,n7201);
and (s1n7200,n6972,n7203);
wire s0n7201,s1n7201,notn7201;
or (n7201,s0n7201,s1n7201);
not(notn7201,n6971);
and (s0n7201,notn7201,1'b0);
and (s1n7201,n6971,n7202);
or (n7203,1'b0,n7204,n7205,n7206,n7207);
and (n7204,n1472,n903);
and (n7205,n2655,n949);
and (n7206,n5233,n901);
and (n7207,n7202,n960);
and (n7208,n7209,n7210);
wire s0n7209,s1n7209,notn7209;
or (n7209,s0n7209,s1n7209);
not(notn7209,n6989);
and (s0n7209,notn7209,1'b0);
and (s1n7209,n6989,n7187);
wire s0n7210,s1n7210,notn7210;
or (n7210,s0n7210,s1n7210);
not(notn7210,n746);
and (s0n7210,notn7210,1'b0);
and (s1n7210,n746,n7164);
or (n7211,n7212,n7229);
and (n7212,n7213,n7226);
xor (n7213,n7214,n7215);
wire s0n7214,s1n7214,notn7214;
or (n7214,s0n7214,s1n7214);
not(notn7214,n6986);
and (s0n7214,notn7214,1'b0);
and (s1n7214,n6986,n7200);
xor (n7215,n7216,n7217);
xor (n7216,n7209,n7210);
wire s0n7217,s1n7217,notn7217;
or (n7217,s0n7217,s1n7217);
not(notn7217,n6841);
and (s0n7217,notn7217,1'b0);
and (s1n7217,n6841,n7218);
wire s0n7218,s1n7218,notn7218;
or (n7218,s0n7218,s1n7218);
not(notn7218,n6972);
and (s0n7218,notn7218,n7219);
and (s1n7218,n6972,n7221);
wire s0n7219,s1n7219,notn7219;
or (n7219,s0n7219,s1n7219);
not(notn7219,n6971);
and (s0n7219,notn7219,1'b0);
and (s1n7219,n6971,n7220);
or (n7221,1'b0,n7222,n7223,n7224,n7225);
and (n7222,n1579,n903);
and (n7223,n2700,n949);
and (n7224,n5304,n901);
and (n7225,n7220,n960);
and (n7226,n7227,n7228);
wire s0n7227,s1n7227,notn7227;
or (n7227,s0n7227,s1n7227);
not(notn7227,n6989);
and (s0n7227,notn7227,1'b0);
and (s1n7227,n6989,n7200);
wire s0n7228,s1n7228,notn7228;
or (n7228,s0n7228,s1n7228);
not(notn7228,n746);
and (s0n7228,notn7228,1'b0);
and (s1n7228,n746,n7187);
and (n7229,n7214,n7215);
not (n7230,n7231);
nand (n7231,n7232,n7286,n7289);
nand (n7232,n7233,n7254,n7283);
or (n7233,n7234,n7235);
xor (n7234,n7213,n7226);
or (n7235,n7236,n7253);
and (n7236,n7237,n7242);
xor (n7237,n7238,n7239);
wire s0n7238,s1n7238,notn7238;
or (n7238,s0n7238,s1n7238);
not(notn7238,n6986);
and (s0n7238,notn7238,1'b0);
and (s1n7238,n6986,n7218);
and (n7239,n7240,n7241);
wire s0n7240,s1n7240,notn7240;
or (n7240,s0n7240,s1n7240);
not(notn7240,n6989);
and (s0n7240,notn7240,1'b0);
and (s1n7240,n6989,n7218);
wire s0n7241,s1n7241,notn7241;
or (n7241,s0n7241,s1n7241);
not(notn7241,n746);
and (s0n7241,notn7241,1'b0);
and (s1n7241,n746,n7200);
xor (n7242,n7243,n7244);
xor (n7243,n7227,n7228);
wire s0n7244,s1n7244,notn7244;
or (n7244,s0n7244,s1n7244);
not(notn7244,n6841);
and (s0n7244,notn7244,1'b0);
and (s1n7244,n6841,n7245);
wire s0n7245,s1n7245,notn7245;
or (n7245,s0n7245,s1n7245);
not(notn7245,n6972);
and (s0n7245,notn7245,n7246);
and (s1n7245,n6972,n7248);
wire s0n7246,s1n7246,notn7246;
or (n7246,s0n7246,s1n7246);
not(notn7246,n6971);
and (s0n7246,notn7246,1'b0);
and (s1n7246,n6971,n7247);
or (n7248,1'b0,n7249,n7250,n7251,n7252);
and (n7249,n1686,n903);
and (n7250,n2745,n949);
and (n7251,n5375,n901);
and (n7252,n7247,n960);
and (n7253,n7238,n7239);
or (n7254,n7255,n7282);
and (n7255,n7256,n7277);
xor (n7256,n7257,n7260);
and (n7257,n7258,n7259);
wire s0n7258,s1n7258,notn7258;
or (n7258,s0n7258,s1n7258);
not(notn7258,n6989);
and (s0n7258,notn7258,1'b0);
and (s1n7258,n6989,n7245);
wire s0n7259,s1n7259,notn7259;
or (n7259,s0n7259,s1n7259);
not(notn7259,n746);
and (s0n7259,notn7259,1'b0);
and (s1n7259,n746,n7218);
or (n7260,n7261,n7276);
and (n7261,n7262,n7275);
xor (n7262,n7263,n7274);
and (n7263,n7264,n7273);
wire s0n7264,s1n7264,notn7264;
or (n7264,s0n7264,s1n7264);
not(notn7264,n6989);
and (s0n7264,notn7264,1'b0);
and (s1n7264,n6989,n7265);
wire s0n7265,s1n7265,notn7265;
or (n7265,s0n7265,s1n7265);
not(notn7265,n6972);
and (s0n7265,notn7265,n7266);
and (s1n7265,n6972,n7268);
wire s0n7266,s1n7266,notn7266;
or (n7266,s0n7266,s1n7266);
not(notn7266,n6971);
and (s0n7266,notn7266,1'b0);
and (s1n7266,n6971,n7267);
or (n7268,1'b0,n7269,n7270,n7271,n7272);
and (n7269,n1792,n903);
and (n7270,n2789,n949);
and (n7271,n5445,n901);
and (n7272,n7267,n960);
wire s0n7273,s1n7273,notn7273;
or (n7273,s0n7273,s1n7273);
not(notn7273,n746);
and (s0n7273,notn7273,1'b0);
and (s1n7273,n746,n7245);
wire s0n7274,s1n7274,notn7274;
or (n7274,s0n7274,s1n7274);
not(notn7274,n6986);
and (s0n7274,notn7274,1'b0);
and (s1n7274,n6986,n7265);
xor (n7275,n7258,n7259);
and (n7276,n7263,n7274);
xor (n7277,n7278,n7281);
xor (n7278,n7279,n7280);
wire s0n7279,s1n7279,notn7279;
or (n7279,s0n7279,s1n7279);
not(notn7279,n6841);
and (s0n7279,notn7279,1'b0);
and (s1n7279,n6841,n7265);
xor (n7280,n7240,n7241);
wire s0n7281,s1n7281,notn7281;
or (n7281,s0n7281,s1n7281);
not(notn7281,n6986);
and (s0n7281,notn7281,1'b0);
and (s1n7281,n6986,n7245);
and (n7282,n7257,n7260);
or (n7283,n7284,n7285);
xor (n7284,n7237,n7242);
and (n7285,n7278,n7281);
nand (n7286,n7287,n7233);
not (n7287,n7288);
nand (n7288,n7284,n7285);
nand (n7289,n7234,n7235);
nand (n7290,n7184,n7211);
or (n7291,n7292,n7299);
xor (n7292,n7293,n7298);
xor (n7293,n7294,n7295);
wire s0n7294,s1n7294,notn7294;
or (n7294,s0n7294,s1n7294);
not(notn7294,n6986);
and (s0n7294,notn7294,1'b0);
and (s1n7294,n6986,n7164);
xor (n7295,n7296,n7297);
xor (n7296,n7173,n7174);
wire s0n7297,s1n7297,notn7297;
or (n7297,s0n7297,s1n7297);
not(notn7297,n6841);
and (s0n7297,notn7297,1'b0);
and (s1n7297,n6841,n7187);
and (n7298,n7197,n7198);
or (n7299,n7300,n7301);
and (n7300,n7185,n7208);
and (n7301,n7186,n7195);
and (n7302,n7292,n7299);
nor (n7303,n7304,n7307);
or (n7304,n7305,n7306);
and (n7305,n7293,n7298);
and (n7306,n7294,n7295);
xor (n7307,n7159,n7172);
nand (n7308,n7304,n7307);
wire s0n7309,s1n7309,notn7309;
or (n7309,s0n7309,s1n7309);
not(notn7309,n7312);
and (s0n7309,notn7309,1'b0);
and (s1n7309,n7312,n7310);
xor (n7310,n7311,n7076);
xor (n7311,n6975,n6987);
xor (n7312,n6894,n6942);
xor (n7313,n7314,n7695);
xor (n7314,n7315,n7679);
or (n7315,n7316,n7678);
and (n7316,n7317,n7536);
xor (n7317,n7318,n7524);
and (n7318,n7319,n7509);
xor (n7319,n7320,n7434);
wire s0n7320,s1n7320,notn7320;
or (n7320,s0n7320,s1n7320);
not(notn7320,n6893);
and (s0n7320,notn7320,1'b0);
and (s1n7320,n6893,n7321);
xor (n7321,n7322,n7409);
xor (n7322,n7323,n7332);
wire s0n7323,s1n7323,notn7323;
or (n7323,s0n7323,s1n7323);
not(notn7323,n6843);
and (s0n7323,notn7323,1'b0);
and (s1n7323,n6843,n7324);
wire s0n7324,s1n7324,notn7324;
or (n7324,s0n7324,s1n7324);
not(notn7324,n6972);
and (s0n7324,notn7324,n7325);
and (s1n7324,n6972,n7327);
wire s0n7325,s1n7325,notn7325;
or (n7325,s0n7325,s1n7325);
not(notn7325,n6971);
and (s0n7325,notn7325,1'b0);
and (s1n7325,n6971,n7326);
or (n7327,1'b0,n7328,n7329,n7330,n7331);
and (n7328,n1360,n903);
and (n7329,n2065,n949);
and (n7330,n3562,n901);
and (n7331,n7326,n960);
xor (n7332,n7333,n7352);
xor (n7333,n7334,n7343);
wire s0n7334,s1n7334,notn7334;
or (n7334,s0n7334,s1n7334);
not(notn7334,n820);
and (s0n7334,notn7334,1'b0);
and (s1n7334,n820,n7335);
wire s0n7335,s1n7335,notn7335;
or (n7335,s0n7335,s1n7335);
not(notn7335,n6972);
and (s0n7335,notn7335,n7336);
and (s1n7335,n6972,n7338);
wire s0n7336,s1n7336,notn7336;
or (n7336,s0n7336,s1n7336);
not(notn7336,n6971);
and (s0n7336,notn7336,1'b0);
and (s1n7336,n6971,n7337);
or (n7338,1'b0,n7339,n7340,n7341,n7342);
and (n7339,n1253,n903);
and (n7340,n2000,n949);
and (n7341,n3437,n901);
and (n7342,n7337,n960);
wire s0n7343,s1n7343,notn7343;
or (n7343,s0n7343,s1n7343);
not(notn7343,n746);
and (s0n7343,notn7343,1'b0);
and (s1n7343,n746,n7344);
wire s0n7344,s1n7344,notn7344;
or (n7344,s0n7344,s1n7344);
not(notn7344,n6972);
and (s0n7344,notn7344,n7345);
and (s1n7344,n6972,n7347);
wire s0n7345,s1n7345,notn7345;
or (n7345,s0n7345,s1n7345);
not(notn7345,n6971);
and (s0n7345,notn7345,1'b0);
and (s1n7345,n6971,n7346);
or (n7347,1'b0,n7348,n7349,n7350,n7351);
and (n7348,n1146,n903);
and (n7349,n1935,n949);
and (n7350,n3312,n901);
and (n7351,n7346,n960);
or (n7352,n7353,n7356,n7408);
and (n7353,n7354,n7355);
wire s0n7354,s1n7354,notn7354;
or (n7354,s0n7354,s1n7354);
not(notn7354,n820);
and (s0n7354,notn7354,1'b0);
and (s1n7354,n820,n7324);
wire s0n7355,s1n7355,notn7355;
or (n7355,s0n7355,s1n7355);
not(notn7355,n746);
and (s0n7355,notn7355,1'b0);
and (s1n7355,n746,n7335);
and (n7356,n7355,n7357);
or (n7357,n7358,n7369,n7407);
and (n7358,n7359,n7368);
wire s0n7359,s1n7359,notn7359;
or (n7359,s0n7359,s1n7359);
not(notn7359,n820);
and (s0n7359,notn7359,1'b0);
and (s1n7359,n820,n7360);
wire s0n7360,s1n7360,notn7360;
or (n7360,s0n7360,s1n7360);
not(notn7360,n6972);
and (s0n7360,notn7360,n7361);
and (s1n7360,n6972,n7363);
wire s0n7361,s1n7361,notn7361;
or (n7361,s0n7361,s1n7361);
not(notn7361,n6971);
and (s0n7361,notn7361,1'b0);
and (s1n7361,n6971,n7362);
or (n7363,1'b0,n7364,n7365,n7366,n7367);
and (n7364,n1467,n903);
and (n7365,n2130,n949);
and (n7366,n3687,n901);
and (n7367,n7362,n960);
wire s0n7368,s1n7368,notn7368;
or (n7368,s0n7368,s1n7368);
not(notn7368,n746);
and (s0n7368,notn7368,1'b0);
and (s1n7368,n746,n7324);
and (n7369,n7368,n7370);
or (n7370,n7371,n7382,n7384);
and (n7371,n7372,n7381);
wire s0n7372,s1n7372,notn7372;
or (n7372,s0n7372,s1n7372);
not(notn7372,n820);
and (s0n7372,notn7372,1'b0);
and (s1n7372,n820,n7373);
wire s0n7373,s1n7373,notn7373;
or (n7373,s0n7373,s1n7373);
not(notn7373,n6972);
and (s0n7373,notn7373,n7374);
and (s1n7373,n6972,n7376);
wire s0n7374,s1n7374,notn7374;
or (n7374,s0n7374,s1n7374);
not(notn7374,n6971);
and (s0n7374,notn7374,1'b0);
and (s1n7374,n6971,n7375);
or (n7376,1'b0,n7377,n7378,n7379,n7380);
and (n7377,n1574,n903);
and (n7378,n2195,n949);
and (n7379,n3812,n901);
and (n7380,n7375,n960);
wire s0n7381,s1n7381,notn7381;
or (n7381,s0n7381,s1n7381);
not(notn7381,n746);
and (s0n7381,notn7381,1'b0);
and (s1n7381,n746,n7360);
and (n7382,n7381,n7383);
or (n7383,n7384,n7395,n7396);
and (n7384,n7385,n7394);
wire s0n7385,s1n7385,notn7385;
or (n7385,s0n7385,s1n7385);
not(notn7385,n820);
and (s0n7385,notn7385,1'b0);
and (s1n7385,n820,n7386);
wire s0n7386,s1n7386,notn7386;
or (n7386,s0n7386,s1n7386);
not(notn7386,n6972);
and (s0n7386,notn7386,n7387);
and (s1n7386,n6972,n7389);
wire s0n7387,s1n7387,notn7387;
or (n7387,s0n7387,s1n7387);
not(notn7387,n6971);
and (s0n7387,notn7387,1'b0);
and (s1n7387,n6971,n7388);
or (n7389,1'b0,n7390,n7391,n7392,n7393);
and (n7390,n1681,n903);
and (n7391,n2260,n949);
and (n7392,n3937,n901);
and (n7393,n7388,n960);
wire s0n7394,s1n7394,notn7394;
or (n7394,s0n7394,s1n7394);
not(notn7394,n746);
and (s0n7394,notn7394,1'b0);
and (s1n7394,n746,n7373);
and (n7395,n7394,n7396);
and (n7396,n7397,n7406);
wire s0n7397,s1n7397,notn7397;
or (n7397,s0n7397,s1n7397);
not(notn7397,n820);
and (s0n7397,notn7397,1'b0);
and (s1n7397,n820,n7398);
wire s0n7398,s1n7398,notn7398;
or (n7398,s0n7398,s1n7398);
not(notn7398,n6972);
and (s0n7398,notn7398,n7399);
and (s1n7398,n6972,n7401);
wire s0n7399,s1n7399,notn7399;
or (n7399,s0n7399,s1n7399);
not(notn7399,n6971);
and (s0n7399,notn7399,1'b0);
and (s1n7399,n6971,n7400);
or (n7401,1'b0,n7402,n7403,n7404,n7405);
and (n7402,n1787,n903);
and (n7403,n2324,n949);
and (n7404,n4061,n901);
and (n7405,n7400,n960);
wire s0n7406,s1n7406,notn7406;
or (n7406,s0n7406,s1n7406);
not(notn7406,n746);
and (s0n7406,notn7406,1'b0);
and (s1n7406,n746,n7386);
and (n7407,n7359,n7370);
and (n7408,n7354,n7357);
or (n7409,n7410,n7414,n7433);
and (n7410,n7411,n7412);
wire s0n7411,s1n7411,notn7411;
or (n7411,s0n7411,s1n7411);
not(notn7411,n6843);
and (s0n7411,notn7411,1'b0);
and (s1n7411,n6843,n7360);
xor (n7412,n7413,n7357);
xor (n7413,n7354,n7355);
and (n7414,n7412,n7415);
or (n7415,n7416,n7420,n7432);
and (n7416,n7417,n7418);
wire s0n7417,s1n7417,notn7417;
or (n7417,s0n7417,s1n7417);
not(notn7417,n6843);
and (s0n7417,notn7417,1'b0);
and (s1n7417,n6843,n7373);
xor (n7418,n7419,n7370);
xor (n7419,n7359,n7368);
and (n7420,n7418,n7421);
or (n7421,n7422,n7426,n7431);
and (n7422,n7423,n7424);
wire s0n7423,s1n7423,notn7423;
or (n7423,s0n7423,s1n7423);
not(notn7423,n6843);
and (s0n7423,notn7423,1'b0);
and (s1n7423,n6843,n7386);
xor (n7424,n7425,n7383);
xor (n7425,n7372,n7381);
and (n7426,n7424,n7427);
and (n7427,n7428,n7429);
wire s0n7428,s1n7428,notn7428;
or (n7428,s0n7428,s1n7428);
not(notn7428,n6843);
and (s0n7428,notn7428,1'b0);
and (s1n7428,n6843,n7398);
xor (n7429,n7430,n7396);
xor (n7430,n7385,n7394);
and (n7431,n7423,n7427);
and (n7432,n7417,n7421);
and (n7433,n7411,n7415);
xor (n7434,n7435,n7470);
xor (n7435,n7436,n7460);
xor (n7436,n7437,n7458);
xor (n7437,n7438,n7448);
and (n7438,n7439,n27);
and (n7439,n6843,n7440);
wire s0n7440,s1n7440,notn7440;
or (n7440,s0n7440,s1n7440);
not(notn7440,n6972);
and (s0n7440,notn7440,n7441);
and (s1n7440,n6972,n7443);
wire s0n7441,s1n7441,notn7441;
or (n7441,s0n7441,s1n7441);
not(notn7441,n6971);
and (s0n7441,notn7441,1'b0);
and (s1n7441,n6971,n7442);
or (n7443,1'b0,n7444,n7445,n7446,n7447);
and (n7444,n1037,n903);
and (n7445,n1871,n949);
and (n7446,n4946,n901);
and (n7447,n7442,n960);
and (n7448,n7449,n27);
wire s0n7449,s1n7449,notn7449;
or (n7449,s0n7449,s1n7449);
not(notn7449,n6843);
and (s0n7449,notn7449,1'b0);
and (s1n7449,n6843,n7450);
wire s0n7450,s1n7450,notn7450;
or (n7450,s0n7450,s1n7450);
not(notn7450,n6972);
and (s0n7450,notn7450,n7451);
and (s1n7450,n6972,n7453);
wire s0n7451,s1n7451,notn7451;
or (n7451,s0n7451,s1n7451);
not(notn7451,n6971);
and (s0n7451,notn7451,1'b0);
and (s1n7451,n6971,n7452);
or (n7453,1'b0,n7454,n7455,n7456,n7457);
and (n7454,n1036,n903);
and (n7455,n1870,n949);
and (n7456,n3187,n901);
and (n7457,n7452,n960);
and (n7458,n7448,n7459);
wire s0n7459,s1n7459,notn7459;
or (n7459,s0n7459,s1n7459);
not(notn7459,n820);
and (s0n7459,notn7459,1'b0);
and (s1n7459,n820,n7344);
and (n7460,n7438,n7461);
wire s0n7461,s1n7461,notn7461;
or (n7461,s0n7461,s1n7461);
not(notn7461,n820);
and (s0n7461,notn7461,1'b0);
and (s1n7461,n820,n7462);
wire s0n7462,s1n7462,notn7462;
or (n7462,s0n7462,s1n7462);
not(notn7462,n6972);
and (s0n7462,notn7462,n7463);
and (s1n7462,n6972,n7465);
wire s0n7463,s1n7463,notn7463;
or (n7463,s0n7463,s1n7463);
not(notn7463,n6971);
and (s0n7463,notn7463,1'b0);
and (s1n7463,n6971,n7464);
or (n7465,1'b0,n7466,n7467,n7468,n7469);
and (n7466,n1147,n903);
and (n7467,n1936,n949);
and (n7468,n5017,n901);
and (n7469,n7464,n960);
or (n7470,n7471,n7508);
and (n7471,n7472,n7488);
xor (n7472,n7473,n7480);
nor (n7473,n7474,n6944);
xnor (n7474,n7475,n7478);
not (n7475,n7476);
not (n7476,n7477);
nand (n7477,n6843,n7462);
not (n7478,n7479);
wire s0n7479,s1n7479,notn7479;
or (n7479,s0n7479,s1n7479);
not(notn7479,n820);
and (s0n7479,notn7479,1'b0);
and (s1n7479,n820,n7440);
and (n7480,n7481,n27);
nand (n7481,n7482,n7486);
or (n7482,n7483,n7485);
not (n7483,n7484);
wire s0n7484,s1n7484,notn7484;
or (n7484,s0n7484,s1n7484);
not(notn7484,n820);
and (s0n7484,notn7484,1'b0);
and (s1n7484,n820,n7450);
wire s0n7485,s1n7485,notn7485;
or (n7485,s0n7485,s1n7485);
not(notn7485,n6843);
and (s0n7485,notn7485,1'b0);
and (s1n7485,n6843,n7344);
or (n7486,n7487,n7484);
not (n7487,n7485);
and (n7488,n7489,n27);
nand (n7489,n7490,n7504);
or (n7490,n7491,n7503);
and (n7491,n7492,n7494);
not (n7492,n7493);
wire s0n7493,s1n7493,notn7493;
or (n7493,s0n7493,s1n7493);
not(notn7493,n746);
and (s0n7493,notn7493,1'b0);
and (s1n7493,n746,n7440);
nand (n7494,n6843,n7495);
wire s0n7495,s1n7495,notn7495;
or (n7495,s0n7495,s1n7495);
not(notn7495,n6972);
and (s0n7495,notn7495,n7496);
and (s1n7495,n6972,n7498);
wire s0n7496,s1n7496,notn7496;
or (n7496,s0n7496,s1n7496);
not(notn7496,n6971);
and (s0n7496,notn7496,1'b0);
and (s1n7496,n6971,n7497);
or (n7498,1'b0,n7499,n7500,n7501,n7502);
and (n7499,n1254,n903);
and (n7500,n2001,n949);
and (n7501,n5088,n901);
and (n7502,n7497,n960);
not (n7503,n7461);
or (n7504,n7505,n7507);
not (n7505,n7506);
wire s0n7506,s1n7506,notn7506;
or (n7506,s0n7506,s1n7506);
not(notn7506,n746);
and (s0n7506,notn7506,1'b0);
and (s1n7506,n746,n7495);
not (n7507,n7439);
and (n7508,n7473,n7480);
wire s0n7509,s1n7509,notn7509;
or (n7509,s0n7509,s1n7509);
not(notn7509,n7312);
and (s0n7509,notn7509,1'b0);
and (s1n7509,n7312,n7510);
xor (n7510,n7511,n7520);
xor (n7511,n7512,n7513);
wire s0n7512,s1n7512,notn7512;
or (n7512,s0n7512,s1n7512);
not(notn7512,n6843);
and (s0n7512,notn7512,1'b0);
and (s1n7512,n6843,n7335);
xor (n7513,n7514,n7516);
xor (n7514,n7459,n7515);
wire s0n7515,s1n7515,notn7515;
or (n7515,s0n7515,s1n7515);
not(notn7515,n746);
and (s0n7515,notn7515,1'b0);
and (s1n7515,n746,n7450);
or (n7516,n7517,n7518,n7519);
and (n7517,n7334,n7343);
and (n7518,n7343,n7352);
and (n7519,n7334,n7352);
or (n7520,n7521,n7522,n7523);
and (n7521,n7323,n7332);
and (n7522,n7332,n7409);
and (n7523,n7323,n7409);
wire s0n7524,s1n7524,notn7524;
or (n7524,s0n7524,s1n7524);
not(notn7524,n7312);
and (s0n7524,notn7524,1'b0);
and (s1n7524,n7312,n7525);
xor (n7525,n7526,n7532);
xor (n7526,n7485,n7527);
xor (n7527,n7484,n7528);
or (n7528,n7529,n7530,n7531);
and (n7529,n7459,n7515);
and (n7530,n7515,n7516);
and (n7531,n7459,n7516);
or (n7532,n7533,n7534,n7535);
and (n7533,n7512,n7513);
and (n7534,n7513,n7520);
and (n7535,n7512,n7520);
wire s0n7536,s1n7536,notn7536;
or (n7536,s0n7536,s1n7536);
not(notn7536,n6895);
and (s0n7536,notn7536,1'b0);
and (s1n7536,n6895,n7537);
xor (n7537,n7538,n7540);
xor (n7538,n7489,n7539);
not (n7539,n7474);
or (n7540,n7541,n7677);
and (n7541,n7542,n7567);
xor (n7542,n7543,n7548);
nor (n7543,n7544,n7546);
and (n7544,n7545,n7461);
xor (n7545,n7492,n7494);
and (n7546,n7547,n7503);
not (n7547,n7545);
nand (n7548,n7549,n7560,n7564);
or (n7549,n7494,n7550);
not (n7550,n7551);
wire s0n7551,s1n7551,notn7551;
or (n7551,s0n7551,s1n7551);
not(notn7551,n820);
and (s0n7551,notn7551,1'b0);
and (s1n7551,n820,n7552);
wire s0n7552,s1n7552,notn7552;
or (n7552,s0n7552,s1n7552);
not(notn7552,n6972);
and (s0n7552,notn7552,n7553);
and (s1n7552,n6972,n7555);
wire s0n7553,s1n7553,notn7553;
or (n7553,s0n7553,s1n7553);
not(notn7553,n6971);
and (s0n7553,notn7553,1'b0);
and (s1n7553,n6971,n7554);
or (n7555,1'b0,n7556,n7557,n7558,n7559);
and (n7556,n1361,n903);
and (n7557,n2066,n949);
and (n7558,n5159,n901);
and (n7559,n7554,n960);
or (n7560,n7561,n7562);
nand (n7561,n6843,n7552);
not (n7562,n7563);
wire s0n7563,s1n7563,notn7563;
or (n7563,s0n7563,s1n7563);
not(notn7563,n746);
and (s0n7563,notn7563,1'b0);
and (s1n7563,n746,n7462);
not (n7564,n7565);
and (n7565,n7566,n7563);
wire s0n7566,s1n7566,notn7566;
or (n7566,s0n7566,s1n7566);
not(notn7566,n820);
and (s0n7566,notn7566,1'b0);
and (s1n7566,n820,n7495);
nand (n7567,n7568,n7676);
or (n7568,n7569,n7595);
not (n7569,n7570);
nand (n7570,n7571,n7575);
xor (n7571,n7572,n7573);
xor (n7572,n7566,n7563);
not (n7573,n7574);
not (n7574,n7561);
not (n7575,n7576);
nand (n7576,n7577,n7590,n7593);
or (n7577,n7578,n7588);
not (n7578,n7579);
wire s0n7579,s1n7579,notn7579;
or (n7579,s0n7579,s1n7579);
not(notn7579,n746);
and (s0n7579,notn7579,1'b0);
and (s1n7579,n746,n7580);
wire s0n7580,s1n7580,notn7580;
or (n7580,s0n7580,s1n7580);
not(notn7580,n6972);
and (s0n7580,notn7580,n7581);
and (s1n7580,n6972,n7583);
wire s0n7581,s1n7581,notn7581;
or (n7581,s0n7581,s1n7581);
not(notn7581,n6971);
and (s0n7581,notn7581,1'b0);
and (s1n7581,n6971,n7582);
or (n7583,1'b0,n7584,n7585,n7586,n7587);
and (n7584,n1468,n903);
and (n7585,n2131,n949);
and (n7586,n5230,n901);
and (n7587,n7582,n960);
not (n7588,n7589);
not (n7589,n7494);
or (n7590,n7573,n7591);
not (n7591,n7592);
wire s0n7592,s1n7592,notn7592;
or (n7592,s0n7592,s1n7592);
not(notn7592,n820);
and (s0n7592,notn7592,1'b0);
and (s1n7592,n820,n7580);
not (n7593,n7594);
and (n7594,n7551,n7506);
not (n7595,n7596);
or (n7596,n7597,n7675);
and (n7597,n7598,n7622);
xor (n7598,n7599,n7618);
nand (n7599,n7600,n7611,n7615);
or (n7600,n7561,n7601);
not (n7601,n7602);
wire s0n7602,s1n7602,notn7602;
or (n7602,s0n7602,s1n7602);
not(notn7602,n746);
and (s0n7602,notn7602,1'b0);
and (s1n7602,n746,n7603);
wire s0n7603,s1n7603,notn7603;
or (n7603,s0n7603,s1n7603);
not(notn7603,n6972);
and (s0n7603,notn7603,n7604);
and (s1n7603,n6972,n7606);
wire s0n7604,s1n7604,notn7604;
or (n7604,s0n7604,s1n7604);
not(notn7604,n6971);
and (s0n7604,notn7604,1'b0);
and (s1n7604,n6971,n7605);
or (n7606,1'b0,n7607,n7608,n7609,n7610);
and (n7607,n1575,n903);
and (n7608,n2196,n949);
and (n7609,n5301,n901);
and (n7610,n7605,n960);
or (n7611,n7612,n7613);
nand (n7612,n6843,n7580);
not (n7613,n7614);
wire s0n7614,s1n7614,notn7614;
or (n7614,s0n7614,s1n7614);
not(notn7614,n820);
and (s0n7614,notn7614,1'b0);
and (s1n7614,n820,n7603);
not (n7615,n7616);
and (n7616,n7592,n7617);
wire s0n7617,s1n7617,notn7617;
or (n7617,s0n7617,s1n7617);
not(notn7617,n746);
and (s0n7617,notn7617,1'b0);
and (s1n7617,n746,n7552);
nand (n7618,n7619,n7621);
or (n7619,n7612,n7620);
xor (n7620,n7551,n7506);
nand (n7621,n7620,n7612);
or (n7622,n7623,n7674);
and (n7623,n7624,n7648);
xor (n7624,n7625,n7645);
nand (n7625,n7626,n7640,n7643);
not (n7626,n7627);
and (n7627,n7628,n7630);
not (n7628,n7629);
nand (n7629,n6843,n7603);
not (n7630,n7631);
nand (n7631,n820,n7632);
wire s0n7632,s1n7632,notn7632;
or (n7632,s0n7632,s1n7632);
not(notn7632,n6972);
and (s0n7632,notn7632,n7633);
and (s1n7632,n6972,n7635);
wire s0n7633,s1n7633,notn7633;
or (n7633,s0n7633,s1n7633);
not(notn7633,n6971);
and (s0n7633,notn7633,1'b0);
and (s1n7633,n6971,n7634);
or (n7635,1'b0,n7636,n7637,n7638,n7639);
and (n7636,n1682,n903);
and (n7637,n2261,n949);
and (n7638,n5372,n901);
and (n7639,n7634,n960);
or (n7640,n7612,n7641);
not (n7641,n7642);
wire s0n7642,s1n7642,notn7642;
or (n7642,s0n7642,s1n7642);
not(notn7642,n746);
and (s0n7642,notn7642,1'b0);
and (s1n7642,n746,n7632);
not (n7643,n7644);
and (n7644,n7614,n7579);
xnor (n7645,n7646,n7647);
not (n7646,n7628);
xor (n7647,n7592,n7617);
or (n7648,n7649,n7673);
and (n7649,n7650,n7667);
xor (n7650,n7651,n7661);
nor (n7651,n7652,n7601);
nand (n7652,n6843,n7653);
wire s0n7653,s1n7653,notn7653;
or (n7653,s0n7653,s1n7653);
not(notn7653,n6972);
and (s0n7653,notn7653,n7654);
and (s1n7653,n6972,n7656);
wire s0n7654,s1n7654,notn7654;
or (n7654,s0n7654,s1n7654);
not(notn7654,n6971);
and (s0n7654,notn7654,1'b0);
and (s1n7654,n6971,n7655);
or (n7656,1'b0,n7657,n7658,n7659,n7660);
and (n7657,n1788,n903);
and (n7658,n2325,n949);
and (n7659,n5442,n901);
and (n7660,n7655,n960);
xnor (n7661,n7662,n7613);
nand (n7662,n7663,n7666);
or (n7663,n7664,n7578);
not (n7664,n7665);
nand (n7665,n6843,n7632);
nand (n7666,n7664,n7578);
nand (n7667,n7668,n7670);
or (n7668,n7669,n7631);
xnor (n7669,n7601,n7652);
not (n7670,n7671);
and (n7671,n7672,n7642);
wire s0n7672,s1n7672,notn7672;
or (n7672,s0n7672,s1n7672);
not(notn7672,n820);
and (s0n7672,notn7672,1'b0);
and (s1n7672,n820,n7653);
and (n7673,n7651,n7661);
and (n7674,n7625,n7645);
and (n7675,n7599,n7618);
or (n7676,n7571,n7575);
and (n7677,n7543,n7548);
and (n7678,n7318,n7524);
xor (n7679,n7680,n7692);
xor (n7680,n7681,n7691);
wire s0n7681,s1n7681,notn7681;
or (n7681,s0n7681,s1n7681);
not(notn7681,n7134);
and (s0n7681,notn7681,1'b0);
and (s1n7681,n7134,n7682);
or (n7682,n7683,n7685,n7690);
and (n7683,n7449,n7684);
and (n7684,n7484,n7528);
and (n7685,n7684,n7686);
or (n7686,n7687,n7688,n7689);
and (n7687,n7485,n7527);
and (n7688,n7527,n7532);
and (n7689,n7485,n7532);
and (n7690,n7449,n7686);
wire s0n7691,s1n7691,notn7691;
or (n7691,s0n7691,s1n7691);
not(notn7691,n6893);
and (s0n7691,notn7691,1'b0);
and (s1n7691,n6893,n7525);
wire s0n7692,s1n7692,notn7692;
or (n7692,s0n7692,s1n7692);
not(notn7692,n7312);
and (s0n7692,notn7692,1'b0);
and (s1n7692,n7312,n7693);
xor (n7693,n7694,n7686);
xor (n7694,n7449,n7684);
wire s0n7695,s1n7695,notn7695;
or (n7695,s0n7695,s1n7695);
not(notn7695,n673);
and (s0n7695,notn7695,1'b0);
and (s1n7695,n673,n7696);
or (n7696,n7697,n7717,n7755);
and (n7697,n7439,n7698);
and (n7698,n7479,n7699);
or (n7699,n7700,n7701,n7716);
and (n7700,n7461,n7493);
and (n7701,n7493,n7702);
or (n7702,n7565,n7703,n7715);
and (n7703,n7563,n7704);
or (n7704,n7594,n7705,n7714);
and (n7705,n7506,n7706);
or (n7706,n7616,n7707,n7713);
and (n7707,n7617,n7708);
or (n7708,n7644,n7709,n7711);
and (n7709,n7579,n7710);
or (n7710,n7711,n7712,n7671);
and (n7711,n7630,n7602);
and (n7712,n7602,n7671);
and (n7713,n7592,n7708);
and (n7714,n7551,n7706);
and (n7715,n7566,n7704);
and (n7716,n7461,n7702);
and (n7717,n7698,n7718);
or (n7718,n7719,n7721,n7754);
and (n7719,n7476,n7720);
xor (n7720,n7479,n7699);
and (n7721,n7720,n7722);
or (n7722,n7723,n7726,n7753);
and (n7723,n7589,n7724);
xor (n7724,n7725,n7702);
xor (n7725,n7461,n7493);
and (n7726,n7724,n7727);
or (n7727,n7728,n7730,n7752);
and (n7728,n7574,n7729);
xor (n7729,n7572,n7704);
and (n7730,n7729,n7731);
or (n7731,n7732,n7735,n7751);
and (n7732,n7733,n7734);
not (n7733,n7612);
xor (n7734,n7620,n7706);
and (n7735,n7734,n7736);
or (n7736,n7737,n7739,n7750);
and (n7737,n7628,n7738);
xor (n7738,n7647,n7708);
and (n7739,n7738,n7740);
or (n7740,n7741,n7744,n7749);
and (n7741,n7664,n7742);
xor (n7742,n7743,n7710);
xor (n7743,n7614,n7579);
and (n7744,n7742,n7745);
and (n7745,n7746,n7747);
not (n7746,n7652);
xor (n7747,n7748,n7671);
xor (n7748,n7630,n7602);
and (n7749,n7664,n7745);
and (n7750,n7628,n7740);
and (n7751,n7733,n7736);
and (n7752,n7574,n7731);
and (n7753,n7589,n7727);
and (n7754,n7476,n7722);
and (n7755,n7439,n7718);
or (n7756,n7757,n7888);
and (n7757,n7758,n7824);
xor (n7758,n7759,n7823);
or (n7759,n7760,n7822);
and (n7760,n7761,n7819);
xor (n7761,n7762,n7815);
wire s0n7762,s1n7762,notn7762;
or (n7762,s0n7762,s1n7762);
not(notn7762,n673);
and (s0n7762,notn7762,1'b0);
and (s1n7762,n673,n7763);
xor (n7763,n7764,n7783);
xor (n7764,n7765,n7766);
xor (n7765,n7163,n7160);
xor (n7766,n7162,n7767);
or (n7767,n7172,n7768,n7782);
and (n7768,n7174,n7769);
or (n7769,n7298,n7770,n7781);
and (n7770,n7198,n7771);
or (n7771,n7208,n7772,n7780);
and (n7772,n7210,n7773);
or (n7773,n7226,n7774,n7779);
and (n7774,n7228,n7775);
or (n7775,n7239,n7776,n7257);
and (n7776,n7241,n7777);
or (n7777,n7257,n7778,n7263);
and (n7778,n7259,n7263);
and (n7779,n7227,n7775);
and (n7780,n7209,n7773);
and (n7781,n7197,n7771);
and (n7782,n7173,n7769);
or (n7783,n7784,n7787,n7814);
and (n7784,n7785,n7786);
xor (n7785,n7297,n7294);
xor (n7786,n7296,n7769);
and (n7787,n7786,n7788);
or (n7788,n7789,n7792,n7813);
and (n7789,n7790,n7791);
xor (n7790,n7199,n7186);
xor (n7791,n7196,n7771);
and (n7792,n7791,n7793);
or (n7793,n7794,n7797,n7812);
and (n7794,n7795,n7796);
xor (n7795,n7217,n7214);
xor (n7796,n7216,n7773);
and (n7797,n7796,n7798);
or (n7798,n7799,n7802,n7811);
and (n7799,n7800,n7801);
xor (n7800,n7244,n7238);
xor (n7801,n7243,n7775);
and (n7802,n7801,n7803);
or (n7803,n7804,n7807,n7810);
and (n7804,n7805,n7806);
xor (n7805,n7279,n7281);
xor (n7806,n7280,n7777);
and (n7807,n7806,n7808);
and (n7808,n7274,n7809);
xor (n7809,n7275,n7263);
and (n7810,n7805,n7808);
and (n7811,n7800,n7803);
and (n7812,n7795,n7798);
and (n7813,n7790,n7793);
and (n7814,n7785,n7788);
wire s0n7815,s1n7815,notn7815;
or (n7815,s0n7815,s1n7815);
not(notn7815,n6895);
and (s0n7815,notn7815,1'b0);
and (s1n7815,n6895,n7816);
xor (n7816,n7817,n7180);
nor (n7817,n7818,n7302);
not (n7818,n7291);
wire s0n7819,s1n7819,notn7819;
or (n7819,s0n7819,s1n7819);
not(notn7819,n7312);
and (s0n7819,notn7819,1'b0);
and (s1n7819,n7312,n7820);
xor (n7820,n7821,n7091);
xor (n7821,n7085,n7088);
and (n7822,n7762,n7815);
xor (n7823,n7317,n7536);
and (n7824,n7825,n7885);
xor (n7825,n7826,n7829);
wire s0n7826,s1n7826,notn7826;
or (n7826,s0n7826,s1n7826);
not(notn7826,n6893);
and (s0n7826,notn7826,1'b0);
and (s1n7826,n6893,n7827);
xor (n7827,n7828,n7099);
xor (n7828,n7093,n7096);
or (n7829,n7830,n7884);
and (n7830,n7831,n7858);
xor (n7831,n7832,n7835);
wire s0n7832,s1n7832,notn7832;
or (n7832,s0n7832,s1n7832);
not(notn7832,n6895);
and (s0n7832,notn7832,1'b0);
and (s1n7832,n6895,n7833);
xor (n7833,n7834,n7731);
xor (n7834,n7574,n7729);
and (n7835,n7836,n7857);
or (n7836,n7837,n7856);
and (n7837,n7838,n7847);
xor (n7838,n7839,n7840);
and (n7839,n7576,n27);
nor (n7840,n6944,n7841);
nor (n7841,n7353,n7842);
nor (n7842,n7843,n7846);
and (n7843,n7844,n7845);
not (n7844,n7355);
not (n7845,n7354);
not (n7846,n7411);
nor (n7847,n7848,n6944);
nor (n7848,n7849,n7854);
and (n7849,n7850,n7334);
not (n7850,n7851);
xor (n7851,n7852,n7853);
not (n7852,n7323);
not (n7853,n7343);
and (n7854,n7851,n7855);
not (n7855,n7334);
and (n7856,n7839,n7840);
and (n7857,n7543,n27);
or (n7858,n7859,n7883);
and (n7859,n7860,n7881);
xor (n7860,n7861,n7864);
wire s0n7861,s1n7861,notn7861;
or (n7861,s0n7861,s1n7861);
not(notn7861,n7312);
and (s0n7861,notn7861,1'b0);
and (s1n7861,n7312,n7862);
xor (n7862,n7863,n7415);
xor (n7863,n7411,n7412);
xor (n7864,n7865,n7873);
xor (n7865,n7866,n7872);
and (n7866,n7867,n27);
nand (n7867,n7868,n7870,n7871);
or (n7868,n7869,n7845);
not (n7869,n7512);
not (n7870,n7517);
or (n7871,n7852,n7853);
and (n7872,n7548,n27);
and (n7873,n7874,n27);
nor (n7874,n7875,n7878);
and (n7875,n7876,n7459);
xor (n7876,n7877,n7869);
not (n7877,n7515);
and (n7878,n7879,n7880);
not (n7879,n7876);
not (n7880,n7459);
wire s0n7881,s1n7881,notn7881;
or (n7881,s0n7881,s1n7881);
not(notn7881,n6895);
and (s0n7881,notn7881,1'b0);
and (s1n7881,n6895,n7882);
xor (n7882,n7598,n7622);
and (n7883,n7861,n7864);
and (n7884,n7832,n7835);
wire s0n7885,s1n7885,notn7885;
or (n7885,s0n7885,s1n7885);
not(notn7885,n7134);
and (s0n7885,notn7885,1'b0);
and (s1n7885,n7134,n7886);
xor (n7886,n7887,n7083);
xor (n7887,n7078,n7081);
and (n7888,n7759,n7823);
xor (n7889,n7890,n7921);
xor (n7890,n7891,n7904);
xor (n7891,n7892,n7901);
xor (n7892,n7893,n7894);
wire s0n7893,s1n7893,notn7893;
or (n7893,s0n7893,s1n7893);
not(notn7893,n6893);
and (s0n7893,notn7893,1'b0);
and (s1n7893,n6893,n7886);
and (n7894,n7895,n7898);
or (n7895,n7896,n7897);
and (n7896,n7435,n7470);
and (n7897,n7436,n7460);
or (n7898,n7899,n7900);
and (n7899,n7437,n7458);
and (n7900,n7438,n7448);
wire s0n7901,s1n7901,notn7901;
or (n7901,s0n7901,s1n7901);
not(notn7901,n6895);
and (s0n7901,notn7901,1'b0);
and (s1n7901,n6895,n7902);
xor (n7902,n7903,n7718);
xor (n7903,n7439,n7698);
or (n7904,n7905,n7920);
and (n7905,n7906,n7919);
xor (n7906,n7907,n7918);
or (n7907,n7908,n7917);
and (n7908,n7909,n7916);
xor (n7909,n7910,n7911);
xor (n7910,n7319,n7509);
and (n7911,n7912,n7915);
xor (n7912,n7913,n7914);
wire s0n7913,s1n7913,notn7913;
or (n7913,s0n7913,s1n7913);
not(notn7913,n6893);
and (s0n7913,notn7913,1'b0);
and (s1n7913,n6893,n7862);
wire s0n7914,s1n7914,notn7914;
or (n7914,s0n7914,s1n7914);
not(notn7914,n7312);
and (s0n7914,notn7914,1'b0);
and (s1n7914,n7312,n7321);
wire s0n7915,s1n7915,notn7915;
or (n7915,s0n7915,s1n7915);
not(notn7915,n7134);
and (s0n7915,notn7915,1'b0);
and (s1n7915,n7134,n7510);
wire s0n7916,s1n7916,notn7916;
or (n7916,s0n7916,s1n7916);
not(notn7916,n673);
and (s0n7916,notn7916,1'b0);
and (s1n7916,n673,n7537);
and (n7917,n7910,n7911);
wire s0n7918,s1n7918,notn7918;
or (n7918,s0n7918,s1n7918);
not(notn7918,n6895);
and (s0n7918,notn7918,1'b0);
and (s1n7918,n6895,n7763);
wire s0n7919,s1n7919,notn7919;
or (n7919,s0n7919,s1n7919);
not(notn7919,n7312);
and (s0n7919,notn7919,1'b0);
and (s1n7919,n7312,n7886);
and (n7920,n7907,n7918);
or (n7921,n7922,n7931);
and (n7922,n7923,n7930);
xor (n7923,n7924,n7925);
wire s0n7924,s1n7924,notn7924;
or (n7924,s0n7924,s1n7924);
not(notn7924,n27);
and (s0n7924,notn7924,1'b0);
and (s1n7924,n27,n6967);
wire s0n7925,s1n7925,notn7925;
or (n7925,s0n7925,s1n7925);
not(notn7925,n27);
and (s0n7925,notn7925,1'b0);
and (s1n7925,n27,n7926);
xor (n7926,n7927,n7928);
wire s0n7927,s1n7927,notn7927;
or (n7927,s0n7927,s1n7927);
not(notn7927,n6841);
and (s0n7927,notn7927,1'b0);
and (s1n7927,n6841,n7149);
or (n7928,n7929,n7175);
and (n7929,n7137,n7176);
wire s0n7930,s1n7930,notn7930;
or (n7930,s0n7930,s1n7930);
not(notn7930,n7134);
and (s0n7930,notn7930,1'b0);
and (s1n7930,n7134,n7310);
and (n7931,n7924,n7925);
or (n7932,n7933,n8103);
and (n7933,n7934,n7974);
xor (n7934,n7935,n7936);
xor (n7935,n7758,n7824);
or (n7936,n7937,n7973);
and (n7937,n7938,n7947);
xor (n7938,n7939,n7940);
xor (n7939,n7825,n7885);
or (n7940,n7941,n7946);
and (n7941,n7942,n7945);
xor (n7942,n7943,n7944);
wire s0n7943,s1n7943,notn7943;
or (n7943,s0n7943,s1n7943);
not(notn7943,n7312);
and (s0n7943,notn7943,1'b0);
and (s1n7943,n7312,n7827);
xor (n7944,n7831,n7858);
wire s0n7945,s1n7945,notn7945;
or (n7945,s0n7945,s1n7945);
not(notn7945,n27);
and (s0n7945,notn7945,1'b0);
and (s1n7945,n27,n7763);
and (n7946,n7943,n7944);
or (n7947,n7948,n7972);
and (n7948,n7949,n7971);
xor (n7949,n7950,n7951);
wire s0n7950,s1n7950,notn7950;
or (n7950,s0n7950,s1n7950);
not(notn7950,n673);
and (s0n7950,notn7950,1'b0);
and (s1n7950,n673,n7816);
or (n7951,n7952,n7970);
and (n7952,n7953,n7967);
xor (n7953,n7954,n7959);
xor (n7954,n7955,n7956);
xor (n7955,n7836,n7857);
wire s0n7956,s1n7956,notn7956;
or (n7956,s0n7956,s1n7956);
not(notn7956,n6893);
and (s0n7956,notn7956,1'b0);
and (s1n7956,n6893,n7957);
xor (n7957,n7958,n7421);
xor (n7958,n7417,n7418);
and (n7959,n7960,n7965);
xor (n7960,n7961,n7962);
xor (n7961,n7838,n7847);
wire s0n7962,s1n7962,notn7962;
or (n7962,s0n7962,s1n7962);
not(notn7962,n6893);
and (s0n7962,notn7962,1'b0);
and (s1n7962,n6893,n7963);
xor (n7963,n7964,n7427);
xor (n7964,n7423,n7424);
wire s0n7965,s1n7965,notn7965;
or (n7965,s0n7965,s1n7965);
not(notn7965,n6895);
and (s0n7965,notn7965,1'b0);
and (s1n7965,n6895,n7966);
xor (n7966,n7624,n7648);
wire s0n7967,s1n7967,notn7967;
or (n7967,s0n7967,s1n7967);
not(notn7967,n6893);
and (s0n7967,notn7967,1'b0);
and (s1n7967,n6893,n7968);
xor (n7968,n7969,n7115);
xor (n7969,n7109,n7112);
and (n7970,n7954,n7959);
wire s0n7971,s1n7971,notn7971;
or (n7971,s0n7971,s1n7971);
not(notn7971,n7134);
and (s0n7971,notn7971,1'b0);
and (s1n7971,n7134,n7820);
and (n7972,n7950,n7951);
and (n7973,n7939,n7940);
or (n7974,n7975,n8102);
and (n7975,n7976,n8079);
xor (n7976,n7977,n8078);
or (n7977,n7978,n8077);
and (n7978,n7979,n8076);
xor (n7979,n7980,n8004);
or (n7980,n7981,n8003);
and (n7981,n7982,n8000);
xor (n7982,n7983,n7984);
xor (n7983,n7860,n7881);
or (n7984,n7985,n7999);
and (n7985,n7986,n7998);
xor (n7986,n7987,n7988);
wire s0n7987,s1n7987,notn7987;
or (n7987,s0n7987,s1n7987);
not(notn7987,n7134);
and (s0n7987,notn7987,1'b0);
and (s1n7987,n7134,n7862);
or (n7988,n7989,n7997);
and (n7989,n7990,n7996);
xor (n7990,n7991,n7992);
and (n7991,n7618,n27);
and (n7992,n7993,n27);
nand (n7993,n7994,n7995);
or (n7994,n7846,n7413);
nand (n7995,n7413,n7846);
wire s0n7996,s1n7996,notn7996;
or (n7996,s0n7996,s1n7996);
not(notn7996,n7312);
and (s0n7996,notn7996,1'b0);
and (s1n7996,n7312,n7963);
and (n7997,n7991,n7992);
wire s0n7998,s1n7998,notn7998;
or (n7998,s0n7998,s1n7998);
not(notn7998,n673);
and (s0n7998,notn7998,1'b0);
and (s1n7998,n673,n7882);
and (n7999,n7987,n7988);
wire s0n8000,s1n8000,notn8000;
or (n8000,s0n8000,s1n8000);
not(notn8000,n6895);
and (s0n8000,notn8000,1'b0);
and (s1n8000,n6895,n8001);
xor (n8001,n8002,n7798);
xor (n8002,n7795,n7796);
and (n8003,n7983,n7984);
or (n8004,n8005,n8075);
and (n8005,n8006,n8072);
xor (n8006,n8007,n8026);
xor (n8007,n8008,n8025);
xor (n8008,n8009,n8010);
wire s0n8009,s1n8009,notn8009;
or (n8009,s0n8009,s1n8009);
not(notn8009,n7134);
and (s0n8009,notn8009,1'b0);
and (s1n8009,n7134,n7321);
or (n8010,n8011,n8024);
and (n8011,n8012,n8023);
xor (n8012,n8013,n8022);
or (n8013,n8014,n8021);
and (n8014,n8015,n27);
nand (n8015,n8016,n8018,n8020);
or (n8016,n7852,n8017);
not (n8017,n7394);
or (n8018,n7846,n8019);
not (n8019,n7372);
not (n8020,n7358);
and (n8021,n7599,n27);
nor (n8022,n7571,n6944);
wire s0n8023,s1n8023,notn8023;
or (n8023,s0n8023,s1n8023);
not(notn8023,n7312);
and (s0n8023,notn8023,1'b0);
and (s1n8023,n7312,n7957);
and (n8024,n8013,n8022);
wire s0n8025,s1n8025,notn8025;
or (n8025,s0n8025,s1n8025);
not(notn8025,n673);
and (s0n8025,notn8025,1'b0);
and (s1n8025,n673,n7833);
and (n8026,n8027,n8071);
xor (n8027,n8028,n8065);
or (n8028,n8029,n8064);
and (n8029,n8030,n8062);
xor (n8030,n8031,n8044);
and (n8031,n8032,n8043);
xor (n8032,n8033,n8041);
and (n8033,n8034,n8038);
nor (n8034,n8035,n7646);
not (n8035,n8036);
wire s0n8036,s1n8036,notn8036;
or (n8036,s0n8036,s1n8036);
not(notn8036,n27);
and (s0n8036,notn8036,1'b0);
and (s1n8036,n27,n8037);
wire s0n8037,s1n8037,notn8037;
or (n8037,s0n8037,s1n8037);
not(notn8037,n746);
and (s0n8037,notn8037,1'b0);
and (s1n8037,n746,n7653);
and (n8038,n8039,n27);
nor (n8039,n8040,n8017);
not (n8040,n7428);
wire s0n8041,s1n8041,notn8041;
or (n8041,s0n8041,s1n8041);
not(notn8041,n6893);
and (s0n8041,notn8041,1'b0);
and (s1n8041,n6893,n8042);
xor (n8042,n7397,n7406);
and (n8043,n7645,n27);
or (n8044,n8045,n8061);
and (n8045,n8046,n8055);
xor (n8046,n8047,n8054);
and (n8047,n8048,n27);
nand (n8048,n8049,n8051,n8053);
or (n8049,n8050,n8019);
not (n8050,n7423);
or (n8051,n7846,n8052);
not (n8052,n7406);
not (n8053,n7371);
and (n8054,n7625,n27);
and (n8055,n8056,n27);
xor (n8056,n8057,n8058);
not (n8057,n7359);
xnor (n8058,n8059,n8060);
not (n8059,n7417);
not (n8060,n7368);
and (n8061,n8047,n8054);
wire s0n8062,s1n8062,notn8062;
or (n8062,s0n8062,s1n8062);
not(notn8062,n6895);
and (s0n8062,notn8062,1'b0);
and (s1n8062,n6895,n8063);
xor (n8063,n7650,n7667);
and (n8064,n8031,n8044);
and (n8065,n8066,n8070);
xor (n8066,n8067,n8068);
wire s0n8067,s1n8067,notn8067;
or (n8067,s0n8067,s1n8067);
not(notn8067,n673);
and (s0n8067,notn8067,1'b0);
and (s1n8067,n673,n7966);
wire s0n8068,s1n8068,notn8068;
or (n8068,s0n8068,s1n8068);
not(notn8068,n6893);
and (s0n8068,notn8068,1'b0);
and (s1n8068,n6893,n8069);
xor (n8069,n7428,n7429);
wire s0n8070,s1n8070,notn8070;
or (n8070,s0n8070,s1n8070);
not(notn8070,n7134);
and (s0n8070,notn8070,1'b0);
and (s1n8070,n7134,n7957);
xor (n8071,n7960,n7965);
wire s0n8072,s1n8072,notn8072;
or (n8072,s0n8072,s1n8072);
not(notn8072,n7312);
and (s0n8072,notn8072,1'b0);
and (s1n8072,n7312,n8073);
xor (n8073,n8074,n7107);
xor (n8074,n7101,n7104);
and (n8075,n8007,n8026);
wire s0n8076,s1n8076,notn8076;
or (n8076,s0n8076,s1n8076);
not(notn8076,n27);
and (s0n8076,notn8076,1'b0);
and (s1n8076,n27,n7886);
and (n8077,n7980,n8004);
xor (n8078,n7761,n7819);
xor (n8079,n8080,n8101);
xor (n8080,n8081,n8082);
and (n8081,n7136,n27);
xor (n8082,n8083,n8099);
xor (n8083,n8084,n8085);
wire s0n8084,s1n8084,notn8084;
or (n8084,s0n8084,s1n8084);
not(notn8084,n7134);
and (s0n8084,notn8084,1'b0);
and (s1n8084,n7134,n7525);
or (n8085,n8086,n8098);
and (n8086,n8087,n8095);
xor (n8087,n8088,n8089);
xor (n8088,n7472,n7488);
and (n8089,n8090,n27);
nand (n8090,n8091,n8093);
or (n8091,n8092,n7880);
and (n8092,n7877,n7869);
or (n8093,n7844,n8094);
not (n8094,n7449);
or (n8095,n8096,n8097);
and (n8096,n7865,n7873);
and (n8097,n7866,n7872);
and (n8098,n8088,n8089);
wire s0n8099,s1n8099,notn8099;
or (n8099,s0n8099,s1n8099);
not(notn8099,n6895);
and (s0n8099,notn8099,1'b0);
and (s1n8099,n6895,n8100);
xor (n8100,n7542,n7567);
wire s0n8101,s1n8101,notn8101;
or (n8101,s0n8101,s1n8101);
not(notn8101,n27);
and (s0n8101,notn8101,1'b0);
and (s1n8101,n27,n7310);
and (n8102,n7977,n8078);
and (n8103,n7935,n7936);
and (n8104,n6962,n7889);
xor (n8105,n8106,n8129);
xor (n8106,n8107,n8110);
or (n8107,n8108,n8109);
and (n8108,n7890,n7921);
and (n8109,n7891,n7904);
and (n8110,n8111,n8122);
xor (n8111,n8112,n8121);
or (n8112,n8113,n8120);
and (n8113,n8114,n8119);
xor (n8114,n8115,n8116);
wire s0n8115,s1n8115,notn8115;
or (n8115,s0n8115,s1n8115);
not(notn8115,n7134);
and (s0n8115,notn8115,1'b0);
and (s1n8115,n7134,n7693);
xor (n8116,n8117,n8118);
xor (n8117,n7895,n7898);
wire s0n8118,s1n8118,notn8118;
or (n8118,s0n8118,s1n8118);
not(notn8118,n6893);
and (s0n8118,notn8118,1'b0);
and (s1n8118,n6893,n7510);
wire s0n8119,s1n8119,notn8119;
or (n8119,s0n8119,s1n8119);
not(notn8119,n673);
and (s0n8119,notn8119,1'b0);
and (s1n8119,n673,n7136);
and (n8120,n8115,n8116);
wire s0n8121,s1n8121,notn8121;
or (n8121,s0n8121,s1n8121);
not(notn8121,n673);
and (s0n8121,notn8121,1'b0);
and (s1n8121,n673,n7926);
and (n8122,n8123,n8128);
xor (n8123,n8124,n8125);
wire s0n8124,s1n8124,notn8124;
or (n8124,s0n8124,s1n8124);
not(notn8124,n6893);
and (s0n8124,notn8124,1'b0);
and (s1n8124,n6893,n7820);
or (n8125,n8126,n8127);
and (n8126,n8083,n8099);
and (n8127,n8084,n8085);
wire s0n8128,s1n8128,notn8128;
or (n8128,s0n8128,s1n8128);
not(notn8128,n673);
and (s0n8128,notn8128,1'b0);
and (s1n8128,n673,n7902);
xor (n8129,n8130,n8133);
xor (n8130,n8131,n8132);
and (n8131,n7892,n7901);
and (n8132,n7680,n7692);
or (n8133,n8134,n8135);
and (n8134,n6965,n7309);
and (n8135,n6966,n7135);
xor (n8136,n8137,n8156);
xor (n8137,n8138,n8141);
or (n8138,n8139,n8140);
and (n8139,n6963,n7756);
and (n8140,n6964,n7313);
xor (n8141,n8142,n8151);
xor (n8142,n8143,n8146);
or (n8143,n8144,n8145);
and (n8144,n7314,n7695);
and (n8145,n7315,n7679);
xor (n8146,n8147,n8150);
xor (n8147,n8148,n8149);
wire s0n8148,s1n8148,notn8148;
or (n8148,s0n8148,s1n8148);
not(notn8148,n6893);
and (s0n8148,notn8148,1'b0);
and (s1n8148,n6893,n7693);
wire s0n8149,s1n8149,notn8149;
or (n8149,s0n8149,s1n8149);
not(notn8149,n7312);
and (s0n8149,notn8149,1'b0);
and (s1n8149,n7312,n7682);
wire s0n8150,s1n8150,notn8150;
or (n8150,s0n8150,s1n8150);
not(notn8150,n6893);
and (s0n8150,notn8150,1'b0);
and (s1n8150,n6893,n7310);
xor (n8151,n8152,n8155);
xor (n8152,n8153,n8154);
wire s0n8153,s1n8153,notn8153;
or (n8153,s0n8153,s1n8153);
not(notn8153,n6895);
and (s0n8153,notn8153,1'b0);
and (s1n8153,n6895,n7926);
wire s0n8154,s1n8154,notn8154;
or (n8154,s0n8154,s1n8154);
not(notn8154,n6895);
and (s0n8154,notn8154,1'b0);
and (s1n8154,n6895,n7696);
wire s0n8155,s1n8155,notn8155;
or (n8155,s0n8155,s1n8155);
not(notn8155,n7312);
and (s0n8155,notn8155,1'b0);
and (s1n8155,n7312,n6967);
or (n8156,n8157,n8198);
and (n8157,n8158,n8169);
xor (n8158,n8159,n8168);
or (n8159,n8160,n8167);
and (n8160,n8161,n8164);
xor (n8161,n8162,n8163);
xor (n8162,n7906,n7919);
xor (n8163,n8114,n8119);
or (n8164,n8165,n8166);
and (n8165,n8080,n8101);
and (n8166,n8081,n8082);
and (n8167,n8162,n8163);
xor (n8168,n8111,n8122);
or (n8169,n8170,n8197);
and (n8170,n8171,n8196);
xor (n8171,n8172,n8173);
xor (n8172,n8123,n8128);
or (n8173,n8174,n8195);
and (n8174,n8175,n8186);
xor (n8175,n8176,n8177);
xor (n8176,n7909,n7916);
or (n8177,n8178,n8185);
and (n8178,n8179,n8184);
xor (n8179,n8180,n8183);
or (n8180,n8181,n8182);
and (n8181,n8008,n8025);
and (n8182,n8009,n8010);
xor (n8183,n8087,n8095);
wire s0n8184,s1n8184,notn8184;
or (n8184,s0n8184,s1n8184);
not(notn8184,n673);
and (s0n8184,notn8184,1'b0);
and (s1n8184,n673,n8100);
and (n8185,n8180,n8183);
or (n8186,n8187,n8194);
and (n8187,n8188,n8191);
xor (n8188,n8189,n8190);
wire s0n8189,s1n8189,notn8189;
or (n8189,s0n8189,s1n8189);
not(notn8189,n6893);
and (s0n8189,notn8189,1'b0);
and (s1n8189,n6893,n8073);
xor (n8190,n7912,n7915);
wire s0n8191,s1n8191,notn8191;
or (n8191,s0n8191,s1n8191);
not(notn8191,n6895);
and (s0n8191,notn8191,1'b0);
and (s1n8191,n6895,n8192);
xnor (n8192,n7231,n8193);
nand (n8193,n7183,n7290);
and (n8194,n8189,n8190);
and (n8195,n8176,n8177);
xor (n8196,n7923,n7930);
and (n8197,n8172,n8173);
and (n8198,n8159,n8168);
or (n8199,n8200,n8271);
and (n8200,n8201,n8270);
xor (n8201,n8202,n8203);
xor (n8202,n8158,n8169);
or (n8203,n8204,n8269);
and (n8204,n8205,n8208);
xor (n8205,n8206,n8207);
xor (n8206,n8171,n8196);
xor (n8207,n8161,n8164);
or (n8208,n8209,n8268);
and (n8209,n8210,n8255);
xor (n8210,n8211,n8254);
or (n8211,n8212,n8253);
and (n8212,n8213,n8216);
xor (n8213,n8214,n8215);
xor (n8214,n8188,n8191);
xor (n8215,n8179,n8184);
or (n8216,n8217,n8252);
and (n8217,n8218,n8251);
xor (n8218,n8219,n8242);
or (n8219,n8220,n8241);
and (n8220,n8221,n8240);
xor (n8221,n8222,n8223);
xor (n8222,n7986,n7998);
or (n8223,n8224,n8239);
and (n8224,n8225,n8231);
xor (n8225,n8226,n8227);
xor (n8226,n7990,n7996);
nand (n8227,n8228,n8013);
or (n8228,n8229,n8230);
not (n8229,n8021);
not (n8230,n8014);
or (n8231,n8232,n8238);
and (n8232,n8233,n8237);
xor (n8233,n8234,n8235);
wire s0n8234,s1n8234,notn8234;
or (n8234,s0n8234,s1n8234);
not(notn8234,n7312);
and (s0n8234,notn8234,1'b0);
and (s1n8234,n7312,n8069);
wire s0n8235,s1n8235,notn8235;
or (n8235,s0n8235,s1n8235);
not(notn8235,n6895);
and (s0n8235,notn8235,1'b0);
and (s1n8235,n6895,n8236);
xor (n8236,n7746,n7747);
wire s0n8237,s1n8237,notn8237;
or (n8237,s0n8237,s1n8237);
not(notn8237,n7134);
and (s0n8237,notn8237,1'b0);
and (s1n8237,n7134,n7963);
and (n8238,n8234,n8235);
and (n8239,n8226,n8227);
wire s0n8240,s1n8240,notn8240;
or (n8240,s0n8240,s1n8240);
not(notn8240,n7312);
and (s0n8240,notn8240,1'b0);
and (s1n8240,n7312,n7968);
and (n8241,n8222,n8223);
and (n8242,n8243,n8248);
xor (n8243,n8244,n8247);
wire s0n8244,s1n8244,notn8244;
or (n8244,s0n8244,s1n8244);
not(notn8244,n6893);
and (s0n8244,notn8244,1'b0);
and (s1n8244,n6893,n8245);
xor (n8245,n8246,n7123);
xor (n8246,n7117,n7120);
xor (n8247,n8012,n8023);
wire s0n8248,s1n8248,notn8248;
or (n8248,s0n8248,s1n8248);
not(notn8248,n6895);
and (s0n8248,notn8248,1'b0);
and (s1n8248,n6895,n8249);
xor (n8249,n8250,n7803);
xor (n8250,n7800,n7801);
and (n8251,n7816,n27);
and (n8252,n8219,n8242);
and (n8253,n8214,n8215);
xor (n8254,n8175,n8186);
or (n8255,n8256,n8267);
and (n8256,n8257,n8266);
xor (n8257,n8258,n8259);
xor (n8258,n7942,n7945);
or (n8259,n8260,n8265);
and (n8260,n8261,n8264);
xor (n8261,n8262,n8263);
wire s0n8262,s1n8262,notn8262;
or (n8262,s0n8262,s1n8262);
not(notn8262,n7134);
and (s0n8262,notn8262,1'b0);
and (s1n8262,n7134,n7827);
wire s0n8263,s1n8263,notn8263;
or (n8263,s0n8263,s1n8263);
not(notn8263,n673);
and (s0n8263,notn8263,1'b0);
and (s1n8263,n673,n8192);
wire s0n8264,s1n8264,notn8264;
or (n8264,s0n8264,s1n8264);
not(notn8264,n27);
and (s0n8264,notn8264,1'b0);
and (s1n8264,n27,n7820);
and (n8265,n8262,n8263);
xor (n8266,n7949,n7971);
and (n8267,n8258,n8259);
and (n8268,n8211,n8254);
and (n8269,n8206,n8207);
xor (n8270,n6961,n7932);
and (n8271,n8202,n8203);
or (n8272,n8273,n8735);
and (n8273,n8274,n8344);
xor (n8274,n8275,n8276);
xor (n8275,n8201,n8270);
or (n8276,n8277,n8343);
and (n8277,n8278,n8342);
xor (n8278,n8279,n8280);
xor (n8279,n7934,n7974);
or (n8280,n8281,n8341);
and (n8281,n8282,n8285);
xor (n8282,n8283,n8284);
xor (n8283,n7938,n7947);
xor (n8284,n7976,n8079);
or (n8285,n8286,n8340);
and (n8286,n8287,n8320);
xor (n8287,n8288,n8289);
xor (n8288,n7979,n8076);
or (n8289,n8290,n8319);
and (n8290,n8291,n8294);
xor (n8291,n8292,n8293);
xor (n8292,n7982,n8000);
xor (n8293,n7953,n7967);
or (n8294,n8295,n8318);
and (n8295,n8296,n8317);
xor (n8296,n8297,n8316);
and (n8297,n8298,n8299);
xor (n8298,n8030,n8062);
or (n8299,n8300,n8315);
and (n8300,n8301,n8314);
xor (n8301,n8302,n8313);
or (n8302,n8303,n8312);
and (n8303,n8304,n8311);
xor (n8304,n8305,n8307);
wire s0n8305,s1n8305,notn8305;
or (n8305,s0n8305,s1n8305);
not(notn8305,n6895);
and (s0n8305,notn8305,1'b0);
and (s1n8305,n6895,n8306);
xor (n8306,n7672,n7642);
and (n8307,n8308,n8309);
wire s0n8308,s1n8308,notn8308;
or (n8308,s0n8308,s1n8308);
not(notn8308,n6895);
and (s0n8308,notn8308,1'b0);
and (s1n8308,n6895,n8037);
wire s0n8309,s1n8309,notn8309;
or (n8309,s0n8309,s1n8309);
not(notn8309,n6895);
and (s0n8309,notn8309,1'b0);
and (s1n8309,n6895,n8310);
wire s0n8310,s1n8310,notn8310;
or (n8310,s0n8310,s1n8310);
not(notn8310,n746);
and (s0n8310,notn8310,1'b0);
and (s1n8310,n746,n7265);
and (n8311,n7661,n27);
and (n8312,n8305,n8307);
xor (n8313,n8046,n8055);
wire s0n8314,s1n8314,notn8314;
or (n8314,s0n8314,s1n8314);
not(notn8314,n673);
and (s0n8314,notn8314,1'b0);
and (s1n8314,n673,n8063);
and (n8315,n8302,n8313);
wire s0n8316,s1n8316,notn8316;
or (n8316,s0n8316,s1n8316);
not(notn8316,n7134);
and (s0n8316,notn8316,1'b0);
and (s1n8316,n7134,n8073);
wire s0n8317,s1n8317,notn8317;
or (n8317,s0n8317,s1n8317);
not(notn8317,n673);
and (s0n8317,notn8317,1'b0);
and (s1n8317,n673,n8001);
and (n8318,n8297,n8316);
and (n8319,n8292,n8293);
or (n8320,n8321,n8339);
and (n8321,n8322,n8338);
xor (n8322,n8323,n8324);
xor (n8323,n8006,n8072);
or (n8324,n8325,n8337);
and (n8325,n8326,n8336);
xor (n8326,n8327,n8335);
or (n8327,n8328,n8334);
and (n8328,n8329,n8333);
xor (n8329,n8330,n8331);
xor (n8330,n8066,n8070);
wire s0n8331,s1n8331,notn8331;
or (n8331,s0n8331,s1n8331);
not(notn8331,n6895);
and (s0n8331,notn8331,1'b0);
and (s1n8331,n6895,n8332);
xor (n8332,n7256,n7277);
wire s0n8333,s1n8333,notn8333;
or (n8333,s0n8333,s1n8333);
not(notn8333,n7312);
and (s0n8333,notn8333,1'b0);
and (s1n8333,n7312,n8245);
and (n8334,n8330,n8331);
xor (n8335,n8027,n8071);
wire s0n8336,s1n8336,notn8336;
or (n8336,s0n8336,s1n8336);
not(notn8336,n27);
and (s0n8336,notn8336,1'b0);
and (s1n8336,n27,n7827);
and (n8337,n8327,n8335);
xor (n8338,n8261,n8264);
and (n8339,n8323,n8324);
and (n8340,n8288,n8289);
and (n8341,n8283,n8284);
xor (n8342,n8205,n8208);
and (n8343,n8279,n8280);
or (n8344,n8345,n8734);
and (n8345,n8346,n8472);
xor (n8346,n8347,n8348);
xor (n8347,n8278,n8342);
or (n8348,n8349,n8471);
and (n8349,n8350,n8470);
xor (n8350,n8351,n8352);
xor (n8351,n8210,n8255);
or (n8352,n8353,n8469);
and (n8353,n8354,n8468);
xor (n8354,n8355,n8356);
xor (n8355,n8213,n8216);
or (n8356,n8357,n8467);
and (n8357,n8358,n8403);
xor (n8358,n8359,n8402);
or (n8359,n8360,n8401);
and (n8360,n8361,n8364);
xor (n8361,n8362,n8363);
xor (n8362,n8243,n8248);
and (n8363,n8192,n27);
or (n8364,n8365,n8400);
and (n8365,n8366,n8399);
xor (n8366,n8367,n8381);
or (n8367,n8368,n8380);
and (n8368,n8369,n8378);
xor (n8369,n8370,n8372);
wire s0n8370,s1n8370,notn8370;
or (n8370,s0n8370,s1n8370);
not(notn8370,n6895);
and (s0n8370,notn8370,1'b0);
and (s1n8370,n6895,n8371);
xor (n8371,n7262,n7275);
and (n8372,n8373,n8377);
xor (n8373,n8374,n8375);
xor (n8374,n8034,n8038);
wire s0n8375,s1n8375,notn8375;
or (n8375,s0n8375,s1n8375);
not(notn8375,n6893);
and (s0n8375,notn8375,1'b0);
and (s1n8375,n6893,n8376);
wire s0n8376,s1n8376,notn8376;
or (n8376,s0n8376,s1n8376);
not(notn8376,n746);
and (s0n8376,notn8376,1'b0);
and (s1n8376,n746,n7398);
wire s0n8377,s1n8377,notn8377;
or (n8377,s0n8377,s1n8377);
not(notn8377,n673);
and (s0n8377,notn8377,1'b0);
and (s1n8377,n673,n8236);
wire s0n8378,s1n8378,notn8378;
or (n8378,s0n8378,s1n8378);
not(notn8378,n7312);
and (s0n8378,notn8378,1'b0);
and (s1n8378,n7312,n8379);
xor (n8379,n7124,n7125);
and (n8380,n8370,n8372);
or (n8381,n8382,n8398);
and (n8382,n8383,n8396);
xor (n8383,n8384,n8385);
xor (n8384,n8032,n8043);
and (n8385,n8386,n8395);
xor (n8386,n8387,n8393);
and (n8387,n8388,n27);
xnor (n8388,n8389,n8019);
nand (n8389,n8390,n8392);
or (n8390,n7423,n8391);
not (n8391,n7381);
nand (n8392,n7423,n8391);
wire s0n8393,s1n8393,notn8393;
or (n8393,s0n8393,s1n8393);
not(notn8393,n6893);
and (s0n8393,notn8393,1'b0);
and (s1n8393,n6893,n8394);
wire s0n8394,s1n8394,notn8394;
or (n8394,s0n8394,s1n8394);
not(notn8394,n746);
and (s0n8394,notn8394,1'b0);
and (s1n8394,n746,n7062);
wire s0n8395,s1n8395,notn8395;
or (n8395,s0n8395,s1n8395);
not(notn8395,n7312);
and (s0n8395,notn8395,1'b0);
and (s1n8395,n7312,n8042);
wire s0n8396,s1n8396,notn8396;
or (n8396,s0n8396,s1n8396);
not(notn8396,n6893);
and (s0n8396,notn8396,1'b0);
and (s1n8396,n6893,n8397);
xor (n8397,n7061,n7070);
and (n8398,n8384,n8385);
wire s0n8399,s1n8399,notn8399;
or (n8399,s0n8399,s1n8399);
not(notn8399,n7134);
and (s0n8399,notn8399,1'b0);
and (s1n8399,n7134,n7968);
and (n8400,n8367,n8381);
and (n8401,n8362,n8363);
xor (n8402,n8218,n8251);
or (n8403,n8404,n8466);
and (n8404,n8405,n8465);
xor (n8405,n8406,n8464);
or (n8406,n8407,n8463);
and (n8407,n8408,n8462);
xor (n8408,n8409,n8410);
xor (n8409,n8225,n8231);
or (n8410,n8411,n8461);
and (n8411,n8412,n8437);
xor (n8412,n8413,n8414);
xor (n8413,n8233,n8237);
or (n8414,n8415,n8436);
and (n8415,n8416,n8435);
xor (n8416,n8417,n8427);
or (n8417,n8418,n8426);
and (n8418,n8419,n8422);
xor (n8419,n8420,n8421);
wire s0n8420,s1n8420,notn8420;
or (n8420,s0n8420,s1n8420);
not(notn8420,n673);
and (s0n8420,notn8420,1'b0);
and (s1n8420,n673,n8306);
xor (n8421,n8308,n8309);
and (n8422,n8423,n27);
nand (n8423,n8424,n8425);
or (n8424,n7394,n8040);
or (n8425,n7428,n8017);
and (n8426,n8420,n8421);
or (n8427,n8428,n8434);
and (n8428,n8429,n8432);
xor (n8429,n8430,n8431);
and (n8430,n7385,n27);
and (n8431,n7630,n27);
and (n8432,n8433,n27);
not (n8433,n7669);
and (n8434,n8430,n8431);
wire s0n8435,s1n8435,notn8435;
or (n8435,s0n8435,s1n8435);
not(notn8435,n7134);
and (s0n8435,notn8435,1'b0);
and (s1n8435,n7134,n8069);
and (n8436,n8417,n8427);
or (n8437,n8438,n8460);
and (n8438,n8439,n8458);
xor (n8439,n8440,n8441);
xor (n8440,n8304,n8311);
or (n8441,n8442,n8457);
and (n8442,n8443,n8456);
xor (n8443,n8444,n8451);
or (n8444,n8445,n8450);
and (n8445,n8446,n8449);
xor (n8446,n8447,n8448);
nor (n8447,n8052,n6944);
wire s0n8448,s1n8448,notn8448;
or (n8448,s0n8448,s1n8448);
not(notn8448,n673);
and (s0n8448,notn8448,1'b0);
and (s1n8448,n673,n8037);
nor (n8449,n7641,n6944);
and (n8450,n8447,n8448);
and (n8451,n8452,n8454);
nor (n8452,n8453,n6944);
not (n8453,n7397);
nor (n8454,n8455,n6944);
not (n8455,n7672);
wire s0n8456,s1n8456,notn8456;
or (n8456,s0n8456,s1n8456);
not(notn8456,n7312);
and (s0n8456,notn8456,1'b0);
and (s1n8456,n7312,n8394);
and (n8457,n8444,n8451);
wire s0n8458,s1n8458,notn8458;
or (n8458,s0n8458,s1n8458);
not(notn8458,n6895);
and (s0n8458,notn8458,1'b0);
and (s1n8458,n6895,n8459);
xor (n8459,n7264,n7273);
and (n8460,n8440,n8441);
and (n8461,n8413,n8414);
wire s0n8462,s1n8462,notn8462;
or (n8462,s0n8462,s1n8462);
not(notn8462,n673);
and (s0n8462,notn8462,1'b0);
and (s1n8462,n673,n8249);
and (n8463,n8409,n8410);
xor (n8464,n8221,n8240);
xor (n8465,n8296,n8317);
and (n8466,n8406,n8464);
and (n8467,n8359,n8402);
xor (n8468,n8257,n8266);
and (n8469,n8355,n8356);
xor (n8470,n8282,n8285);
and (n8471,n8351,n8352);
or (n8472,n8473,n8733);
and (n8473,n8474,n8533);
xor (n8474,n8475,n8476);
xor (n8475,n8350,n8470);
or (n8476,n8477,n8532);
and (n8477,n8478,n8531);
xor (n8478,n8479,n8480);
xor (n8479,n8287,n8320);
or (n8480,n8481,n8530);
and (n8481,n8482,n8529);
xor (n8482,n8483,n8484);
xor (n8483,n8291,n8294);
or (n8484,n8485,n8528);
and (n8485,n8486,n8527);
xor (n8486,n8487,n8496);
or (n8487,n8488,n8495);
and (n8488,n8489,n8494);
xor (n8489,n8490,n8493);
xor (n8490,n8491,n8492);
xor (n8491,n8298,n8299);
wire s0n8492,s1n8492,notn8492;
or (n8492,s0n8492,s1n8492);
not(notn8492,n6893);
and (s0n8492,notn8492,1'b0);
and (s1n8492,n6893,n8379);
wire s0n8493,s1n8493,notn8493;
or (n8493,s0n8493,s1n8493);
not(notn8493,n27);
and (s0n8493,notn8493,1'b0);
and (s1n8493,n27,n8073);
wire s0n8494,s1n8494,notn8494;
or (n8494,s0n8494,s1n8494);
not(notn8494,n27);
and (s0n8494,notn8494,1'b0);
and (s1n8494,n27,n8001);
and (n8495,n8490,n8493);
or (n8496,n8497,n8526);
and (n8497,n8498,n8519);
xor (n8498,n8499,n8518);
or (n8499,n8500,n8517);
and (n8500,n8501,n8516);
xor (n8501,n8502,n8503);
xor (n8502,n8383,n8396);
or (n8503,n8504,n8515);
and (n8504,n8505,n8514);
xor (n8505,n8506,n8507);
wire s0n8506,s1n8506,notn8506;
or (n8506,s0n8506,s1n8506);
not(notn8506,n7312);
and (s0n8506,notn8506,1'b0);
and (s1n8506,n7312,n8397);
or (n8507,n8508,n8513);
and (n8508,n8509,n8512);
xor (n8509,n8510,n8511);
xor (n8510,n8429,n8432);
wire s0n8511,s1n8511,notn8511;
or (n8511,s0n8511,s1n8511);
not(notn8511,n7134);
and (s0n8511,notn8511,1'b0);
and (s1n8511,n7134,n8042);
wire s0n8512,s1n8512,notn8512;
or (n8512,s0n8512,s1n8512);
not(notn8512,n7312);
and (s0n8512,notn8512,1'b0);
and (s1n8512,n7312,n8376);
and (n8513,n8510,n8511);
xor (n8514,n8373,n8377);
and (n8515,n8506,n8507);
wire s0n8516,s1n8516,notn8516;
or (n8516,s0n8516,s1n8516);
not(notn8516,n7134);
and (s0n8516,notn8516,1'b0);
and (s1n8516,n7134,n8245);
and (n8517,n8502,n8503);
xor (n8518,n8329,n8333);
or (n8519,n8520,n8525);
and (n8520,n8521,n8524);
xor (n8521,n8522,n8523);
wire s0n8522,s1n8522,notn8522;
or (n8522,s0n8522,s1n8522);
not(notn8522,n673);
and (s0n8522,notn8522,1'b0);
and (s1n8522,n673,n8332);
xor (n8523,n8301,n8314);
wire s0n8524,s1n8524,notn8524;
or (n8524,s0n8524,s1n8524);
not(notn8524,n27);
and (s0n8524,notn8524,1'b0);
and (s1n8524,n27,n7968);
and (n8525,n8522,n8523);
and (n8526,n8499,n8518);
xor (n8527,n8326,n8336);
and (n8528,n8487,n8496);
xor (n8529,n8322,n8338);
and (n8530,n8483,n8484);
xor (n8531,n8354,n8468);
and (n8532,n8479,n8480);
or (n8533,n8534,n8732);
and (n8534,n8535,n8568);
xor (n8535,n8536,n8567);
or (n8536,n8537,n8566);
and (n8537,n8538,n8565);
xor (n8538,n8539,n8564);
or (n8539,n8540,n8563);
and (n8540,n8541,n8562);
xor (n8541,n8542,n8561);
or (n8542,n8543,n8560);
and (n8543,n8544,n8547);
xor (n8544,n8545,n8546);
xor (n8545,n8366,n8399);
xor (n8546,n8408,n8462);
or (n8547,n8548,n8559);
and (n8548,n8549,n8558);
xor (n8549,n8550,n8551);
xor (n8550,n8369,n8378);
or (n8551,n8552,n8557);
and (n8552,n8553,n8556);
xor (n8553,n8554,n8555);
xor (n8554,n8386,n8395);
wire s0n8555,s1n8555,notn8555;
or (n8555,s0n8555,s1n8555);
not(notn8555,n673);
and (s0n8555,notn8555,1'b0);
and (s1n8555,n673,n8371);
wire s0n8556,s1n8556,notn8556;
or (n8556,s0n8556,s1n8556);
not(notn8556,n7134);
and (s0n8556,notn8556,1'b0);
and (s1n8556,n7134,n8379);
and (n8557,n8554,n8555);
wire s0n8558,s1n8558,notn8558;
or (n8558,s0n8558,s1n8558);
not(notn8558,n27);
and (s0n8558,notn8558,1'b0);
and (s1n8558,n27,n8249);
and (n8559,n8550,n8551);
and (n8560,n8545,n8546);
xor (n8561,n8361,n8364);
xor (n8562,n8405,n8465);
and (n8563,n8542,n8561);
xor (n8564,n8358,n8403);
xor (n8565,n8482,n8529);
and (n8566,n8539,n8564);
xor (n8567,n8478,n8531);
or (n8568,n8569,n8731);
and (n8569,n8570,n8635);
xor (n8570,n8571,n8634);
or (n8571,n8572,n8633);
and (n8572,n8573,n8632);
xor (n8573,n8574,n8631);
or (n8574,n8575,n8630);
and (n8575,n8576,n8623);
xor (n8576,n8577,n8622);
or (n8577,n8578,n8621);
and (n8578,n8579,n8602);
xor (n8579,n8580,n8601);
or (n8580,n8581,n8600);
and (n8581,n8582,n8599);
xor (n8582,n8583,n8598);
or (n8583,n8584,n8597);
and (n8584,n8585,n8596);
xor (n8585,n8586,n8587);
xor (n8586,n8419,n8422);
or (n8587,n8588,n8595);
and (n8588,n8589,n8594);
xor (n8589,n8590,n8593);
and (n8590,n8591,n8592);
wire s0n8591,s1n8591,notn8591;
or (n8591,s0n8591,s1n8591);
not(notn8591,n27);
and (s0n8591,notn8591,1'b0);
and (s1n8591,n27,n8376);
wire s0n8592,s1n8592,notn8592;
or (n8592,s0n8592,s1n8592);
not(notn8592,n27);
and (s0n8592,notn8592,1'b0);
and (s1n8592,n27,n8310);
wire s0n8593,s1n8593,notn8593;
or (n8593,s0n8593,s1n8593);
not(notn8593,n673);
and (s0n8593,notn8593,1'b0);
and (s1n8593,n673,n8310);
xor (n8594,n8452,n8454);
and (n8595,n8590,n8593);
wire s0n8596,s1n8596,notn8596;
or (n8596,s0n8596,s1n8596);
not(notn8596,n7134);
and (s0n8596,notn8596,1'b0);
and (s1n8596,n7134,n8397);
and (n8597,n8586,n8587);
xor (n8598,n8416,n8435);
xor (n8599,n8439,n8458);
and (n8600,n8583,n8598);
xor (n8601,n8412,n8437);
or (n8602,n8603,n8620);
and (n8603,n8604,n8619);
xor (n8604,n8605,n8618);
or (n8605,n8606,n8617);
and (n8606,n8607,n8616);
xor (n8607,n8608,n8609);
wire s0n8608,s1n8608,notn8608;
or (n8608,s0n8608,s1n8608);
not(notn8608,n673);
and (s0n8608,notn8608,1'b0);
and (s1n8608,n673,n8459);
or (n8609,n8610,n8615);
and (n8610,n8611,n8614);
xor (n8611,n8612,n8613);
wire s0n8612,s1n8612,notn8612;
or (n8612,s0n8612,s1n8612);
not(notn8612,n7134);
and (s0n8612,notn8612,1'b0);
and (s1n8612,n7134,n8394);
xor (n8613,n8446,n8449);
wire s0n8614,s1n8614,notn8614;
or (n8614,s0n8614,s1n8614);
not(notn8614,n7134);
and (s0n8614,notn8614,1'b0);
and (s1n8614,n7134,n8376);
and (n8615,n8612,n8613);
xor (n8616,n8509,n8512);
and (n8617,n8608,n8609);
and (n8618,n8332,n27);
wire s0n8619,s1n8619,notn8619;
or (n8619,s0n8619,s1n8619);
not(notn8619,n27);
and (s0n8619,notn8619,1'b0);
and (s1n8619,n27,n8245);
and (n8620,n8605,n8618);
and (n8621,n8580,n8601);
xor (n8622,n8489,n8494);
or (n8623,n8624,n8629);
and (n8624,n8625,n8628);
xor (n8625,n8626,n8627);
xor (n8626,n8501,n8516);
xor (n8627,n8521,n8524);
xor (n8628,n8549,n8558);
and (n8629,n8626,n8627);
and (n8630,n8577,n8622);
xor (n8631,n8486,n8527);
xor (n8632,n8541,n8562);
and (n8633,n8574,n8631);
xor (n8634,n8538,n8565);
or (n8635,n8636,n8730);
and (n8636,n8637,n8729);
xor (n8637,n8638,n8681);
or (n8638,n8639,n8680);
and (n8639,n8640,n8679);
xor (n8640,n8641,n8678);
or (n8641,n8642,n8677);
and (n8642,n8643,n8658);
xor (n8643,n8644,n8657);
or (n8644,n8645,n8656);
and (n8645,n8646,n8655);
xor (n8646,n8647,n8654);
or (n8647,n8648,n8653);
and (n8648,n8649,n8652);
xor (n8649,n8650,n8651);
and (n8650,n8371,n27);
xor (n8651,n8443,n8456);
wire s0n8652,s1n8652,notn8652;
or (n8652,s0n8652,s1n8652);
not(notn8652,n27);
and (s0n8652,notn8652,1'b0);
and (s1n8652,n27,n8379);
and (n8653,n8650,n8651);
xor (n8654,n8505,n8514);
xor (n8655,n8553,n8556);
and (n8656,n8647,n8654);
xor (n8657,n8579,n8602);
or (n8658,n8659,n8676);
and (n8659,n8660,n8675);
xor (n8660,n8661,n8662);
xor (n8661,n8582,n8599);
or (n8662,n8663,n8674);
and (n8663,n8664,n8673);
xor (n8664,n8665,n8672);
or (n8665,n8666,n8671);
and (n8666,n8667,n8670);
xor (n8667,n8668,n8669);
wire s0n8668,s1n8668,notn8668;
or (n8668,s0n8668,s1n8668);
not(notn8668,n27);
and (s0n8668,notn8668,1'b0);
and (s1n8668,n27,n8397);
xor (n8669,n8589,n8594);
wire s0n8670,s1n8670,notn8670;
or (n8670,s0n8670,s1n8670);
not(notn8670,n27);
and (s0n8670,notn8670,1'b0);
and (s1n8670,n27,n8459);
and (n8671,n8668,n8669);
xor (n8672,n8585,n8596);
xor (n8673,n8607,n8616);
and (n8674,n8665,n8672);
xor (n8675,n8604,n8619);
and (n8676,n8661,n8662);
and (n8677,n8644,n8657);
xor (n8678,n8498,n8519);
xor (n8679,n8544,n8547);
and (n8680,n8641,n8678);
nand (n8681,n8682,n8725);
or (n8682,n8683,n8723);
not (n8683,n8684);
nand (n8684,n8685,n8687,n8722);
not (n8685,n8686);
xor (n8686,n8576,n8623);
nand (n8687,n8688,n8721);
or (n8688,n8689,n8690);
xor (n8689,n8643,n8658);
nand (n8690,n8691,n8718);
or (n8691,n8692,n8716);
not (n8692,n8693);
nand (n8693,n8694,n8713);
or (n8694,n8695,n8711);
not (n8695,n8696);
nand (n8696,n8697,n8708);
or (n8697,n8698,n8706);
not (n8698,n8699);
nand (n8699,n8700,n8703);
or (n8700,n8035,n8701);
not (n8701,n8702);
wire s0n8702,s1n8702,notn8702;
or (n8702,s0n8702,s1n8702);
not(notn8702,n27);
and (s0n8702,notn8702,1'b0);
and (s1n8702,n27,n8394);
nand (n8703,n8704,n8705);
or (n8704,n8702,n8036);
xor (n8705,n8591,n8592);
not (n8706,n8707);
xor (n8707,n8611,n8614);
nand (n8708,n8709,n8710);
or (n8709,n8707,n8699);
xor (n8710,n8667,n8670);
not (n8711,n8712);
xor (n8712,n8649,n8652);
nand (n8713,n8714,n8715);
or (n8714,n8712,n8696);
xor (n8715,n8664,n8673);
not (n8716,n8717);
xor (n8717,n8646,n8655);
nand (n8718,n8719,n8720);
or (n8719,n8717,n8693);
xor (n8720,n8660,n8675);
xor (n8721,n8625,n8628);
nand (n8722,n8689,n8690);
not (n8723,n8724);
xor (n8724,n8640,n8679);
nand (n8725,n8726,n8686);
or (n8726,n8727,n8728);
not (n8727,n8722);
not (n8728,n8687);
xor (n8729,n8573,n8632);
and (n8730,n8638,n8681);
and (n8731,n8571,n8634);
and (n8732,n8536,n8567);
and (n8733,n8475,n8476);
and (n8734,n8347,n8348);
and (n8735,n8275,n8276);
and (n8736,n6957,n8199);
nor (n8737,n8738,n8763);
not (n8738,n8739);
nor (n8739,n8740,n8760);
not (n8740,n8741);
nor (n8741,n8742,n8757);
not (n8742,n8743);
nor (n8743,n8744,n8754);
not (n8744,n8745);
nor (n8745,n8746,n8747);
and (n8746,n8152,n8155);
not (n8747,n8748);
nor (n8748,n8749,n8750);
and (n8749,n8147,n8150);
not (n8750,n8751);
xnor (n8751,n8752,n8753);
wire s0n8752,s1n8752,notn8752;
or (n8752,s0n8752,s1n8752);
not(notn8752,n6893);
and (s0n8752,notn8752,1'b0);
and (s1n8752,n6893,n6967);
wire s0n8753,s1n8753,notn8753;
or (n8753,s0n8753,s1n8753);
not(notn8753,n6893);
and (s0n8753,notn8753,1'b0);
and (s1n8753,n6893,n7682);
or (n8754,n8755,n8756);
and (n8755,n8142,n8151);
and (n8756,n8143,n8146);
or (n8757,n8758,n8759);
and (n8758,n8106,n8129);
and (n8759,n8107,n8110);
or (n8760,n8761,n8762);
and (n8761,n8137,n8156);
and (n8762,n8138,n8141);
or (n8763,n8764,n8765);
and (n8764,n6958,n8136);
and (n8765,n6959,n8105);
nor (n8766,n8767,n6839);
not (n8767,n8768);
and (n8768,n66,n21);
wire s0n8769,s1n8769,notn8769;
or (n8769,s0n8769,s1n8769);
not(notn8769,n9514);
and (s0n8769,notn8769,n8770);
and (s1n8769,n9514,n9510);
wire s0n8770,s1n8770,notn8770;
or (n8770,s0n8770,s1n8770);
not(notn8770,n6839);
and (s0n8770,notn8770,n8771);
and (s1n8770,n6839,n6829);
xor (n8771,n8772,n9487);
xor (n8772,n8773,n9388);
xor (n8773,n8774,n9091);
xor (n8774,n8775,n8998);
xor (n8775,n8776,n8883);
xor (n8776,n8752,n8777);
or (n8777,n8778,n8816,n8882);
and (n8778,n8779,n8780);
xor (n8779,n8150,n8155);
and (n8780,n6966,n8781);
or (n8781,n8782,n8783,n8815);
and (n8782,n7930,n7924);
and (n8783,n7924,n8784);
or (n8784,n8785,n8786,n8814);
and (n8785,n7885,n8101);
and (n8786,n8101,n8787);
or (n8787,n8788,n8789,n8813);
and (n8788,n7971,n8076);
and (n8789,n8076,n8790);
or (n8790,n8791,n8792,n8812);
and (n8791,n8262,n8264);
and (n8792,n8264,n8793);
or (n8793,n8794,n8795,n8811);
and (n8794,n8316,n8336);
and (n8795,n8336,n8796);
or (n8796,n8797,n8798,n8810);
and (n8797,n8399,n8493);
and (n8798,n8493,n8799);
or (n8799,n8800,n8801,n8809);
and (n8800,n8516,n8524);
and (n8801,n8524,n8802);
or (n8802,n8803,n8804,n8806);
and (n8803,n8556,n8619);
and (n8804,n8619,n8805);
or (n8805,n8806,n8807,n8808);
and (n8806,n8596,n8652);
and (n8807,n8652,n8808);
and (n8808,n8612,n8668);
and (n8809,n8516,n8802);
and (n8810,n8399,n8799);
and (n8811,n8316,n8796);
and (n8812,n8262,n8793);
and (n8813,n7971,n8790);
and (n8814,n7885,n8787);
and (n8815,n7930,n8784);
and (n8816,n8780,n8817);
or (n8817,n8818,n8821,n8881);
and (n8818,n8819,n8820);
xor (n8819,n7893,n7309);
xor (n8820,n6966,n8781);
and (n8821,n8820,n8822);
or (n8822,n8823,n8827,n8880);
and (n8823,n8824,n8825);
xor (n8824,n8124,n7919);
xor (n8825,n8826,n8784);
xor (n8826,n7930,n7924);
and (n8827,n8825,n8828);
or (n8828,n8829,n8833,n8879);
and (n8829,n8830,n8831);
xor (n8830,n7826,n7819);
xor (n8831,n8832,n8787);
xor (n8832,n7885,n8101);
and (n8833,n8831,n8834);
or (n8834,n8835,n8839,n8878);
and (n8835,n8836,n8837);
xor (n8836,n8189,n7943);
xor (n8837,n8838,n8790);
xor (n8838,n7971,n8076);
and (n8839,n8837,n8840);
or (n8840,n8841,n8845,n8877);
and (n8841,n8842,n8843);
xor (n8842,n7967,n8072);
xor (n8843,n8844,n8793);
xor (n8844,n8262,n8264);
and (n8845,n8843,n8846);
or (n8846,n8847,n8851,n8876);
and (n8847,n8848,n8849);
xor (n8848,n8244,n8240);
xor (n8849,n8850,n8796);
xor (n8850,n8316,n8336);
and (n8851,n8849,n8852);
or (n8852,n8853,n8857,n8875);
and (n8853,n8854,n8855);
xor (n8854,n8492,n8333);
xor (n8855,n8856,n8799);
xor (n8856,n8399,n8493);
and (n8857,n8855,n8858);
or (n8858,n8859,n8863,n8874);
and (n8859,n8860,n8861);
xor (n8860,n8396,n8378);
xor (n8861,n8862,n8802);
xor (n8862,n8516,n8524);
and (n8863,n8861,n8864);
or (n8864,n8865,n8869,n8873);
and (n8865,n8866,n8867);
xor (n8866,n8393,n8506);
xor (n8867,n8868,n8805);
xor (n8868,n8556,n8619);
and (n8869,n8867,n8870);
and (n8870,n8456,n8871);
xor (n8871,n8872,n8808);
xor (n8872,n8596,n8652);
and (n8873,n8866,n8870);
and (n8874,n8860,n8864);
and (n8875,n8854,n8858);
and (n8876,n8848,n8852);
and (n8877,n8842,n8846);
and (n8878,n8836,n8840);
and (n8879,n8830,n8834);
and (n8880,n8824,n8828);
and (n8881,n8819,n8822);
and (n8882,n8779,n8817);
xor (n8883,n8753,n8884);
or (n8884,n8885,n8932,n8997);
and (n8885,n8147,n8886);
and (n8886,n7681,n8887);
or (n8887,n8888,n8890,n8931);
and (n8888,n8115,n8889);
wire s0n8889,s1n8889,notn8889;
or (n8889,s0n8889,s1n8889);
not(notn8889,n27);
and (s0n8889,notn8889,1'b0);
and (s1n8889,n27,n7682);
and (n8890,n8889,n8891);
or (n8891,n8892,n8894,n8930);
and (n8892,n8084,n8893);
wire s0n8893,s1n8893,notn8893;
or (n8893,s0n8893,s1n8893);
not(notn8893,n27);
and (s0n8893,notn8893,1'b0);
and (s1n8893,n27,n7693);
and (n8894,n8893,n8895);
or (n8895,n8896,n8898,n8929);
and (n8896,n7915,n8897);
wire s0n8897,s1n8897,notn8897;
or (n8897,s0n8897,s1n8897);
not(notn8897,n27);
and (s0n8897,notn8897,1'b0);
and (s1n8897,n27,n7525);
and (n8898,n8897,n8899);
or (n8899,n8900,n8902,n8928);
and (n8900,n8009,n8901);
wire s0n8901,s1n8901,notn8901;
or (n8901,s0n8901,s1n8901);
not(notn8901,n27);
and (s0n8901,notn8901,1'b0);
and (s1n8901,n27,n7510);
and (n8902,n8901,n8903);
or (n8903,n8904,n8906,n8927);
and (n8904,n7987,n8905);
wire s0n8905,s1n8905,notn8905;
or (n8905,s0n8905,s1n8905);
not(notn8905,n27);
and (s0n8905,notn8905,1'b0);
and (s1n8905,n27,n7321);
and (n8906,n8905,n8907);
or (n8907,n8908,n8910,n8926);
and (n8908,n8070,n8909);
wire s0n8909,s1n8909,notn8909;
or (n8909,s0n8909,s1n8909);
not(notn8909,n27);
and (s0n8909,notn8909,1'b0);
and (s1n8909,n27,n7862);
and (n8910,n8909,n8911);
or (n8911,n8912,n8914,n8925);
and (n8912,n8237,n8913);
wire s0n8913,s1n8913,notn8913;
or (n8913,s0n8913,s1n8913);
not(notn8913,n27);
and (s0n8913,notn8913,1'b0);
and (s1n8913,n27,n7957);
and (n8914,n8913,n8915);
or (n8915,n8916,n8918,n8920);
and (n8916,n8435,n8917);
wire s0n8917,s1n8917,notn8917;
or (n8917,s0n8917,s1n8917);
not(notn8917,n27);
and (s0n8917,notn8917,1'b0);
and (s1n8917,n27,n7963);
and (n8918,n8917,n8919);
or (n8919,n8920,n8922,n8923);
and (n8920,n8511,n8921);
wire s0n8921,s1n8921,notn8921;
or (n8921,s0n8921,s1n8921);
not(notn8921,n27);
and (s0n8921,notn8921,1'b0);
and (s1n8921,n27,n8069);
and (n8922,n8921,n8923);
and (n8923,n8614,n8924);
wire s0n8924,s1n8924,notn8924;
or (n8924,s0n8924,s1n8924);
not(notn8924,n27);
and (s0n8924,notn8924,1'b0);
and (s1n8924,n27,n8042);
and (n8925,n8237,n8915);
and (n8926,n8070,n8911);
and (n8927,n7987,n8907);
and (n8928,n8009,n8903);
and (n8929,n7915,n8899);
and (n8930,n8084,n8895);
and (n8931,n8115,n8891);
and (n8932,n8886,n8933);
or (n8933,n8934,n8937,n8996);
and (n8934,n8935,n8936);
xor (n8935,n7691,n7692);
xor (n8936,n7681,n8887);
and (n8937,n8936,n8938);
or (n8938,n8939,n8943,n8995);
and (n8939,n8940,n8941);
xor (n8940,n8118,n7524);
xor (n8941,n8942,n8891);
xor (n8942,n8115,n8889);
and (n8943,n8941,n8944);
or (n8944,n8945,n8949,n8994);
and (n8945,n8946,n8947);
xor (n8946,n7320,n7509);
xor (n8947,n8948,n8895);
xor (n8948,n8084,n8893);
and (n8949,n8947,n8950);
or (n8950,n8951,n8954,n8993);
and (n8951,n7912,n8952);
xor (n8952,n8953,n8899);
xor (n8953,n7915,n8897);
and (n8954,n8952,n8955);
or (n8955,n8956,n8960,n8992);
and (n8956,n8957,n8958);
xor (n8957,n7956,n7861);
xor (n8958,n8959,n8903);
xor (n8959,n8009,n8901);
and (n8960,n8958,n8961);
or (n8961,n8962,n8966,n8991);
and (n8962,n8963,n8964);
xor (n8963,n7962,n8023);
xor (n8964,n8965,n8907);
xor (n8965,n7987,n8905);
and (n8966,n8964,n8967);
or (n8967,n8968,n8972,n8990);
and (n8968,n8969,n8970);
xor (n8969,n8068,n7996);
xor (n8970,n8971,n8911);
xor (n8971,n8070,n8909);
and (n8972,n8970,n8973);
or (n8973,n8974,n8978,n8989);
and (n8974,n8975,n8976);
xor (n8975,n8041,n8234);
xor (n8976,n8977,n8915);
xor (n8977,n8237,n8913);
and (n8978,n8976,n8979);
or (n8979,n8980,n8984,n8988);
and (n8980,n8981,n8982);
xor (n8981,n8375,n8395);
xor (n8982,n8983,n8919);
xor (n8983,n8435,n8917);
and (n8984,n8982,n8985);
and (n8985,n8512,n8986);
xor (n8986,n8987,n8923);
xor (n8987,n8511,n8921);
and (n8988,n8981,n8985);
and (n8989,n8975,n8979);
and (n8990,n8969,n8973);
and (n8991,n8963,n8967);
and (n8992,n8957,n8961);
and (n8993,n7912,n8955);
and (n8994,n8946,n8950);
and (n8995,n8940,n8944);
and (n8996,n8935,n8938);
and (n8997,n8147,n8933);
or (n8998,n8999,n9004,n9090);
and (n8999,n9000,n9002);
xor (n9000,n9001,n8817);
xor (n9001,n8779,n8780);
xor (n9002,n9003,n8933);
xor (n9003,n8147,n8886);
and (n9004,n9002,n9005);
or (n9005,n9006,n9011,n9089);
and (n9006,n9007,n9009);
xor (n9007,n9008,n8822);
xor (n9008,n8819,n8820);
xor (n9009,n9010,n8938);
xor (n9010,n8935,n8936);
and (n9011,n9009,n9012);
or (n9012,n9013,n9018,n9088);
and (n9013,n9014,n9016);
xor (n9014,n9015,n8828);
xor (n9015,n8824,n8825);
xor (n9016,n9017,n8944);
xor (n9017,n8940,n8941);
and (n9018,n9016,n9019);
or (n9019,n9020,n9025,n9087);
and (n9020,n9021,n9023);
xor (n9021,n9022,n8834);
xor (n9022,n8830,n8831);
xor (n9023,n9024,n8950);
xor (n9024,n8946,n8947);
and (n9025,n9023,n9026);
or (n9026,n9027,n9032,n9086);
and (n9027,n9028,n9030);
xor (n9028,n9029,n8840);
xor (n9029,n8836,n8837);
xor (n9030,n9031,n8955);
xor (n9031,n7912,n8952);
and (n9032,n9030,n9033);
or (n9033,n9034,n9039,n9085);
and (n9034,n9035,n9037);
xor (n9035,n9036,n8846);
xor (n9036,n8842,n8843);
xor (n9037,n9038,n8961);
xor (n9038,n8957,n8958);
and (n9039,n9037,n9040);
or (n9040,n9041,n9046,n9084);
and (n9041,n9042,n9044);
xor (n9042,n9043,n8852);
xor (n9043,n8848,n8849);
xor (n9044,n9045,n8967);
xor (n9045,n8963,n8964);
and (n9046,n9044,n9047);
or (n9047,n9048,n9053,n9083);
and (n9048,n9049,n9051);
xor (n9049,n9050,n8858);
xor (n9050,n8854,n8855);
xor (n9051,n9052,n8973);
xor (n9052,n8969,n8970);
and (n9053,n9051,n9054);
or (n9054,n9055,n9060,n9082);
and (n9055,n9056,n9058);
xor (n9056,n9057,n8864);
xor (n9057,n8860,n8861);
xor (n9058,n9059,n8979);
xor (n9059,n8975,n8976);
and (n9060,n9058,n9061);
or (n9061,n9062,n9067,n9081);
and (n9062,n9063,n9065);
xor (n9063,n9064,n8870);
xor (n9064,n8866,n8867);
xor (n9065,n9066,n8985);
xor (n9066,n8981,n8982);
and (n9067,n9065,n9068);
or (n9068,n9069,n9072,n9080);
and (n9069,n9070,n9071);
xor (n9070,n8456,n8871);
xor (n9071,n8512,n8986);
and (n9072,n9071,n9073);
or (n9073,n9074,n9077,n9079);
and (n9074,n9075,n9076);
xor (n9075,n8612,n8668);
xor (n9076,n8614,n8924);
and (n9077,n9076,n9078);
and (n9078,n8702,n8591);
and (n9079,n9075,n9078);
and (n9080,n9070,n9073);
and (n9081,n9063,n9068);
and (n9082,n9056,n9061);
and (n9083,n9049,n9054);
and (n9084,n9042,n9047);
and (n9085,n9035,n9040);
and (n9086,n9028,n9033);
and (n9087,n9021,n9026);
and (n9088,n9014,n9019);
and (n9089,n9007,n9012);
and (n9090,n9000,n9005);
xor (n9091,n9092,n9295);
xor (n9092,n9093,n9189);
or (n9093,n9094,n9131,n9188);
and (n9094,n8153,n9095);
and (n9095,n8121,n9096);
or (n9096,n9097,n9098,n9130);
and (n9097,n8119,n7925);
and (n9098,n7925,n9099);
or (n9099,n9100,n9101,n9129);
and (n9100,n7762,n8081);
and (n9101,n8081,n9102);
or (n9102,n9103,n9104,n9128);
and (n9103,n7950,n7945);
and (n9104,n7945,n9105);
or (n9105,n9106,n9107,n9127);
and (n9106,n8263,n8251);
and (n9107,n8251,n9108);
or (n9108,n9109,n9110,n9126);
and (n9109,n8317,n8363);
and (n9110,n8363,n9111);
or (n9111,n9112,n9113,n9125);
and (n9112,n8462,n8494);
and (n9113,n8494,n9114);
or (n9114,n9115,n9116,n9124);
and (n9115,n8522,n8558);
and (n9116,n8558,n9117);
or (n9117,n9118,n9119,n9121);
and (n9118,n8555,n8618);
and (n9119,n8618,n9120);
or (n9120,n9121,n9122,n9123);
and (n9121,n8608,n8650);
and (n9122,n8650,n9123);
and (n9123,n8593,n8670);
and (n9124,n8522,n9117);
and (n9125,n8462,n9114);
and (n9126,n8317,n9111);
and (n9127,n8263,n9108);
and (n9128,n7950,n9105);
and (n9129,n7762,n9102);
and (n9130,n8119,n9099);
and (n9131,n9095,n9132);
or (n9132,n9133,n9135,n9187);
and (n9133,n7135,n9134);
xor (n9134,n8121,n9096);
and (n9135,n9134,n9136);
or (n9136,n9137,n9140,n9186);
and (n9137,n7918,n9138);
xor (n9138,n9139,n9099);
xor (n9139,n8119,n7925);
and (n9140,n9138,n9141);
or (n9141,n9142,n9145,n9185);
and (n9142,n7815,n9143);
xor (n9143,n9144,n9102);
xor (n9144,n7762,n8081);
and (n9145,n9143,n9146);
or (n9146,n9147,n9150,n9184);
and (n9147,n8191,n9148);
xor (n9148,n9149,n9105);
xor (n9149,n7950,n7945);
and (n9150,n9148,n9151);
or (n9151,n9152,n9155,n9183);
and (n9152,n8000,n9153);
xor (n9153,n9154,n9108);
xor (n9154,n8263,n8251);
and (n9155,n9153,n9156);
or (n9156,n9157,n9160,n9182);
and (n9157,n8248,n9158);
xor (n9158,n9159,n9111);
xor (n9159,n8317,n8363);
and (n9160,n9158,n9161);
or (n9161,n9162,n9165,n9181);
and (n9162,n8331,n9163);
xor (n9163,n9164,n9114);
xor (n9164,n8462,n8494);
and (n9165,n9163,n9166);
or (n9166,n9167,n9170,n9180);
and (n9167,n8370,n9168);
xor (n9168,n9169,n9117);
xor (n9169,n8522,n8558);
and (n9170,n9168,n9171);
or (n9171,n9172,n9175,n9179);
and (n9172,n8458,n9173);
xor (n9173,n9174,n9120);
xor (n9174,n8555,n8618);
and (n9175,n9173,n9176);
and (n9176,n8309,n9177);
xor (n9177,n9178,n9123);
xor (n9178,n8608,n8650);
and (n9179,n8458,n9176);
and (n9180,n8370,n9171);
and (n9181,n8331,n9166);
and (n9182,n8248,n9161);
and (n9183,n8000,n9156);
and (n9184,n8191,n9151);
and (n9185,n7815,n9146);
and (n9186,n7918,n9141);
and (n9187,n7135,n9136);
and (n9188,n8153,n9132);
or (n9189,n9190,n9237,n9294);
and (n9190,n8154,n9191);
and (n9191,n7695,n9192);
or (n9192,n9193,n9195,n9236);
and (n9193,n8128,n9194);
wire s0n9194,s1n9194,notn9194;
or (n9194,s0n9194,s1n9194);
not(notn9194,n27);
and (s0n9194,notn9194,1'b0);
and (s1n9194,n27,n7696);
and (n9195,n9194,n9196);
or (n9196,n9197,n9199,n9235);
and (n9197,n7916,n9198);
wire s0n9198,s1n9198,notn9198;
or (n9198,s0n9198,s1n9198);
not(notn9198,n27);
and (s0n9198,notn9198,1'b0);
and (s1n9198,n27,n7902);
and (n9199,n9198,n9200);
or (n9200,n9201,n9203,n9234);
and (n9201,n8184,n9202);
wire s0n9202,s1n9202,notn9202;
or (n9202,s0n9202,s1n9202);
not(notn9202,n27);
and (s0n9202,notn9202,1'b0);
and (s1n9202,n27,n7537);
and (n9203,n9202,n9204);
or (n9204,n9205,n9207,n9233);
and (n9205,n8025,n9206);
wire s0n9206,s1n9206,notn9206;
or (n9206,s0n9206,s1n9206);
not(notn9206,n27);
and (s0n9206,notn9206,1'b0);
and (s1n9206,n27,n8100);
and (n9207,n9206,n9208);
or (n9208,n9209,n9211,n9232);
and (n9209,n7998,n9210);
wire s0n9210,s1n9210,notn9210;
or (n9210,s0n9210,s1n9210);
not(notn9210,n27);
and (s0n9210,notn9210,1'b0);
and (s1n9210,n27,n7833);
and (n9211,n9210,n9212);
or (n9212,n9213,n9215,n9231);
and (n9213,n8067,n9214);
wire s0n9214,s1n9214,notn9214;
or (n9214,s0n9214,s1n9214);
not(notn9214,n27);
and (s0n9214,notn9214,1'b0);
and (s1n9214,n27,n7882);
and (n9215,n9214,n9216);
or (n9216,n9217,n9219,n9230);
and (n9217,n8314,n9218);
wire s0n9218,s1n9218,notn9218;
or (n9218,s0n9218,s1n9218);
not(notn9218,n27);
and (s0n9218,notn9218,1'b0);
and (s1n9218,n27,n7966);
and (n9219,n9218,n9220);
or (n9220,n9221,n9223,n9225);
and (n9221,n8377,n9222);
wire s0n9222,s1n9222,notn9222;
or (n9222,s0n9222,s1n9222);
not(notn9222,n27);
and (s0n9222,notn9222,1'b0);
and (s1n9222,n27,n8063);
and (n9223,n9222,n9224);
or (n9224,n9225,n9227,n9228);
and (n9225,n8420,n9226);
wire s0n9226,s1n9226,notn9226;
or (n9226,s0n9226,s1n9226);
not(notn9226,n27);
and (s0n9226,notn9226,1'b0);
and (s1n9226,n27,n8236);
and (n9227,n9226,n9228);
and (n9228,n8448,n9229);
wire s0n9229,s1n9229,notn9229;
or (n9229,s0n9229,s1n9229);
not(notn9229,n27);
and (s0n9229,notn9229,1'b0);
and (s1n9229,n27,n8306);
and (n9230,n8314,n9220);
and (n9231,n8067,n9216);
and (n9232,n7998,n9212);
and (n9233,n8025,n9208);
and (n9234,n8184,n9204);
and (n9235,n7916,n9200);
and (n9236,n8128,n9196);
and (n9237,n9191,n9238);
or (n9238,n9239,n9241,n9293);
and (n9239,n7901,n9240);
xor (n9240,n7695,n9192);
and (n9241,n9240,n9242);
or (n9242,n9243,n9246,n9292);
and (n9243,n7536,n9244);
xor (n9244,n9245,n9196);
xor (n9245,n8128,n9194);
and (n9246,n9244,n9247);
or (n9247,n9248,n9251,n9291);
and (n9248,n8099,n9249);
xor (n9249,n9250,n9200);
xor (n9250,n7916,n9198);
and (n9251,n9249,n9252);
or (n9252,n9253,n9256,n9290);
and (n9253,n7832,n9254);
xor (n9254,n9255,n9204);
xor (n9255,n8184,n9202);
and (n9256,n9254,n9257);
or (n9257,n9258,n9261,n9289);
and (n9258,n7881,n9259);
xor (n9259,n9260,n9208);
xor (n9260,n8025,n9206);
and (n9261,n9259,n9262);
or (n9262,n9263,n9266,n9288);
and (n9263,n7965,n9264);
xor (n9264,n9265,n9212);
xor (n9265,n7998,n9210);
and (n9266,n9264,n9267);
or (n9267,n9268,n9271,n9287);
and (n9268,n8062,n9269);
xor (n9269,n9270,n9216);
xor (n9270,n8067,n9214);
and (n9271,n9269,n9272);
or (n9272,n9273,n9276,n9286);
and (n9273,n8235,n9274);
xor (n9274,n9275,n9220);
xor (n9275,n8314,n9218);
and (n9276,n9274,n9277);
or (n9277,n9278,n9281,n9285);
and (n9278,n8305,n9279);
xor (n9279,n9280,n9224);
xor (n9280,n8377,n9222);
and (n9281,n9279,n9282);
and (n9282,n8308,n9283);
xor (n9283,n9284,n9228);
xor (n9284,n8420,n9226);
and (n9285,n8305,n9282);
and (n9286,n8235,n9277);
and (n9287,n8062,n9272);
and (n9288,n7965,n9267);
and (n9289,n7881,n9262);
and (n9290,n7832,n9257);
and (n9291,n8099,n9252);
and (n9292,n7536,n9247);
and (n9293,n7901,n9242);
and (n9294,n8154,n9238);
or (n9295,n9296,n9301,n9387);
and (n9296,n9297,n9299);
xor (n9297,n9298,n9132);
xor (n9298,n8153,n9095);
xor (n9299,n9300,n9238);
xor (n9300,n8154,n9191);
and (n9301,n9299,n9302);
or (n9302,n9303,n9308,n9386);
and (n9303,n9304,n9306);
xor (n9304,n9305,n9136);
xor (n9305,n7135,n9134);
xor (n9306,n9307,n9242);
xor (n9307,n7901,n9240);
and (n9308,n9306,n9309);
or (n9309,n9310,n9315,n9385);
and (n9310,n9311,n9313);
xor (n9311,n9312,n9141);
xor (n9312,n7918,n9138);
xor (n9313,n9314,n9247);
xor (n9314,n7536,n9244);
and (n9315,n9313,n9316);
or (n9316,n9317,n9322,n9384);
and (n9317,n9318,n9320);
xor (n9318,n9319,n9146);
xor (n9319,n7815,n9143);
xor (n9320,n9321,n9252);
xor (n9321,n8099,n9249);
and (n9322,n9320,n9323);
or (n9323,n9324,n9329,n9383);
and (n9324,n9325,n9327);
xor (n9325,n9326,n9151);
xor (n9326,n8191,n9148);
xor (n9327,n9328,n9257);
xor (n9328,n7832,n9254);
and (n9329,n9327,n9330);
or (n9330,n9331,n9336,n9382);
and (n9331,n9332,n9334);
xor (n9332,n9333,n9156);
xor (n9333,n8000,n9153);
xor (n9334,n9335,n9262);
xor (n9335,n7881,n9259);
and (n9336,n9334,n9337);
or (n9337,n9338,n9343,n9381);
and (n9338,n9339,n9341);
xor (n9339,n9340,n9161);
xor (n9340,n8248,n9158);
xor (n9341,n9342,n9267);
xor (n9342,n7965,n9264);
and (n9343,n9341,n9344);
or (n9344,n9345,n9350,n9380);
and (n9345,n9346,n9348);
xor (n9346,n9347,n9166);
xor (n9347,n8331,n9163);
xor (n9348,n9349,n9272);
xor (n9349,n8062,n9269);
and (n9350,n9348,n9351);
or (n9351,n9352,n9357,n9379);
and (n9352,n9353,n9355);
xor (n9353,n9354,n9171);
xor (n9354,n8370,n9168);
xor (n9355,n9356,n9277);
xor (n9356,n8235,n9274);
and (n9357,n9355,n9358);
or (n9358,n9359,n9364,n9378);
and (n9359,n9360,n9362);
xor (n9360,n9361,n9176);
xor (n9361,n8458,n9173);
xor (n9362,n9363,n9282);
xor (n9363,n8305,n9279);
and (n9364,n9362,n9365);
or (n9365,n9366,n9369,n9377);
and (n9366,n9367,n9368);
xor (n9367,n8309,n9177);
xor (n9368,n8308,n9283);
and (n9369,n9368,n9370);
or (n9370,n9371,n9374,n9376);
and (n9371,n9372,n9373);
xor (n9372,n8593,n8670);
xor (n9373,n8448,n9229);
and (n9374,n9373,n9375);
and (n9375,n8592,n8036);
and (n9376,n9372,n9375);
and (n9377,n9367,n9370);
and (n9378,n9360,n9365);
and (n9379,n9353,n9358);
and (n9380,n9346,n9351);
and (n9381,n9339,n9344);
and (n9382,n9332,n9337);
and (n9383,n9325,n9330);
and (n9384,n9318,n9323);
and (n9385,n9311,n9316);
and (n9386,n9304,n9309);
and (n9387,n9297,n9302);
or (n9388,n9389,n9394,n9486);
and (n9389,n9390,n9392);
xor (n9390,n9391,n9005);
xor (n9391,n9000,n9002);
xor (n9392,n9393,n9302);
xor (n9393,n9297,n9299);
and (n9394,n9392,n9395);
or (n9395,n9396,n9401,n9485);
and (n9396,n9397,n9399);
xor (n9397,n9398,n9012);
xor (n9398,n9007,n9009);
xor (n9399,n9400,n9309);
xor (n9400,n9304,n9306);
and (n9401,n9399,n9402);
or (n9402,n9403,n9408,n9484);
and (n9403,n9404,n9406);
xor (n9404,n9405,n9019);
xor (n9405,n9014,n9016);
xor (n9406,n9407,n9316);
xor (n9407,n9311,n9313);
and (n9408,n9406,n9409);
or (n9409,n9410,n9415,n9483);
and (n9410,n9411,n9413);
xor (n9411,n9412,n9026);
xor (n9412,n9021,n9023);
xor (n9413,n9414,n9323);
xor (n9414,n9318,n9320);
and (n9415,n9413,n9416);
or (n9416,n9417,n9422,n9482);
and (n9417,n9418,n9420);
xor (n9418,n9419,n9033);
xor (n9419,n9028,n9030);
xor (n9420,n9421,n9330);
xor (n9421,n9325,n9327);
and (n9422,n9420,n9423);
or (n9423,n9424,n9429,n9481);
and (n9424,n9425,n9427);
xor (n9425,n9426,n9040);
xor (n9426,n9035,n9037);
xor (n9427,n9428,n9337);
xor (n9428,n9332,n9334);
and (n9429,n9427,n9430);
or (n9430,n9431,n9436,n9480);
and (n9431,n9432,n9434);
xor (n9432,n9433,n9047);
xor (n9433,n9042,n9044);
xor (n9434,n9435,n9344);
xor (n9435,n9339,n9341);
and (n9436,n9434,n9437);
or (n9437,n9438,n9443,n9479);
and (n9438,n9439,n9441);
xor (n9439,n9440,n9054);
xor (n9440,n9049,n9051);
xor (n9441,n9442,n9351);
xor (n9442,n9346,n9348);
and (n9443,n9441,n9444);
or (n9444,n9445,n9450,n9478);
and (n9445,n9446,n9448);
xor (n9446,n9447,n9061);
xor (n9447,n9056,n9058);
xor (n9448,n9449,n9358);
xor (n9449,n9353,n9355);
and (n9450,n9448,n9451);
or (n9451,n9452,n9457,n9477);
and (n9452,n9453,n9455);
xor (n9453,n9454,n9068);
xor (n9454,n9063,n9065);
xor (n9455,n9456,n9365);
xor (n9456,n9360,n9362);
and (n9457,n9455,n9458);
or (n9458,n9459,n9464,n9476);
and (n9459,n9460,n9462);
xor (n9460,n9461,n9073);
xor (n9461,n9070,n9071);
xor (n9462,n9463,n9370);
xor (n9463,n9367,n9368);
and (n9464,n9462,n9465);
or (n9465,n9466,n9471,n9475);
and (n9466,n9467,n9469);
xor (n9467,n9468,n9078);
xor (n9468,n9075,n9076);
xor (n9469,n9470,n9375);
xor (n9470,n9372,n9373);
and (n9471,n9469,n9472);
and (n9472,n9473,n9474);
xor (n9473,n8702,n8591);
xor (n9474,n8592,n8036);
and (n9475,n9467,n9472);
and (n9476,n9460,n9465);
and (n9477,n9453,n9458);
and (n9478,n9446,n9451);
and (n9479,n9439,n9444);
and (n9480,n9432,n9437);
and (n9481,n9425,n9430);
and (n9482,n9418,n9423);
and (n9483,n9411,n9416);
and (n9484,n9404,n9409);
and (n9485,n9397,n9402);
and (n9486,n9390,n9395);
and (n9487,n9488,n9490);
xor (n9488,n9489,n9395);
xor (n9489,n9390,n9392);
and (n9490,n9491,n9493);
xor (n9491,n9492,n9402);
xor (n9492,n9397,n9399);
and (n9493,n9494,n9496);
xor (n9494,n9495,n9409);
xor (n9495,n9404,n9406);
and (n9496,n9497,n9499);
xor (n9497,n9498,n9416);
xor (n9498,n9411,n9413);
and (n9499,n9500,n9502);
xor (n9500,n9501,n9423);
xor (n9501,n9418,n9420);
and (n9502,n9503,n9505);
xor (n9503,n9504,n9430);
xor (n9504,n9425,n9427);
and (n9505,n9506,n9508);
xor (n9506,n9507,n9437);
xor (n9507,n9432,n9434);
xor (n9508,n9509,n9444);
xor (n9509,n9439,n9441);
or (n9510,n9511,n4,n6829);
and (n9511,n9512,n9513);
wire s0n9512,s1n9512,notn9512;
or (n9512,s0n9512,s1n9512);
not(notn9512,n3077);
and (s0n9512,notn9512,1'b0);
and (s1n9512,n3077,n2);
nor (n9513,n2955,n905,n906);
and (n9514,n594,n21);
endmodule
