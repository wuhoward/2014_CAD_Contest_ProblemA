module top (out,n20,n21,n25,n27,n29,n30,n31,n35,n36
        ,n37,n46,n47,n48,n55,n56,n60,n62,n64,n65
        ,n68,n70,n72,n74,n75,n76,n77,n78,n79,n80
        ,n81,n82,n83,n84,n85,n86,n87,n88,n89,n90
        ,n91,n92,n93,n94,n95,n96,n97,n98,n99,n100
        ,n101,n102,n109,n110,n111,n120,n121,n122,n127,n128
        ,n129,n132,n133,n134,n140,n141,n142,n160,n161,n162
        ,n169,n170,n171,n174,n175,n176,n189,n190,n191,n201
        ,n202,n203,n209,n210,n211,n219,n220,n221,n225,n226
        ,n227,n235,n236,n237,n241,n242,n243,n255,n256,n257
        ,n268,n269,n270,n279,n280,n281,n284,n285,n286,n294
        ,n295,n296,n313,n314,n315,n324,n325,n326,n333,n334
        ,n335,n348,n349,n350,n361,n362,n363,n371,n372,n373
        ,n380,n381,n382,n392,n393,n394,n401,n402,n403,n410
        ,n411,n412,n1260,n1261,n1265,n1267,n1269,n1272,n1273,n1277
        ,n1279,n1281,n1282,n1285,n1287,n1289,n1291,n1292,n1293,n1294
        ,n1295,n1296,n1297,n1298,n1299,n1300,n1301,n1302,n1303,n1304
        ,n1305,n1306,n1307,n1308,n1309,n1310,n1311,n1312,n1313,n1314
        ,n1315,n1316,n1317,n1318,n1319,n1322,n1323,n1326,n1327,n1328
        ,n1333,n1334,n1338,n1339,n1340);
output out;
input n20;
input n21;
input n25;
input n27;
input n29;
input n30;
input n31;
input n35;
input n36;
input n37;
input n46;
input n47;
input n48;
input n55;
input n56;
input n60;
input n62;
input n64;
input n65;
input n68;
input n70;
input n72;
input n74;
input n75;
input n76;
input n77;
input n78;
input n79;
input n80;
input n81;
input n82;
input n83;
input n84;
input n85;
input n86;
input n87;
input n88;
input n89;
input n90;
input n91;
input n92;
input n93;
input n94;
input n95;
input n96;
input n97;
input n98;
input n99;
input n100;
input n101;
input n102;
input n109;
input n110;
input n111;
input n120;
input n121;
input n122;
input n127;
input n128;
input n129;
input n132;
input n133;
input n134;
input n140;
input n141;
input n142;
input n160;
input n161;
input n162;
input n169;
input n170;
input n171;
input n174;
input n175;
input n176;
input n189;
input n190;
input n191;
input n201;
input n202;
input n203;
input n209;
input n210;
input n211;
input n219;
input n220;
input n221;
input n225;
input n226;
input n227;
input n235;
input n236;
input n237;
input n241;
input n242;
input n243;
input n255;
input n256;
input n257;
input n268;
input n269;
input n270;
input n279;
input n280;
input n281;
input n284;
input n285;
input n286;
input n294;
input n295;
input n296;
input n313;
input n314;
input n315;
input n324;
input n325;
input n326;
input n333;
input n334;
input n335;
input n348;
input n349;
input n350;
input n361;
input n362;
input n363;
input n371;
input n372;
input n373;
input n380;
input n381;
input n382;
input n392;
input n393;
input n394;
input n401;
input n402;
input n403;
input n410;
input n411;
input n412;
input n1260;
input n1261;
input n1265;
input n1267;
input n1269;
input n1272;
input n1273;
input n1277;
input n1279;
input n1281;
input n1282;
input n1285;
input n1287;
input n1289;
input n1291;
input n1292;
input n1293;
input n1294;
input n1295;
input n1296;
input n1297;
input n1298;
input n1299;
input n1300;
input n1301;
input n1302;
input n1303;
input n1304;
input n1305;
input n1306;
input n1307;
input n1308;
input n1309;
input n1310;
input n1311;
input n1312;
input n1313;
input n1314;
input n1315;
input n1316;
input n1317;
input n1318;
input n1319;
input n1322;
input n1323;
input n1326;
input n1327;
input n1328;
input n1333;
input n1334;
input n1338;
input n1339;
input n1340;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n22;
wire n23;
wire n24;
wire n26;
wire n28;
wire n32;
wire n33;
wire n34;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n57;
wire n58;
wire n59;
wire n61;
wire n63;
wire n66;
wire n67;
wire n69;
wire n71;
wire n73;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n123;
wire n124;
wire n125;
wire n126;
wire n130;
wire n131;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n172;
wire n173;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n222;
wire n223;
wire n224;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n238;
wire n239;
wire n240;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n282;
wire n283;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1262;
wire n1263;
wire n1264;
wire n1266;
wire n1268;
wire n1270;
wire n1271;
wire n1274;
wire n1275;
wire n1276;
wire n1278;
wire n1280;
wire n1283;
wire n1284;
wire n1286;
wire n1288;
wire n1290;
wire n1320;
wire n1321;
wire n1324;
wire n1325;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1335;
wire n1336;
wire n1337;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
xnor (out,n0,n1364);
nand (n0,n1,n1252);
nand (n1,n2,n1251);
or (n2,n3,n702);
nand (n3,n4,n701);
nand (n4,n5,n639);
not (n5,n6);
xor (n6,n7,n590);
xor (n7,n8,n416);
xor (n8,n9,n303);
xor (n9,n10,n194);
xor (n10,n11,n152);
xor (n11,n12,n114);
nand (n12,n13,n104);
or (n13,n14,n50);
nand (n14,n15,n41);
or (n15,n16,n38);
not (n16,n17);
nand (n17,n18,n32);
wire s0n18,s1n18,notn18;
or (n18,s0n18,s1n18);
not(notn18,n31);
and (s0n18,notn18,n19);
and (s1n18,n31,n30);
wire s0n19,s1n19,notn19;
or (n19,s0n19,s1n19);
not(notn19,n22);
and (s0n19,notn19,n20);
and (s1n19,n22,n21);
and (n22,n23,n28);
and (n23,n24,n26);
not (n24,n25);
not (n26,n27);
not (n28,n29);
not (n32,n33);
wire s0n33,s1n33,notn33;
or (n33,s0n33,s1n33);
not(notn33,n31);
and (s0n33,notn33,n34);
and (s1n33,n31,n37);
wire s0n34,s1n34,notn34;
or (n34,s0n34,s1n34);
not(notn34,n22);
and (s0n34,notn34,n35);
and (s1n34,n22,n36);
not (n38,n39);
nand (n39,n40,n33);
not (n40,n18);
nor (n41,n42,n49);
and (n42,n43,n33);
not (n43,n44);
wire s0n44,s1n44,notn44;
or (n44,s0n44,s1n44);
not(notn44,n31);
and (s0n44,notn44,n45);
and (s1n44,n31,n48);
wire s0n45,s1n45,notn45;
or (n45,s0n45,s1n45);
not(notn45,n22);
and (s0n45,notn45,n46);
and (s1n45,n22,n47);
and (n49,n44,n32);
not (n50,n51);
nand (n51,n52,n103);
or (n52,n40,n53);
wire s0n53,s1n53,notn53;
or (n53,s0n53,s1n53);
not(notn53,n66);
and (s0n53,notn53,n54);
and (s1n53,n66,n65);
wire s0n54,s1n54,notn54;
or (n54,s0n54,s1n54);
not(notn54,n57);
and (s0n54,notn54,n55);
and (s1n54,n57,n56);
and (n57,n58,n63);
and (n58,n59,n61);
not (n59,n60);
not (n61,n62);
not (n63,n64);
and (n66,n67,n69);
not (n67,n68);
or (n69,n70,n71);
and (n71,n72,n73);
or (n73,n74,n75,n76,n77,n78,n79,n80,n81,n82,n83,n84,n85,n86,n87,n88,n89,n90,n91,n92,n93,n94,n95,n96,n97,n98,n99,n100,n101,n102);
nand (n103,n53,n40);
nand (n104,n105,n113);
nand (n105,n106,n112);
or (n106,n40,n107);
wire s0n107,s1n107,notn107;
or (n107,s0n107,s1n107);
not(notn107,n66);
and (s0n107,notn107,n108);
and (s1n107,n66,n111);
wire s0n108,s1n108,notn108;
or (n108,s0n108,s1n108);
not(notn108,n57);
and (s0n108,notn108,n109);
and (s1n108,n57,n110);
nand (n112,n107,n40);
not (n113,n41);
nand (n114,n115,n135);
or (n115,n116,n124);
nor (n116,n117,n123);
and (n117,n118,n43);
wire s0n118,s1n118,notn118;
or (n118,s0n118,s1n118);
not(notn118,n66);
and (s0n118,notn118,n119);
and (s1n118,n66,n122);
wire s0n119,s1n119,notn119;
or (n119,s0n119,s1n119);
not(notn119,n57);
and (s0n119,notn119,n120);
and (s1n119,n57,n121);
nor (n123,n118,n43);
xnor (n124,n125,n130);
wire s0n125,s1n125,notn125;
or (n125,s0n125,s1n125);
not(notn125,n31);
and (s0n125,notn125,n126);
and (s1n125,n31,n129);
wire s0n126,s1n126,notn126;
or (n126,s0n126,s1n126);
not(notn126,n22);
and (s0n126,notn126,n127);
and (s1n126,n22,n128);
wire s0n130,s1n130,notn130;
or (n130,s0n130,s1n130);
not(notn130,n31);
and (s0n130,notn130,n131);
and (s1n130,n31,n134);
wire s0n131,s1n131,notn131;
or (n131,s0n131,s1n131);
not(notn131,n22);
and (s0n131,notn131,n132);
and (s1n131,n22,n133);
nand (n135,n136,n144);
nand (n136,n137,n143);
or (n137,n43,n138);
wire s0n138,s1n138,notn138;
or (n138,s0n138,s1n138);
not(notn138,n66);
and (s0n138,notn138,n139);
and (s1n138,n66,n142);
wire s0n139,s1n139,notn139;
or (n139,s0n139,s1n139);
not(notn139,n57);
and (s0n139,notn139,n140);
and (s1n139,n57,n141);
nand (n143,n138,n43);
not (n144,n145);
nand (n145,n146,n124);
or (n146,n147,n150);
not (n147,n148);
nand (n148,n44,n149);
not (n149,n130);
not (n150,n151);
nand (n151,n43,n130);
nand (n152,n153,n180);
or (n153,n154,n164);
not (n154,n155);
nand (n155,n156,n163);
or (n156,n157,n18);
not (n157,n158);
wire s0n158,s1n158,notn158;
or (n158,s0n158,s1n158);
not(notn158,n31);
and (s0n158,notn158,n159);
and (s1n158,n31,n162);
wire s0n159,s1n159,notn159;
or (n159,s0n159,s1n159);
not(notn159,n22);
and (s0n159,notn159,n160);
and (s1n159,n22,n161);
nand (n163,n18,n157);
not (n164,n165);
nor (n165,n166,n177);
and (n166,n167,n172);
wire s0n167,s1n167,notn167;
or (n167,s0n167,s1n167);
not(notn167,n66);
and (s0n167,notn167,n168);
and (s1n167,n66,n171);
wire s0n168,s1n168,notn168;
or (n168,s0n168,s1n168);
not(notn168,n57);
and (s0n168,notn168,n169);
and (s1n168,n57,n170);
wire s0n172,s1n172,notn172;
or (n172,s0n172,s1n172);
not(notn172,n31);
and (s0n172,notn172,n173);
and (s1n172,n31,n176);
wire s0n173,s1n173,notn173;
or (n173,s0n173,s1n173);
not(notn173,n22);
and (s0n173,notn173,n174);
and (s1n173,n22,n175);
and (n177,n178,n179);
not (n178,n172);
not (n179,n167);
nand (n180,n181,n185);
nor (n181,n155,n182);
nor (n182,n183,n184);
and (n183,n158,n178);
and (n184,n157,n172);
nor (n185,n186,n192);
and (n186,n187,n172);
wire s0n187,s1n187,notn187;
or (n187,s0n187,s1n187);
not(notn187,n66);
and (s0n187,notn187,n188);
and (s1n187,n66,n191);
wire s0n188,s1n188,notn188;
or (n188,s0n188,s1n188);
not(notn188,n57);
and (s0n188,notn188,n189);
and (s1n188,n57,n190);
and (n192,n178,n193);
not (n193,n187);
xor (n194,n195,n260);
xor (n195,n196,n212);
nor (n196,n197,n206);
nor (n197,n198,n204);
and (n198,n199,n178);
wire s0n199,s1n199,notn199;
or (n199,s0n199,s1n199);
not(notn199,n31);
and (s0n199,notn199,n200);
and (s1n199,n31,n203);
wire s0n200,s1n200,notn200;
or (n200,s0n200,s1n200);
not(notn200,n22);
and (s0n200,notn200,n201);
and (s1n200,n22,n202);
and (n204,n205,n172);
not (n205,n199);
not (n206,n207);
wire s0n207,s1n207,notn207;
or (n207,s0n207,s1n207);
not(notn207,n66);
and (s0n207,notn207,n208);
and (s1n207,n66,n211);
wire s0n208,s1n208,notn208;
or (n208,s0n208,s1n208);
not(notn208,n57);
and (s0n208,notn208,n209);
and (s1n208,n57,n210);
nand (n212,n213,n248);
or (n213,n214,n229);
not (n214,n215);
nand (n215,n216,n228);
or (n216,n217,n222);
wire s0n217,s1n217,notn217;
or (n217,s0n217,s1n217);
not(notn217,n31);
and (s0n217,notn217,n218);
and (s1n217,n31,n221);
wire s0n218,s1n218,notn218;
or (n218,s0n218,s1n218);
not(notn218,n22);
and (s0n218,notn218,n219);
and (s1n218,n22,n220);
not (n222,n223);
wire s0n223,s1n223,notn223;
or (n223,s0n223,s1n223);
not(notn223,n66);
and (s0n223,notn223,n224);
and (s1n223,n66,n227);
wire s0n224,s1n224,notn224;
or (n224,s0n224,s1n224);
not(notn224,n57);
and (s0n224,notn224,n225);
and (s1n224,n57,n226);
nand (n228,n222,n217);
nand (n229,n230,n245);
not (n230,n231);
nand (n231,n232,n244);
or (n232,n233,n238);
wire s0n233,s1n233,notn233;
or (n233,s0n233,s1n233);
not(notn233,n31);
and (s0n233,notn233,n234);
and (s1n233,n31,n237);
wire s0n234,s1n234,notn234;
or (n234,s0n234,s1n234);
not(notn234,n22);
and (s0n234,notn234,n235);
and (s1n234,n22,n236);
not (n238,n239);
wire s0n239,s1n239,notn239;
or (n239,s0n239,s1n239);
not(notn239,n31);
and (s0n239,notn239,n240);
and (s1n239,n31,n243);
wire s0n240,s1n240,notn240;
or (n240,s0n240,s1n240);
not(notn240,n22);
and (s0n240,notn240,n241);
and (s1n240,n22,n242);
nand (n244,n238,n233);
nand (n245,n246,n247);
or (n246,n238,n217);
nand (n247,n217,n238);
nand (n248,n249,n231);
not (n249,n250);
nor (n250,n251,n258);
and (n251,n217,n252);
not (n252,n253);
wire s0n253,s1n253,notn253;
or (n253,s0n253,s1n253);
not(notn253,n66);
and (s0n253,notn253,n254);
and (s1n253,n66,n257);
wire s0n254,s1n254,notn254;
or (n254,s0n254,s1n254);
not(notn254,n57);
and (s0n254,notn254,n255);
and (s1n254,n57,n256);
and (n258,n259,n253);
not (n259,n217);
nand (n260,n261,n288);
or (n261,n262,n273);
not (n262,n263);
nand (n263,n264,n271);
or (n264,n265,n233);
not (n265,n266);
wire s0n266,s1n266,notn266;
or (n266,s0n266,s1n266);
not(notn266,n66);
and (s0n266,notn266,n267);
and (s1n266,n66,n270);
wire s0n267,s1n267,notn267;
or (n267,s0n267,s1n267);
not(notn267,n57);
and (s0n267,notn267,n268);
and (s1n267,n57,n269);
or (n271,n266,n272);
not (n272,n233);
not (n273,n274);
nand (n274,n275,n287);
or (n275,n276,n282);
not (n276,n277);
wire s0n277,s1n277,notn277;
or (n277,s0n277,s1n277);
not(notn277,n31);
and (s0n277,notn277,n278);
and (s1n277,n31,n281);
wire s0n278,s1n278,notn278;
or (n278,s0n278,s1n278);
not(notn278,n22);
and (s0n278,notn278,n279);
and (s1n278,n22,n280);
wire s0n282,s1n282,notn282;
or (n282,s0n282,s1n282);
not(notn282,n31);
and (s0n282,notn282,n283);
and (s1n282,n31,n286);
wire s0n283,s1n283,notn283;
or (n283,s0n283,s1n283);
not(notn283,n22);
and (s0n283,notn283,n284);
and (s1n283,n22,n285);
nand (n287,n282,n276);
nand (n288,n289,n298);
nor (n289,n290,n297);
and (n290,n272,n291);
not (n291,n292);
wire s0n292,s1n292,notn292;
or (n292,s0n292,s1n292);
not(notn292,n66);
and (s0n292,notn292,n293);
and (s1n292,n66,n296);
wire s0n293,s1n293,notn293;
or (n293,s0n293,s1n293);
not(notn293,n57);
and (s0n293,notn293,n294);
and (s1n293,n57,n295);
and (n297,n292,n233);
not (n298,n299);
nand (n299,n273,n300);
nand (n300,n301,n302);
or (n301,n272,n277);
nand (n302,n272,n277);
xor (n303,n304,n385);
xor (n304,n305,n341);
nand (n305,n306,n328);
or (n306,n307,n317);
not (n307,n308);
nand (n308,n309,n316);
or (n309,n310,n217);
not (n310,n311);
wire s0n311,s1n311,notn311;
or (n311,s0n311,s1n311);
not(notn311,n31);
and (s0n311,notn311,n312);
and (s1n311,n31,n315);
wire s0n312,s1n312,notn312;
or (n312,s0n312,s1n312);
not(notn312,n22);
and (s0n312,notn312,n313);
and (s1n312,n22,n314);
nand (n316,n217,n310);
not (n317,n318);
nor (n318,n319,n327);
and (n319,n320,n321);
not (n320,n125);
not (n321,n322);
wire s0n322,s1n322,notn322;
or (n322,s0n322,s1n322);
not(notn322,n66);
and (s0n322,notn322,n323);
and (s1n322,n66,n326);
wire s0n323,s1n323,notn323;
or (n323,s0n323,s1n323);
not(notn323,n57);
and (s0n323,notn323,n324);
and (s1n323,n57,n325);
and (n327,n322,n125);
nand (n328,n329,n337);
nand (n329,n330,n336);
or (n330,n320,n331);
wire s0n331,s1n331,notn331;
or (n331,s0n331,s1n331);
not(notn331,n66);
and (s0n331,notn331,n332);
and (s1n331,n66,n335);
wire s0n332,s1n332,notn332;
or (n332,s0n332,s1n332);
not(notn332,n57);
and (s0n332,notn332,n333);
and (s1n332,n57,n334);
nand (n336,n331,n320);
nor (n337,n338,n308);
nor (n338,n339,n340);
and (n339,n320,n311);
and (n340,n125,n310);
nand (n341,n342,n375);
or (n342,n343,n354);
not (n343,n344);
nor (n344,n345,n351);
and (n345,n346,n282);
wire s0n346,s1n346,notn346;
or (n346,s0n346,s1n346);
not(notn346,n66);
and (s0n346,notn346,n347);
and (s1n346,n66,n350);
wire s0n347,s1n347,notn347;
or (n347,s0n347,s1n347);
not(notn347,n57);
and (s0n347,notn347,n348);
and (s1n347,n57,n349);
and (n351,n352,n353);
not (n352,n282);
not (n353,n346);
nand (n354,n355,n366);
or (n355,n356,n364);
not (n356,n357);
nand (n357,n282,n358);
not (n358,n359);
wire s0n359,s1n359,notn359;
or (n359,s0n359,s1n359);
not(notn359,n31);
and (s0n359,notn359,n360);
and (s1n359,n31,n363);
wire s0n360,s1n360,notn360;
or (n360,s0n360,s1n360);
not(notn360,n22);
and (s0n360,notn360,n361);
and (s1n360,n22,n362);
not (n364,n365);
nand (n365,n352,n359);
not (n366,n367);
nand (n367,n368,n374);
or (n368,n369,n358);
wire s0n369,s1n369,notn369;
or (n369,s0n369,s1n369);
not(notn369,n31);
and (s0n369,notn369,n370);
and (s1n369,n31,n373);
wire s0n370,s1n370,notn370;
or (n370,s0n370,s1n370);
not(notn370,n22);
and (s0n370,notn370,n371);
and (s1n370,n22,n372);
nand (n374,n358,n369);
nand (n375,n367,n376);
nor (n376,n377,n383);
and (n377,n378,n282);
wire s0n378,s1n378,notn378;
or (n378,s0n378,s1n378);
not(notn378,n66);
and (s0n378,notn378,n379);
and (s1n378,n66,n382);
wire s0n379,s1n379,notn379;
or (n379,s0n379,s1n379);
not(notn379,n57);
and (s0n379,notn379,n380);
and (s1n379,n57,n381);
and (n383,n352,n384);
not (n384,n378);
nand (n385,n386,n405);
or (n386,n387,n395);
not (n387,n388);
nor (n388,n389,n390);
not (n389,n369);
wire s0n390,s1n390,notn390;
or (n390,s0n390,s1n390);
not(notn390,n31);
and (s0n390,notn390,n391);
and (s1n390,n31,n394);
wire s0n391,s1n391,notn391;
or (n391,s0n391,s1n391);
not(notn391,n22);
and (s0n391,notn391,n392);
and (s1n391,n22,n393);
not (n395,n396);
nand (n396,n397,n404);
or (n397,n369,n398);
not (n398,n399);
wire s0n399,s1n399,notn399;
or (n399,s0n399,s1n399);
not(notn399,n66);
and (s0n399,notn399,n400);
and (s1n399,n66,n403);
wire s0n400,s1n400,notn400;
or (n400,s0n400,s1n400);
not(notn400,n57);
and (s0n400,notn400,n401);
and (s1n400,n57,n402);
nand (n404,n398,n369);
or (n405,n406,n415);
nor (n406,n407,n413);
and (n407,n408,n389);
wire s0n408,s1n408,notn408;
or (n408,s0n408,s1n408);
not(notn408,n66);
and (s0n408,notn408,n409);
and (s1n408,n66,n412);
wire s0n409,s1n409,notn409;
or (n409,s0n409,s1n409);
not(notn409,n57);
and (s0n409,notn409,n410);
and (s1n409,n57,n411);
and (n413,n414,n369);
not (n414,n408);
not (n415,n390);
or (n416,n417,n589);
and (n417,n418,n520);
xor (n418,n419,n461);
or (n419,n420,n460);
and (n420,n421,n442);
xor (n421,n422,n432);
nand (n422,n423,n428);
or (n423,n424,n14);
not (n424,n425);
nand (n425,n426,n427);
or (n426,n40,n187);
nand (n427,n187,n40);
nand (n428,n429,n113);
nand (n429,n430,n431);
or (n430,n40,n167);
nand (n431,n167,n40);
nand (n432,n433,n438);
or (n433,n434,n354);
not (n434,n435);
nand (n435,n436,n437);
or (n436,n352,n292);
nand (n437,n292,n352);
nand (n438,n439,n367);
nand (n439,n440,n441);
or (n440,n282,n265);
nand (n441,n265,n282);
and (n442,n443,n449);
nor (n443,n444,n40);
and (n444,n445,n448);
nand (n445,n446,n43);
not (n446,n447);
and (n447,n207,n33);
nand (n448,n206,n32);
nand (n449,n450,n455);
or (n450,n229,n451);
not (n451,n452);
nand (n452,n453,n454);
or (n453,n259,n118);
nand (n454,n118,n259);
nand (n455,n456,n231);
nand (n456,n457,n459);
or (n457,n217,n458);
not (n458,n331);
nand (n459,n458,n217);
and (n460,n422,n432);
xor (n461,n462,n484);
xor (n462,n463,n470);
nand (n463,n464,n466);
or (n464,n154,n465);
not (n465,n185);
nand (n466,n467,n181);
nor (n467,n468,n469);
and (n468,n207,n172);
and (n469,n178,n206);
xor (n470,n471,n477);
nor (n471,n472,n178);
and (n472,n473,n476);
nand (n473,n474,n40);
not (n474,n475);
and (n475,n207,n158);
nand (n476,n206,n157);
nand (n477,n478,n483);
or (n478,n479,n229);
not (n479,n480);
nand (n480,n481,n482);
or (n481,n259,n322);
nand (n482,n322,n259);
nand (n483,n215,n231);
or (n484,n485,n519);
and (n485,n486,n508);
xor (n486,n487,n497);
nand (n487,n488,n493);
or (n488,n489,n299);
not (n489,n490);
nand (n490,n491,n492);
or (n491,n233,n222);
nand (n492,n222,n233);
nand (n493,n494,n274);
nand (n494,n495,n496);
or (n495,n233,n252);
nand (n496,n252,n233);
nand (n497,n498,n504);
or (n498,n499,n500);
not (n499,n337);
not (n500,n501);
nand (n501,n502,n503);
or (n502,n320,n138);
nand (n503,n138,n320);
nand (n504,n505,n308);
nand (n505,n506,n507);
or (n506,n320,n118);
nand (n507,n118,n320);
nand (n508,n509,n514);
or (n509,n145,n510);
not (n510,n511);
nand (n511,n512,n513);
or (n512,n43,n53);
nand (n513,n53,n43);
nand (n514,n515,n518);
nand (n515,n516,n517);
or (n516,n43,n107);
nand (n517,n107,n43);
not (n518,n124);
and (n519,n487,n497);
or (n520,n521,n588);
and (n521,n522,n574);
xor (n522,n523,n547);
or (n523,n524,n546);
and (n524,n525,n539);
xor (n525,n526,n533);
nand (n526,n527,n532);
or (n527,n528,n145);
not (n528,n529);
nand (n529,n530,n531);
or (n530,n43,n167);
nand (n531,n167,n43);
nand (n532,n518,n511);
nand (n533,n534,n538);
or (n534,n535,n14);
nor (n535,n536,n537);
and (n536,n18,n206);
and (n537,n40,n207);
nand (n538,n425,n113);
nand (n539,n540,n545);
or (n540,n541,n354);
not (n541,n542);
nand (n542,n543,n544);
or (n543,n352,n253);
nand (n544,n253,n352);
nand (n545,n435,n367);
and (n546,n526,n533);
or (n547,n548,n573);
and (n548,n549,n566);
xor (n549,n550,n560);
nand (n550,n551,n556);
or (n551,n552,n387);
not (n552,n553);
nand (n553,n554,n555);
or (n554,n389,n266);
nand (n555,n266,n389);
nand (n556,n557,n390);
nand (n557,n558,n559);
or (n558,n389,n346);
nand (n559,n346,n389);
nand (n560,n561,n565);
nand (n561,n298,n562);
nand (n562,n563,n564);
or (n563,n233,n321);
nand (n564,n321,n233);
nand (n565,n274,n490);
nand (n566,n567,n572);
or (n567,n499,n568);
not (n568,n569);
nand (n569,n570,n571);
or (n570,n320,n107);
nand (n571,n107,n320);
nand (n572,n501,n308);
and (n573,n550,n560);
xor (n574,n575,n581);
xor (n575,n576,n577);
and (n576,n155,n207);
nand (n577,n578,n580);
or (n578,n579,n229);
not (n579,n456);
nand (n580,n480,n231);
nand (n581,n582,n584);
or (n582,n583,n387);
not (n583,n557);
nand (n584,n585,n390);
nor (n585,n586,n587);
and (n586,n389,n384);
and (n587,n378,n369);
and (n588,n523,n547);
and (n589,n419,n461);
xor (n590,n591,n630);
xor (n591,n592,n595);
or (n592,n593,n594);
and (n593,n462,n484);
and (n594,n463,n470);
xor (n595,n596,n614);
xor (n596,n597,n598);
and (n597,n471,n477);
or (n598,n599,n613);
and (n599,n600,n609);
xor (n600,n601,n605);
nand (n601,n602,n604);
or (n602,n603,n387);
not (n603,n585);
nand (n604,n396,n390);
nand (n605,n606,n607);
or (n606,n41,n50);
nand (n607,n608,n429);
not (n608,n14);
nand (n609,n610,n612);
or (n610,n145,n611);
not (n611,n515);
nand (n612,n136,n518);
and (n613,n601,n605);
or (n614,n615,n629);
and (n615,n616,n625);
xor (n616,n617,n621);
nand (n617,n618,n620);
or (n618,n619,n299);
not (n619,n494);
nand (n620,n289,n274);
nand (n621,n622,n624);
or (n622,n499,n623);
not (n623,n505);
nand (n624,n329,n308);
nand (n625,n626,n628);
or (n626,n627,n354);
not (n627,n439);
nand (n628,n367,n344);
and (n629,n617,n621);
or (n630,n631,n638);
and (n631,n632,n637);
xor (n632,n633,n636);
or (n633,n634,n635);
and (n634,n575,n581);
and (n635,n576,n577);
xor (n636,n600,n609);
xor (n637,n616,n625);
and (n638,n633,n636);
not (n639,n640);
or (n640,n641,n700);
and (n641,n642,n699);
xor (n642,n643,n644);
xor (n643,n632,n637);
or (n644,n645,n698);
and (n645,n646,n649);
xor (n646,n647,n648);
xor (n647,n486,n508);
xor (n648,n421,n442);
or (n649,n650,n697);
and (n650,n651,n673);
xor (n651,n652,n653);
xor (n652,n443,n449);
or (n653,n654,n672);
and (n654,n655,n664);
xor (n655,n656,n657);
nor (n656,n206,n41);
nand (n657,n658,n663);
or (n658,n659,n299);
not (n659,n660);
nand (n660,n661,n662);
or (n661,n272,n331);
nand (n662,n331,n272);
nand (n663,n562,n274);
nand (n664,n665,n671);
or (n665,n666,n229);
not (n666,n667);
nand (n667,n668,n670);
or (n668,n217,n669);
not (n669,n138);
nand (n670,n669,n217);
nand (n671,n452,n231);
and (n672,n656,n657);
or (n673,n674,n696);
and (n674,n675,n689);
xor (n675,n676,n683);
nand (n676,n677,n682);
or (n677,n678,n145);
not (n678,n679);
nand (n679,n680,n681);
or (n680,n43,n187);
nand (n681,n43,n187);
nand (n682,n529,n518);
nand (n683,n684,n685);
or (n684,n307,n568);
nand (n685,n686,n337);
nand (n686,n687,n688);
or (n687,n320,n53);
nand (n688,n53,n320);
nand (n689,n690,n695);
or (n690,n387,n691);
not (n691,n692);
nand (n692,n693,n694);
or (n693,n369,n291);
nand (n694,n291,n369);
nand (n695,n553,n390);
and (n696,n676,n683);
and (n697,n652,n653);
and (n698,n647,n648);
xor (n699,n418,n520);
and (n700,n643,n644);
nand (n701,n6,n640);
nand (n702,n703,n934);
nor (n703,n704,n926);
and (n704,n705,n813);
and (n705,n706,n776);
nand (n706,n707,n709);
not (n707,n708);
xor (n708,n642,n699);
not (n709,n710);
or (n710,n711,n775);
and (n711,n712,n715);
xor (n712,n713,n714);
xor (n713,n522,n574);
xor (n714,n646,n649);
or (n715,n716,n774);
and (n716,n717,n720);
xor (n717,n718,n719);
xor (n718,n525,n539);
xor (n719,n549,n566);
or (n720,n721,n773);
and (n721,n722,n748);
xor (n722,n723,n730);
nand (n723,n724,n729);
or (n724,n725,n354);
not (n725,n726);
nand (n726,n727,n728);
or (n727,n352,n223);
nand (n728,n223,n352);
nand (n729,n542,n367);
nor (n730,n731,n740);
not (n731,n732);
nand (n732,n733,n739);
or (n733,n734,n299);
not (n734,n735);
nand (n735,n736,n738);
or (n736,n233,n737);
not (n737,n118);
nand (n738,n737,n233);
nand (n739,n660,n274);
nand (n740,n741,n44);
or (n741,n742,n744);
not (n742,n743);
nand (n743,n206,n149);
not (n744,n745);
nand (n745,n746,n320);
not (n746,n747);
and (n747,n207,n130);
or (n748,n749,n772);
and (n749,n750,n765);
xor (n750,n751,n758);
nand (n751,n752,n753);
or (n752,n230,n666);
nand (n753,n754,n757);
nand (n754,n755,n756);
or (n755,n259,n107);
nand (n756,n107,n259);
not (n757,n229);
nand (n758,n759,n764);
or (n759,n760,n145);
not (n760,n761);
nor (n761,n762,n763);
and (n762,n43,n206);
and (n763,n207,n44);
nand (n764,n679,n518);
nand (n765,n766,n768);
or (n766,n307,n767);
not (n767,n686);
nand (n768,n769,n337);
nand (n769,n770,n771);
or (n770,n320,n167);
nand (n771,n167,n320);
and (n772,n751,n758);
and (n773,n723,n730);
and (n774,n718,n719);
and (n775,n713,n714);
not (n776,n777);
nor (n777,n778,n779);
xor (n778,n712,n715);
or (n779,n780,n812);
and (n780,n781,n811);
xor (n781,n782,n783);
xor (n782,n651,n673);
or (n783,n784,n810);
and (n784,n785,n788);
xor (n785,n786,n787);
xor (n786,n675,n689);
xor (n787,n655,n664);
or (n788,n789,n809);
and (n789,n790,n805);
xor (n790,n791,n798);
nand (n791,n792,n797);
or (n792,n793,n354);
not (n793,n794);
nand (n794,n795,n796);
or (n795,n352,n322);
nand (n796,n322,n352);
nand (n797,n367,n726);
nand (n798,n799,n804);
or (n799,n800,n387);
not (n800,n801);
nand (n801,n802,n803);
or (n802,n369,n252);
nand (n803,n252,n369);
nand (n804,n692,n390);
nand (n805,n806,n808);
or (n806,n807,n731);
not (n807,n740);
or (n808,n740,n732);
and (n809,n791,n798);
and (n810,n786,n787);
xor (n811,n717,n720);
and (n812,n782,n783);
nand (n813,n814,n925);
or (n814,n815,n873);
nor (n815,n816,n817);
xor (n816,n781,n811);
or (n817,n818,n872);
and (n818,n819,n871);
xor (n819,n820,n821);
xor (n820,n722,n748);
or (n821,n822,n870);
and (n822,n823,n869);
xor (n823,n824,n850);
or (n824,n825,n849);
and (n825,n826,n842);
xor (n826,n827,n834);
nand (n827,n828,n833);
or (n828,n829,n499);
not (n829,n830);
nand (n830,n831,n832);
or (n831,n125,n193);
nand (n832,n193,n125);
nand (n833,n769,n308);
nand (n834,n835,n837);
or (n835,n230,n836);
not (n836,n754);
nand (n837,n757,n838);
nand (n838,n839,n841);
or (n839,n217,n840);
not (n840,n53);
nand (n841,n840,n217);
nand (n842,n843,n848);
or (n843,n844,n354);
not (n844,n845);
nor (n845,n846,n847);
and (n846,n331,n282);
and (n847,n352,n458);
nand (n848,n794,n367);
and (n849,n827,n834);
or (n850,n851,n868);
and (n851,n852,n861);
xor (n852,n853,n854);
nor (n853,n206,n124);
nand (n854,n855,n860);
or (n855,n299,n856);
not (n856,n857);
nand (n857,n858,n859);
or (n858,n233,n669);
nand (n859,n669,n233);
nand (n860,n735,n274);
nand (n861,n862,n867);
or (n862,n863,n387);
not (n863,n864);
nand (n864,n865,n866);
or (n865,n369,n222);
nand (n866,n222,n369);
nand (n867,n801,n390);
and (n868,n853,n854);
xor (n869,n750,n765);
and (n870,n824,n850);
xor (n871,n785,n788);
and (n872,n820,n821);
nand (n873,n874,n875);
xor (n874,n819,n871);
or (n875,n876,n924);
and (n876,n877,n880);
xor (n877,n878,n879);
xor (n878,n790,n805);
xor (n879,n823,n869);
or (n880,n881,n923);
and (n881,n882,n922);
xor (n882,n883,n897);
and (n883,n884,n890);
nor (n884,n885,n320);
and (n885,n886,n889);
nand (n886,n887,n259);
not (n887,n888);
and (n888,n207,n311);
nand (n889,n206,n310);
nand (n890,n891,n896);
or (n891,n299,n892);
not (n892,n893);
nand (n893,n894,n895);
or (n894,n272,n107);
nand (n895,n107,n272);
nand (n896,n857,n274);
or (n897,n898,n921);
and (n898,n899,n914);
xor (n899,n900,n907);
nand (n900,n901,n906);
or (n901,n387,n902);
not (n902,n903);
nand (n903,n904,n905);
or (n904,n369,n321);
nand (n905,n321,n369);
nand (n906,n864,n390);
nand (n907,n908,n913);
or (n908,n909,n354);
not (n909,n910);
nand (n910,n911,n912);
or (n911,n352,n118);
nand (n912,n118,n352);
nand (n913,n845,n367);
nand (n914,n915,n920);
or (n915,n916,n229);
not (n916,n917);
nand (n917,n918,n919);
or (n918,n259,n167);
nand (n919,n167,n259);
nand (n920,n838,n231);
and (n921,n900,n907);
xor (n922,n852,n861);
and (n923,n883,n897);
and (n924,n878,n879);
nand (n925,n816,n817);
nand (n926,n927,n933);
or (n927,n928,n932);
not (n928,n929);
nor (n929,n930,n931);
not (n930,n778);
not (n931,n779);
not (n932,n706);
nand (n933,n708,n710);
nand (n934,n706,n935,n1247,n776);
nand (n935,n936,n1231,n1237);
nand (n936,n937,n978,n1085);
nand (n937,n938,n940);
not (n938,n939);
xor (n939,n877,n880);
not (n940,n941);
or (n941,n942,n977);
and (n942,n943,n976);
xor (n943,n944,n945);
xor (n944,n826,n842);
or (n945,n946,n975);
and (n946,n947,n956);
xor (n947,n948,n955);
nand (n948,n949,n954);
or (n949,n499,n950);
not (n950,n951);
nor (n951,n952,n953);
and (n952,n207,n125);
and (n953,n320,n206);
nand (n954,n308,n830);
xor (n955,n884,n890);
or (n956,n957,n974);
and (n957,n958,n967);
xor (n958,n959,n960);
and (n959,n308,n207);
nand (n960,n961,n966);
or (n961,n354,n962);
not (n962,n963);
nand (n963,n964,n965);
or (n964,n282,n669);
nand (n965,n669,n282);
nand (n966,n910,n367);
nand (n967,n968,n973);
or (n968,n387,n969);
not (n969,n970);
nor (n970,n971,n972);
and (n971,n331,n369);
and (n972,n389,n458);
nand (n973,n903,n390);
and (n974,n959,n960);
and (n975,n948,n955);
xor (n976,n882,n922);
and (n977,n944,n945);
not (n978,n979);
nand (n979,n980,n1078);
nor (n980,n981,n1048);
nor (n981,n982,n1018);
xor (n982,n983,n1017);
xor (n983,n984,n985);
xor (n984,n899,n914);
or (n985,n986,n1016);
and (n986,n987,n1002);
xor (n987,n988,n995);
nand (n988,n989,n994);
or (n989,n990,n229);
not (n990,n991);
nand (n991,n992,n993);
or (n992,n259,n187);
nand (n993,n187,n259);
nand (n994,n917,n231);
nand (n995,n996,n1001);
or (n996,n997,n299);
not (n997,n998);
nand (n998,n999,n1000);
or (n999,n272,n53);
nand (n1000,n53,n272);
nand (n1001,n893,n274);
and (n1002,n1003,n1010);
nand (n1003,n1004,n1009);
or (n1004,n1005,n354);
not (n1005,n1006);
nand (n1006,n1007,n1008);
or (n1007,n352,n107);
nand (n1008,n107,n352);
nand (n1009,n963,n367);
nor (n1010,n1011,n259);
and (n1011,n1012,n1015);
nand (n1012,n1013,n272);
not (n1013,n1014);
and (n1014,n207,n239);
nand (n1015,n206,n238);
and (n1016,n988,n995);
xor (n1017,n947,n956);
or (n1018,n1019,n1047);
and (n1019,n1020,n1046);
xor (n1020,n1021,n1045);
or (n1021,n1022,n1044);
and (n1022,n1023,n1037);
xor (n1023,n1024,n1030);
nand (n1024,n1025,n1029);
nand (n1025,n1026,n388);
nand (n1026,n1027,n1028);
or (n1027,n389,n118);
nand (n1028,n118,n389);
nand (n1029,n970,n390);
nand (n1030,n1031,n1036);
or (n1031,n1032,n229);
not (n1032,n1033);
nand (n1033,n1034,n1035);
or (n1034,n217,n206);
or (n1035,n207,n259);
nand (n1036,n991,n231);
nand (n1037,n1038,n1043);
or (n1038,n1039,n299);
not (n1039,n1040);
nand (n1040,n1041,n1042);
or (n1041,n272,n167);
nand (n1042,n167,n272);
nand (n1043,n998,n274);
and (n1044,n1024,n1030);
xor (n1045,n958,n967);
xor (n1046,n987,n1002);
and (n1047,n1021,n1045);
nor (n1048,n1049,n1050);
xor (n1049,n1020,n1046);
or (n1050,n1051,n1077);
and (n1051,n1052,n1076);
xor (n1052,n1053,n1057);
nand (n1053,n1054,n1056);
or (n1054,n1010,n1055);
not (n1055,n1003);
nand (n1056,n1055,n1010);
or (n1057,n1058,n1075);
and (n1058,n1059,n1068);
xor (n1059,n1060,n1061);
nor (n1060,n206,n230);
nand (n1061,n1062,n1067);
or (n1062,n1063,n354);
not (n1063,n1064);
nand (n1064,n1065,n1066);
or (n1065,n282,n840);
nand (n1066,n840,n282);
nand (n1067,n1006,n367);
nand (n1068,n1069,n1074);
or (n1069,n1070,n299);
not (n1070,n1071);
nand (n1071,n1072,n1073);
or (n1072,n272,n187);
nand (n1073,n187,n272);
nand (n1074,n1040,n274);
and (n1075,n1060,n1061);
xor (n1076,n1023,n1037);
and (n1077,n1053,n1057);
nand (n1078,n1079,n1081);
not (n1079,n1080);
xor (n1080,n943,n976);
not (n1081,n1082);
or (n1082,n1083,n1084);
and (n1083,n983,n1017);
and (n1084,n984,n985);
nand (n1085,n1086,n1230);
or (n1086,n1087,n1118);
not (n1087,n1088);
nand (n1088,n1089,n1091);
not (n1089,n1090);
xor (n1090,n1052,n1076);
not (n1091,n1092);
or (n1092,n1093,n1117);
and (n1093,n1094,n1116);
xor (n1094,n1095,n1102);
nand (n1095,n1096,n1101);
or (n1096,n387,n1097);
not (n1097,n1098);
nand (n1098,n1099,n1100);
or (n1099,n369,n669);
nand (n1100,n369,n669);
nand (n1101,n1026,n390);
and (n1102,n1103,n1110);
nand (n1103,n1104,n1105);
or (n1104,n366,n1063);
nand (n1105,n1106,n1107);
not (n1106,n354);
nand (n1107,n1108,n1109);
or (n1108,n352,n167);
nand (n1109,n167,n352);
nor (n1110,n1111,n272);
and (n1111,n1112,n1115);
nand (n1112,n1113,n352);
not (n1113,n1114);
and (n1114,n207,n277);
nand (n1115,n206,n276);
xor (n1116,n1059,n1068);
and (n1117,n1095,n1102);
not (n1118,n1119);
nand (n1119,n1120,n1229);
or (n1120,n1121,n1148);
not (n1121,n1122);
nand (n1122,n1123,n1125);
not (n1123,n1124);
xor (n1124,n1094,n1116);
not (n1125,n1126);
or (n1126,n1127,n1147);
and (n1127,n1128,n1143);
xor (n1128,n1129,n1136);
nand (n1129,n1130,n1135);
or (n1130,n1131,n299);
not (n1131,n1132);
nor (n1132,n1133,n1134);
and (n1133,n272,n206);
and (n1134,n207,n233);
nand (n1135,n274,n1071);
nand (n1136,n1137,n1138);
or (n1137,n415,n1097);
nand (n1138,n1139,n388);
nand (n1139,n1140,n1142);
or (n1140,n369,n1141);
not (n1141,n107);
nand (n1142,n369,n1141);
nand (n1143,n1144,n1146);
or (n1144,n1110,n1145);
not (n1145,n1103);
nand (n1146,n1145,n1110);
and (n1147,n1129,n1136);
not (n1148,n1149);
nand (n1149,n1150,n1228);
or (n1150,n1151,n1223);
nor (n1151,n1152,n1222);
and (n1152,n1153,n1189);
nand (n1153,n1154,n1172);
not (n1154,n1155);
xor (n1155,n1156,n1165);
xor (n1156,n1157,n1158);
and (n1157,n274,n207);
nand (n1158,n1159,n1161);
or (n1159,n415,n1160);
not (n1160,n1139);
nand (n1161,n1162,n388);
nand (n1162,n1163,n1164);
or (n1163,n369,n840);
nand (n1164,n840,n369);
nand (n1165,n1166,n1171);
or (n1166,n1167,n354);
not (n1167,n1168);
nand (n1168,n1169,n1170);
or (n1169,n352,n187);
nand (n1170,n187,n352);
nand (n1171,n1107,n367);
nand (n1172,n1173,n1182);
not (n1173,n1174);
nand (n1174,n1175,n282);
or (n1175,n1176,n1178);
not (n1176,n1177);
nand (n1177,n358,n206);
not (n1178,n1179);
nand (n1179,n1180,n389);
not (n1180,n1181);
and (n1181,n207,n359);
nand (n1182,n1183,n1185);
or (n1183,n415,n1184);
not (n1184,n1162);
nand (n1185,n1186,n388);
nand (n1186,n1187,n1188);
or (n1187,n389,n167);
nand (n1188,n167,n389);
nand (n1189,n1190,n1221);
nand (n1190,n1191,n1202);
or (n1191,n1192,n1195);
nand (n1192,n1193,n1194);
or (n1193,n1174,n1182);
nand (n1194,n1182,n1174);
nand (n1195,n1196,n1201);
or (n1196,n1197,n354);
not (n1197,n1198);
nor (n1198,n1199,n1200);
and (n1199,n352,n206);
and (n1200,n207,n282);
nand (n1201,n367,n1168);
or (n1202,n1203,n1220);
and (n1203,n1204,n1213);
xor (n1204,n1205,n1206);
and (n1205,n207,n367);
nand (n1206,n1207,n1209);
or (n1207,n415,n1208);
not (n1208,n1186);
nand (n1209,n1210,n388);
nand (n1210,n1211,n1212);
or (n1211,n389,n187);
nand (n1212,n187,n389);
nor (n1213,n1214,n1217);
nor (n1214,n1215,n1216);
and (n1215,n388,n206);
and (n1216,n1210,n390);
nand (n1217,n1218,n369);
not (n1218,n1219);
and (n1219,n207,n390);
and (n1220,n1205,n1206);
nand (n1221,n1192,n1195);
nor (n1222,n1154,n1172);
nor (n1223,n1224,n1225);
xor (n1224,n1128,n1143);
or (n1225,n1226,n1227);
and (n1226,n1156,n1165);
and (n1227,n1157,n1158);
nand (n1228,n1224,n1225);
nand (n1229,n1124,n1126);
nand (n1230,n1090,n1092);
nand (n1231,n1232,n937);
or (n1232,n1233,n1235);
not (n1233,n1234);
nand (n1234,n1080,n1082);
not (n1235,n1236);
nand (n1236,n939,n941);
nand (n1237,n937,n1238);
nor (n1238,n1239,n1246);
nand (n1239,n1240,n1245);
or (n1240,n1241,n1243);
not (n1241,n1242);
nand (n1242,n1049,n1050);
not (n1243,n1244);
nand (n1244,n982,n1018);
not (n1245,n981);
not (n1246,n1078);
not (n1247,n1248);
nand (n1248,n1249,n1250);
not (n1249,n815);
or (n1250,n874,n875);
nand (n1251,n702,n3);
not (n1252,n1253);
or (n1253,n1254,n1351,n1363);
and (n1254,n1255,n1341);
xor (n1255,n1256,n1335);
xor (n1256,n1257,n1329);
xor (n1257,n1258,n1320);
and (n1258,n1259,n1270);
wire s0n1259,s1n1259,notn1259;
or (n1259,s0n1259,s1n1259);
not(notn1259,n1262);
and (s0n1259,notn1259,n1260);
and (s1n1259,n1262,n1261);
and (n1262,n1263,n1268);
and (n1263,n1264,n1266);
not (n1264,n1265);
not (n1266,n1267);
not (n1268,n1269);
wire s0n1270,s1n1270,notn1270;
or (n1270,s0n1270,s1n1270);
not(notn1270,n1283);
and (s0n1270,notn1270,n1271);
and (s1n1270,n1283,n1282);
wire s0n1271,s1n1271,notn1271;
or (n1271,s0n1271,s1n1271);
not(notn1271,n1274);
and (s0n1271,notn1271,n1272);
and (s1n1271,n1274,n1273);
and (n1274,n1275,n1280);
and (n1275,n1276,n1278);
not (n1276,n1277);
not (n1278,n1279);
not (n1280,n1281);
and (n1283,n1284,n1286);
not (n1284,n1285);
or (n1286,n1287,n1288);
and (n1288,n1289,n1290);
or (n1290,n1291,n1292,n1293,n1294,n1295,n1296,n1297,n1298,n1299,n1300,n1301,n1302,n1303,n1304,n1305,n1306,n1307,n1308,n1309,n1310,n1311,n1312,n1313,n1314,n1315,n1316,n1317,n1318,n1319);
and (n1320,n1321,n1324);
wire s0n1321,s1n1321,notn1321;
or (n1321,s0n1321,s1n1321);
not(notn1321,n1262);
and (s0n1321,notn1321,n1322);
and (s1n1321,n1262,n1323);
wire s0n1324,s1n1324,notn1324;
or (n1324,s0n1324,s1n1324);
not(notn1324,n1283);
and (s0n1324,notn1324,n1325);
and (s1n1324,n1283,n1328);
wire s0n1325,s1n1325,notn1325;
or (n1325,s0n1325,s1n1325);
not(notn1325,n1274);
and (s0n1325,notn1325,n1326);
and (s1n1325,n1274,n1327);
and (n1329,n1330,n1331);
and (n1330,n1321,n1270);
and (n1331,n1332,n1324);
wire s0n1332,s1n1332,notn1332;
or (n1332,s0n1332,s1n1332);
not(notn1332,n1262);
and (s0n1332,notn1332,n1333);
and (s1n1332,n1262,n1334);
and (n1335,n1332,n1336);
wire s0n1336,s1n1336,notn1336;
or (n1336,s0n1336,s1n1336);
not(notn1336,n1283);
and (s0n1336,notn1336,n1337);
and (s1n1336,n1283,n1340);
wire s0n1337,s1n1337,notn1337;
or (n1337,s0n1337,s1n1337);
not(notn1337,n1274);
and (s0n1337,notn1337,n1338);
and (s1n1337,n1274,n1339);
not (n1341,n1342);
xor (n1342,n1343,n1350);
xor (n1343,n1344,n1347);
xor (n1344,n1345,n1346);
and (n1345,n360,n207);
and (n1346,n370,n187);
and (n1347,n1348,n1349);
and (n1348,n370,n207);
and (n1349,n391,n187);
and (n1350,n391,n167);
and (n1351,n1341,n1352);
or (n1352,n1353,n1357,n1362);
and (n1353,n1354,n1355);
xor (n1354,n1330,n1331);
not (n1355,n1356);
xor (n1356,n1348,n1349);
and (n1357,n1355,n1358);
or (n1358,n1359,n1360);
and (n1359,n1332,n1270);
not (n1360,n1361);
and (n1361,n391,n207);
and (n1362,n1354,n1358);
and (n1363,n1255,n1352);
and (n1364,n1365,n2578);
xor (n1365,n1366,n2558);
xor (n1366,n1367,n2474);
xor (n1367,n1368,n2449);
xor (n1368,n1369,n2370);
xor (n1369,n1370,n2340);
xor (n1370,n1371,n2266);
xor (n1371,n1372,n2231);
xor (n1372,n1373,n2164);
xor (n1373,n1374,n2124);
xor (n1374,n1375,n2063);
xor (n1375,n1376,n2018);
xor (n1376,n1377,n1964);
xor (n1377,n1378,n1914);
xor (n1378,n1379,n1865);
xor (n1379,n1380,n1810);
xor (n1380,n1381,n1768);
xor (n1381,n1382,n1708);
xor (n1382,n1383,n1669);
xor (n1383,n1384,n1604);
xor (n1384,n1385,n1572);
xor (n1385,n1386,n1468);
xor (n1386,n1387,n1443);
xor (n1387,n1388,n1442);
xor (n1388,n1389,n1423);
xor (n1389,n1390,n1422);
xor (n1390,n1391,n1409);
xor (n1391,n1392,n1408);
xor (n1392,n1393,n1401);
xor (n1393,n1394,n1400);
xor (n1394,n1395,n1396);
and (n1395,n1252,n1219);
and (n1396,n1252,n1397);
xor (n1397,n1398,n1399);
and (n1398,n187,n390);
and (n1399,n207,n369);
and (n1400,n1395,n1396);
and (n1401,n1252,n1402);
xor (n1402,n1403,n1181);
xor (n1403,n1404,n1407);
xor (n1404,n1405,n1406);
and (n1405,n167,n390);
and (n1406,n187,n369);
and (n1407,n1398,n1399);
and (n1408,n1393,n1401);
and (n1409,n1252,n1410);
xor (n1410,n1411,n1200);
xor (n1411,n1412,n1421);
xor (n1412,n1413,n1420);
xor (n1413,n1414,n1417);
xor (n1414,n1415,n1416);
and (n1415,n53,n390);
and (n1416,n167,n369);
or (n1417,n1418,n1419);
and (n1418,n1405,n1406);
and (n1419,n1404,n1407);
and (n1420,n187,n359);
and (n1421,n1403,n1181);
and (n1422,n1391,n1409);
and (n1423,n1252,n1424);
xor (n1424,n1425,n1114);
xor (n1425,n1426,n1441);
xor (n1426,n1427,n1440);
xor (n1427,n1428,n1437);
xor (n1428,n1429,n1436);
xor (n1429,n1430,n1433);
xor (n1430,n1431,n1432);
and (n1431,n107,n390);
and (n1432,n53,n369);
or (n1433,n1434,n1435);
and (n1434,n1415,n1416);
and (n1435,n1414,n1417);
and (n1436,n167,n359);
or (n1437,n1438,n1439);
and (n1438,n1413,n1420);
and (n1439,n1412,n1421);
and (n1440,n187,n282);
and (n1441,n1411,n1200);
and (n1442,n1389,n1423);
and (n1443,n1252,n1444);
xor (n1444,n1445,n1134);
xor (n1445,n1446,n1467);
xor (n1446,n1447,n1466);
xor (n1447,n1448,n1463);
xor (n1448,n1449,n1462);
xor (n1449,n1450,n1459);
xor (n1450,n1451,n1458);
xor (n1451,n1452,n1455);
xor (n1452,n1453,n1454);
and (n1453,n138,n390);
and (n1454,n107,n369);
or (n1455,n1456,n1457);
and (n1456,n1431,n1432);
and (n1457,n1430,n1433);
and (n1458,n53,n359);
or (n1459,n1460,n1461);
and (n1460,n1429,n1436);
and (n1461,n1428,n1437);
and (n1462,n167,n282);
or (n1463,n1464,n1465);
and (n1464,n1427,n1440);
and (n1465,n1426,n1441);
and (n1466,n187,n277);
and (n1467,n1425,n1114);
or (n1468,n1469,n1470);
and (n1469,n1387,n1443);
and (n1470,n1386,n1471);
or (n1471,n1469,n1472);
and (n1472,n1386,n1473);
or (n1473,n1469,n1474);
and (n1474,n1386,n1475);
or (n1475,n1469,n1476);
and (n1476,n1386,n1477);
or (n1477,n1469,n1478);
and (n1478,n1386,n1479);
or (n1479,n1469,n1480);
and (n1480,n1386,n1481);
or (n1481,n1469,n1482);
and (n1482,n1386,n1483);
or (n1483,n1469,n1484);
and (n1484,n1386,n1485);
or (n1485,n1469,n1486);
and (n1486,n1386,n1487);
or (n1487,n1469,n1488);
and (n1488,n1386,n1489);
or (n1489,n1469,n1490);
and (n1490,n1386,n1491);
or (n1491,n1492,n1561);
and (n1492,n1493,n1560);
xor (n1493,n1388,n1494);
or (n1494,n1495,n1549);
and (n1495,n1496,n1548);
xor (n1496,n1390,n1497);
or (n1497,n1498,n1536);
and (n1498,n1499,n1535);
xor (n1499,n1392,n1500);
or (n1500,n1501,n1523);
and (n1501,n1502,n1522);
xor (n1502,n1394,n1503);
or (n1503,n1504,n1508);
and (n1504,n1395,n1505);
and (n1505,n1506,n1397);
xor (n1506,n1507,n1352);
xor (n1507,n1255,n1341);
and (n1508,n1509,n1510);
xor (n1509,n1395,n1505);
or (n1510,n1511,n1516);
and (n1511,n1512,n1513);
and (n1512,n1506,n1219);
and (n1513,n1514,n1397);
xor (n1514,n1515,n1358);
xor (n1515,n1354,n1355);
and (n1516,n1517,n1518);
xor (n1517,n1512,n1513);
and (n1518,n1519,n1520);
and (n1519,n1514,n1219);
and (n1520,n1521,n1397);
xor (n1521,n1359,n1361);
and (n1522,n1506,n1402);
and (n1523,n1524,n1525);
xor (n1524,n1502,n1522);
or (n1525,n1526,n1529);
and (n1526,n1527,n1528);
xor (n1527,n1509,n1510);
and (n1528,n1514,n1402);
and (n1529,n1530,n1531);
xor (n1530,n1527,n1528);
and (n1531,n1532,n1533);
xor (n1532,n1517,n1518);
not (n1533,n1534);
nand (n1534,n1402,n1521);
and (n1535,n1506,n1410);
and (n1536,n1537,n1538);
xor (n1537,n1499,n1535);
or (n1538,n1539,n1542);
and (n1539,n1540,n1541);
xor (n1540,n1524,n1525);
and (n1541,n1514,n1410);
and (n1542,n1543,n1544);
xor (n1543,n1540,n1541);
and (n1544,n1545,n1546);
xor (n1545,n1530,n1531);
not (n1546,n1547);
nand (n1547,n1410,n1521);
and (n1548,n1506,n1424);
and (n1549,n1550,n1551);
xor (n1550,n1496,n1548);
or (n1551,n1552,n1555);
and (n1552,n1553,n1554);
xor (n1553,n1537,n1538);
and (n1554,n1514,n1424);
and (n1555,n1556,n1557);
xor (n1556,n1553,n1554);
and (n1557,n1558,n1559);
xor (n1558,n1543,n1544);
and (n1559,n1424,n1521);
and (n1560,n1506,n1444);
and (n1561,n1562,n1563);
xor (n1562,n1493,n1560);
or (n1563,n1564,n1567);
and (n1564,n1565,n1566);
xor (n1565,n1550,n1551);
and (n1566,n1444,n1514);
and (n1567,n1568,n1569);
xor (n1568,n1565,n1566);
and (n1569,n1570,n1571);
xor (n1570,n1556,n1557);
and (n1571,n1444,n1521);
not (n1572,n1573);
nand (n1573,n1574,n1252);
xor (n1574,n1575,n1014);
xor (n1575,n1576,n1603);
xor (n1576,n1577,n1602);
xor (n1577,n1578,n1599);
xor (n1578,n1579,n1598);
xor (n1579,n1580,n1595);
xor (n1580,n1581,n1594);
xor (n1581,n1582,n1591);
xor (n1582,n1583,n1590);
xor (n1583,n1584,n1587);
xor (n1584,n1585,n1586);
and (n1585,n118,n390);
and (n1586,n138,n369);
or (n1587,n1588,n1589);
and (n1588,n1453,n1454);
and (n1589,n1452,n1455);
and (n1590,n107,n359);
or (n1591,n1592,n1593);
and (n1592,n1451,n1458);
and (n1593,n1450,n1459);
and (n1594,n53,n282);
or (n1595,n1596,n1597);
and (n1596,n1449,n1462);
and (n1597,n1448,n1463);
and (n1598,n167,n277);
or (n1599,n1600,n1601);
and (n1600,n1447,n1466);
and (n1601,n1446,n1467);
and (n1602,n187,n233);
and (n1603,n1445,n1134);
or (n1604,n1605,n1607);
and (n1605,n1606,n1572);
xor (n1606,n1386,n1471);
and (n1607,n1608,n1609);
xor (n1608,n1606,n1572);
or (n1609,n1610,n1612);
and (n1610,n1611,n1572);
xor (n1611,n1386,n1473);
and (n1612,n1613,n1614);
xor (n1613,n1611,n1572);
or (n1614,n1615,n1617);
and (n1615,n1616,n1572);
xor (n1616,n1386,n1475);
and (n1617,n1618,n1619);
xor (n1618,n1616,n1572);
or (n1619,n1620,n1622);
and (n1620,n1621,n1572);
xor (n1621,n1386,n1477);
and (n1622,n1623,n1624);
xor (n1623,n1621,n1572);
or (n1624,n1625,n1627);
and (n1625,n1626,n1572);
xor (n1626,n1386,n1479);
and (n1627,n1628,n1629);
xor (n1628,n1626,n1572);
or (n1629,n1630,n1632);
and (n1630,n1631,n1572);
xor (n1631,n1386,n1481);
and (n1632,n1633,n1634);
xor (n1633,n1631,n1572);
or (n1634,n1635,n1637);
and (n1635,n1636,n1572);
xor (n1636,n1386,n1483);
and (n1637,n1638,n1639);
xor (n1638,n1636,n1572);
or (n1639,n1640,n1642);
and (n1640,n1641,n1572);
xor (n1641,n1386,n1485);
and (n1642,n1643,n1644);
xor (n1643,n1641,n1572);
or (n1644,n1645,n1647);
and (n1645,n1646,n1572);
xor (n1646,n1386,n1487);
and (n1647,n1648,n1649);
xor (n1648,n1646,n1572);
or (n1649,n1650,n1652);
and (n1650,n1651,n1572);
xor (n1651,n1386,n1489);
and (n1652,n1653,n1654);
xor (n1653,n1651,n1572);
or (n1654,n1655,n1658);
and (n1655,n1656,n1657);
xor (n1656,n1386,n1491);
and (n1657,n1574,n1506);
and (n1658,n1659,n1660);
xor (n1659,n1656,n1657);
or (n1660,n1661,n1664);
and (n1661,n1662,n1663);
xor (n1662,n1562,n1563);
and (n1663,n1514,n1574);
and (n1664,n1665,n1666);
xor (n1665,n1662,n1663);
and (n1666,n1667,n1668);
xor (n1667,n1568,n1569);
and (n1668,n1574,n1521);
not (n1669,n1670);
nand (n1670,n1671,n1252);
xor (n1671,n1672,n1707);
xor (n1672,n1673,n1706);
xor (n1673,n1674,n1705);
xor (n1674,n1675,n1702);
xor (n1675,n1676,n1701);
xor (n1676,n1677,n1698);
xor (n1677,n1678,n1697);
xor (n1678,n1679,n1694);
xor (n1679,n1680,n1693);
xor (n1680,n1681,n1690);
xor (n1681,n1682,n1689);
xor (n1682,n1683,n1686);
xor (n1683,n1684,n1685);
and (n1684,n331,n390);
and (n1685,n118,n369);
or (n1686,n1687,n1688);
and (n1687,n1585,n1586);
and (n1688,n1584,n1587);
and (n1689,n138,n359);
or (n1690,n1691,n1692);
and (n1691,n1583,n1590);
and (n1692,n1582,n1591);
and (n1693,n107,n282);
or (n1694,n1695,n1696);
and (n1695,n1581,n1594);
and (n1696,n1580,n1595);
and (n1697,n53,n277);
or (n1698,n1699,n1700);
and (n1699,n1579,n1598);
and (n1700,n1578,n1599);
and (n1701,n167,n233);
or (n1702,n1703,n1704);
and (n1703,n1577,n1602);
and (n1704,n1576,n1603);
and (n1705,n187,n239);
and (n1706,n1575,n1014);
and (n1707,n207,n217);
or (n1708,n1709,n1711);
and (n1709,n1710,n1669);
xor (n1710,n1608,n1609);
and (n1711,n1712,n1713);
xor (n1712,n1710,n1669);
or (n1713,n1714,n1716);
and (n1714,n1715,n1669);
xor (n1715,n1613,n1614);
and (n1716,n1717,n1718);
xor (n1717,n1715,n1669);
or (n1718,n1719,n1721);
and (n1719,n1720,n1669);
xor (n1720,n1618,n1619);
and (n1721,n1722,n1723);
xor (n1722,n1720,n1669);
or (n1723,n1724,n1726);
and (n1724,n1725,n1669);
xor (n1725,n1623,n1624);
and (n1726,n1727,n1728);
xor (n1727,n1725,n1669);
or (n1728,n1729,n1731);
and (n1729,n1730,n1669);
xor (n1730,n1628,n1629);
and (n1731,n1732,n1733);
xor (n1732,n1730,n1669);
or (n1733,n1734,n1736);
and (n1734,n1735,n1669);
xor (n1735,n1633,n1634);
and (n1736,n1737,n1738);
xor (n1737,n1735,n1669);
or (n1738,n1739,n1741);
and (n1739,n1740,n1669);
xor (n1740,n1638,n1639);
and (n1741,n1742,n1743);
xor (n1742,n1740,n1669);
or (n1743,n1744,n1746);
and (n1744,n1745,n1669);
xor (n1745,n1643,n1644);
and (n1746,n1747,n1748);
xor (n1747,n1745,n1669);
or (n1748,n1749,n1751);
and (n1749,n1750,n1669);
xor (n1750,n1648,n1649);
and (n1751,n1752,n1753);
xor (n1752,n1750,n1669);
or (n1753,n1754,n1757);
and (n1754,n1755,n1756);
xor (n1755,n1653,n1654);
and (n1756,n1671,n1506);
and (n1757,n1758,n1759);
xor (n1758,n1755,n1756);
or (n1759,n1760,n1763);
and (n1760,n1761,n1762);
xor (n1761,n1659,n1660);
and (n1762,n1514,n1671);
and (n1763,n1764,n1765);
xor (n1764,n1761,n1762);
and (n1765,n1766,n1767);
xor (n1766,n1665,n1666);
and (n1767,n1521,n1671);
and (n1768,n1252,n1769);
xor (n1769,n1770,n888);
xor (n1770,n1771,n1809);
xor (n1771,n1772,n1808);
xor (n1772,n1773,n1805);
xor (n1773,n1774,n1804);
xor (n1774,n1775,n1801);
xor (n1775,n1776,n1800);
xor (n1776,n1777,n1797);
xor (n1777,n1778,n1796);
xor (n1778,n1779,n1793);
xor (n1779,n1780,n1792);
xor (n1780,n1781,n1789);
xor (n1781,n1782,n1788);
xor (n1782,n1783,n1785);
xor (n1783,n1784,n971);
and (n1784,n322,n390);
or (n1785,n1786,n1787);
and (n1786,n1684,n1685);
and (n1787,n1683,n1686);
and (n1788,n118,n359);
or (n1789,n1790,n1791);
and (n1790,n1682,n1689);
and (n1791,n1681,n1690);
and (n1792,n138,n282);
or (n1793,n1794,n1795);
and (n1794,n1680,n1693);
and (n1795,n1679,n1694);
and (n1796,n107,n277);
or (n1797,n1798,n1799);
and (n1798,n1678,n1697);
and (n1799,n1677,n1698);
and (n1800,n53,n233);
or (n1801,n1802,n1803);
and (n1802,n1676,n1701);
and (n1803,n1675,n1702);
and (n1804,n167,n239);
or (n1805,n1806,n1807);
and (n1806,n1674,n1705);
and (n1807,n1673,n1706);
and (n1808,n187,n217);
and (n1809,n1672,n1707);
or (n1810,n1811,n1813);
and (n1811,n1812,n1768);
xor (n1812,n1712,n1713);
and (n1813,n1814,n1815);
xor (n1814,n1812,n1768);
or (n1815,n1816,n1818);
and (n1816,n1817,n1768);
xor (n1817,n1717,n1718);
and (n1818,n1819,n1820);
xor (n1819,n1817,n1768);
or (n1820,n1821,n1823);
and (n1821,n1822,n1768);
xor (n1822,n1722,n1723);
and (n1823,n1824,n1825);
xor (n1824,n1822,n1768);
or (n1825,n1826,n1828);
and (n1826,n1827,n1768);
xor (n1827,n1727,n1728);
and (n1828,n1829,n1830);
xor (n1829,n1827,n1768);
or (n1830,n1831,n1833);
and (n1831,n1832,n1768);
xor (n1832,n1732,n1733);
and (n1833,n1834,n1835);
xor (n1834,n1832,n1768);
or (n1835,n1836,n1838);
and (n1836,n1837,n1768);
xor (n1837,n1737,n1738);
and (n1838,n1839,n1840);
xor (n1839,n1837,n1768);
or (n1840,n1841,n1843);
and (n1841,n1842,n1768);
xor (n1842,n1742,n1743);
and (n1843,n1844,n1845);
xor (n1844,n1842,n1768);
or (n1845,n1846,n1848);
and (n1846,n1847,n1768);
xor (n1847,n1747,n1748);
and (n1848,n1849,n1850);
xor (n1849,n1847,n1768);
or (n1850,n1851,n1854);
and (n1851,n1852,n1853);
xor (n1852,n1752,n1753);
and (n1853,n1769,n1506);
and (n1854,n1855,n1856);
xor (n1855,n1852,n1853);
or (n1856,n1857,n1860);
and (n1857,n1858,n1859);
xor (n1858,n1758,n1759);
and (n1859,n1769,n1514);
and (n1860,n1861,n1862);
xor (n1861,n1858,n1859);
and (n1862,n1863,n1864);
xor (n1863,n1764,n1765);
and (n1864,n1769,n1521);
and (n1865,n1252,n1866);
xor (n1866,n1867,n952);
xor (n1867,n1868,n1913);
xor (n1868,n1869,n1912);
xor (n1869,n1870,n1909);
xor (n1870,n1871,n1908);
xor (n1871,n1872,n1905);
xor (n1872,n1873,n1904);
xor (n1873,n1874,n1901);
xor (n1874,n1875,n1900);
xor (n1875,n1876,n1897);
xor (n1876,n1877,n1896);
xor (n1877,n1878,n1893);
xor (n1878,n1879,n1892);
xor (n1879,n1880,n1889);
xor (n1880,n1881,n1888);
xor (n1881,n1882,n1885);
xor (n1882,n1883,n1884);
and (n1883,n223,n390);
and (n1884,n322,n369);
or (n1885,n1886,n1887);
and (n1886,n1784,n971);
and (n1887,n1783,n1785);
and (n1888,n331,n359);
or (n1889,n1890,n1891);
and (n1890,n1782,n1788);
and (n1891,n1781,n1789);
and (n1892,n118,n282);
or (n1893,n1894,n1895);
and (n1894,n1780,n1792);
and (n1895,n1779,n1793);
and (n1896,n138,n277);
or (n1897,n1898,n1899);
and (n1898,n1778,n1796);
and (n1899,n1777,n1797);
and (n1900,n107,n233);
or (n1901,n1902,n1903);
and (n1902,n1776,n1800);
and (n1903,n1775,n1801);
and (n1904,n53,n239);
or (n1905,n1906,n1907);
and (n1906,n1774,n1804);
and (n1907,n1773,n1805);
and (n1908,n167,n217);
or (n1909,n1910,n1911);
and (n1910,n1772,n1808);
and (n1911,n1771,n1809);
and (n1912,n187,n311);
and (n1913,n1770,n888);
or (n1914,n1915,n1917);
and (n1915,n1916,n1865);
xor (n1916,n1814,n1815);
and (n1917,n1918,n1919);
xor (n1918,n1916,n1865);
or (n1919,n1920,n1922);
and (n1920,n1921,n1865);
xor (n1921,n1819,n1820);
and (n1922,n1923,n1924);
xor (n1923,n1921,n1865);
or (n1924,n1925,n1927);
and (n1925,n1926,n1865);
xor (n1926,n1824,n1825);
and (n1927,n1928,n1929);
xor (n1928,n1926,n1865);
or (n1929,n1930,n1932);
and (n1930,n1931,n1865);
xor (n1931,n1829,n1830);
and (n1932,n1933,n1934);
xor (n1933,n1931,n1865);
or (n1934,n1935,n1937);
and (n1935,n1936,n1865);
xor (n1936,n1834,n1835);
and (n1937,n1938,n1939);
xor (n1938,n1936,n1865);
or (n1939,n1940,n1942);
and (n1940,n1941,n1865);
xor (n1941,n1839,n1840);
and (n1942,n1943,n1944);
xor (n1943,n1941,n1865);
or (n1944,n1945,n1947);
and (n1945,n1946,n1865);
xor (n1946,n1844,n1845);
and (n1947,n1948,n1949);
xor (n1948,n1946,n1865);
or (n1949,n1950,n1953);
and (n1950,n1951,n1952);
xor (n1951,n1849,n1850);
and (n1952,n1506,n1866);
and (n1953,n1954,n1955);
xor (n1954,n1951,n1952);
or (n1955,n1956,n1959);
and (n1956,n1957,n1958);
xor (n1957,n1855,n1856);
and (n1958,n1514,n1866);
and (n1959,n1960,n1961);
xor (n1960,n1957,n1958);
and (n1961,n1962,n1963);
xor (n1962,n1861,n1862);
and (n1963,n1521,n1866);
and (n1964,n1252,n1965);
xor (n1965,n1966,n747);
xor (n1966,n1967,n2017);
xor (n1967,n1968,n2016);
xor (n1968,n1969,n2013);
xor (n1969,n1970,n2012);
xor (n1970,n1971,n2009);
xor (n1971,n1972,n2008);
xor (n1972,n1973,n2005);
xor (n1973,n1974,n2004);
xor (n1974,n1975,n2001);
xor (n1975,n1976,n2000);
xor (n1976,n1977,n1997);
xor (n1977,n1978,n1996);
xor (n1978,n1979,n1993);
xor (n1979,n1980,n846);
xor (n1980,n1981,n1990);
xor (n1981,n1982,n1989);
xor (n1982,n1983,n1986);
xor (n1983,n1984,n1985);
and (n1984,n253,n390);
and (n1985,n223,n369);
or (n1986,n1987,n1988);
and (n1987,n1883,n1884);
and (n1988,n1882,n1885);
and (n1989,n322,n359);
or (n1990,n1991,n1992);
and (n1991,n1881,n1888);
and (n1992,n1880,n1889);
or (n1993,n1994,n1995);
and (n1994,n1879,n1892);
and (n1995,n1878,n1893);
and (n1996,n118,n277);
or (n1997,n1998,n1999);
and (n1998,n1877,n1896);
and (n1999,n1876,n1897);
and (n2000,n138,n233);
or (n2001,n2002,n2003);
and (n2002,n1875,n1900);
and (n2003,n1874,n1901);
and (n2004,n107,n239);
or (n2005,n2006,n2007);
and (n2006,n1873,n1904);
and (n2007,n1872,n1905);
and (n2008,n53,n217);
or (n2009,n2010,n2011);
and (n2010,n1871,n1908);
and (n2011,n1870,n1909);
and (n2012,n167,n311);
or (n2013,n2014,n2015);
and (n2014,n1869,n1912);
and (n2015,n1868,n1913);
and (n2016,n187,n125);
and (n2017,n1867,n952);
or (n2018,n2019,n2021);
and (n2019,n2020,n1964);
xor (n2020,n1918,n1919);
and (n2021,n2022,n2023);
xor (n2022,n2020,n1964);
or (n2023,n2024,n2026);
and (n2024,n2025,n1964);
xor (n2025,n1923,n1924);
and (n2026,n2027,n2028);
xor (n2027,n2025,n1964);
or (n2028,n2029,n2031);
and (n2029,n2030,n1964);
xor (n2030,n1928,n1929);
and (n2031,n2032,n2033);
xor (n2032,n2030,n1964);
or (n2033,n2034,n2036);
and (n2034,n2035,n1964);
xor (n2035,n1933,n1934);
and (n2036,n2037,n2038);
xor (n2037,n2035,n1964);
or (n2038,n2039,n2041);
and (n2039,n2040,n1964);
xor (n2040,n1938,n1939);
and (n2041,n2042,n2043);
xor (n2042,n2040,n1964);
or (n2043,n2044,n2046);
and (n2044,n2045,n1964);
xor (n2045,n1943,n1944);
and (n2046,n2047,n2048);
xor (n2047,n2045,n1964);
or (n2048,n2049,n2052);
and (n2049,n2050,n2051);
xor (n2050,n1948,n1949);
and (n2051,n1506,n1965);
and (n2052,n2053,n2054);
xor (n2053,n2050,n2051);
or (n2054,n2055,n2058);
and (n2055,n2056,n2057);
xor (n2056,n1954,n1955);
and (n2057,n1514,n1965);
and (n2058,n2059,n2060);
xor (n2059,n2056,n2057);
and (n2060,n2061,n2062);
xor (n2061,n1960,n1961);
and (n2062,n1521,n1965);
and (n2063,n1252,n2064);
xor (n2064,n2065,n763);
xor (n2065,n2066,n2123);
xor (n2066,n2067,n2122);
xor (n2067,n2068,n2119);
xor (n2068,n2069,n2118);
xor (n2069,n2070,n2115);
xor (n2070,n2071,n2114);
xor (n2071,n2072,n2111);
xor (n2072,n2073,n2110);
xor (n2073,n2074,n2107);
xor (n2074,n2075,n2106);
xor (n2075,n2076,n2103);
xor (n2076,n2077,n2102);
xor (n2077,n2078,n2099);
xor (n2078,n2079,n2098);
xor (n2079,n2080,n2095);
xor (n2080,n2081,n2094);
xor (n2081,n2082,n2091);
xor (n2082,n2083,n2090);
xor (n2083,n2084,n2087);
xor (n2084,n2085,n2086);
and (n2085,n292,n390);
and (n2086,n253,n369);
or (n2087,n2088,n2089);
and (n2088,n1984,n1985);
and (n2089,n1983,n1986);
and (n2090,n223,n359);
or (n2091,n2092,n2093);
and (n2092,n1982,n1989);
and (n2093,n1981,n1990);
and (n2094,n322,n282);
or (n2095,n2096,n2097);
and (n2096,n1980,n846);
and (n2097,n1979,n1993);
and (n2098,n331,n277);
or (n2099,n2100,n2101);
and (n2100,n1978,n1996);
and (n2101,n1977,n1997);
and (n2102,n118,n233);
or (n2103,n2104,n2105);
and (n2104,n1976,n2000);
and (n2105,n1975,n2001);
and (n2106,n138,n239);
or (n2107,n2108,n2109);
and (n2108,n1974,n2004);
and (n2109,n1973,n2005);
and (n2110,n107,n217);
or (n2111,n2112,n2113);
and (n2112,n1972,n2008);
and (n2113,n1971,n2009);
and (n2114,n53,n311);
or (n2115,n2116,n2117);
and (n2116,n1970,n2012);
and (n2117,n1969,n2013);
and (n2118,n167,n125);
or (n2119,n2120,n2121);
and (n2120,n1968,n2016);
and (n2121,n1967,n2017);
and (n2122,n187,n130);
and (n2123,n1966,n747);
or (n2124,n2125,n2127);
and (n2125,n2126,n2063);
xor (n2126,n2022,n2023);
and (n2127,n2128,n2129);
xor (n2128,n2126,n2063);
or (n2129,n2130,n2132);
and (n2130,n2131,n2063);
xor (n2131,n2027,n2028);
and (n2132,n2133,n2134);
xor (n2133,n2131,n2063);
or (n2134,n2135,n2137);
and (n2135,n2136,n2063);
xor (n2136,n2032,n2033);
and (n2137,n2138,n2139);
xor (n2138,n2136,n2063);
or (n2139,n2140,n2142);
and (n2140,n2141,n2063);
xor (n2141,n2037,n2038);
and (n2142,n2143,n2144);
xor (n2143,n2141,n2063);
or (n2144,n2145,n2147);
and (n2145,n2146,n2063);
xor (n2146,n2042,n2043);
and (n2147,n2148,n2149);
xor (n2148,n2146,n2063);
or (n2149,n2150,n2153);
and (n2150,n2151,n2152);
xor (n2151,n2047,n2048);
and (n2152,n1506,n2064);
and (n2153,n2154,n2155);
xor (n2154,n2151,n2152);
or (n2155,n2156,n2159);
and (n2156,n2157,n2158);
xor (n2157,n2053,n2054);
and (n2158,n1514,n2064);
and (n2159,n2160,n2161);
xor (n2160,n2157,n2158);
and (n2161,n2162,n2163);
xor (n2162,n2059,n2060);
and (n2163,n1521,n2064);
and (n2164,n1252,n2165);
xor (n2165,n2166,n447);
xor (n2166,n2167,n2230);
xor (n2167,n2168,n2229);
xor (n2168,n2169,n2226);
xor (n2169,n2170,n2225);
xor (n2170,n2171,n2222);
xor (n2171,n2172,n2221);
xor (n2172,n2173,n2218);
xor (n2173,n2174,n2217);
xor (n2174,n2175,n2214);
xor (n2175,n2176,n2213);
xor (n2176,n2177,n2210);
xor (n2177,n2178,n2209);
xor (n2178,n2179,n2206);
xor (n2179,n2180,n2205);
xor (n2180,n2181,n2202);
xor (n2181,n2182,n2201);
xor (n2182,n2183,n2198);
xor (n2183,n2184,n2197);
xor (n2184,n2185,n2194);
xor (n2185,n2186,n2193);
xor (n2186,n2187,n2190);
xor (n2187,n2188,n2189);
and (n2188,n266,n390);
and (n2189,n292,n369);
or (n2190,n2191,n2192);
and (n2191,n2085,n2086);
and (n2192,n2084,n2087);
and (n2193,n253,n359);
or (n2194,n2195,n2196);
and (n2195,n2083,n2090);
and (n2196,n2082,n2091);
and (n2197,n223,n282);
or (n2198,n2199,n2200);
and (n2199,n2081,n2094);
and (n2200,n2080,n2095);
and (n2201,n322,n277);
or (n2202,n2203,n2204);
and (n2203,n2079,n2098);
and (n2204,n2078,n2099);
and (n2205,n331,n233);
or (n2206,n2207,n2208);
and (n2207,n2077,n2102);
and (n2208,n2076,n2103);
and (n2209,n118,n239);
or (n2210,n2211,n2212);
and (n2211,n2075,n2106);
and (n2212,n2074,n2107);
and (n2213,n138,n217);
or (n2214,n2215,n2216);
and (n2215,n2073,n2110);
and (n2216,n2072,n2111);
and (n2217,n107,n311);
or (n2218,n2219,n2220);
and (n2219,n2071,n2114);
and (n2220,n2070,n2115);
and (n2221,n53,n125);
or (n2222,n2223,n2224);
and (n2223,n2069,n2118);
and (n2224,n2068,n2119);
and (n2225,n167,n130);
or (n2226,n2227,n2228);
and (n2227,n2067,n2122);
and (n2228,n2066,n2123);
and (n2229,n187,n44);
and (n2230,n2065,n763);
or (n2231,n2232,n2234);
and (n2232,n2233,n2164);
xor (n2233,n2128,n2129);
and (n2234,n2235,n2236);
xor (n2235,n2233,n2164);
or (n2236,n2237,n2239);
and (n2237,n2238,n2164);
xor (n2238,n2133,n2134);
and (n2239,n2240,n2241);
xor (n2240,n2238,n2164);
or (n2241,n2242,n2244);
and (n2242,n2243,n2164);
xor (n2243,n2138,n2139);
and (n2244,n2245,n2246);
xor (n2245,n2243,n2164);
or (n2246,n2247,n2249);
and (n2247,n2248,n2164);
xor (n2248,n2143,n2144);
and (n2249,n2250,n2251);
xor (n2250,n2248,n2164);
or (n2251,n2252,n2255);
and (n2252,n2253,n2254);
xor (n2253,n2148,n2149);
and (n2254,n1506,n2165);
and (n2255,n2256,n2257);
xor (n2256,n2253,n2254);
or (n2257,n2258,n2261);
and (n2258,n2259,n2260);
xor (n2259,n2154,n2155);
and (n2260,n1514,n2165);
and (n2261,n2262,n2263);
xor (n2262,n2259,n2260);
and (n2263,n2264,n2265);
xor (n2264,n2160,n2161);
and (n2265,n1521,n2165);
and (n2266,n1252,n2267);
xor (n2267,n2268,n2339);
xor (n2268,n2269,n2338);
xor (n2269,n2270,n2337);
xor (n2270,n2271,n2334);
xor (n2271,n2272,n2333);
xor (n2272,n2273,n2330);
xor (n2273,n2274,n2329);
xor (n2274,n2275,n2326);
xor (n2275,n2276,n2325);
xor (n2276,n2277,n2322);
xor (n2277,n2278,n2321);
xor (n2278,n2279,n2318);
xor (n2279,n2280,n2317);
xor (n2280,n2281,n2314);
xor (n2281,n2282,n2313);
xor (n2282,n2283,n2310);
xor (n2283,n2284,n2309);
xor (n2284,n2285,n2306);
xor (n2285,n2286,n2305);
xor (n2286,n2287,n2302);
xor (n2287,n2288,n2301);
xor (n2288,n2289,n2298);
xor (n2289,n2290,n2297);
xor (n2290,n2291,n2294);
xor (n2291,n2292,n2293);
and (n2292,n346,n390);
and (n2293,n266,n369);
or (n2294,n2295,n2296);
and (n2295,n2188,n2189);
and (n2296,n2187,n2190);
and (n2297,n292,n359);
or (n2298,n2299,n2300);
and (n2299,n2186,n2193);
and (n2300,n2185,n2194);
and (n2301,n253,n282);
or (n2302,n2303,n2304);
and (n2303,n2184,n2197);
and (n2304,n2183,n2198);
and (n2305,n223,n277);
or (n2306,n2307,n2308);
and (n2307,n2182,n2201);
and (n2308,n2181,n2202);
and (n2309,n322,n233);
or (n2310,n2311,n2312);
and (n2311,n2180,n2205);
and (n2312,n2179,n2206);
and (n2313,n331,n239);
or (n2314,n2315,n2316);
and (n2315,n2178,n2209);
and (n2316,n2177,n2210);
and (n2317,n118,n217);
or (n2318,n2319,n2320);
and (n2319,n2176,n2213);
and (n2320,n2175,n2214);
and (n2321,n138,n311);
or (n2322,n2323,n2324);
and (n2323,n2174,n2217);
and (n2324,n2173,n2218);
and (n2325,n107,n125);
or (n2326,n2327,n2328);
and (n2327,n2172,n2221);
and (n2328,n2171,n2222);
and (n2329,n53,n130);
or (n2330,n2331,n2332);
and (n2331,n2170,n2225);
and (n2332,n2169,n2226);
and (n2333,n167,n44);
or (n2334,n2335,n2336);
and (n2335,n2168,n2229);
and (n2336,n2167,n2230);
and (n2337,n187,n33);
and (n2338,n2166,n447);
and (n2339,n207,n18);
or (n2340,n2341,n2343);
and (n2341,n2342,n2266);
xor (n2342,n2235,n2236);
and (n2343,n2344,n2345);
xor (n2344,n2342,n2266);
or (n2345,n2346,n2348);
and (n2346,n2347,n2266);
xor (n2347,n2240,n2241);
and (n2348,n2349,n2350);
xor (n2349,n2347,n2266);
or (n2350,n2351,n2353);
and (n2351,n2352,n2266);
xor (n2352,n2245,n2246);
and (n2353,n2354,n2355);
xor (n2354,n2352,n2266);
or (n2355,n2356,n2359);
and (n2356,n2357,n2358);
xor (n2357,n2250,n2251);
and (n2358,n1506,n2267);
and (n2359,n2360,n2361);
xor (n2360,n2357,n2358);
or (n2361,n2362,n2365);
and (n2362,n2363,n2364);
xor (n2363,n2256,n2257);
and (n2364,n1514,n2267);
and (n2365,n2366,n2367);
xor (n2366,n2363,n2364);
and (n2367,n2368,n2369);
xor (n2368,n2262,n2263);
and (n2369,n1521,n2267);
and (n2370,n1252,n2371);
xor (n2371,n2372,n475);
xor (n2372,n2373,n2448);
xor (n2373,n2374,n2447);
xor (n2374,n2375,n2444);
xor (n2375,n2376,n2443);
xor (n2376,n2377,n2440);
xor (n2377,n2378,n2439);
xor (n2378,n2379,n2436);
xor (n2379,n2380,n2435);
xor (n2380,n2381,n2432);
xor (n2381,n2382,n2431);
xor (n2382,n2383,n2428);
xor (n2383,n2384,n2427);
xor (n2384,n2385,n2424);
xor (n2385,n2386,n2423);
xor (n2386,n2387,n2420);
xor (n2387,n2388,n2419);
xor (n2388,n2389,n2416);
xor (n2389,n2390,n2415);
xor (n2390,n2391,n2412);
xor (n2391,n2392,n2411);
xor (n2392,n2393,n2408);
xor (n2393,n2394,n2407);
xor (n2394,n2395,n2404);
xor (n2395,n2396,n2403);
xor (n2396,n2397,n2400);
xor (n2397,n2398,n2399);
and (n2398,n378,n390);
and (n2399,n346,n369);
or (n2400,n2401,n2402);
and (n2401,n2292,n2293);
and (n2402,n2291,n2294);
and (n2403,n266,n359);
or (n2404,n2405,n2406);
and (n2405,n2290,n2297);
and (n2406,n2289,n2298);
and (n2407,n292,n282);
or (n2408,n2409,n2410);
and (n2409,n2288,n2301);
and (n2410,n2287,n2302);
and (n2411,n253,n277);
or (n2412,n2413,n2414);
and (n2413,n2286,n2305);
and (n2414,n2285,n2306);
and (n2415,n223,n233);
or (n2416,n2417,n2418);
and (n2417,n2284,n2309);
and (n2418,n2283,n2310);
and (n2419,n322,n239);
or (n2420,n2421,n2422);
and (n2421,n2282,n2313);
and (n2422,n2281,n2314);
and (n2423,n331,n217);
or (n2424,n2425,n2426);
and (n2425,n2280,n2317);
and (n2426,n2279,n2318);
and (n2427,n118,n311);
or (n2428,n2429,n2430);
and (n2429,n2278,n2321);
and (n2430,n2277,n2322);
and (n2431,n138,n125);
or (n2432,n2433,n2434);
and (n2433,n2276,n2325);
and (n2434,n2275,n2326);
and (n2435,n107,n130);
or (n2436,n2437,n2438);
and (n2437,n2274,n2329);
and (n2438,n2273,n2330);
and (n2439,n53,n44);
or (n2440,n2441,n2442);
and (n2441,n2272,n2333);
and (n2442,n2271,n2334);
and (n2443,n167,n33);
or (n2444,n2445,n2446);
and (n2445,n2270,n2337);
and (n2446,n2269,n2338);
and (n2447,n187,n18);
and (n2448,n2268,n2339);
or (n2449,n2450,n2452);
and (n2450,n2451,n2370);
xor (n2451,n2344,n2345);
and (n2452,n2453,n2454);
xor (n2453,n2451,n2370);
or (n2454,n2455,n2457);
and (n2455,n2456,n2370);
xor (n2456,n2349,n2350);
and (n2457,n2458,n2459);
xor (n2458,n2456,n2370);
or (n2459,n2460,n2463);
and (n2460,n2461,n2462);
xor (n2461,n2354,n2355);
and (n2462,n1506,n2371);
and (n2463,n2464,n2465);
xor (n2464,n2461,n2462);
or (n2465,n2466,n2469);
and (n2466,n2467,n2468);
xor (n2467,n2360,n2361);
and (n2468,n1514,n2371);
and (n2469,n2470,n2471);
xor (n2470,n2467,n2468);
and (n2471,n2472,n2473);
xor (n2472,n2366,n2367);
and (n2473,n1521,n2371);
and (n2474,n1252,n2475);
xor (n2475,n2476,n468);
xor (n2476,n2477,n2557);
xor (n2477,n2478,n2556);
xor (n2478,n2479,n2553);
xor (n2479,n2480,n2552);
xor (n2480,n2481,n2549);
xor (n2481,n2482,n2548);
xor (n2482,n2483,n2545);
xor (n2483,n2484,n2544);
xor (n2484,n2485,n2541);
xor (n2485,n2486,n2540);
xor (n2486,n2487,n2537);
xor (n2487,n2488,n2536);
xor (n2488,n2489,n2533);
xor (n2489,n2490,n2532);
xor (n2490,n2491,n2529);
xor (n2491,n2492,n2528);
xor (n2492,n2493,n2525);
xor (n2493,n2494,n2524);
xor (n2494,n2495,n2521);
xor (n2495,n2496,n2520);
xor (n2496,n2497,n2517);
xor (n2497,n2498,n2516);
xor (n2498,n2499,n2513);
xor (n2499,n2500,n2512);
xor (n2500,n2501,n2509);
xor (n2501,n2502,n2508);
xor (n2502,n2503,n2505);
xor (n2503,n2504,n587);
and (n2504,n399,n390);
or (n2505,n2506,n2507);
and (n2506,n2398,n2399);
and (n2507,n2397,n2400);
and (n2508,n346,n359);
or (n2509,n2510,n2511);
and (n2510,n2396,n2403);
and (n2511,n2395,n2404);
and (n2512,n266,n282);
or (n2513,n2514,n2515);
and (n2514,n2394,n2407);
and (n2515,n2393,n2408);
and (n2516,n292,n277);
or (n2517,n2518,n2519);
and (n2518,n2392,n2411);
and (n2519,n2391,n2412);
and (n2520,n253,n233);
or (n2521,n2522,n2523);
and (n2522,n2390,n2415);
and (n2523,n2389,n2416);
and (n2524,n223,n239);
or (n2525,n2526,n2527);
and (n2526,n2388,n2419);
and (n2527,n2387,n2420);
and (n2528,n322,n217);
or (n2529,n2530,n2531);
and (n2530,n2386,n2423);
and (n2531,n2385,n2424);
and (n2532,n331,n311);
or (n2533,n2534,n2535);
and (n2534,n2384,n2427);
and (n2535,n2383,n2428);
and (n2536,n118,n125);
or (n2537,n2538,n2539);
and (n2538,n2382,n2431);
and (n2539,n2381,n2432);
and (n2540,n138,n130);
or (n2541,n2542,n2543);
and (n2542,n2380,n2435);
and (n2543,n2379,n2436);
and (n2544,n107,n44);
or (n2545,n2546,n2547);
and (n2546,n2378,n2439);
and (n2547,n2377,n2440);
and (n2548,n53,n33);
or (n2549,n2550,n2551);
and (n2550,n2376,n2443);
and (n2551,n2375,n2444);
and (n2552,n167,n18);
or (n2553,n2554,n2555);
and (n2554,n2374,n2447);
and (n2555,n2373,n2448);
and (n2556,n187,n158);
and (n2557,n2372,n475);
or (n2558,n2559,n2561);
and (n2559,n2560,n2474);
xor (n2560,n2453,n2454);
and (n2561,n2562,n2563);
xor (n2562,n2560,n2474);
or (n2563,n2564,n2567);
and (n2564,n2565,n2566);
xor (n2565,n2458,n2459);
and (n2566,n1506,n2475);
and (n2567,n2568,n2569);
xor (n2568,n2565,n2566);
or (n2569,n2570,n2573);
and (n2570,n2571,n2572);
xor (n2571,n2464,n2465);
and (n2572,n1514,n2475);
and (n2573,n2574,n2575);
xor (n2574,n2571,n2572);
and (n2575,n2576,n2577);
xor (n2576,n2470,n2471);
and (n2577,n1521,n2475);
and (n2578,n1252,n2579);
xor (n2579,n2580,n2666);
xor (n2580,n2581,n2665);
xor (n2581,n2582,n186);
xor (n2582,n2583,n2662);
xor (n2583,n2584,n2661);
xor (n2584,n2585,n2658);
xor (n2585,n2586,n2657);
xor (n2586,n2587,n2654);
xor (n2587,n2588,n2653);
xor (n2588,n2589,n2650);
xor (n2589,n2590,n2649);
xor (n2590,n2591,n2646);
xor (n2591,n2592,n2645);
xor (n2592,n2593,n2642);
xor (n2593,n2594,n2641);
xor (n2594,n2595,n2638);
xor (n2595,n2596,n2637);
xor (n2596,n2597,n2634);
xor (n2597,n2598,n2633);
xor (n2598,n2599,n2630);
xor (n2599,n2600,n2629);
xor (n2600,n2601,n2626);
xor (n2601,n2602,n297);
xor (n2602,n2603,n2623);
xor (n2603,n2604,n2622);
xor (n2604,n2605,n2619);
xor (n2605,n2606,n345);
xor (n2606,n2607,n2616);
xor (n2607,n2608,n2615);
xor (n2608,n2609,n2612);
xor (n2609,n2610,n2611);
and (n2610,n408,n390);
and (n2611,n399,n369);
or (n2612,n2613,n2614);
and (n2613,n2504,n587);
and (n2614,n2503,n2505);
and (n2615,n378,n359);
or (n2616,n2617,n2618);
and (n2617,n2502,n2508);
and (n2618,n2501,n2509);
or (n2619,n2620,n2621);
and (n2620,n2500,n2512);
and (n2621,n2499,n2513);
and (n2622,n266,n277);
or (n2623,n2624,n2625);
and (n2624,n2498,n2516);
and (n2625,n2497,n2517);
or (n2626,n2627,n2628);
and (n2627,n2496,n2520);
and (n2628,n2495,n2521);
and (n2629,n253,n239);
or (n2630,n2631,n2632);
and (n2631,n2494,n2524);
and (n2632,n2493,n2525);
and (n2633,n223,n217);
or (n2634,n2635,n2636);
and (n2635,n2492,n2528);
and (n2636,n2491,n2529);
and (n2637,n322,n311);
or (n2638,n2639,n2640);
and (n2639,n2490,n2532);
and (n2640,n2489,n2533);
and (n2641,n331,n125);
or (n2642,n2643,n2644);
and (n2643,n2488,n2536);
and (n2644,n2487,n2537);
and (n2645,n118,n130);
or (n2646,n2647,n2648);
and (n2647,n2486,n2540);
and (n2648,n2485,n2541);
and (n2649,n138,n44);
or (n2650,n2651,n2652);
and (n2651,n2484,n2544);
and (n2652,n2483,n2545);
and (n2653,n107,n33);
or (n2654,n2655,n2656);
and (n2655,n2482,n2548);
and (n2656,n2481,n2549);
and (n2657,n53,n18);
or (n2658,n2659,n2660);
and (n2659,n2480,n2552);
and (n2660,n2479,n2553);
and (n2661,n167,n158);
or (n2662,n2663,n2664);
and (n2663,n2478,n2556);
and (n2664,n2477,n2557);
and (n2665,n2476,n468);
and (n2666,n207,n199);
endmodule
