module top (out,n15,n16,n25,n26,n35,n42,n43,n48,n53
        ,n60,n61,n69,n74,n79,n90,n102,n112,n123,n138
        ,n150,n175,n195);
output out;
input n15;
input n16;
input n25;
input n26;
input n35;
input n42;
input n43;
input n48;
input n53;
input n60;
input n61;
input n69;
input n74;
input n79;
input n90;
input n102;
input n112;
input n123;
input n138;
input n150;
input n175;
input n195;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n24;
wire n27;
wire n28;
wire n29;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n44;
wire n45;
wire n46;
wire n47;
wire n49;
wire n50;
wire n51;
wire n52;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n70;
wire n71;
wire n72;
wire n73;
wire n75;
wire n76;
wire n77;
wire n78;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
xor (out,n0,n455);
nand (n0,n1,n454);
or (n1,n2,n249);
not (n2,n3);
and (n3,n4,n248);
not (n4,n5);
nor (n5,n6,n212);
xor (n6,n7,n164);
xor (n7,n8,n83);
xor (n8,n9,n55);
xor (n9,n10,n37);
nand (n10,n11,n31);
or (n11,n12,n20);
not (n12,n13);
nor (n13,n14,n17);
and (n14,n15,n16);
and (n17,n18,n19);
not (n18,n16);
not (n19,n15);
nand (n20,n21,n28);
not (n21,n22);
nand (n22,n23,n27);
or (n23,n24,n26);
not (n24,n25);
nand (n27,n26,n24);
nand (n28,n29,n30);
or (n29,n26,n19);
nand (n30,n19,n26);
nand (n31,n22,n32);
nor (n32,n33,n36);
and (n33,n34,n19);
not (n34,n35);
and (n36,n15,n35);
nand (n37,n38,n49);
or (n38,n39,n46);
nor (n39,n40,n44);
and (n40,n41,n43);
not (n41,n42);
and (n44,n42,n45);
not (n45,n43);
nand (n46,n42,n47);
not (n47,n48);
or (n49,n50,n47);
nor (n50,n51,n54);
and (n51,n52,n42);
not (n52,n53);
and (n54,n53,n41);
nand (n55,n56,n76);
or (n56,n57,n64);
nor (n57,n58,n62);
and (n58,n59,n61);
not (n59,n60);
and (n62,n60,n63);
not (n63,n61);
not (n64,n65);
nor (n65,n66,n71);
nor (n66,n67,n70);
and (n67,n68,n60);
not (n68,n69);
nor (n70,n60,n68);
nand (n71,n72,n75);
or (n72,n73,n69);
not (n73,n74);
nand (n75,n73,n69);
or (n76,n77,n82);
nor (n77,n78,n80);
and (n78,n59,n79);
and (n80,n60,n81);
not (n81,n79);
not (n82,n71);
or (n83,n84,n163);
and (n84,n85,n125);
xor (n85,n86,n94);
nand (n86,n87,n93);
or (n87,n64,n88);
nor (n88,n89,n91);
and (n89,n59,n90);
and (n91,n60,n92);
not (n92,n90);
or (n93,n82,n57);
xor (n94,n95,n103);
and (n95,n96,n15);
nand (n96,n97,n98);
or (n97,n25,n26);
nand (n98,n99,n101);
or (n99,n100,n24);
not (n100,n26);
not (n101,n102);
nand (n103,n104,n118);
or (n104,n105,n109);
not (n105,n106);
nand (n106,n107,n108);
or (n107,n74,n81);
or (n108,n73,n79);
nand (n109,n110,n115);
nor (n110,n111,n113);
and (n111,n41,n112);
and (n113,n42,n114);
not (n114,n112);
nand (n115,n116,n117);
or (n116,n114,n74);
nand (n117,n74,n114);
nand (n118,n119,n120);
not (n119,n110);
nor (n120,n121,n124);
and (n121,n122,n73);
not (n122,n123);
and (n124,n74,n123);
or (n125,n126,n162);
and (n126,n127,n141);
xor (n127,n128,n129);
and (n128,n22,n102);
nand (n129,n130,n135);
or (n130,n46,n131);
not (n131,n132);
nor (n132,n133,n134);
and (n133,n122,n41);
and (n134,n42,n123);
or (n135,n136,n47);
nor (n136,n137,n139);
and (n137,n41,n138);
and (n139,n42,n140);
not (n140,n138);
nand (n141,n142,n152);
or (n142,n143,n147);
not (n143,n144);
nor (n144,n145,n146);
and (n145,n34,n24);
and (n146,n25,n35);
not (n147,n148);
nand (n148,n149,n151);
or (n149,n59,n150);
nand (n151,n59,n150);
or (n152,n153,n159);
not (n153,n154);
nor (n154,n155,n148);
nor (n155,n156,n157);
and (n156,n150,n24);
and (n157,n25,n158);
not (n158,n150);
nor (n159,n160,n161);
and (n160,n16,n24);
and (n161,n18,n25);
and (n162,n128,n129);
and (n163,n86,n94);
xor (n164,n165,n189);
xor (n165,n166,n167);
and (n166,n95,n103);
or (n167,n168,n188);
and (n168,n169,n185);
xor (n169,n170,n178);
nand (n170,n171,n172);
or (n171,n143,n153);
nand (n172,n148,n173);
nor (n173,n174,n176);
and (n174,n25,n175);
and (n176,n177,n24);
not (n177,n175);
nand (n178,n179,n184);
or (n179,n180,n20);
not (n180,n181);
nand (n181,n182,n183);
or (n182,n15,n101);
or (n183,n19,n102);
nand (n184,n22,n13);
nand (n185,n186,n187);
or (n186,n46,n136);
or (n187,n39,n47);
and (n188,n170,n178);
xor (n189,n190,n204);
xor (n190,n191,n197);
and (n191,n192,n102);
nand (n192,n193,n196);
or (n193,n194,n15);
not (n194,n195);
or (n196,n19,n195);
nand (n197,n198,n200);
or (n198,n199,n109);
not (n199,n120);
nand (n200,n119,n201);
nor (n201,n202,n203);
and (n202,n140,n73);
and (n203,n74,n138);
nand (n204,n205,n207);
or (n205,n206,n153);
not (n206,n173);
nand (n207,n208,n148);
not (n208,n209);
nor (n209,n210,n211);
and (n210,n24,n90);
and (n211,n25,n92);
or (n212,n213,n247);
and (n213,n214,n246);
xor (n214,n215,n216);
xor (n215,n169,n185);
or (n216,n217,n245);
and (n217,n218,n232);
xor (n218,n219,n226);
nand (n219,n220,n225);
or (n220,n221,n109);
not (n221,n222);
nand (n222,n223,n224);
or (n223,n74,n63);
or (n224,n73,n61);
nand (n225,n119,n106);
nand (n226,n227,n231);
or (n227,n64,n228);
nor (n228,n229,n230);
and (n229,n59,n175);
and (n230,n60,n177);
or (n231,n88,n82);
and (n232,n233,n238);
nor (n233,n234,n24);
nor (n234,n235,n237);
and (n235,n236,n101);
nand (n236,n60,n150);
and (n237,n59,n158);
nand (n238,n239,n244);
or (n239,n46,n240);
not (n240,n241);
nor (n241,n242,n243);
and (n242,n81,n41);
and (n243,n42,n79);
or (n244,n131,n47);
and (n245,n219,n226);
xor (n246,n85,n125);
and (n247,n215,n216);
nand (n248,n6,n212);
not (n249,n250);
nor (n250,n251,n450);
and (n251,n252,n431);
or (n252,n253,n430);
and (n253,n254,n322);
xor (n254,n255,n300);
or (n255,n256,n299);
and (n256,n257,n283);
xor (n257,n258,n267);
nand (n258,n259,n263);
or (n259,n64,n260);
nor (n260,n261,n262);
and (n261,n59,n16);
and (n262,n60,n18);
or (n263,n264,n82);
nor (n264,n265,n266);
and (n265,n59,n35);
and (n266,n60,n34);
and (n267,n268,n273);
and (n268,n269,n60);
nand (n269,n270,n271);
or (n270,n74,n69);
nand (n271,n272,n101);
or (n272,n68,n73);
nand (n273,n274,n279);
or (n274,n46,n275);
not (n275,n276);
nor (n276,n277,n278);
and (n277,n92,n41);
and (n278,n42,n90);
nand (n279,n280,n48);
nand (n280,n281,n282);
or (n281,n63,n42);
nand (n282,n42,n63);
xor (n283,n284,n290);
xor (n284,n285,n286);
and (n285,n148,n102);
nand (n286,n287,n288);
or (n287,n47,n240);
or (n288,n289,n46);
not (n289,n280);
nand (n290,n291,n295);
or (n291,n109,n292);
nor (n292,n293,n294);
and (n293,n73,n175);
and (n294,n74,n177);
or (n295,n110,n296);
nor (n296,n297,n298);
and (n297,n92,n74);
and (n298,n90,n73);
and (n299,n258,n267);
xor (n300,n301,n306);
xor (n301,n302,n303);
xor (n302,n233,n238);
or (n303,n304,n305);
and (n304,n284,n290);
and (n305,n285,n286);
xor (n306,n307,n319);
xor (n307,n308,n316);
nand (n308,n309,n314);
or (n309,n310,n153);
not (n310,n311);
nand (n311,n312,n313);
or (n312,n25,n101);
or (n313,n24,n102);
nand (n314,n315,n148);
not (n315,n159);
nand (n316,n317,n318);
or (n317,n296,n109);
nand (n318,n119,n222);
nand (n319,n320,n321);
or (n320,n64,n264);
or (n321,n228,n82);
or (n322,n323,n429);
and (n323,n324,n347);
xor (n324,n325,n346);
or (n325,n326,n345);
and (n326,n327,n344);
xor (n327,n328,n336);
nand (n328,n329,n334);
or (n329,n330,n109);
not (n330,n331);
nor (n331,n332,n333);
and (n332,n34,n73);
and (n333,n74,n35);
nand (n334,n335,n119);
not (n335,n292);
nand (n336,n337,n342);
or (n337,n338,n64);
not (n338,n339);
nand (n339,n340,n341);
or (n340,n60,n101);
or (n341,n59,n102);
nand (n342,n343,n71);
not (n343,n260);
xor (n344,n268,n273);
and (n345,n328,n336);
xor (n346,n257,n283);
nand (n347,n348,n428);
or (n348,n349,n423);
nor (n349,n350,n422);
and (n350,n351,n384);
nand (n351,n352,n370);
not (n352,n353);
xor (n353,n354,n363);
xor (n354,n355,n356);
and (n355,n71,n102);
nand (n356,n357,n362);
or (n357,n358,n109);
not (n358,n359);
nor (n359,n360,n361);
and (n360,n74,n16);
and (n361,n18,n73);
nand (n362,n119,n331);
nand (n363,n364,n365);
or (n364,n47,n275);
or (n365,n46,n366);
not (n366,n367);
nor (n367,n368,n369);
and (n368,n177,n41);
and (n369,n42,n175);
nand (n370,n371,n378);
nand (n371,n372,n373);
or (n372,n47,n366);
nand (n373,n374,n377);
nand (n374,n375,n376);
or (n375,n35,n41);
nand (n376,n41,n35);
not (n377,n46);
not (n378,n379);
nand (n379,n380,n74);
nand (n380,n381,n383);
or (n381,n382,n102);
nor (n382,n41,n114);
or (n383,n42,n112);
or (n384,n385,n421);
and (n385,n386,n398);
xor (n386,n387,n394);
nand (n387,n388,n393);
or (n388,n389,n109);
not (n389,n390);
nand (n390,n391,n392);
or (n391,n74,n101);
or (n392,n73,n102);
nand (n393,n119,n359);
nand (n394,n395,n397);
or (n395,n378,n396);
not (n396,n371);
nand (n397,n396,n378);
or (n398,n399,n420);
and (n399,n400,n410);
xor (n400,n401,n402);
nor (n401,n110,n101);
nand (n402,n403,n408);
or (n403,n46,n404);
not (n404,n405);
nand (n405,n406,n407);
or (n406,n16,n41);
nand (n407,n41,n16);
or (n408,n409,n47);
not (n409,n374);
nor (n410,n411,n418);
nor (n411,n412,n417);
and (n412,n413,n377);
not (n413,n414);
nor (n414,n415,n416);
and (n415,n41,n102);
and (n416,n42,n101);
and (n417,n405,n48);
or (n418,n419,n41);
nor (n419,n101,n47);
and (n420,n401,n402);
and (n421,n387,n394);
nor (n422,n352,n370);
nor (n423,n424,n425);
xor (n424,n327,n344);
or (n425,n426,n427);
and (n426,n354,n363);
and (n427,n355,n356);
nand (n428,n424,n425);
and (n429,n325,n346);
and (n430,n255,n300);
not (n431,n432);
nand (n432,n433,n445);
not (n433,n434);
nor (n434,n435,n436);
xor (n435,n214,n246);
or (n436,n437,n444);
and (n437,n438,n443);
xor (n438,n439,n442);
or (n439,n440,n441);
and (n440,n307,n319);
and (n441,n308,n316);
xor (n442,n127,n141);
xor (n443,n218,n232);
and (n444,n439,n442);
or (n445,n446,n447);
xor (n446,n438,n443);
or (n447,n448,n449);
and (n448,n301,n306);
and (n449,n302,n303);
nand (n450,n451,n453);
or (n451,n434,n452);
nand (n452,n446,n447);
nand (n453,n435,n436);
or (n454,n250,n3);
xor (n455,n456,n717);
xor (n456,n457,n714);
xor (n457,n458,n713);
xor (n458,n459,n704);
xor (n459,n460,n703);
xor (n460,n461,n689);
xor (n461,n462,n124);
xor (n462,n463,n669);
xor (n463,n464,n668);
xor (n464,n465,n641);
xor (n465,n466,n640);
xor (n466,n467,n608);
xor (n467,n468,n607);
xor (n468,n469,n569);
xor (n469,n470,n174);
xor (n470,n471,n526);
xor (n471,n472,n525);
xor (n472,n473,n475);
xor (n473,n474,n14);
and (n474,n195,n102);
or (n475,n476,n479);
and (n476,n477,n478);
and (n477,n15,n102);
and (n478,n26,n16);
and (n479,n480,n481);
xor (n480,n477,n478);
or (n481,n482,n485);
and (n482,n483,n484);
and (n483,n26,n102);
and (n484,n25,n16);
and (n485,n486,n487);
xor (n486,n483,n484);
or (n487,n488,n491);
and (n488,n489,n490);
and (n489,n25,n102);
and (n490,n150,n16);
and (n491,n492,n493);
xor (n492,n489,n490);
or (n493,n494,n497);
and (n494,n495,n496);
and (n495,n150,n102);
and (n496,n60,n16);
and (n497,n498,n499);
xor (n498,n495,n496);
or (n499,n500,n503);
and (n500,n501,n502);
and (n501,n60,n102);
and (n502,n69,n16);
and (n503,n504,n505);
xor (n504,n501,n502);
or (n505,n506,n508);
and (n506,n507,n360);
and (n507,n69,n102);
and (n508,n509,n510);
xor (n509,n507,n360);
or (n510,n511,n514);
and (n511,n512,n513);
and (n512,n74,n102);
and (n513,n112,n16);
and (n514,n515,n516);
xor (n515,n512,n513);
or (n516,n517,n520);
and (n517,n518,n519);
and (n518,n112,n102);
and (n519,n42,n16);
and (n520,n521,n522);
xor (n521,n518,n519);
and (n522,n523,n524);
and (n523,n42,n102);
and (n524,n48,n16);
and (n525,n26,n35);
or (n526,n527,n529);
and (n527,n528,n146);
xor (n528,n480,n481);
and (n529,n530,n531);
xor (n530,n528,n146);
or (n531,n532,n535);
and (n532,n533,n534);
xor (n533,n486,n487);
and (n534,n150,n35);
and (n535,n536,n537);
xor (n536,n533,n534);
or (n537,n538,n541);
and (n538,n539,n540);
xor (n539,n492,n493);
and (n540,n60,n35);
and (n541,n542,n543);
xor (n542,n539,n540);
or (n543,n544,n547);
and (n544,n545,n546);
xor (n545,n498,n499);
and (n546,n69,n35);
and (n547,n548,n549);
xor (n548,n545,n546);
or (n549,n550,n552);
and (n550,n551,n333);
xor (n551,n504,n505);
and (n552,n553,n554);
xor (n553,n551,n333);
or (n554,n555,n558);
and (n555,n556,n557);
xor (n556,n509,n510);
and (n557,n112,n35);
and (n558,n559,n560);
xor (n559,n556,n557);
or (n560,n561,n564);
and (n561,n562,n563);
xor (n562,n515,n516);
and (n563,n42,n35);
and (n564,n565,n566);
xor (n565,n562,n563);
and (n566,n567,n568);
xor (n567,n521,n522);
and (n568,n48,n35);
or (n569,n570,n573);
and (n570,n571,n572);
xor (n571,n530,n531);
and (n572,n150,n175);
and (n573,n574,n575);
xor (n574,n571,n572);
or (n575,n576,n579);
and (n576,n577,n578);
xor (n577,n536,n537);
and (n578,n60,n175);
and (n579,n580,n581);
xor (n580,n577,n578);
or (n581,n582,n585);
and (n582,n583,n584);
xor (n583,n542,n543);
and (n584,n69,n175);
and (n585,n586,n587);
xor (n586,n583,n584);
or (n587,n588,n591);
and (n588,n589,n590);
xor (n589,n548,n549);
and (n590,n74,n175);
and (n591,n592,n593);
xor (n592,n589,n590);
or (n593,n594,n597);
and (n594,n595,n596);
xor (n595,n553,n554);
and (n596,n112,n175);
and (n597,n598,n599);
xor (n598,n595,n596);
or (n599,n600,n602);
and (n600,n601,n369);
xor (n601,n559,n560);
and (n602,n603,n604);
xor (n603,n601,n369);
and (n604,n605,n606);
xor (n605,n565,n566);
and (n606,n48,n175);
and (n607,n150,n90);
or (n608,n609,n612);
and (n609,n610,n611);
xor (n610,n574,n575);
and (n611,n60,n90);
and (n612,n613,n614);
xor (n613,n610,n611);
or (n614,n615,n618);
and (n615,n616,n617);
xor (n616,n580,n581);
and (n617,n69,n90);
and (n618,n619,n620);
xor (n619,n616,n617);
or (n620,n621,n624);
and (n621,n622,n623);
xor (n622,n586,n587);
and (n623,n74,n90);
and (n624,n625,n626);
xor (n625,n622,n623);
or (n626,n627,n630);
and (n627,n628,n629);
xor (n628,n592,n593);
and (n629,n112,n90);
and (n630,n631,n632);
xor (n631,n628,n629);
or (n632,n633,n635);
and (n633,n634,n278);
xor (n634,n598,n599);
and (n635,n636,n637);
xor (n636,n634,n278);
and (n637,n638,n639);
xor (n638,n603,n604);
and (n639,n48,n90);
and (n640,n60,n61);
or (n641,n642,n645);
and (n642,n643,n644);
xor (n643,n613,n614);
and (n644,n69,n61);
and (n645,n646,n647);
xor (n646,n643,n644);
or (n647,n648,n651);
and (n648,n649,n650);
xor (n649,n619,n620);
and (n650,n74,n61);
and (n651,n652,n653);
xor (n652,n649,n650);
or (n653,n654,n657);
and (n654,n655,n656);
xor (n655,n625,n626);
and (n656,n112,n61);
and (n657,n658,n659);
xor (n658,n655,n656);
or (n659,n660,n663);
and (n660,n661,n662);
xor (n661,n631,n632);
and (n662,n42,n61);
and (n663,n664,n665);
xor (n664,n661,n662);
and (n665,n666,n667);
xor (n666,n636,n637);
and (n667,n48,n61);
and (n668,n69,n79);
or (n669,n670,n673);
and (n670,n671,n672);
xor (n671,n646,n647);
and (n672,n74,n79);
and (n673,n674,n675);
xor (n674,n671,n672);
or (n675,n676,n679);
and (n676,n677,n678);
xor (n677,n652,n653);
and (n678,n112,n79);
and (n679,n680,n681);
xor (n680,n677,n678);
or (n681,n682,n684);
and (n682,n683,n243);
xor (n683,n658,n659);
and (n684,n685,n686);
xor (n685,n683,n243);
and (n686,n687,n688);
xor (n687,n664,n665);
and (n688,n48,n79);
or (n689,n690,n693);
and (n690,n691,n692);
xor (n691,n674,n675);
and (n692,n112,n123);
and (n693,n694,n695);
xor (n694,n691,n692);
or (n695,n696,n698);
and (n696,n697,n134);
xor (n697,n680,n681);
and (n698,n699,n700);
xor (n699,n697,n134);
and (n700,n701,n702);
xor (n701,n685,n686);
and (n702,n48,n123);
and (n703,n112,n138);
or (n704,n705,n708);
and (n705,n706,n707);
xor (n706,n694,n695);
and (n707,n42,n138);
and (n708,n709,n710);
xor (n709,n706,n707);
and (n710,n711,n712);
xor (n711,n699,n700);
and (n712,n48,n138);
and (n713,n42,n43);
and (n714,n715,n716);
xor (n715,n709,n710);
and (n716,n48,n43);
and (n717,n48,n53);
endmodule
