module top (out,n19,n24,n25,n26,n28,n29,n40,n43,n45
        ,n48,n51,n61,n71,n76,n79,n82,n85,n88,n91
        ,n93,n95,n103,n116,n121,n137,n149,n154,n157,n160
        ,n167,n177,n358,n371);
output out;
input n19;
input n24;
input n25;
input n26;
input n28;
input n29;
input n40;
input n43;
input n45;
input n48;
input n51;
input n61;
input n71;
input n76;
input n79;
input n82;
input n85;
input n88;
input n91;
input n93;
input n95;
input n103;
input n116;
input n121;
input n137;
input n149;
input n154;
input n157;
input n160;
input n167;
input n177;
input n358;
input n371;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n20;
wire n21;
wire n22;
wire n23;
wire n27;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n41;
wire n42;
wire n44;
wire n46;
wire n47;
wire n49;
wire n50;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n72;
wire n73;
wire n74;
wire n75;
wire n77;
wire n78;
wire n80;
wire n81;
wire n83;
wire n84;
wire n86;
wire n87;
wire n89;
wire n90;
wire n92;
wire n94;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n117;
wire n118;
wire n119;
wire n120;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n150;
wire n151;
wire n152;
wire n153;
wire n155;
wire n156;
wire n158;
wire n159;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
xor (out,n0,n724);
nand (n0,n1,n722);
or (n1,n2,n453);
not (n2,n3);
and (n3,n4,n452);
or (n4,n5,n407);
xor (n5,n6,n348);
xor (n6,n7,n270);
xor (n7,n8,n181);
xor (n8,n9,n109);
nand (n9,n10,n98);
or (n10,n11,n67);
nand (n11,n12,n56);
not (n12,n13);
nand (n13,n14,n55);
or (n14,n15,n49);
not (n15,n16);
wire s0n16,s1n16,notn16;
or (n16,s0n16,s1n16);
not(notn16,n46);
and (s0n16,notn16,n17);
and (s1n16,n46,n36);
wire s0n17,s1n17,notn17;
or (n17,s0n17,s1n17);
not(notn17,n20);
and (s0n17,notn17,1'b0);
and (s1n17,n20,n19);
or (n20,n21,n32);
or (n21,n22,n30);
nor (n22,n23,n25,n26,n27,n29);
not (n23,n24);
not (n27,n28);
nor (n30,n24,n31,n26,n27,n29);
not (n31,n25);
or (n32,n33,n35);
and (n33,n23,n25,n26,n27,n34);
not (n34,n29);
nor (n35,n23,n31,n26,n27,n29);
xor (n36,n37,n38);
not (n37,n19);
and (n38,n39,n41);
not (n39,n40);
and (n41,n42,n44);
not (n42,n43);
not (n44,n45);
and (n46,n47,n48);
or (n47,n22,n33);
wire s0n49,s1n49,notn49;
or (n49,s0n49,s1n49);
not(notn49,n46);
and (s0n49,notn49,n50);
and (s1n49,n46,n52);
wire s0n50,s1n50,notn50;
or (n50,s0n50,s1n50);
not(notn50,n20);
and (s0n50,notn50,1'b0);
and (s1n50,n20,n51);
xor (n52,n53,n54);
not (n53,n51);
and (n54,n37,n38);
nand (n55,n49,n15);
nor (n56,n57,n66);
and (n57,n58,n65);
not (n58,n59);
wire s0n59,s1n59,notn59;
or (n59,s0n59,s1n59);
not(notn59,n46);
and (s0n59,notn59,n60);
and (s1n59,n46,n62);
wire s0n60,s1n60,notn60;
or (n60,s0n60,s1n60);
not(notn60,n20);
and (s0n60,notn60,1'b0);
and (s1n60,n20,n61);
xor (n62,n63,n64);
not (n63,n61);
and (n64,n53,n54);
not (n65,n49);
and (n66,n59,n49);
nor (n67,n68,n96);
and (n68,n69,n58);
wire s0n69,s1n69,notn69;
or (n69,s0n69,s1n69);
not(notn69,n94);
and (s0n69,notn69,n70);
and (s1n69,n94,n72);
wire s0n70,s1n70,notn70;
or (n70,s0n70,s1n70);
not(notn70,n20);
and (s0n70,notn70,1'b0);
and (s1n70,n20,n71);
xor (n72,n73,n74);
not (n73,n71);
and (n74,n75,n77);
not (n75,n76);
and (n77,n78,n80);
not (n78,n79);
and (n80,n81,n83);
not (n81,n82);
and (n83,n84,n86);
not (n84,n85);
and (n86,n87,n89);
not (n87,n88);
and (n89,n90,n92);
not (n90,n91);
not (n92,n93);
and (n94,n47,n95);
and (n96,n97,n59);
not (n97,n69);
or (n98,n12,n99);
nor (n99,n100,n107);
and (n100,n101,n58);
wire s0n101,s1n101,notn101;
or (n101,s0n101,s1n101);
not(notn101,n94);
and (s0n101,notn101,n102);
and (s1n101,n94,n104);
wire s0n102,s1n102,notn102;
or (n102,s0n102,s1n102);
not(notn102,n20);
and (s0n102,notn102,1'b0);
and (s1n102,n20,n103);
xor (n104,n105,n106);
not (n105,n103);
and (n106,n73,n74);
and (n107,n108,n59);
not (n108,n101);
and (n109,n110,n143);
nand (n110,n111,n132);
or (n111,n112,n129);
nor (n112,n113,n127);
and (n113,n114,n123);
wire s0n114,s1n114,notn114;
or (n114,s0n114,s1n114);
not(notn114,n94);
and (s0n114,notn114,n115);
and (s1n114,n94,n117);
wire s0n115,s1n115,notn115;
or (n115,s0n115,s1n115);
not(notn115,n20);
and (s0n115,notn115,1'b0);
and (s1n115,n20,n116);
xor (n117,n118,n119);
not (n118,n116);
and (n119,n120,n122);
not (n120,n121);
and (n122,n105,n106);
not (n123,n124);
wire s0n124,s1n124,notn124;
or (n124,s0n124,s1n124);
not(notn124,n46);
and (s0n124,notn124,n125);
and (s1n124,n46,n126);
wire s0n125,s1n125,notn125;
or (n125,s0n125,s1n125);
not(notn125,n20);
and (s0n125,notn125,1'b0);
and (s1n125,n20,n43);
xor (n126,n42,n44);
and (n127,n128,n124);
not (n128,n114);
nand (n129,n124,n130);
not (n130,n131);
wire s0n131,s1n131,notn131;
or (n131,s0n131,s1n131);
not(notn131,n20);
and (s0n131,notn131,1'b0);
and (s1n131,n20,n45);
or (n132,n133,n130);
nor (n133,n134,n141);
and (n134,n123,n135);
wire s0n135,s1n135,notn135;
or (n135,s0n135,s1n135);
not(notn135,n94);
and (s0n135,notn135,n136);
and (s1n135,n94,n138);
wire s0n136,s1n136,notn136;
or (n136,s0n136,s1n136);
not(notn136,n20);
and (s0n136,notn136,1'b0);
and (s1n136,n20,n137);
xor (n138,n139,n140);
not (n139,n137);
and (n140,n118,n119);
and (n141,n142,n124);
not (n142,n135);
nor (n143,n144,n174);
nor (n144,n145,n171);
and (n145,n146,n162);
not (n146,n147);
wire s0n147,s1n147,notn147;
or (n147,s0n147,s1n147);
not(notn147,n46);
and (s0n147,notn147,n148);
and (s1n147,n46,n150);
wire s0n148,s1n148,notn148;
or (n148,s0n148,s1n148);
not(notn148,n20);
and (s0n148,notn148,1'b0);
and (s1n148,n20,n149);
xor (n150,n151,n152);
not (n151,n149);
and (n152,n153,n155);
not (n153,n154);
and (n155,n156,n158);
not (n156,n157);
and (n158,n159,n161);
not (n159,n160);
and (n161,n63,n64);
not (n162,n163);
and (n163,n164,n165);
wire s0n164,s1n164,notn164;
or (n164,s0n164,s1n164);
not(notn164,n20);
and (s0n164,notn164,1'b0);
and (s1n164,n20,n93);
wire s0n165,s1n165,notn165;
or (n165,s0n165,s1n165);
not(notn165,n46);
and (s0n165,notn165,n166);
and (s1n165,n46,n168);
wire s0n166,s1n166,notn166;
or (n166,s0n166,s1n166);
not(notn166,n20);
and (s0n166,notn166,1'b0);
and (s1n166,n20,n167);
xor (n168,n169,n170);
not (n169,n167);
and (n170,n151,n152);
and (n171,n172,n173);
not (n172,n165);
not (n173,n164);
not (n174,n175);
wire s0n175,s1n175,notn175;
or (n175,s0n175,s1n175);
not(notn175,n46);
and (s0n175,notn175,n176);
and (s1n175,n46,n178);
wire s0n176,s1n176,notn176;
or (n176,s0n176,s1n176);
not(notn176,n20);
and (s0n176,notn176,1'b0);
and (s1n176,n20,n177);
xor (n178,n179,n180);
not (n179,n177);
and (n180,n169,n170);
or (n181,n182,n269);
and (n182,n183,n240);
xor (n183,n184,n208);
nand (n184,n185,n200);
or (n185,n186,n197);
nand (n186,n187,n194);
nor (n187,n188,n192);
and (n188,n123,n189);
wire s0n189,s1n189,notn189;
or (n189,s0n189,s1n189);
not(notn189,n46);
and (s0n189,notn189,n190);
and (s1n189,n46,n191);
wire s0n190,s1n190,notn190;
or (n190,s0n190,s1n190);
not(notn190,n20);
and (s0n190,notn190,1'b0);
and (s1n190,n20,n40);
xor (n191,n39,n41);
and (n192,n124,n193);
not (n193,n189);
nand (n194,n195,n196);
or (n195,n15,n189);
nand (n196,n15,n189);
nor (n197,n198,n199);
and (n198,n101,n15);
and (n199,n108,n16);
or (n200,n187,n201);
nor (n201,n202,n206);
and (n202,n203,n15);
wire s0n203,s1n203,notn203;
or (n203,s0n203,s1n203);
not(notn203,n94);
and (s0n203,notn203,n204);
and (s1n203,n94,n205);
wire s0n204,s1n204,notn204;
or (n204,s0n204,s1n204);
not(notn204,n20);
and (s0n204,notn204,1'b0);
and (s1n204,n20,n121);
xor (n205,n120,n122);
and (n206,n207,n16);
not (n207,n203);
nand (n208,n209,n232);
or (n209,n210,n225);
nand (n210,n211,n218);
or (n211,n212,n216);
and (n212,n59,n213);
wire s0n213,s1n213,notn213;
or (n213,s0n213,s1n213);
not(notn213,n46);
and (s0n213,notn213,n214);
and (s1n213,n46,n215);
wire s0n214,s1n214,notn214;
or (n214,s0n214,s1n214);
not(notn214,n20);
and (s0n214,notn214,1'b0);
and (s1n214,n20,n160);
xor (n215,n159,n161);
and (n216,n58,n217);
not (n217,n213);
nor (n218,n219,n223);
and (n219,n220,n213);
wire s0n220,s1n220,notn220;
or (n220,s0n220,s1n220);
not(notn220,n46);
and (s0n220,notn220,n221);
and (s1n220,n46,n222);
wire s0n221,s1n221,notn221;
or (n221,s0n221,s1n221);
not(notn221,n20);
and (s0n221,notn221,1'b0);
and (s1n221,n20,n157);
xor (n222,n156,n158);
and (n223,n224,n217);
not (n224,n220);
nor (n225,n226,n230);
and (n226,n227,n224);
wire s0n227,s1n227,notn227;
or (n227,s0n227,s1n227);
not(notn227,n94);
and (s0n227,notn227,n228);
and (s1n227,n94,n229);
wire s0n228,s1n228,notn228;
or (n228,s0n228,s1n228);
not(notn228,n20);
and (s0n228,notn228,1'b0);
and (s1n228,n20,n82);
xor (n229,n81,n83);
and (n230,n231,n220);
not (n231,n227);
or (n232,n233,n211);
nor (n233,n234,n238);
and (n234,n235,n224);
wire s0n235,s1n235,notn235;
or (n235,s0n235,s1n235);
not(notn235,n94);
and (s0n235,notn235,n236);
and (s1n235,n94,n237);
wire s0n236,s1n236,notn236;
or (n236,s0n236,s1n236);
not(notn236,n20);
and (s0n236,notn236,1'b0);
and (s1n236,n20,n79);
xor (n237,n78,n80);
and (n238,n239,n220);
not (n239,n235);
nand (n240,n241,n261);
or (n241,n242,n254);
nand (n242,n243,n250);
nor (n243,n244,n248);
and (n244,n245,n147);
wire s0n245,s1n245,notn245;
or (n245,s0n245,s1n245);
not(notn245,n46);
and (s0n245,notn245,n246);
and (s1n245,n46,n247);
wire s0n246,s1n246,notn246;
or (n246,s0n246,s1n246);
not(notn246,n20);
and (s0n246,notn246,1'b0);
and (s1n246,n20,n154);
xor (n247,n153,n155);
and (n248,n249,n146);
not (n249,n245);
not (n250,n251);
nor (n251,n252,n253);
and (n252,n220,n245);
and (n253,n224,n249);
nor (n254,n255,n259);
and (n255,n256,n146);
wire s0n256,s1n256,notn256;
or (n256,s0n256,s1n256);
not(notn256,n94);
and (s0n256,notn256,n257);
and (s1n256,n94,n258);
wire s0n257,s1n257,notn257;
or (n257,s0n257,s1n257);
not(notn257,n20);
and (s0n257,notn257,1'b0);
and (s1n257,n20,n88);
xor (n258,n87,n89);
and (n259,n260,n147);
not (n260,n256);
or (n261,n262,n250);
nor (n262,n263,n267);
and (n263,n146,n264);
wire s0n264,s1n264,notn264;
or (n264,s0n264,s1n264);
not(notn264,n94);
and (s0n264,notn264,n265);
and (s1n264,n94,n266);
wire s0n265,s1n265,notn265;
or (n265,s0n265,s1n265);
not(notn265,n20);
and (s0n265,notn265,1'b0);
and (s1n265,n20,n85);
xor (n266,n84,n86);
and (n267,n147,n268);
not (n268,n264);
and (n269,n184,n208);
or (n270,n271,n347);
and (n271,n272,n328);
xor (n272,n273,n293);
or (n273,n274,n292);
and (n274,n275,n286);
xor (n275,n276,n280);
nor (n276,n277,n173);
or (n277,n278,n279);
and (n278,n165,n147);
and (n279,n172,n146);
nand (n280,n281,n285);
or (n281,n282,n129);
nor (n282,n283,n284);
and (n283,n123,n203);
and (n284,n207,n124);
or (n285,n112,n130);
nand (n286,n287,n291);
or (n287,n186,n288);
nor (n288,n289,n290);
and (n289,n69,n15);
and (n290,n97,n16);
or (n291,n187,n197);
and (n292,n276,n280);
or (n293,n294,n327);
and (n294,n295,n314);
xor (n295,n296,n303);
nand (n296,n297,n302);
or (n297,n210,n298);
not (n298,n299);
nor (n299,n300,n301);
and (n300,n224,n268);
and (n301,n264,n220);
or (n302,n225,n211);
nand (n303,n304,n313);
or (n304,n305,n242);
not (n305,n306);
nand (n306,n307,n312);
or (n307,n308,n147);
not (n308,n309);
wire s0n309,s1n309,notn309;
or (n309,s0n309,s1n309);
not(notn309,n94);
and (s0n309,notn309,n310);
and (s1n309,n94,n311);
wire s0n310,s1n310,notn310;
or (n310,s0n310,s1n310);
not(notn310,n20);
and (s0n310,notn310,1'b0);
and (s1n310,n20,n91);
xor (n311,n90,n92);
or (n312,n309,n146);
or (n313,n254,n250);
nand (n314,n315,n319);
or (n315,n11,n316);
nor (n316,n317,n318);
and (n317,n235,n58);
and (n318,n239,n59);
or (n319,n12,n320);
nor (n320,n321,n325);
and (n321,n322,n58);
wire s0n322,s1n322,notn322;
or (n322,s0n322,s1n322);
not(notn322,n94);
and (s0n322,notn322,n323);
and (s1n322,n94,n324);
wire s0n323,s1n323,notn323;
or (n323,s0n323,s1n323);
not(notn323,n20);
and (s0n323,notn323,1'b0);
and (s1n323,n20,n76);
xor (n324,n75,n77);
and (n325,n326,n59);
not (n326,n322);
and (n327,n296,n303);
xor (n328,n329,n346);
xor (n329,n330,n343);
nand (n330,n331,n339);
or (n331,n332,n336);
nand (n332,n277,n333);
nand (n333,n334,n335);
or (n334,n172,n175);
or (n335,n174,n165);
nor (n336,n337,n338);
and (n337,n175,n173);
and (n338,n174,n164);
or (n339,n340,n277);
nor (n340,n341,n342);
and (n341,n309,n174);
and (n342,n308,n175);
nand (n343,n344,n345);
or (n344,n11,n320);
or (n345,n67,n12);
xor (n346,n110,n143);
and (n347,n273,n293);
xor (n348,n349,n404);
xor (n349,n350,n383);
xor (n350,n351,n377);
xor (n351,n352,n364);
nor (n352,n353,n173);
not (n353,n354);
nor (n354,n355,n362);
and (n355,n356,n175);
wire s0n356,s1n356,notn356;
or (n356,s0n356,s1n356);
not(notn356,n46);
and (s0n356,notn356,n357);
and (s1n356,n46,n359);
wire s0n357,s1n357,notn357;
or (n357,s0n357,s1n357);
not(notn357,n20);
and (s0n357,notn357,1'b0);
and (s1n357,n20,n358);
xor (n359,n360,n361);
not (n360,n358);
and (n361,n179,n180);
and (n362,n363,n174);
not (n363,n356);
nand (n364,n365,n366);
or (n365,n133,n129);
or (n366,n367,n130);
nor (n367,n368,n375);
and (n368,n123,n369);
wire s0n369,s1n369,notn369;
or (n369,s0n369,s1n369);
not(notn369,n94);
and (s0n369,notn369,n370);
and (s1n369,n94,n372);
wire s0n370,s1n370,notn370;
or (n370,s0n370,s1n370);
not(notn370,n20);
and (s0n370,notn370,1'b0);
and (s1n370,n20,n371);
xor (n372,n373,n374);
not (n373,n371);
and (n374,n139,n140);
and (n375,n376,n124);
not (n376,n369);
nand (n377,n378,n382);
or (n378,n187,n379);
nor (n379,n380,n381);
and (n380,n15,n114);
and (n381,n128,n16);
or (n382,n186,n201);
xor (n383,n384,n398);
xor (n384,n385,n391);
nand (n385,n386,n387);
or (n386,n210,n233);
or (n387,n388,n211);
nor (n388,n389,n390);
and (n389,n322,n224);
and (n390,n326,n220);
nand (n391,n392,n397);
or (n392,n250,n393);
not (n393,n394);
nand (n394,n395,n396);
or (n395,n147,n231);
or (n396,n146,n227);
or (n397,n242,n262);
nand (n398,n399,n403);
or (n399,n277,n400);
nor (n400,n401,n402);
and (n401,n256,n174);
and (n402,n260,n175);
or (n403,n332,n340);
or (n404,n405,n406);
and (n405,n329,n346);
and (n406,n330,n343);
or (n407,n408,n451);
and (n408,n409,n450);
xor (n409,n410,n411);
xor (n410,n183,n240);
or (n411,n412,n449);
and (n412,n413,n427);
xor (n413,n414,n426);
and (n414,n415,n421);
nor (n415,n416,n146);
nor (n416,n417,n420);
and (n417,n418,n224);
not (n418,n419);
and (n419,n164,n245);
and (n420,n249,n173);
nand (n421,n422,n425);
or (n422,n129,n423);
not (n423,n424);
xnor (n424,n101,n123);
or (n425,n282,n130);
xor (n426,n275,n286);
or (n427,n428,n448);
and (n428,n429,n442);
xor (n429,n430,n436);
nand (n430,n431,n435);
or (n431,n186,n432);
nor (n432,n433,n434);
and (n433,n15,n322);
and (n434,n326,n16);
or (n435,n288,n187);
nand (n436,n437,n438);
or (n437,n211,n298);
or (n438,n439,n210);
nor (n439,n440,n441);
and (n440,n256,n224);
and (n441,n260,n220);
nand (n442,n443,n444);
or (n443,n250,n305);
or (n444,n242,n445);
nor (n445,n446,n447);
and (n446,n147,n173);
and (n447,n146,n164);
and (n448,n430,n436);
and (n449,n414,n426);
xor (n450,n272,n328);
and (n451,n410,n411);
nand (n452,n5,n407);
or (n453,n454,n721);
and (n454,n455,n491);
xor (n455,n456,n490);
or (n456,n457,n489);
and (n457,n458,n488);
xor (n458,n459,n460);
xor (n459,n295,n314);
or (n460,n461,n487);
and (n461,n462,n470);
xor (n462,n463,n469);
nand (n463,n464,n468);
or (n464,n11,n465);
nor (n465,n466,n467);
and (n466,n227,n58);
and (n467,n231,n59);
or (n468,n316,n12);
xor (n469,n415,n421);
or (n470,n471,n486);
and (n471,n472,n480);
xor (n472,n473,n474);
nor (n473,n250,n173);
nand (n474,n475,n476);
or (n475,n130,n423);
or (n476,n477,n129);
nor (n477,n478,n479);
and (n478,n123,n69);
and (n479,n97,n124);
nand (n480,n481,n485);
or (n481,n210,n482);
nor (n482,n483,n484);
and (n483,n309,n224);
and (n484,n308,n220);
or (n485,n439,n211);
and (n486,n473,n474);
and (n487,n463,n469);
xor (n488,n413,n427);
and (n489,n459,n460);
xor (n490,n409,n450);
or (n491,n492,n720);
and (n492,n493,n530);
xor (n493,n494,n529);
or (n494,n495,n528);
and (n495,n496,n527);
xor (n496,n497,n526);
or (n497,n498,n525);
and (n498,n499,n512);
xor (n499,n500,n506);
nand (n500,n501,n505);
or (n501,n186,n502);
nor (n502,n503,n504);
and (n503,n235,n15);
and (n504,n16,n239);
or (n505,n432,n187);
nand (n506,n507,n511);
or (n507,n11,n508);
nor (n508,n509,n510);
and (n509,n264,n58);
and (n510,n268,n59);
or (n511,n465,n12);
and (n512,n513,n519);
nor (n513,n514,n224);
nor (n514,n515,n518);
and (n515,n516,n58);
not (n516,n517);
and (n517,n164,n213);
and (n518,n217,n173);
nand (n519,n520,n524);
or (n520,n521,n129);
nor (n521,n522,n523);
and (n522,n123,n322);
and (n523,n326,n124);
or (n524,n477,n130);
and (n525,n500,n506);
xor (n526,n429,n442);
xor (n527,n462,n470);
and (n528,n497,n526);
xor (n529,n458,n488);
nand (n530,n531,n717,n719);
or (n531,n532,n590);
nand (n532,n533,n585);
not (n533,n534);
nor (n534,n535,n561);
xor (n535,n536,n560);
xor (n536,n537,n559);
or (n537,n538,n558);
and (n538,n539,n552);
xor (n539,n540,n546);
nand (n540,n541,n545);
or (n541,n210,n542);
nor (n542,n543,n544);
and (n543,n220,n173);
and (n544,n224,n164);
or (n545,n482,n211);
nand (n546,n547,n551);
or (n547,n548,n186);
nor (n548,n549,n550);
and (n549,n16,n231);
and (n550,n15,n227);
or (n551,n502,n187);
nand (n552,n553,n557);
or (n553,n11,n554);
nor (n554,n555,n556);
and (n555,n256,n58);
and (n556,n260,n59);
or (n557,n508,n12);
and (n558,n540,n546);
xor (n559,n472,n480);
xor (n560,n499,n512);
or (n561,n562,n584);
and (n562,n563,n583);
xor (n563,n564,n565);
xor (n564,n513,n519);
or (n565,n566,n582);
and (n566,n567,n576);
xor (n567,n568,n569);
nor (n568,n211,n173);
nand (n569,n570,n575);
or (n570,n571,n129);
not (n571,n572);
nand (n572,n573,n574);
or (n573,n124,n239);
nand (n574,n239,n124);
or (n575,n521,n130);
nand (n576,n577,n581);
or (n577,n186,n578);
nor (n578,n579,n580);
and (n579,n15,n264);
and (n580,n16,n268);
or (n581,n548,n187);
and (n582,n568,n569);
xor (n583,n539,n552);
and (n584,n564,n565);
or (n585,n586,n587);
xor (n586,n496,n527);
or (n587,n588,n589);
and (n588,n536,n560);
and (n589,n537,n559);
nor (n590,n591,n716);
and (n591,n592,n711);
or (n592,n593,n710);
and (n593,n594,n635);
xor (n594,n595,n628);
or (n595,n596,n627);
and (n596,n597,n613);
xor (n597,n598,n604);
nand (n598,n599,n603);
or (n599,n186,n600);
nor (n600,n601,n602);
and (n601,n16,n260);
and (n602,n15,n256);
or (n603,n578,n187);
or (n604,n605,n609);
nor (n605,n606,n12);
nor (n606,n607,n608);
and (n607,n58,n309);
and (n608,n59,n308);
nor (n609,n11,n610);
nor (n610,n611,n612);
and (n611,n59,n173);
and (n612,n58,n164);
xor (n613,n614,n620);
nor (n614,n615,n58);
nor (n615,n616,n619);
and (n616,n617,n15);
not (n617,n618);
and (n618,n164,n49);
and (n619,n65,n173);
nand (n620,n621,n626);
or (n621,n129,n622);
not (n622,n623);
nand (n623,n624,n625);
or (n624,n123,n227);
nand (n625,n227,n123);
nand (n626,n572,n131);
and (n627,n598,n604);
xor (n628,n629,n634);
xor (n629,n630,n633);
nand (n630,n631,n632);
or (n631,n11,n606);
or (n632,n554,n12);
and (n633,n614,n620);
xor (n634,n567,n576);
or (n635,n636,n709);
and (n636,n637,n657);
xor (n637,n638,n656);
or (n638,n639,n655);
and (n639,n640,n649);
xor (n640,n641,n642);
and (n641,n13,n164);
nand (n642,n643,n648);
or (n643,n129,n644);
not (n644,n645);
nand (n645,n646,n647);
or (n646,n124,n268);
nand (n647,n268,n124);
nand (n648,n623,n131);
nand (n649,n650,n654);
or (n650,n186,n651);
nor (n651,n652,n653);
and (n652,n15,n309);
and (n653,n16,n308);
or (n654,n600,n187);
and (n655,n641,n642);
xor (n656,n597,n613);
or (n657,n658,n708);
and (n658,n659,n676);
xor (n659,n660,n675);
and (n660,n661,n667);
and (n661,n662,n16);
nand (n662,n663,n666);
nand (n663,n664,n123);
not (n664,n665);
and (n665,n164,n189);
nand (n666,n193,n173);
nand (n667,n668,n669);
or (n668,n130,n644);
nand (n669,n670,n674);
not (n670,n671);
nor (n671,n672,n673);
and (n672,n260,n124);
and (n673,n256,n123);
not (n674,n129);
xor (n675,n640,n649);
or (n676,n677,n707);
and (n677,n678,n686);
xor (n678,n679,n685);
nand (n679,n680,n684);
or (n680,n186,n681);
nor (n681,n682,n683);
and (n682,n16,n173);
and (n683,n15,n164);
or (n684,n651,n187);
xor (n685,n661,n667);
or (n686,n687,n706);
and (n687,n688,n696);
xor (n688,n689,n690);
nor (n689,n187,n173);
nand (n690,n691,n695);
or (n691,n692,n129);
or (n692,n693,n694);
and (n693,n123,n308);
and (n694,n309,n124);
or (n695,n671,n130);
nor (n696,n697,n704);
nor (n697,n698,n700);
and (n698,n699,n131);
not (n699,n692);
and (n700,n701,n674);
nand (n701,n702,n703);
or (n702,n123,n164);
or (n703,n124,n173);
or (n704,n123,n705);
and (n705,n164,n131);
and (n706,n689,n690);
and (n707,n679,n685);
and (n708,n660,n675);
and (n709,n638,n656);
and (n710,n595,n628);
or (n711,n712,n713);
xor (n712,n563,n583);
or (n713,n714,n715);
and (n714,n629,n634);
and (n715,n630,n633);
and (n716,n712,n713);
nand (n717,n585,n718);
and (n718,n535,n561);
nand (n719,n586,n587);
and (n720,n494,n529);
and (n721,n456,n490);
or (n722,n723,n3);
not (n723,n453);
xor (n724,n725,n1115);
xor (n725,n726,n1112);
xor (n726,n727,n1111);
xor (n727,n728,n1103);
xor (n728,n729,n1102);
xor (n729,n730,n1087);
xor (n730,n731,n1086);
xor (n731,n732,n1066);
xor (n732,n733,n1065);
xor (n733,n734,n1039);
xor (n734,n735,n1038);
xor (n735,n736,n1006);
xor (n736,n737,n1005);
xor (n737,n738,n966);
xor (n738,n739,n965);
xor (n739,n740,n921);
xor (n740,n741,n920);
xor (n741,n742,n869);
xor (n742,n743,n868);
xor (n743,n744,n812);
xor (n744,n745,n811);
xor (n745,n746,n749);
xor (n746,n747,n748);
and (n747,n369,n131);
and (n748,n135,n124);
or (n749,n750,n753);
and (n750,n751,n752);
and (n751,n135,n131);
and (n752,n114,n124);
and (n753,n754,n755);
xor (n754,n751,n752);
or (n755,n756,n759);
and (n756,n757,n758);
and (n757,n114,n131);
and (n758,n203,n124);
and (n759,n760,n761);
xor (n760,n757,n758);
or (n761,n762,n765);
and (n762,n763,n764);
and (n763,n203,n131);
and (n764,n101,n124);
and (n765,n766,n767);
xor (n766,n763,n764);
or (n767,n768,n771);
and (n768,n769,n770);
and (n769,n101,n131);
and (n770,n69,n124);
and (n771,n772,n773);
xor (n772,n769,n770);
or (n773,n774,n777);
and (n774,n775,n776);
and (n775,n69,n131);
and (n776,n322,n124);
and (n777,n778,n779);
xor (n778,n775,n776);
or (n779,n780,n783);
and (n780,n781,n782);
and (n781,n322,n131);
and (n782,n235,n124);
and (n783,n784,n785);
xor (n784,n781,n782);
or (n785,n786,n789);
and (n786,n787,n788);
and (n787,n235,n131);
and (n788,n227,n124);
and (n789,n790,n791);
xor (n790,n787,n788);
or (n791,n792,n795);
and (n792,n793,n794);
and (n793,n227,n131);
and (n794,n264,n124);
and (n795,n796,n797);
xor (n796,n793,n794);
or (n797,n798,n801);
and (n798,n799,n800);
and (n799,n264,n131);
and (n800,n256,n124);
and (n801,n802,n803);
xor (n802,n799,n800);
or (n803,n804,n806);
and (n804,n805,n694);
and (n805,n256,n131);
and (n806,n807,n808);
xor (n807,n805,n694);
and (n808,n809,n810);
and (n809,n309,n131);
and (n810,n164,n124);
and (n811,n114,n189);
or (n812,n813,n816);
and (n813,n814,n815);
xor (n814,n754,n755);
and (n815,n203,n189);
and (n816,n817,n818);
xor (n817,n814,n815);
or (n818,n819,n822);
and (n819,n820,n821);
xor (n820,n760,n761);
and (n821,n101,n189);
and (n822,n823,n824);
xor (n823,n820,n821);
or (n824,n825,n828);
and (n825,n826,n827);
xor (n826,n766,n767);
and (n827,n69,n189);
and (n828,n829,n830);
xor (n829,n826,n827);
or (n830,n831,n834);
and (n831,n832,n833);
xor (n832,n772,n773);
and (n833,n322,n189);
and (n834,n835,n836);
xor (n835,n832,n833);
or (n836,n837,n840);
and (n837,n838,n839);
xor (n838,n778,n779);
and (n839,n235,n189);
and (n840,n841,n842);
xor (n841,n838,n839);
or (n842,n843,n846);
and (n843,n844,n845);
xor (n844,n784,n785);
and (n845,n227,n189);
and (n846,n847,n848);
xor (n847,n844,n845);
or (n848,n849,n852);
and (n849,n850,n851);
xor (n850,n790,n791);
and (n851,n264,n189);
and (n852,n853,n854);
xor (n853,n850,n851);
or (n854,n855,n858);
and (n855,n856,n857);
xor (n856,n796,n797);
and (n857,n256,n189);
and (n858,n859,n860);
xor (n859,n856,n857);
or (n860,n861,n864);
and (n861,n862,n863);
xor (n862,n802,n803);
and (n863,n309,n189);
and (n864,n865,n866);
xor (n865,n862,n863);
and (n866,n867,n665);
xor (n867,n807,n808);
and (n868,n203,n16);
or (n869,n870,n873);
and (n870,n871,n872);
xor (n871,n817,n818);
and (n872,n101,n16);
and (n873,n874,n875);
xor (n874,n871,n872);
or (n875,n876,n879);
and (n876,n877,n878);
xor (n877,n823,n824);
and (n878,n69,n16);
and (n879,n880,n881);
xor (n880,n877,n878);
or (n881,n882,n885);
and (n882,n883,n884);
xor (n883,n829,n830);
and (n884,n322,n16);
and (n885,n886,n887);
xor (n886,n883,n884);
or (n887,n888,n891);
and (n888,n889,n890);
xor (n889,n835,n836);
and (n890,n235,n16);
and (n891,n892,n893);
xor (n892,n889,n890);
or (n893,n894,n897);
and (n894,n895,n896);
xor (n895,n841,n842);
and (n896,n227,n16);
and (n897,n898,n899);
xor (n898,n895,n896);
or (n899,n900,n903);
and (n900,n901,n902);
xor (n901,n847,n848);
and (n902,n264,n16);
and (n903,n904,n905);
xor (n904,n901,n902);
or (n905,n906,n909);
and (n906,n907,n908);
xor (n907,n853,n854);
and (n908,n256,n16);
and (n909,n910,n911);
xor (n910,n907,n908);
or (n911,n912,n915);
and (n912,n913,n914);
xor (n913,n859,n860);
and (n914,n309,n16);
and (n915,n916,n917);
xor (n916,n913,n914);
and (n917,n918,n919);
xor (n918,n865,n866);
and (n919,n164,n16);
and (n920,n101,n49);
or (n921,n922,n925);
and (n922,n923,n924);
xor (n923,n874,n875);
and (n924,n69,n49);
and (n925,n926,n927);
xor (n926,n923,n924);
or (n927,n928,n931);
and (n928,n929,n930);
xor (n929,n880,n881);
and (n930,n322,n49);
and (n931,n932,n933);
xor (n932,n929,n930);
or (n933,n934,n937);
and (n934,n935,n936);
xor (n935,n886,n887);
and (n936,n235,n49);
and (n937,n938,n939);
xor (n938,n935,n936);
or (n939,n940,n943);
and (n940,n941,n942);
xor (n941,n892,n893);
and (n942,n227,n49);
and (n943,n944,n945);
xor (n944,n941,n942);
or (n945,n946,n949);
and (n946,n947,n948);
xor (n947,n898,n899);
and (n948,n264,n49);
and (n949,n950,n951);
xor (n950,n947,n948);
or (n951,n952,n955);
and (n952,n953,n954);
xor (n953,n904,n905);
and (n954,n256,n49);
and (n955,n956,n957);
xor (n956,n953,n954);
or (n957,n958,n961);
and (n958,n959,n960);
xor (n959,n910,n911);
and (n960,n309,n49);
and (n961,n962,n963);
xor (n962,n959,n960);
and (n963,n964,n618);
xor (n964,n916,n917);
and (n965,n69,n59);
or (n966,n967,n970);
and (n967,n968,n969);
xor (n968,n926,n927);
and (n969,n322,n59);
and (n970,n971,n972);
xor (n971,n968,n969);
or (n972,n973,n976);
and (n973,n974,n975);
xor (n974,n932,n933);
and (n975,n235,n59);
and (n976,n977,n978);
xor (n977,n974,n975);
or (n978,n979,n982);
and (n979,n980,n981);
xor (n980,n938,n939);
and (n981,n227,n59);
and (n982,n983,n984);
xor (n983,n980,n981);
or (n984,n985,n988);
and (n985,n986,n987);
xor (n986,n944,n945);
and (n987,n264,n59);
and (n988,n989,n990);
xor (n989,n986,n987);
or (n990,n991,n994);
and (n991,n992,n993);
xor (n992,n950,n951);
and (n993,n256,n59);
and (n994,n995,n996);
xor (n995,n992,n993);
or (n996,n997,n1000);
and (n997,n998,n999);
xor (n998,n956,n957);
and (n999,n309,n59);
and (n1000,n1001,n1002);
xor (n1001,n998,n999);
and (n1002,n1003,n1004);
xor (n1003,n962,n963);
and (n1004,n164,n59);
and (n1005,n322,n213);
or (n1006,n1007,n1010);
and (n1007,n1008,n1009);
xor (n1008,n971,n972);
and (n1009,n235,n213);
and (n1010,n1011,n1012);
xor (n1011,n1008,n1009);
or (n1012,n1013,n1016);
and (n1013,n1014,n1015);
xor (n1014,n977,n978);
and (n1015,n227,n213);
and (n1016,n1017,n1018);
xor (n1017,n1014,n1015);
or (n1018,n1019,n1022);
and (n1019,n1020,n1021);
xor (n1020,n983,n984);
and (n1021,n264,n213);
and (n1022,n1023,n1024);
xor (n1023,n1020,n1021);
or (n1024,n1025,n1028);
and (n1025,n1026,n1027);
xor (n1026,n989,n990);
and (n1027,n256,n213);
and (n1028,n1029,n1030);
xor (n1029,n1026,n1027);
or (n1030,n1031,n1034);
and (n1031,n1032,n1033);
xor (n1032,n995,n996);
and (n1033,n309,n213);
and (n1034,n1035,n1036);
xor (n1035,n1032,n1033);
and (n1036,n1037,n517);
xor (n1037,n1001,n1002);
and (n1038,n235,n220);
or (n1039,n1040,n1043);
and (n1040,n1041,n1042);
xor (n1041,n1011,n1012);
and (n1042,n227,n220);
and (n1043,n1044,n1045);
xor (n1044,n1041,n1042);
or (n1045,n1046,n1048);
and (n1046,n1047,n301);
xor (n1047,n1017,n1018);
and (n1048,n1049,n1050);
xor (n1049,n1047,n301);
or (n1050,n1051,n1054);
and (n1051,n1052,n1053);
xor (n1052,n1023,n1024);
and (n1053,n256,n220);
and (n1054,n1055,n1056);
xor (n1055,n1052,n1053);
or (n1056,n1057,n1060);
and (n1057,n1058,n1059);
xor (n1058,n1029,n1030);
and (n1059,n309,n220);
and (n1060,n1061,n1062);
xor (n1061,n1058,n1059);
and (n1062,n1063,n1064);
xor (n1063,n1035,n1036);
and (n1064,n164,n220);
and (n1065,n227,n245);
or (n1066,n1067,n1070);
and (n1067,n1068,n1069);
xor (n1068,n1044,n1045);
and (n1069,n264,n245);
and (n1070,n1071,n1072);
xor (n1071,n1068,n1069);
or (n1072,n1073,n1076);
and (n1073,n1074,n1075);
xor (n1074,n1049,n1050);
and (n1075,n256,n245);
and (n1076,n1077,n1078);
xor (n1077,n1074,n1075);
or (n1078,n1079,n1082);
and (n1079,n1080,n1081);
xor (n1080,n1055,n1056);
and (n1081,n309,n245);
and (n1082,n1083,n1084);
xor (n1083,n1080,n1081);
and (n1084,n1085,n419);
xor (n1085,n1061,n1062);
and (n1086,n264,n147);
or (n1087,n1088,n1091);
and (n1088,n1089,n1090);
xor (n1089,n1071,n1072);
and (n1090,n256,n147);
and (n1091,n1092,n1093);
xor (n1092,n1089,n1090);
or (n1093,n1094,n1097);
and (n1094,n1095,n1096);
xor (n1095,n1077,n1078);
and (n1096,n309,n147);
and (n1097,n1098,n1099);
xor (n1098,n1095,n1096);
and (n1099,n1100,n1101);
xor (n1100,n1083,n1084);
and (n1101,n164,n147);
and (n1102,n256,n165);
or (n1103,n1104,n1107);
and (n1104,n1105,n1106);
xor (n1105,n1092,n1093);
and (n1106,n309,n165);
and (n1107,n1108,n1109);
xor (n1108,n1105,n1106);
and (n1109,n1110,n163);
xor (n1110,n1098,n1099);
and (n1111,n309,n175);
and (n1112,n1113,n1114);
xor (n1113,n1108,n1109);
and (n1114,n164,n175);
and (n1115,n164,n356);
endmodule
