module top (out,n12,n14,n15,n17,n20,n24,n26,n28,n31
        ,n39,n41,n42,n46,n51,n53,n56,n61,n63,n64
        ,n66,n69,n74,n81,n83,n89,n95,n97,n100,n112
        ,n117,n119,n158,n160,n162,n203,n277,n299,n300,n455
        ,n540,n557,n558,n653,n657,n659,n670,n682,n696);
output out;
input n12;
input n14;
input n15;
input n17;
input n20;
input n24;
input n26;
input n28;
input n31;
input n39;
input n41;
input n42;
input n46;
input n51;
input n53;
input n56;
input n61;
input n63;
input n64;
input n66;
input n69;
input n74;
input n81;
input n83;
input n89;
input n95;
input n97;
input n100;
input n112;
input n117;
input n119;
input n158;
input n160;
input n162;
input n203;
input n277;
input n299;
input n300;
input n455;
input n540;
input n557;
input n558;
input n653;
input n657;
input n659;
input n670;
input n682;
input n696;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n13;
wire n16;
wire n18;
wire n19;
wire n21;
wire n22;
wire n23;
wire n25;
wire n27;
wire n29;
wire n30;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n40;
wire n43;
wire n44;
wire n45;
wire n47;
wire n48;
wire n49;
wire n50;
wire n52;
wire n54;
wire n55;
wire n57;
wire n58;
wire n59;
wire n60;
wire n62;
wire n65;
wire n67;
wire n68;
wire n70;
wire n71;
wire n72;
wire n73;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n82;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n96;
wire n98;
wire n99;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n113;
wire n114;
wire n115;
wire n116;
wire n118;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n159;
wire n161;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n654;
wire n655;
wire n656;
wire n658;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2988;
wire n2989;
wire n2990;
wire n2991;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2996;
wire n2997;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3003;
wire n3004;
wire n3005;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3010;
wire n3011;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3038;
wire n3039;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
wire n3056;
wire n3057;
wire n3058;
wire n3059;
wire n3060;
wire n3061;
wire n3062;
wire n3063;
wire n3064;
wire n3065;
wire n3066;
wire n3067;
wire n3068;
wire n3069;
wire n3070;
wire n3071;
wire n3072;
wire n3073;
wire n3074;
wire n3075;
wire n3076;
wire n3077;
wire n3078;
wire n3079;
wire n3080;
wire n3081;
wire n3082;
wire n3083;
wire n3084;
wire n3085;
wire n3086;
wire n3087;
wire n3088;
wire n3089;
wire n3090;
wire n3091;
wire n3092;
wire n3093;
wire n3094;
wire n3095;
wire n3096;
wire n3097;
wire n3098;
wire n3099;
wire n3100;
wire n3101;
wire n3102;
wire n3103;
wire n3104;
wire n3105;
wire n3106;
wire n3107;
wire n3108;
wire n3109;
wire n3110;
wire n3111;
wire n3112;
wire n3113;
wire n3114;
wire n3115;
wire n3116;
wire n3117;
wire n3118;
wire n3119;
wire n3120;
wire n3121;
wire n3122;
wire n3123;
wire n3124;
wire n3125;
wire n3126;
wire n3127;
wire n3128;
wire n3129;
wire n3130;
wire n3131;
wire n3132;
wire n3133;
wire n3134;
wire n3135;
wire n3136;
wire n3137;
wire n3138;
wire n3139;
wire n3140;
wire n3141;
wire n3142;
wire n3143;
wire n3144;
wire n3145;
wire n3146;
wire n3147;
wire n3148;
wire n3149;
wire n3150;
wire n3151;
wire n3152;
wire n3153;
wire n3154;
wire n3155;
wire n3156;
wire n3157;
wire n3158;
wire n3159;
wire n3160;
wire n3161;
wire n3162;
xor (out,n0,n2665);
xnor (n0,n1,n2594);
nand (n1,n2,n390);
nand (n2,n3,n322);
nand (n3,n4,n266,n321);
nand (n4,n5,n145);
xor (n5,n6,n125);
xor (n6,n7,n72);
nand (n7,n8,n32,n71);
nand (n8,n9,n21);
xor (n9,n10,n20);
or (n10,n11,n16);
and (n11,n12,n13);
xor (n13,n14,n15);
and (n16,n17,n18);
nor (n18,n13,n19);
xnor (n19,n20,n14);
xor (n21,n22,n31);
or (n22,n23,n27);
and (n23,n24,n25);
xor (n25,n26,n20);
and (n27,n28,n29);
nor (n29,n25,n30);
xnor (n30,n31,n26);
nand (n32,n33,n21);
nand (n33,n34,n57,n70);
nand (n34,n35,n47);
not (n35,n36);
xor (n36,n37,n46);
or (n37,n38,n43);
and (n38,n39,n40);
xor (n40,n41,n42);
and (n43,n39,n44);
nor (n44,n40,n45);
xnor (n45,n46,n41);
xor (n47,n48,n56);
or (n48,n49,n52);
and (n49,n39,n50);
xor (n50,n51,n46);
and (n52,n53,n54);
nor (n54,n50,n55);
xnor (n55,n56,n51);
nand (n57,n58,n47);
xor (n58,n59,n69);
or (n59,n60,n65);
and (n60,n61,n62);
xor (n62,n63,n64);
and (n65,n66,n67);
nor (n67,n62,n68);
xnor (n68,n69,n63);
nand (n70,n35,n58);
nand (n71,n9,n33);
nand (n72,n73,n101,n124);
nand (n73,n74,n75);
xor (n75,n76,n91);
xor (n76,n77,n86);
xor (n77,n78,n64);
or (n78,n79,n82);
and (n79,n53,n80);
xor (n80,n81,n56);
and (n82,n83,n84);
nor (n84,n80,n85);
xnor (n85,n64,n81);
xor (n86,n87,n69);
or (n87,n88,n90);
and (n88,n89,n62);
and (n90,n61,n67);
xor (n91,n92,n100);
or (n92,n93,n96);
and (n93,n66,n94);
xor (n94,n95,n69);
and (n96,n97,n98);
nor (n98,n94,n99);
xnor (n99,n100,n95);
nand (n101,n102,n75);
nand (n102,n103,n113,n123);
nand (n103,n104,n108);
xor (n104,n105,n64);
or (n105,n106,n107);
and (n106,n83,n80);
and (n107,n89,n84);
xor (n108,n109,n100);
or (n109,n110,n111);
and (n110,n97,n94);
and (n111,n112,n98);
nand (n113,n114,n108);
xor (n114,n115,n15);
or (n115,n116,n120);
and (n116,n117,n118);
xor (n118,n119,n100);
and (n120,n12,n121);
nor (n121,n118,n122);
xnor (n122,n15,n119);
nand (n123,n104,n114);
nand (n124,n74,n102);
xor (n125,n126,n141);
xor (n126,n74,n127);
xor (n127,n128,n137);
xor (n128,n129,n133);
not (n129,n130);
xor (n130,n131,n56);
or (n131,n49,n132);
and (n132,n39,n54);
xor (n133,n134,n64);
or (n134,n135,n136);
and (n135,n39,n80);
and (n136,n53,n84);
xor (n137,n138,n69);
or (n138,n139,n140);
and (n139,n83,n62);
and (n140,n89,n67);
nand (n141,n142,n143,n144);
nand (n142,n77,n86);
nand (n143,n91,n86);
nand (n144,n77,n91);
xor (n145,n146,n212);
xor (n146,n147,n191);
xor (n147,n148,n181);
xor (n148,n149,n167);
nand (n149,n150,n165,n166);
nand (n150,n151,n155);
xor (n151,n152,n15);
or (n152,n153,n154);
and (n153,n112,n118);
and (n154,n117,n121);
xor (n155,n156,n74);
or (n156,n157,n161);
and (n157,n158,n159);
xor (n159,n160,n31);
and (n161,n162,n163);
nor (n163,n159,n164);
xnor (n164,n74,n160);
nand (n165,n129,n155);
nand (n166,n151,n129);
xor (n167,n168,n177);
xor (n168,n169,n173);
xor (n169,n170,n100);
or (n170,n171,n172);
and (n171,n61,n94);
and (n172,n66,n98);
xor (n173,n174,n15);
or (n174,n175,n176);
and (n175,n97,n118);
and (n176,n112,n121);
xor (n177,n178,n74);
or (n178,n179,n180);
and (n179,n28,n159);
and (n180,n158,n163);
xor (n181,n182,n187);
xor (n182,n130,n183);
xor (n183,n184,n20);
or (n184,n185,n186);
and (n185,n117,n13);
and (n186,n12,n18);
xor (n187,n188,n31);
or (n188,n189,n190);
and (n189,n17,n25);
and (n190,n24,n29);
nand (n191,n192,n208,n211);
nand (n192,n193,n206);
nand (n193,n194,n204,n205);
nand (n194,n195,n199);
xor (n195,n196,n31);
or (n196,n197,n198);
and (n197,n28,n25);
and (n198,n158,n29);
xor (n199,n200,n74);
or (n200,n201,n202);
and (n201,n162,n159);
and (n202,n203,n163);
nand (n204,n36,n199);
nand (n205,n195,n36);
xor (n206,n207,n33);
xor (n207,n9,n21);
nand (n208,n209,n206);
xor (n209,n210,n129);
xor (n210,n151,n155);
nand (n211,n193,n209);
nand (n212,n213,n240,n265);
nand (n213,n214,n238);
nand (n214,n215,n220,n237);
nand (n215,n216,n74);
xor (n216,n217,n20);
or (n217,n218,n219);
and (n218,n17,n13);
and (n219,n24,n18);
nand (n220,n221,n74);
nand (n221,n222,n231,n236);
nand (n222,n223,n227);
xor (n223,n224,n69);
or (n224,n225,n226);
and (n225,n66,n62);
and (n226,n97,n67);
xor (n227,n228,n56);
or (n228,n229,n230);
and (n229,n53,n50);
and (n230,n83,n54);
nand (n231,n232,n227);
xor (n232,n233,n64);
or (n233,n234,n235);
and (n234,n89,n80);
and (n235,n61,n84);
nand (n236,n223,n232);
nand (n237,n216,n221);
xor (n238,n239,n102);
xor (n239,n74,n75);
nand (n240,n241,n238);
nand (n241,n242,n247,n264);
nand (n242,n243,n245);
xor (n243,n244,n58);
xor (n244,n35,n47);
xor (n245,n246,n114);
xor (n246,n104,n108);
nand (n247,n248,n245);
nand (n248,n249,n258,n263);
nand (n249,n250,n254);
xor (n250,n251,n100);
or (n251,n252,n253);
and (n252,n112,n94);
and (n253,n117,n98);
xor (n254,n255,n15);
or (n255,n256,n257);
and (n256,n12,n118);
and (n257,n17,n121);
nand (n258,n259,n254);
xor (n259,n260,n31);
or (n260,n261,n262);
and (n261,n158,n25);
and (n262,n162,n29);
nand (n263,n250,n259);
nand (n264,n243,n248);
nand (n265,n214,n241);
nand (n266,n267,n145);
nand (n267,n268,n317,n320);
nand (n268,n269,n315);
nand (n269,n270,n286,n314);
nand (n270,n271,n284);
nand (n271,n272,n278,n283);
nand (n272,n273,n35);
xor (n273,n274,n74);
or (n274,n275,n276);
and (n275,n203,n159);
and (n276,n277,n163);
nand (n278,n279,n35);
xor (n279,n280,n20);
or (n280,n281,n282);
and (n281,n24,n13);
and (n282,n28,n18);
nand (n283,n273,n279);
xor (n284,n285,n36);
xor (n285,n195,n199);
nand (n286,n287,n284);
nand (n287,n288,n310,n313);
nand (n288,n74,n289);
nand (n289,n290,n304,n309);
nand (n290,n291,n294);
xor (n291,n292,n46);
or (n292,n38,n293);
and (n293,n53,n44);
not (n294,n295);
xor (n295,n296,n42);
or (n296,n297,n301);
and (n297,n39,n298);
xor (n298,n299,n300);
and (n301,n39,n302);
nor (n302,n298,n303);
xnor (n303,n42,n299);
nand (n304,n305,n294);
xor (n305,n306,n64);
or (n306,n307,n308);
and (n307,n61,n80);
and (n308,n66,n84);
nand (n309,n291,n305);
nand (n310,n311,n289);
xor (n311,n312,n232);
xor (n312,n223,n227);
nand (n313,n74,n311);
nand (n314,n271,n287);
xor (n315,n316,n209);
xor (n316,n193,n206);
nand (n317,n318,n315);
xor (n318,n319,n241);
xor (n319,n214,n238);
nand (n320,n269,n318);
nand (n321,n5,n267);
xor (n322,n323,n386);
xor (n323,n324,n352);
xor (n324,n325,n348);
xor (n325,n326,n340);
xor (n326,n327,n336);
xor (n327,n328,n332);
not (n328,n329);
xor (n329,n330,n64);
or (n330,n135,n331);
and (n331,n39,n84);
xor (n332,n333,n20);
or (n333,n334,n335);
and (n334,n112,n13);
and (n335,n117,n18);
xor (n336,n337,n31);
or (n337,n338,n339);
and (n338,n12,n25);
and (n339,n17,n29);
xor (n340,n341,n344);
or (n341,n342,n343);
and (n342,n24,n159);
and (n343,n28,n163);
nand (n344,n345,n346,n347);
nand (n345,n129,n133);
nand (n346,n137,n133);
nand (n347,n129,n137);
nand (n348,n349,n350,n351);
nand (n349,n74,n127);
nand (n350,n141,n127);
nand (n351,n74,n141);
xor (n352,n353,n382);
xor (n353,n354,n378);
xor (n354,n355,n374);
xor (n355,n356,n370);
xor (n356,n357,n366);
xor (n357,n358,n362);
xor (n358,n359,n69);
or (n359,n360,n361);
and (n360,n53,n62);
and (n361,n83,n67);
xor (n362,n363,n15);
or (n363,n364,n365);
and (n364,n66,n118);
and (n365,n97,n121);
xor (n366,n367,n100);
or (n367,n368,n369);
and (n368,n89,n94);
and (n369,n61,n98);
nand (n370,n371,n372,n373);
nand (n371,n169,n173);
nand (n372,n177,n173);
nand (n373,n169,n177);
nand (n374,n375,n376,n377);
nand (n375,n130,n183);
nand (n376,n187,n183);
nand (n377,n130,n187);
nand (n378,n379,n380,n381);
nand (n379,n149,n167);
nand (n380,n181,n167);
nand (n381,n149,n181);
nand (n382,n383,n384,n385);
nand (n383,n7,n72);
nand (n384,n125,n72);
nand (n385,n7,n125);
nand (n386,n387,n388,n389);
nand (n387,n147,n191);
nand (n388,n212,n191);
nand (n389,n147,n212);
nand (n390,n391,n2592);
nand (n391,n392,n632);
nor (n392,n393,n630);
nor (n393,n394,n623);
nand (n394,n395,n611);
nand (n395,n396,n527,n610);
nand (n396,n397,n441);
xor (n397,n398,n439);
xor (n398,n399,n401);
xor (n399,n400,n221);
xor (n400,n216,n74);
nand (n401,n402,n421,n438);
nand (n402,n403,n419);
nand (n403,n404,n413,n418);
nand (n404,n405,n409);
xor (n405,n406,n69);
or (n406,n407,n408);
and (n407,n97,n62);
and (n408,n112,n67);
xor (n409,n410,n56);
or (n410,n411,n412);
and (n411,n83,n50);
and (n412,n89,n54);
nand (n413,n414,n409);
xor (n414,n415,n100);
or (n415,n416,n417);
and (n416,n117,n94);
and (n417,n12,n98);
nand (n418,n405,n414);
xor (n419,n420,n259);
xor (n420,n250,n254);
nand (n421,n422,n419);
nand (n422,n423,n432,n437);
nand (n423,n424,n428);
xor (n424,n425,n46);
or (n425,n426,n427);
and (n426,n53,n40);
and (n427,n83,n44);
xor (n428,n429,n15);
or (n429,n430,n431);
and (n430,n17,n118);
and (n431,n24,n121);
nand (n432,n433,n428);
xor (n433,n434,n20);
or (n434,n435,n436);
and (n435,n28,n13);
and (n436,n158,n18);
nand (n437,n424,n433);
nand (n438,n403,n422);
xor (n439,n440,n248);
xor (n440,n243,n245);
xor (n441,n442,n466);
xor (n442,n443,n464);
nand (n443,n444,n460,n463);
nand (n444,n445,n458);
nand (n445,n446,n456,n457);
nand (n446,n447,n451);
xor (n447,n448,n31);
or (n448,n449,n450);
and (n449,n162,n25);
and (n450,n203,n29);
xor (n451,n452,n74);
or (n452,n453,n454);
and (n453,n277,n159);
and (n454,n455,n163);
nand (n456,n74,n451);
nand (n457,n447,n74);
xor (n458,n459,n279);
xor (n459,n273,n35);
nand (n460,n461,n458);
xor (n461,n462,n311);
xor (n462,n74,n289);
nand (n463,n445,n461);
xor (n464,n465,n287);
xor (n465,n271,n284);
nand (n466,n467,n523,n526);
nand (n467,n468,n488);
nand (n468,n469,n484,n487);
nand (n469,n470,n482);
nand (n470,n471,n476,n481);
nand (n471,n295,n472);
xor (n472,n473,n64);
or (n473,n474,n475);
and (n474,n66,n80);
and (n475,n97,n84);
nand (n476,n477,n472);
xor (n477,n478,n69);
or (n478,n479,n480);
and (n479,n112,n62);
and (n480,n117,n67);
nand (n481,n295,n477);
xor (n482,n483,n414);
xor (n483,n405,n409);
nand (n484,n485,n482);
xor (n485,n486,n305);
xor (n486,n291,n294);
nand (n487,n470,n485);
nand (n488,n489,n519,n522);
nand (n489,n490,n503);
nand (n490,n491,n497,n502);
nand (n491,n492,n496);
xor (n492,n493,n56);
or (n493,n494,n495);
and (n494,n89,n50);
and (n495,n61,n54);
not (n496,n424);
nand (n497,n498,n496);
xor (n498,n499,n100);
or (n499,n500,n501);
and (n500,n12,n94);
and (n501,n17,n98);
nand (n502,n492,n498);
nand (n503,n504,n513,n518);
nand (n504,n505,n509);
xor (n505,n506,n15);
or (n506,n507,n508);
and (n507,n24,n118);
and (n508,n28,n121);
xor (n509,n510,n20);
or (n510,n511,n512);
and (n511,n158,n13);
and (n512,n162,n18);
nand (n513,n514,n509);
xor (n514,n515,n31);
or (n515,n516,n517);
and (n516,n203,n25);
and (n517,n277,n29);
nand (n518,n505,n514);
nand (n519,n520,n503);
xor (n520,n521,n433);
xor (n521,n424,n428);
nand (n522,n490,n520);
nand (n523,n524,n488);
xor (n524,n525,n422);
xor (n525,n403,n419);
nand (n526,n468,n524);
nand (n527,n528,n441);
nand (n528,n529,n606,n609);
nand (n529,n530,n532);
xor (n530,n531,n461);
xor (n531,n445,n458);
nand (n532,n533,n566,n605);
nand (n533,n534,n564);
nand (n534,n535,n541,n563);
nand (n535,n536,n74);
xor (n536,n537,n74);
or (n537,n538,n539);
and (n538,n455,n159);
and (n539,n540,n163);
nand (n541,n542,n74);
nand (n542,n543,n551,n562);
nand (n543,n544,n547);
xor (n544,n545,n42);
or (n545,n297,n546);
and (n546,n53,n302);
xor (n547,n548,n46);
or (n548,n549,n550);
and (n549,n83,n40);
and (n550,n89,n44);
nand (n551,n552,n547);
not (n552,n553);
xor (n553,n554,n300);
or (n554,n555,n559);
and (n555,n39,n556);
xor (n556,n557,n558);
and (n559,n39,n560);
nor (n560,n556,n561);
xnor (n561,n300,n557);
nand (n562,n544,n552);
nand (n563,n536,n542);
xor (n564,n565,n74);
xor (n565,n447,n451);
nand (n566,n567,n564);
nand (n567,n568,n587,n604);
nand (n568,n569,n585);
nand (n569,n570,n579,n584);
nand (n570,n571,n575);
xor (n571,n572,n56);
or (n572,n573,n574);
and (n573,n61,n50);
and (n574,n66,n54);
xor (n575,n576,n64);
or (n576,n577,n578);
and (n577,n97,n80);
and (n578,n112,n84);
nand (n579,n580,n575);
xor (n580,n581,n69);
or (n581,n582,n583);
and (n582,n117,n62);
and (n583,n12,n67);
nand (n584,n571,n580);
xor (n585,n586,n477);
xor (n586,n295,n472);
nand (n587,n588,n585);
nand (n588,n589,n598,n603);
nand (n589,n590,n594);
xor (n590,n591,n15);
or (n591,n592,n593);
and (n592,n28,n118);
and (n593,n158,n121);
xor (n594,n595,n42);
or (n595,n596,n597);
and (n596,n53,n298);
and (n597,n83,n302);
nand (n598,n599,n594);
xor (n599,n600,n100);
or (n600,n601,n602);
and (n601,n17,n94);
and (n602,n24,n98);
nand (n603,n590,n599);
nand (n604,n569,n588);
nand (n605,n534,n567);
nand (n606,n607,n532);
xor (n607,n608,n524);
xor (n608,n468,n488);
nand (n609,n530,n607);
nand (n610,n397,n528);
xor (n611,n612,n619);
xor (n612,n613,n617);
nand (n613,n614,n615,n616);
nand (n614,n399,n401);
nand (n615,n439,n401);
nand (n616,n399,n439);
xor (n617,n618,n318);
xor (n618,n269,n315);
nand (n619,n620,n621,n622);
nand (n620,n443,n464);
nand (n621,n466,n464);
nand (n622,n443,n466);
nor (n623,n624,n628);
nand (n624,n625,n626,n627);
nand (n625,n613,n617);
nand (n626,n619,n617);
nand (n627,n613,n619);
xor (n628,n629,n267);
xor (n629,n5,n145);
not (n630,n631);
nand (n631,n624,n628);
nand (n632,n633,n635);
nor (n633,n634,n623);
nor (n634,n395,n611);
nand (n635,n636,n2166);
nor (n636,n637,n2134);
nor (n637,n638,n1607);
nor (n638,n639,n1592);
nor (n639,n640,n1313);
nand (n640,n641,n1096);
nor (n641,n642,n995);
nor (n642,n643,n905);
nand (n643,n644,n820,n904);
nand (n644,n645,n722);
xor (n645,n646,n698);
xor (n646,n647,n672);
xor (n647,n648,n660);
xor (n648,n649,n654);
xor (n649,n650,n100);
or (n650,n651,n652);
and (n651,n540,n94);
and (n652,n653,n98);
xor (n654,n655,n15);
or (n655,n656,n658);
and (n656,n657,n118);
and (n658,n659,n121);
xor (n660,n661,n665);
xor (n661,n662,n300);
or (n662,n663,n664);
and (n663,n97,n556);
and (n664,n112,n560);
xnor (n665,n666,n558);
nor (n666,n667,n671);
and (n667,n66,n668);
and (n668,n669,n558);
not (n669,n670);
and (n671,n61,n670);
nand (n672,n673,n683,n697);
nand (n673,n674,n678);
xor (n674,n675,n100);
or (n675,n676,n677);
and (n676,n653,n94);
and (n677,n657,n98);
xor (n678,n679,n15);
or (n679,n680,n681);
and (n680,n659,n118);
and (n681,n682,n121);
nand (n683,n684,n678);
xor (n684,n685,n694);
xor (n685,n686,n690);
xor (n686,n687,n300);
or (n687,n688,n689);
and (n688,n112,n556);
and (n689,n117,n560);
xor (n690,n691,n46);
or (n691,n692,n693);
and (n692,n24,n40);
and (n693,n28,n44);
xnor (n694,n695,n20);
nand (n695,n696,n13);
nand (n697,n674,n684);
xor (n698,n699,n708);
xor (n699,n700,n704);
xor (n700,n701,n20);
or (n701,n702,n703);
and (n702,n682,n13);
and (n703,n696,n18);
nand (n704,n705,n706,n707);
nand (n705,n686,n690);
nand (n706,n694,n690);
nand (n707,n686,n694);
xor (n708,n709,n718);
xor (n709,n710,n714);
xor (n710,n711,n46);
or (n711,n712,n713);
and (n712,n17,n40);
and (n713,n24,n44);
xor (n714,n715,n42);
or (n715,n716,n717);
and (n716,n117,n298);
and (n717,n12,n302);
xor (n718,n719,n56);
or (n719,n720,n721);
and (n720,n28,n50);
and (n721,n158,n54);
nand (n722,n723,n777,n819);
nand (n723,n724,n726);
xor (n724,n725,n684);
xor (n725,n674,n678);
xor (n726,n727,n766);
xor (n727,n728,n744);
nand (n728,n729,n738,n743);
nand (n729,n730,n734);
xor (n730,n731,n46);
or (n731,n732,n733);
and (n732,n28,n40);
and (n733,n158,n44);
xor (n734,n735,n42);
or (n735,n736,n737);
and (n736,n17,n298);
and (n737,n24,n302);
nand (n738,n739,n734);
xor (n739,n740,n56);
or (n740,n741,n742);
and (n741,n162,n50);
and (n742,n203,n54);
nand (n743,n730,n739);
nand (n744,n745,n760,n765);
nand (n745,n746,n755);
xor (n746,n747,n751);
xnor (n747,n748,n558);
nor (n748,n749,n750);
and (n749,n112,n668);
and (n750,n97,n670);
xor (n751,n752,n300);
or (n752,n753,n754);
and (n753,n117,n556);
and (n754,n12,n560);
and (n755,n756,n15);
xnor (n756,n757,n558);
nor (n757,n758,n759);
and (n758,n117,n668);
and (n759,n112,n670);
nand (n760,n761,n755);
xor (n761,n762,n64);
or (n762,n763,n764);
and (n763,n277,n80);
and (n764,n455,n84);
nand (n765,n746,n761);
xor (n766,n767,n773);
xor (n767,n768,n772);
xor (n768,n769,n64);
or (n769,n770,n771);
and (n770,n203,n80);
and (n771,n277,n84);
and (n772,n747,n751);
xor (n773,n774,n69);
or (n774,n775,n776);
and (n775,n455,n62);
and (n776,n540,n67);
nand (n777,n778,n726);
nand (n778,n779,n803,n818);
nand (n779,n780,n801);
nand (n780,n781,n795,n800);
nand (n781,n782,n791);
and (n782,n783,n787);
xnor (n783,n784,n558);
nor (n784,n785,n786);
and (n785,n12,n668);
and (n786,n117,n670);
xor (n787,n788,n300);
or (n788,n789,n790);
and (n789,n17,n556);
and (n790,n24,n560);
xor (n791,n792,n64);
or (n792,n793,n794);
and (n793,n455,n80);
and (n794,n540,n84);
nand (n795,n796,n791);
xor (n796,n797,n69);
or (n797,n798,n799);
and (n798,n653,n62);
and (n799,n657,n67);
nand (n800,n782,n796);
xor (n801,n802,n761);
xor (n802,n746,n755);
nand (n803,n804,n801);
xor (n804,n805,n814);
xor (n805,n806,n810);
xor (n806,n807,n69);
or (n807,n808,n809);
and (n808,n540,n62);
and (n809,n653,n67);
xor (n810,n811,n100);
or (n811,n812,n813);
and (n812,n657,n94);
and (n813,n659,n98);
xor (n814,n815,n15);
or (n815,n816,n817);
and (n816,n682,n118);
and (n817,n696,n121);
nand (n818,n780,n804);
nand (n819,n724,n778);
nand (n820,n821,n722);
xor (n821,n822,n861);
xor (n822,n823,n827);
nand (n823,n824,n825,n826);
nand (n824,n728,n744);
nand (n825,n766,n744);
nand (n826,n728,n766);
xor (n827,n828,n850);
xor (n828,n829,n846);
nand (n829,n830,n840,n845);
nand (n830,n831,n835);
xor (n831,n832,n42);
or (n832,n833,n834);
and (n833,n12,n298);
and (n834,n17,n302);
xor (n835,n836,n20);
xnor (n836,n837,n558);
nor (n837,n838,n839);
and (n838,n97,n668);
and (n839,n66,n670);
nand (n840,n841,n835);
xor (n841,n842,n56);
or (n842,n843,n844);
and (n843,n158,n50);
and (n844,n162,n54);
nand (n845,n831,n841);
nand (n846,n847,n848,n849);
nand (n847,n768,n772);
nand (n848,n773,n772);
nand (n849,n768,n773);
xor (n850,n851,n857);
xor (n851,n852,n853);
and (n852,n836,n20);
xor (n853,n854,n64);
or (n854,n855,n856);
and (n855,n162,n80);
and (n856,n203,n84);
xor (n857,n858,n69);
or (n858,n859,n860);
and (n859,n277,n62);
and (n860,n455,n67);
nand (n861,n862,n869,n903);
nand (n862,n863,n867);
nand (n863,n864,n865,n866);
nand (n864,n806,n810);
nand (n865,n814,n810);
nand (n866,n806,n814);
xor (n867,n868,n841);
xor (n868,n831,n835);
nand (n869,n870,n867);
nand (n870,n871,n888,n902);
nand (n871,n872,n886);
nand (n872,n873,n882,n885);
nand (n873,n874,n878);
xor (n874,n875,n300);
or (n875,n876,n877);
and (n876,n12,n556);
and (n877,n17,n560);
xor (n878,n879,n46);
or (n879,n880,n881);
and (n880,n158,n40);
and (n881,n162,n44);
nand (n882,n883,n878);
xnor (n883,n884,n15);
nand (n884,n696,n118);
nand (n885,n874,n883);
xor (n886,n887,n739);
xor (n887,n730,n734);
nand (n888,n889,n886);
nand (n889,n890,n896,n901);
nand (n890,n891,n895);
xor (n891,n892,n42);
or (n892,n893,n894);
and (n893,n24,n298);
and (n894,n28,n302);
xor (n895,n756,n15);
nand (n896,n897,n895);
xor (n897,n898,n56);
or (n898,n899,n900);
and (n899,n203,n50);
and (n900,n277,n54);
nand (n901,n891,n897);
nand (n902,n872,n889);
nand (n903,n863,n870);
nand (n904,n645,n821);
xor (n905,n906,n991);
xor (n906,n907,n928);
xor (n907,n908,n924);
xor (n908,n909,n920);
xor (n909,n910,n916);
xor (n910,n911,n915);
xor (n911,n912,n15);
or (n912,n913,n914);
and (n913,n653,n118);
and (n914,n657,n121);
and (n915,n661,n665);
xor (n916,n917,n20);
or (n917,n918,n919);
and (n918,n659,n13);
and (n919,n682,n18);
nand (n920,n921,n922,n923);
nand (n921,n700,n704);
nand (n922,n708,n704);
nand (n923,n700,n708);
nand (n924,n925,n926,n927);
nand (n925,n829,n846);
nand (n926,n850,n846);
nand (n927,n829,n850);
xor (n928,n929,n987);
xor (n929,n930,n954);
xor (n930,n931,n950);
xor (n931,n932,n936);
nand (n932,n933,n934,n935);
nand (n933,n852,n853);
nand (n934,n857,n853);
nand (n935,n852,n857);
xor (n936,n937,n946);
xor (n937,n938,n942);
xnor (n938,n939,n558);
nor (n939,n940,n941);
and (n940,n61,n668);
and (n941,n89,n670);
xor (n942,n943,n46);
or (n943,n944,n945);
and (n944,n12,n40);
and (n945,n17,n44);
xor (n946,n947,n42);
or (n947,n948,n949);
and (n948,n112,n298);
and (n949,n117,n302);
nand (n950,n951,n952,n953);
nand (n951,n710,n714);
nand (n952,n718,n714);
nand (n953,n710,n718);
xor (n954,n955,n973);
xor (n955,n956,n960);
nand (n956,n957,n958,n959);
nand (n957,n649,n654);
nand (n958,n660,n654);
nand (n959,n649,n660);
xor (n960,n961,n971);
xor (n961,n962,n966);
xor (n962,n963,n56);
or (n963,n964,n965);
and (n964,n24,n50);
and (n965,n28,n54);
xor (n966,n31,n967);
xor (n967,n968,n300);
or (n968,n969,n970);
and (n969,n66,n556);
and (n970,n97,n560);
xnor (n971,n972,n31);
nand (n972,n696,n25);
xor (n973,n974,n983);
xor (n974,n975,n979);
xor (n975,n976,n64);
or (n976,n977,n978);
and (n977,n158,n80);
and (n978,n162,n84);
xor (n979,n980,n69);
or (n980,n981,n982);
and (n981,n203,n62);
and (n982,n277,n67);
xor (n983,n984,n100);
or (n984,n985,n986);
and (n985,n455,n94);
and (n986,n540,n98);
nand (n987,n988,n989,n990);
nand (n988,n647,n672);
nand (n989,n698,n672);
nand (n990,n647,n698);
nand (n991,n992,n993,n994);
nand (n992,n823,n827);
nand (n993,n861,n827);
nand (n994,n823,n861);
nor (n995,n996,n1000);
nand (n996,n997,n998,n999);
nand (n997,n907,n928);
nand (n998,n991,n928);
nand (n999,n907,n991);
xor (n1000,n1001,n1010);
xor (n1001,n1002,n1006);
nand (n1002,n1003,n1004,n1005);
nand (n1003,n909,n920);
nand (n1004,n924,n920);
nand (n1005,n909,n924);
nand (n1006,n1007,n1008,n1009);
nand (n1007,n930,n954);
nand (n1008,n987,n954);
nand (n1009,n930,n987);
xor (n1010,n1011,n1072);
xor (n1011,n1012,n1043);
xor (n1012,n1013,n1032);
xor (n1013,n1014,n1028);
xor (n1014,n1015,n1024);
xor (n1015,n1016,n1020);
xor (n1016,n1017,n46);
or (n1017,n1018,n1019);
and (n1018,n117,n40);
and (n1019,n12,n44);
xor (n1020,n1021,n42);
or (n1021,n1022,n1023);
and (n1022,n97,n298);
and (n1023,n112,n302);
xor (n1024,n1025,n56);
or (n1025,n1026,n1027);
and (n1026,n17,n50);
and (n1027,n24,n54);
nand (n1028,n1029,n1030,n1031);
nand (n1029,n962,n966);
nand (n1030,n971,n966);
nand (n1031,n962,n971);
xor (n1032,n1033,n1039);
xor (n1033,n1034,n1038);
xor (n1034,n1035,n64);
or (n1035,n1036,n1037);
and (n1036,n28,n80);
and (n1037,n158,n84);
and (n1038,n31,n967);
xor (n1039,n1040,n69);
or (n1040,n1041,n1042);
and (n1041,n162,n62);
and (n1042,n203,n67);
xor (n1043,n1044,n1068);
xor (n1044,n1045,n1049);
nand (n1045,n1046,n1047,n1048);
nand (n1046,n975,n979);
nand (n1047,n983,n979);
nand (n1048,n975,n983);
xor (n1049,n1050,n1059);
xor (n1050,n1051,n1055);
xor (n1051,n1052,n100);
or (n1052,n1053,n1054);
and (n1053,n277,n94);
and (n1054,n455,n98);
xor (n1055,n1056,n15);
or (n1056,n1057,n1058);
and (n1057,n540,n118);
and (n1058,n653,n121);
xor (n1059,n1060,n1064);
xnor (n1060,n1061,n558);
nor (n1061,n1062,n1063);
and (n1062,n89,n668);
and (n1063,n83,n670);
xor (n1064,n1065,n300);
or (n1065,n1066,n1067);
and (n1066,n61,n556);
and (n1067,n66,n560);
nand (n1068,n1069,n1070,n1071);
nand (n1069,n911,n915);
nand (n1070,n916,n915);
nand (n1071,n911,n916);
xor (n1072,n1073,n1092);
xor (n1073,n1074,n1088);
xor (n1074,n1075,n1084);
xor (n1075,n1076,n1080);
xor (n1076,n1077,n20);
or (n1077,n1078,n1079);
and (n1078,n657,n13);
and (n1079,n659,n18);
xor (n1080,n1081,n31);
or (n1081,n1082,n1083);
and (n1082,n682,n25);
and (n1083,n696,n29);
nand (n1084,n1085,n1086,n1087);
nand (n1085,n938,n942);
nand (n1086,n946,n942);
nand (n1087,n938,n946);
nand (n1088,n1089,n1090,n1091);
nand (n1089,n932,n936);
nand (n1090,n950,n936);
nand (n1091,n932,n950);
nand (n1092,n1093,n1094,n1095);
nand (n1093,n956,n960);
nand (n1094,n973,n960);
nand (n1095,n956,n973);
nor (n1096,n1097,n1202);
nor (n1097,n1098,n1102);
nand (n1098,n1099,n1100,n1101);
nand (n1099,n1002,n1006);
nand (n1100,n1010,n1006);
nand (n1101,n1002,n1010);
xor (n1102,n1103,n1198);
xor (n1103,n1104,n1138);
xor (n1104,n1105,n1134);
xor (n1105,n1106,n1110);
nand (n1106,n1107,n1108,n1109);
nand (n1107,n1014,n1028);
nand (n1108,n1032,n1028);
nand (n1109,n1014,n1032);
xor (n1110,n1111,n1120);
xor (n1111,n1112,n1116);
xor (n1112,n1113,n31);
or (n1113,n1114,n1115);
and (n1114,n659,n25);
and (n1115,n682,n29);
nand (n1116,n1117,n1118,n1119);
nand (n1117,n1034,n1038);
nand (n1118,n1039,n1038);
nand (n1119,n1034,n1039);
xor (n1120,n1121,n1130);
xor (n1121,n1122,n1126);
xor (n1122,n1123,n46);
or (n1123,n1124,n1125);
and (n1124,n112,n40);
and (n1125,n117,n44);
xnor (n1126,n1127,n558);
nor (n1127,n1128,n1129);
and (n1128,n83,n668);
and (n1129,n53,n670);
xor (n1130,n1131,n42);
or (n1131,n1132,n1133);
and (n1132,n66,n298);
and (n1133,n97,n302);
nand (n1134,n1135,n1136,n1137);
nand (n1135,n1045,n1049);
nand (n1136,n1068,n1049);
nand (n1137,n1045,n1068);
xor (n1138,n1139,n1194);
xor (n1139,n1140,n1162);
xor (n1140,n1141,n1150);
xor (n1141,n1142,n1146);
nand (n1142,n1143,n1144,n1145);
nand (n1143,n1016,n1020);
nand (n1144,n1024,n1020);
nand (n1145,n1016,n1024);
nand (n1146,n1147,n1148,n1149);
nand (n1147,n1051,n1055);
nand (n1148,n1059,n1055);
nand (n1149,n1051,n1059);
xor (n1150,n1151,n1158);
xor (n1151,n1152,n1156);
xor (n1152,n1153,n56);
or (n1153,n1154,n1155);
and (n1154,n12,n50);
and (n1155,n17,n54);
xnor (n1156,n1157,n74);
nand (n1157,n696,n159);
xor (n1158,n1159,n64);
or (n1159,n1160,n1161);
and (n1160,n24,n80);
and (n1161,n28,n84);
xor (n1162,n1163,n1182);
xor (n1163,n1164,n1168);
nand (n1164,n1165,n1166,n1167);
nand (n1165,n1076,n1080);
nand (n1166,n1084,n1080);
nand (n1167,n1076,n1084);
xor (n1168,n1169,n1178);
xor (n1169,n1170,n1174);
xor (n1170,n1171,n69);
or (n1171,n1172,n1173);
and (n1172,n158,n62);
and (n1173,n162,n67);
xor (n1174,n1175,n100);
or (n1175,n1176,n1177);
and (n1176,n203,n94);
and (n1177,n277,n98);
xor (n1178,n1179,n15);
or (n1179,n1180,n1181);
and (n1180,n455,n118);
and (n1181,n540,n121);
xor (n1182,n1183,n1190);
xor (n1183,n1184,n1189);
xor (n1184,n74,n1185);
xor (n1185,n1186,n300);
or (n1186,n1187,n1188);
and (n1187,n89,n556);
and (n1188,n61,n560);
and (n1189,n1060,n1064);
xor (n1190,n1191,n20);
or (n1191,n1192,n1193);
and (n1192,n653,n13);
and (n1193,n657,n18);
nand (n1194,n1195,n1196,n1197);
nand (n1195,n1074,n1088);
nand (n1196,n1092,n1088);
nand (n1197,n1074,n1092);
nand (n1198,n1199,n1200,n1201);
nand (n1199,n1012,n1043);
nand (n1200,n1072,n1043);
nand (n1201,n1012,n1072);
nor (n1202,n1203,n1207);
nand (n1203,n1204,n1205,n1206);
nand (n1204,n1104,n1138);
nand (n1205,n1198,n1138);
nand (n1206,n1104,n1198);
xor (n1207,n1208,n1217);
xor (n1208,n1209,n1213);
nand (n1209,n1210,n1211,n1212);
nand (n1210,n1106,n1110);
nand (n1211,n1134,n1110);
nand (n1212,n1106,n1134);
nand (n1213,n1214,n1215,n1216);
nand (n1214,n1140,n1162);
nand (n1215,n1194,n1162);
nand (n1216,n1140,n1194);
xor (n1217,n1218,n1279);
xor (n1218,n1219,n1243);
xor (n1219,n1220,n1239);
xor (n1220,n1221,n1225);
nand (n1221,n1222,n1223,n1224);
nand (n1222,n1170,n1174);
nand (n1223,n1178,n1174);
nand (n1224,n1170,n1178);
xor (n1225,n1226,n1235);
xor (n1226,n1227,n1231);
xor (n1227,n1228,n64);
or (n1228,n1229,n1230);
and (n1229,n17,n80);
and (n1230,n24,n84);
xor (n1231,n1232,n69);
or (n1232,n1233,n1234);
and (n1233,n28,n62);
and (n1234,n158,n67);
xor (n1235,n1236,n100);
or (n1236,n1237,n1238);
and (n1237,n162,n94);
and (n1238,n203,n98);
nand (n1239,n1240,n1241,n1242);
nand (n1240,n1184,n1189);
nand (n1241,n1190,n1189);
nand (n1242,n1184,n1190);
xor (n1243,n1244,n1265);
xor (n1244,n1245,n1261);
xor (n1245,n1246,n1260);
xor (n1246,n1247,n1251);
xor (n1247,n1248,n15);
or (n1248,n1249,n1250);
and (n1249,n277,n118);
and (n1250,n455,n121);
xor (n1251,n1252,n1256);
xnor (n1252,n1253,n558);
nor (n1253,n1254,n1255);
and (n1254,n53,n668);
and (n1255,n39,n670);
xor (n1256,n1257,n300);
or (n1257,n1258,n1259);
and (n1258,n83,n556);
and (n1259,n89,n560);
and (n1260,n74,n1185);
nand (n1261,n1262,n1263,n1264);
nand (n1262,n1112,n1116);
nand (n1263,n1120,n1116);
nand (n1264,n1112,n1120);
xor (n1265,n1266,n1275);
xor (n1266,n1267,n1271);
xor (n1267,n1268,n20);
or (n1268,n1269,n1270);
and (n1269,n540,n13);
and (n1270,n653,n18);
xor (n1271,n1272,n74);
or (n1272,n1273,n1274);
and (n1273,n682,n159);
and (n1274,n696,n163);
xor (n1275,n1276,n31);
or (n1276,n1277,n1278);
and (n1277,n657,n25);
and (n1278,n659,n29);
xor (n1279,n1280,n1309);
xor (n1280,n1281,n1305);
xor (n1281,n1282,n1301);
xor (n1282,n1283,n1287);
nand (n1283,n1284,n1285,n1286);
nand (n1284,n1122,n1126);
nand (n1285,n1130,n1126);
nand (n1286,n1122,n1130);
xor (n1287,n1288,n1297);
xor (n1288,n1289,n1293);
xor (n1289,n1290,n46);
or (n1290,n1291,n1292);
and (n1291,n97,n40);
and (n1292,n112,n44);
xor (n1293,n1294,n42);
or (n1294,n1295,n1296);
and (n1295,n61,n298);
and (n1296,n66,n302);
xor (n1297,n1298,n56);
or (n1298,n1299,n1300);
and (n1299,n117,n50);
and (n1300,n12,n54);
nand (n1301,n1302,n1303,n1304);
nand (n1302,n1152,n1156);
nand (n1303,n1158,n1156);
nand (n1304,n1152,n1158);
nand (n1305,n1306,n1307,n1308);
nand (n1306,n1142,n1146);
nand (n1307,n1150,n1146);
nand (n1308,n1142,n1150);
nand (n1309,n1310,n1311,n1312);
nand (n1310,n1164,n1168);
nand (n1311,n1182,n1168);
nand (n1312,n1164,n1182);
nor (n1313,n1314,n1586);
nor (n1314,n1315,n1562);
nor (n1315,n1316,n1560);
nor (n1316,n1317,n1535);
nand (n1317,n1318,n1497);
nand (n1318,n1319,n1444,n1496);
nand (n1319,n1320,n1371);
xor (n1320,n1321,n1358);
xor (n1321,n1322,n1343);
nand (n1322,n1323,n1337,n1342);
nand (n1323,n1324,n1333);
and (n1324,n1325,n1329);
xnor (n1325,n1326,n558);
nor (n1326,n1327,n1328);
and (n1327,n24,n668);
and (n1328,n17,n670);
xor (n1329,n1330,n300);
or (n1330,n1331,n1332);
and (n1331,n28,n556);
and (n1332,n158,n560);
xor (n1333,n1334,n64);
or (n1334,n1335,n1336);
and (n1335,n653,n80);
and (n1336,n657,n84);
nand (n1337,n1338,n1333);
xor (n1338,n1339,n69);
or (n1339,n1340,n1341);
and (n1340,n659,n62);
and (n1341,n682,n67);
nand (n1342,n1324,n1338);
xor (n1343,n1344,n1353);
xor (n1344,n1345,n1349);
xor (n1345,n1346,n46);
or (n1346,n1347,n1348);
and (n1347,n162,n40);
and (n1348,n203,n44);
xor (n1349,n1350,n42);
or (n1350,n1351,n1352);
and (n1351,n28,n298);
and (n1352,n158,n302);
and (n1353,n1354,n100);
xnor (n1354,n1355,n558);
nor (n1355,n1356,n1357);
and (n1356,n17,n668);
and (n1357,n12,n670);
nand (n1358,n1359,n1365,n1370);
nand (n1359,n1360,n1364);
xor (n1360,n1361,n42);
or (n1361,n1362,n1363);
and (n1362,n158,n298);
and (n1363,n162,n302);
xor (n1364,n1354,n100);
nand (n1365,n1366,n1364);
xor (n1366,n1367,n56);
or (n1367,n1368,n1369);
and (n1368,n455,n50);
and (n1369,n540,n54);
nand (n1370,n1360,n1366);
xor (n1371,n1372,n1408);
xor (n1372,n1373,n1384);
xor (n1373,n1374,n1380);
xor (n1374,n1375,n1379);
xor (n1375,n1376,n56);
or (n1376,n1377,n1378);
and (n1377,n277,n50);
and (n1378,n455,n54);
xor (n1379,n783,n787);
xor (n1380,n1381,n64);
or (n1381,n1382,n1383);
and (n1382,n540,n80);
and (n1383,n653,n84);
xor (n1384,n1385,n1394);
xor (n1385,n1386,n1390);
xor (n1386,n1387,n69);
or (n1387,n1388,n1389);
and (n1388,n657,n62);
and (n1389,n659,n67);
xor (n1390,n1391,n100);
or (n1391,n1392,n1393);
and (n1392,n682,n94);
and (n1393,n696,n98);
nand (n1394,n1395,n1402,n1407);
nand (n1395,n1396,n1400);
xor (n1396,n1397,n300);
or (n1397,n1398,n1399);
and (n1398,n24,n556);
and (n1399,n28,n560);
xnor (n1400,n1401,n100);
nand (n1401,n696,n94);
nand (n1402,n1403,n1400);
xor (n1403,n1404,n46);
or (n1404,n1405,n1406);
and (n1405,n203,n40);
and (n1406,n277,n44);
nand (n1407,n1396,n1403);
nand (n1408,n1409,n1429,n1443);
nand (n1409,n1410,n1412);
xor (n1410,n1411,n1403);
xor (n1411,n1396,n1400);
nand (n1412,n1413,n1422,n1428);
nand (n1413,n1414,n1418);
xor (n1414,n1415,n46);
or (n1415,n1416,n1417);
and (n1416,n277,n40);
and (n1417,n455,n44);
xor (n1418,n1419,n42);
or (n1419,n1420,n1421);
and (n1420,n162,n298);
and (n1421,n203,n302);
nand (n1422,n1423,n1418);
and (n1423,n1424,n69);
xnor (n1424,n1425,n558);
nor (n1425,n1426,n1427);
and (n1426,n28,n668);
and (n1427,n24,n670);
nand (n1428,n1414,n1423);
nand (n1429,n1430,n1412);
nand (n1430,n1431,n1437,n1442);
nand (n1431,n1432,n1436);
xor (n1432,n1433,n56);
or (n1433,n1434,n1435);
and (n1434,n540,n50);
and (n1435,n653,n54);
xor (n1436,n1325,n1329);
nand (n1437,n1438,n1436);
xor (n1438,n1439,n64);
or (n1439,n1440,n1441);
and (n1440,n657,n80);
and (n1441,n659,n84);
nand (n1442,n1432,n1438);
nand (n1443,n1410,n1430);
nand (n1444,n1445,n1371);
nand (n1445,n1446,n1451,n1495);
nand (n1446,n1447,n1449);
xor (n1447,n1448,n1338);
xor (n1448,n1324,n1333);
xor (n1449,n1450,n1366);
xor (n1450,n1360,n1364);
nand (n1451,n1452,n1449);
nand (n1452,n1453,n1472,n1494);
nand (n1453,n1454,n1458);
xor (n1454,n1455,n69);
or (n1455,n1456,n1457);
and (n1456,n682,n62);
and (n1457,n696,n67);
nand (n1458,n1459,n1466,n1471);
nand (n1459,n1460,n1464);
xor (n1460,n1461,n300);
or (n1461,n1462,n1463);
and (n1462,n158,n556);
and (n1463,n162,n560);
xnor (n1464,n1465,n69);
nand (n1465,n696,n62);
nand (n1466,n1467,n1464);
xor (n1467,n1468,n46);
or (n1468,n1469,n1470);
and (n1469,n455,n40);
and (n1470,n540,n44);
nand (n1471,n1460,n1467);
nand (n1472,n1473,n1458);
nand (n1473,n1474,n1488,n1493);
nand (n1474,n1475,n1479);
xor (n1475,n1476,n42);
or (n1476,n1477,n1478);
and (n1477,n203,n298);
and (n1478,n277,n302);
and (n1479,n1480,n1484);
xnor (n1480,n1481,n558);
nor (n1481,n1482,n1483);
and (n1482,n158,n668);
and (n1483,n28,n670);
xor (n1484,n1485,n300);
or (n1485,n1486,n1487);
and (n1486,n162,n556);
and (n1487,n203,n560);
nand (n1488,n1489,n1479);
xor (n1489,n1490,n56);
or (n1490,n1491,n1492);
and (n1491,n653,n50);
and (n1492,n657,n54);
nand (n1493,n1475,n1489);
nand (n1494,n1454,n1473);
nand (n1495,n1447,n1452);
nand (n1496,n1320,n1445);
xor (n1497,n1498,n1513);
xor (n1498,n1499,n1509);
xor (n1499,n1500,n1507);
xor (n1500,n1501,n1505);
nand (n1501,n1502,n1503,n1504);
nand (n1502,n1345,n1349);
nand (n1503,n1353,n1349);
nand (n1504,n1345,n1353);
xor (n1505,n1506,n796);
xor (n1506,n782,n791);
xor (n1507,n1508,n897);
xor (n1508,n891,n895);
nand (n1509,n1510,n1511,n1512);
nand (n1510,n1373,n1384);
nand (n1511,n1408,n1384);
nand (n1512,n1373,n1408);
xor (n1513,n1514,n1523);
xor (n1514,n1515,n1519);
nand (n1515,n1516,n1517,n1518);
nand (n1516,n1386,n1390);
nand (n1517,n1394,n1390);
nand (n1518,n1386,n1394);
nand (n1519,n1520,n1521,n1522);
nand (n1520,n1322,n1343);
nand (n1521,n1358,n1343);
nand (n1522,n1322,n1358);
xor (n1523,n1524,n1533);
xor (n1524,n1525,n1529);
xor (n1525,n1526,n100);
or (n1526,n1527,n1528);
and (n1527,n659,n94);
and (n1528,n682,n98);
nand (n1529,n1530,n1531,n1532);
nand (n1530,n1375,n1379);
nand (n1531,n1380,n1379);
nand (n1532,n1375,n1380);
xor (n1533,n1534,n883);
xor (n1534,n874,n878);
nor (n1535,n1536,n1540);
nand (n1536,n1537,n1538,n1539);
nand (n1537,n1499,n1509);
nand (n1538,n1513,n1509);
nand (n1539,n1499,n1513);
xor (n1540,n1541,n1548);
xor (n1541,n1542,n1544);
xor (n1542,n1543,n804);
xor (n1543,n780,n801);
nand (n1544,n1545,n1546,n1547);
nand (n1545,n1515,n1519);
nand (n1546,n1523,n1519);
nand (n1547,n1515,n1523);
xor (n1548,n1549,n1558);
xor (n1549,n1550,n1554);
nand (n1550,n1551,n1552,n1553);
nand (n1551,n1525,n1529);
nand (n1552,n1533,n1529);
nand (n1553,n1525,n1533);
nand (n1554,n1555,n1556,n1557);
nand (n1555,n1501,n1505);
nand (n1556,n1507,n1505);
nand (n1557,n1501,n1507);
xor (n1558,n1559,n889);
xor (n1559,n872,n886);
not (n1560,n1561);
nand (n1561,n1536,n1540);
not (n1562,n1563);
nor (n1563,n1564,n1579);
nor (n1564,n1565,n1569);
nand (n1565,n1566,n1567,n1568);
nand (n1566,n1542,n1544);
nand (n1567,n1548,n1544);
nand (n1568,n1542,n1548);
xor (n1569,n1570,n1577);
xor (n1570,n1571,n1573);
xor (n1571,n1572,n870);
xor (n1572,n863,n867);
nand (n1573,n1574,n1575,n1576);
nand (n1574,n1550,n1554);
nand (n1575,n1558,n1554);
nand (n1576,n1550,n1558);
xor (n1577,n1578,n778);
xor (n1578,n724,n726);
nor (n1579,n1580,n1584);
nand (n1580,n1581,n1582,n1583);
nand (n1581,n1571,n1573);
nand (n1582,n1577,n1573);
nand (n1583,n1571,n1577);
xor (n1584,n1585,n821);
xor (n1585,n645,n722);
not (n1586,n1587);
nor (n1587,n1588,n1590);
nor (n1588,n1589,n1579);
nand (n1589,n1565,n1569);
not (n1590,n1591);
nand (n1591,n1580,n1584);
not (n1592,n1593);
nor (n1593,n1594,n1601);
nor (n1594,n1595,n1600);
nor (n1595,n1596,n1598);
nor (n1596,n1597,n995);
nand (n1597,n643,n905);
not (n1598,n1599);
nand (n1599,n996,n1000);
not (n1600,n1096);
not (n1601,n1602);
nor (n1602,n1603,n1605);
nor (n1603,n1604,n1202);
nand (n1604,n1098,n1102);
not (n1605,n1606);
nand (n1606,n1203,n1207);
not (n1607,n1608);
nor (n1608,n1609,n2024);
nand (n1609,n1610,n1837);
nor (n1610,n1611,n1723);
nor (n1611,n1612,n1616);
nand (n1612,n1613,n1614,n1615);
nand (n1613,n1209,n1213);
nand (n1614,n1217,n1213);
nand (n1615,n1209,n1217);
xor (n1616,n1617,n1719);
xor (n1617,n1618,n1651);
xor (n1618,n1619,n1647);
xor (n1619,n1620,n1643);
xor (n1620,n1621,n1639);
xor (n1621,n1622,n1635);
xor (n1622,n1623,n1632);
xor (n1623,n1624,n1628);
xor (n1624,n1625,n300);
or (n1625,n1626,n1627);
and (n1626,n53,n556);
and (n1627,n83,n560);
xor (n1628,n1629,n42);
or (n1629,n1630,n1631);
and (n1630,n89,n298);
and (n1631,n61,n302);
xnor (n1632,n1633,n558);
nor (n1633,n1634,n1255);
and (n1634,n39,n668);
nand (n1635,n1636,n1637,n1638);
nand (n1636,n1227,n1231);
nand (n1637,n1235,n1231);
nand (n1638,n1227,n1235);
nand (n1639,n1640,n1641,n1642);
nand (n1640,n1247,n1251);
nand (n1641,n1260,n1251);
nand (n1642,n1247,n1260);
nand (n1643,n1644,n1645,n1646);
nand (n1644,n1221,n1225);
nand (n1645,n1239,n1225);
nand (n1646,n1221,n1239);
nand (n1647,n1648,n1649,n1650);
nand (n1648,n1245,n1261);
nand (n1649,n1265,n1261);
nand (n1650,n1245,n1265);
xor (n1651,n1652,n1715);
xor (n1652,n1653,n1691);
xor (n1653,n1654,n1676);
xor (n1654,n1655,n1669);
xor (n1655,n1656,n1665);
xor (n1656,n1657,n1661);
xor (n1657,n1658,n56);
or (n1658,n1659,n1660);
and (n1659,n112,n50);
and (n1660,n117,n54);
xor (n1661,n1662,n64);
or (n1662,n1663,n1664);
and (n1663,n12,n80);
and (n1664,n17,n84);
xor (n1665,n1666,n69);
or (n1666,n1667,n1668);
and (n1667,n24,n62);
and (n1668,n28,n67);
xor (n1669,n1670,n1672);
xor (n1670,n74,n1671);
and (n1671,n1252,n1256);
xor (n1672,n1673,n20);
or (n1673,n1674,n1675);
and (n1674,n455,n13);
and (n1675,n540,n18);
xor (n1676,n1677,n1686);
xor (n1677,n1678,n1682);
xor (n1678,n1679,n100);
or (n1679,n1680,n1681);
and (n1680,n158,n94);
and (n1681,n162,n98);
xor (n1682,n1683,n15);
or (n1683,n1684,n1685);
and (n1684,n203,n118);
and (n1685,n277,n121);
xor (n1686,n74,n1687);
xor (n1687,n1688,n46);
or (n1688,n1689,n1690);
and (n1689,n66,n40);
and (n1690,n97,n44);
xor (n1691,n1692,n1701);
xor (n1692,n1693,n1697);
nand (n1693,n1694,n1695,n1696);
nand (n1694,n1267,n1271);
nand (n1695,n1275,n1271);
nand (n1696,n1267,n1275);
nand (n1697,n1698,n1699,n1700);
nand (n1698,n1283,n1287);
nand (n1699,n1301,n1287);
nand (n1700,n1283,n1301);
xor (n1701,n1702,n1711);
xor (n1702,n1703,n1707);
xor (n1703,n1704,n31);
or (n1704,n1705,n1706);
and (n1705,n653,n25);
and (n1706,n657,n29);
xor (n1707,n1708,n74);
or (n1708,n1709,n1710);
and (n1709,n659,n159);
and (n1710,n682,n163);
nand (n1711,n1712,n1713,n1714);
nand (n1712,n1289,n1293);
nand (n1713,n1297,n1293);
nand (n1714,n1289,n1297);
nand (n1715,n1716,n1717,n1718);
nand (n1716,n1281,n1305);
nand (n1717,n1309,n1305);
nand (n1718,n1281,n1309);
nand (n1719,n1720,n1721,n1722);
nand (n1720,n1219,n1243);
nand (n1721,n1279,n1243);
nand (n1722,n1219,n1279);
nor (n1723,n1724,n1728);
nand (n1724,n1725,n1726,n1727);
nand (n1725,n1618,n1651);
nand (n1726,n1719,n1651);
nand (n1727,n1618,n1719);
xor (n1728,n1729,n1738);
xor (n1729,n1730,n1734);
nand (n1730,n1731,n1732,n1733);
nand (n1731,n1620,n1643);
nand (n1732,n1647,n1643);
nand (n1733,n1620,n1647);
nand (n1734,n1735,n1736,n1737);
nand (n1735,n1653,n1691);
nand (n1736,n1715,n1691);
nand (n1737,n1653,n1715);
xor (n1738,n1739,n1796);
xor (n1739,n1740,n1771);
xor (n1740,n1741,n1757);
xor (n1741,n1742,n1746);
nand (n1742,n1743,n1744,n1745);
nand (n1743,n74,n1671);
nand (n1744,n1672,n1671);
nand (n1745,n74,n1672);
xor (n1746,n1747,n1753);
xor (n1747,n1748,n1752);
xor (n1748,n1749,n15);
or (n1749,n1750,n1751);
and (n1750,n162,n118);
and (n1751,n203,n121);
and (n1752,n74,n1687);
xor (n1753,n1754,n20);
or (n1754,n1755,n1756);
and (n1755,n277,n13);
and (n1756,n455,n18);
xor (n1757,n1758,n1767);
xor (n1758,n1759,n1763);
xor (n1759,n1760,n31);
or (n1760,n1761,n1762);
and (n1761,n540,n25);
and (n1762,n653,n29);
xor (n1763,n1764,n74);
or (n1764,n1765,n1766);
and (n1765,n657,n159);
and (n1766,n659,n163);
nand (n1767,n1768,n1769,n1770);
nand (n1768,n1624,n1628);
nand (n1769,n1632,n1628);
nand (n1770,n1624,n1632);
xor (n1771,n1772,n1781);
xor (n1772,n1773,n1777);
nand (n1773,n1774,n1775,n1776);
nand (n1774,n1703,n1707);
nand (n1775,n1711,n1707);
nand (n1776,n1703,n1711);
nand (n1777,n1778,n1779,n1780);
nand (n1778,n1622,n1635);
nand (n1779,n1639,n1635);
nand (n1780,n1622,n1639);
xor (n1781,n1782,n74);
xor (n1782,n1783,n1787);
nand (n1783,n1784,n1785,n1786);
nand (n1784,n1657,n1661);
nand (n1785,n1665,n1661);
nand (n1786,n1657,n1665);
xor (n1787,n1788,n1793);
not (n1788,n1789);
xor (n1789,n1790,n46);
or (n1790,n1791,n1792);
and (n1791,n61,n40);
and (n1792,n66,n44);
xor (n1793,n1794,n300);
or (n1794,n555,n1795);
and (n1795,n53,n560);
xor (n1796,n1797,n1833);
xor (n1797,n1798,n1802);
nand (n1798,n1799,n1800,n1801);
nand (n1799,n1655,n1669);
nand (n1800,n1676,n1669);
nand (n1801,n1655,n1676);
xor (n1802,n1803,n1822);
xor (n1803,n1804,n1808);
nand (n1804,n1805,n1806,n1807);
nand (n1805,n1678,n1682);
nand (n1806,n1686,n1682);
nand (n1807,n1678,n1686);
xor (n1808,n1809,n1818);
xor (n1809,n1810,n1814);
xor (n1810,n1811,n64);
or (n1811,n1812,n1813);
and (n1812,n117,n80);
and (n1813,n12,n84);
xor (n1814,n1815,n69);
or (n1815,n1816,n1817);
and (n1816,n17,n62);
and (n1817,n24,n67);
xor (n1818,n1819,n100);
or (n1819,n1820,n1821);
and (n1820,n28,n94);
and (n1821,n158,n98);
xor (n1822,n1823,n1829);
xor (n1823,n1824,n1828);
xor (n1824,n1825,n42);
or (n1825,n1826,n1827);
and (n1826,n83,n298);
and (n1827,n89,n302);
not (n1828,n1632);
xor (n1829,n1830,n56);
or (n1830,n1831,n1832);
and (n1831,n97,n50);
and (n1832,n112,n54);
nand (n1833,n1834,n1835,n1836);
nand (n1834,n1693,n1697);
nand (n1835,n1701,n1697);
nand (n1836,n1693,n1701);
nor (n1837,n1838,n1945);
nor (n1838,n1839,n1843);
nand (n1839,n1840,n1841,n1842);
nand (n1840,n1730,n1734);
nand (n1841,n1738,n1734);
nand (n1842,n1730,n1738);
xor (n1843,n1844,n1941);
xor (n1844,n1845,n1885);
xor (n1845,n1846,n1881);
xor (n1846,n1847,n1877);
xor (n1847,n1848,n1873);
xor (n1848,n1849,n1863);
xor (n1849,n1850,n1859);
xor (n1850,n1851,n1855);
xor (n1851,n1852,n64);
or (n1852,n1853,n1854);
and (n1853,n112,n80);
and (n1854,n117,n84);
xor (n1855,n1856,n69);
or (n1856,n1857,n1858);
and (n1857,n12,n62);
and (n1858,n17,n67);
xor (n1859,n1860,n15);
or (n1860,n1861,n1862);
and (n1861,n158,n118);
and (n1862,n162,n121);
xor (n1863,n1864,n1869);
xor (n1864,n1865,n553);
xor (n1865,n1866,n46);
or (n1866,n1867,n1868);
and (n1867,n89,n40);
and (n1868,n61,n44);
xor (n1869,n1870,n56);
or (n1870,n1871,n1872);
and (n1871,n66,n50);
and (n1872,n97,n54);
nand (n1873,n1874,n1875,n1876);
nand (n1874,n1748,n1752);
nand (n1875,n1753,n1752);
nand (n1876,n1748,n1753);
nand (n1877,n1878,n1879,n1880);
nand (n1878,n1742,n1746);
nand (n1879,n1757,n1746);
nand (n1880,n1742,n1757);
nand (n1881,n1882,n1883,n1884);
nand (n1882,n1773,n1777);
nand (n1883,n1781,n1777);
nand (n1884,n1773,n1781);
xor (n1885,n1886,n1937);
xor (n1886,n1887,n1908);
xor (n1887,n1888,n1904);
xor (n1888,n1889,n1900);
xor (n1889,n1890,n1896);
xor (n1890,n1891,n1892);
not (n1891,n594);
xor (n1892,n1893,n100);
or (n1893,n1894,n1895);
and (n1894,n24,n94);
and (n1895,n28,n98);
xor (n1896,n1897,n20);
or (n1897,n1898,n1899);
and (n1898,n203,n13);
and (n1899,n277,n18);
nand (n1900,n1901,n1902,n1903);
nand (n1901,n1759,n1763);
nand (n1902,n1767,n1763);
nand (n1903,n1759,n1767);
nand (n1904,n1905,n1906,n1907);
nand (n1905,n1783,n1787);
nand (n1906,n74,n1787);
nand (n1907,n1783,n74);
xor (n1908,n1909,n1933);
xor (n1909,n1910,n1923);
xor (n1910,n1911,n1920);
xor (n1911,n1912,n1916);
xor (n1912,n1913,n31);
or (n1913,n1914,n1915);
and (n1914,n455,n25);
and (n1915,n540,n29);
xor (n1916,n1917,n74);
or (n1917,n1918,n1919);
and (n1918,n653,n159);
and (n1919,n657,n163);
nand (n1920,n1788,n1921,n1922);
nand (n1921,n1793,n1789);
not (n1922,n1793);
xor (n1923,n1924,n1929);
xor (n1924,n74,n1925);
nand (n1925,n1926,n1927,n1928);
nand (n1926,n1824,n1828);
nand (n1927,n1829,n1828);
nand (n1928,n1824,n1829);
nand (n1929,n1930,n1931,n1932);
nand (n1930,n1810,n1814);
nand (n1931,n1818,n1814);
nand (n1932,n1810,n1818);
nand (n1933,n1934,n1935,n1936);
nand (n1934,n1804,n1808);
nand (n1935,n1822,n1808);
nand (n1936,n1804,n1822);
nand (n1937,n1938,n1939,n1940);
nand (n1938,n1798,n1802);
nand (n1939,n1833,n1802);
nand (n1940,n1798,n1833);
nand (n1941,n1942,n1943,n1944);
nand (n1942,n1740,n1771);
nand (n1943,n1796,n1771);
nand (n1944,n1740,n1796);
nor (n1945,n1946,n1950);
nand (n1946,n1947,n1948,n1949);
nand (n1947,n1845,n1885);
nand (n1948,n1941,n1885);
nand (n1949,n1845,n1941);
xor (n1950,n1951,n1960);
xor (n1951,n1952,n1956);
nand (n1952,n1953,n1954,n1955);
nand (n1953,n1847,n1877);
nand (n1954,n1881,n1877);
nand (n1955,n1847,n1881);
nand (n1956,n1957,n1958,n1959);
nand (n1957,n1887,n1908);
nand (n1958,n1937,n1908);
nand (n1959,n1887,n1937);
xor (n1960,n1961,n1992);
xor (n1961,n1962,n1966);
nand (n1962,n1963,n1964,n1965);
nand (n1963,n1910,n1923);
nand (n1964,n1933,n1923);
nand (n1965,n1910,n1933);
xor (n1966,n1967,n1980);
xor (n1967,n1968,n1972);
nand (n1968,n1969,n1970,n1971);
nand (n1969,n74,n1925);
nand (n1970,n1929,n1925);
nand (n1971,n74,n1929);
xor (n1972,n1973,n1976);
xor (n1973,n1974,n74);
xor (n1974,n1975,n552);
xor (n1975,n544,n547);
nand (n1976,n1977,n1978,n1979);
nand (n1977,n1865,n553);
nand (n1978,n1869,n553);
nand (n1979,n1865,n1869);
xor (n1980,n1981,n1988);
xor (n1981,n1982,n1984);
xor (n1982,n1983,n580);
xor (n1983,n571,n575);
nand (n1984,n1985,n1986,n1987);
nand (n1985,n1851,n1855);
nand (n1986,n1859,n1855);
nand (n1987,n1851,n1859);
nand (n1988,n1989,n1990,n1991);
nand (n1989,n1912,n1916);
nand (n1990,n1920,n1916);
nand (n1991,n1912,n1920);
xor (n1992,n1993,n2002);
xor (n1993,n1994,n1998);
nand (n1994,n1995,n1996,n1997);
nand (n1995,n1849,n1863);
nand (n1996,n1873,n1863);
nand (n1997,n1849,n1873);
nand (n1998,n1999,n2000,n2001);
nand (n1999,n1889,n1900);
nand (n2000,n1904,n1900);
nand (n2001,n1889,n1904);
xor (n2002,n2003,n2010);
xor (n2003,n2004,n2008);
nand (n2004,n2005,n2006,n2007);
nand (n2005,n1891,n1892);
nand (n2006,n1896,n1892);
nand (n2007,n1891,n1896);
xor (n2008,n2009,n599);
xor (n2009,n590,n594);
xor (n2010,n2011,n2020);
xor (n2011,n2012,n2016);
xor (n2012,n2013,n20);
or (n2013,n2014,n2015);
and (n2014,n162,n13);
and (n2015,n203,n18);
xor (n2016,n2017,n31);
or (n2017,n2018,n2019);
and (n2018,n277,n25);
and (n2019,n455,n29);
xor (n2020,n2021,n74);
or (n2021,n2022,n2023);
and (n2022,n540,n159);
and (n2023,n653,n163);
nand (n2024,n2025,n2109);
nor (n2025,n2026,n2076);
nor (n2026,n2027,n2031);
nand (n2027,n2028,n2029,n2030);
nand (n2028,n1952,n1956);
nand (n2029,n1960,n1956);
nand (n2030,n1952,n1960);
xor (n2031,n2032,n2072);
xor (n2032,n2033,n2053);
xor (n2033,n2034,n2041);
xor (n2034,n2035,n2037);
xor (n2035,n2036,n588);
xor (n2036,n569,n585);
nand (n2037,n2038,n2039,n2040);
nand (n2038,n2004,n2008);
nand (n2039,n2010,n2008);
nand (n2040,n2004,n2010);
xor (n2041,n2042,n2049);
xor (n2042,n2043,n2047);
nand (n2043,n2044,n2045,n2046);
nand (n2044,n2012,n2016);
nand (n2045,n2020,n2016);
nand (n2046,n2012,n2020);
xor (n2047,n2048,n498);
xor (n2048,n492,n496);
nand (n2049,n2050,n2051,n2052);
nand (n2050,n1974,n74);
nand (n2051,n1976,n74);
nand (n2052,n1974,n1976);
xor (n2053,n2054,n2068);
xor (n2054,n2055,n2059);
nand (n2055,n2056,n2057,n2058);
nand (n2056,n1968,n1972);
nand (n2057,n1980,n1972);
nand (n2058,n1968,n1980);
xor (n2059,n2060,n2064);
xor (n2060,n2061,n2063);
xor (n2061,n2062,n514);
xor (n2062,n505,n509);
xor (n2063,n537,n542);
nand (n2064,n2065,n2066,n2067);
nand (n2065,n1982,n1984);
nand (n2066,n1988,n1984);
nand (n2067,n1982,n1988);
nand (n2068,n2069,n2070,n2071);
nand (n2069,n1994,n1998);
nand (n2070,n2002,n1998);
nand (n2071,n1994,n2002);
nand (n2072,n2073,n2074,n2075);
nand (n2073,n1962,n1966);
nand (n2074,n1992,n1966);
nand (n2075,n1962,n1992);
nor (n2076,n2077,n2081);
nand (n2077,n2078,n2079,n2080);
nand (n2078,n2033,n2053);
nand (n2079,n2072,n2053);
nand (n2080,n2033,n2072);
xor (n2081,n2082,n2105);
xor (n2082,n2083,n2093);
xor (n2083,n2084,n2091);
xor (n2084,n2085,n2087);
xor (n2085,n2086,n485);
xor (n2086,n470,n482);
nand (n2087,n2088,n2089,n2090);
nand (n2088,n2043,n2047);
nand (n2089,n2049,n2047);
nand (n2090,n2043,n2049);
xor (n2091,n2092,n520);
xor (n2092,n490,n503);
xor (n2093,n2094,n2101);
xor (n2094,n2095,n2097);
xor (n2095,n2096,n567);
xor (n2096,n534,n564);
nand (n2097,n2098,n2099,n2100);
nand (n2098,n2061,n2063);
nand (n2099,n2064,n2063);
nand (n2100,n2061,n2064);
nand (n2101,n2102,n2103,n2104);
nand (n2102,n2035,n2037);
nand (n2103,n2041,n2037);
nand (n2104,n2035,n2041);
nand (n2105,n2106,n2107,n2108);
nand (n2106,n2055,n2059);
nand (n2107,n2068,n2059);
nand (n2108,n2055,n2068);
nor (n2109,n2110,n2127);
nor (n2110,n2111,n2115);
nand (n2111,n2112,n2113,n2114);
nand (n2112,n2083,n2093);
nand (n2113,n2105,n2093);
nand (n2114,n2083,n2105);
xor (n2115,n2116,n2123);
xor (n2116,n2117,n2121);
nand (n2117,n2118,n2119,n2120);
nand (n2118,n2085,n2087);
nand (n2119,n2091,n2087);
nand (n2120,n2085,n2091);
xor (n2121,n2122,n607);
xor (n2122,n530,n532);
nand (n2123,n2124,n2125,n2126);
nand (n2124,n2095,n2097);
nand (n2125,n2101,n2097);
nand (n2126,n2095,n2101);
nor (n2127,n2128,n2132);
nand (n2128,n2129,n2130,n2131);
nand (n2129,n2117,n2121);
nand (n2130,n2123,n2121);
nand (n2131,n2117,n2123);
xor (n2132,n2133,n528);
xor (n2133,n397,n441);
not (n2134,n2135);
nor (n2135,n2136,n2151);
nor (n2136,n2024,n2137);
nor (n2137,n2138,n2145);
nor (n2138,n2139,n2144);
nor (n2139,n2140,n2142);
nor (n2140,n2141,n1723);
nand (n2141,n1612,n1616);
not (n2142,n2143);
nand (n2143,n1724,n1728);
not (n2144,n1837);
not (n2145,n2146);
nor (n2146,n2147,n2149);
nor (n2147,n2148,n1945);
nand (n2148,n1839,n1843);
not (n2149,n2150);
nand (n2150,n1946,n1950);
not (n2151,n2152);
nor (n2152,n2153,n2160);
nor (n2153,n2154,n2159);
nor (n2154,n2155,n2157);
nor (n2155,n2156,n2076);
nand (n2156,n2027,n2031);
not (n2157,n2158);
nand (n2158,n2077,n2081);
not (n2159,n2109);
not (n2160,n2161);
nor (n2161,n2162,n2164);
nor (n2162,n2163,n2127);
nand (n2163,n2111,n2115);
not (n2164,n2165);
nand (n2165,n2128,n2132);
nand (n2166,n2167,n2586);
nand (n2167,n2168,n2479);
nor (n2168,n2169,n2464);
nor (n2169,n2170,n2335);
nand (n2170,n2171,n2312);
nor (n2171,n2172,n2289);
nor (n2172,n2173,n2262);
nand (n2173,n2174,n2219,n2261);
nand (n2174,n2175,n2187);
xor (n2175,n2176,n2182);
xor (n2176,n2177,n2178);
xor (n2177,n1480,n1484);
xor (n2178,n2179,n64);
or (n2179,n2180,n2181);
and (n2180,n682,n80);
and (n2181,n696,n84);
and (n2182,n64,n2183);
xor (n2183,n2184,n300);
or (n2184,n2185,n2186);
and (n2185,n203,n556);
and (n2186,n277,n560);
nand (n2187,n2188,n2205,n2218);
nand (n2188,n2189,n2190);
xor (n2189,n64,n2183);
nand (n2190,n2191,n2200,n2204);
nand (n2191,n2192,n2196);
xor (n2192,n2193,n46);
or (n2193,n2194,n2195);
and (n2194,n657,n40);
and (n2195,n659,n44);
xor (n2196,n2197,n42);
or (n2197,n2198,n2199);
and (n2198,n540,n298);
and (n2199,n653,n302);
nand (n2200,n2201,n2196);
and (n2201,n56,n2202);
xnor (n2202,n2203,n56);
nand (n2203,n696,n50);
nand (n2204,n2192,n2201);
nand (n2205,n2206,n2190);
xor (n2206,n2207,n2214);
xor (n2207,n2208,n2212);
xnor (n2208,n2209,n558);
nor (n2209,n2210,n2211);
and (n2210,n162,n668);
and (n2211,n158,n670);
xnor (n2212,n2213,n64);
nand (n2213,n696,n80);
xor (n2214,n2215,n46);
or (n2215,n2216,n2217);
and (n2216,n653,n40);
and (n2217,n657,n44);
nand (n2218,n2189,n2206);
nand (n2219,n2220,n2187);
xor (n2220,n2221,n2240);
xor (n2221,n2222,n2226);
nand (n2222,n2223,n2224,n2225);
nand (n2223,n2208,n2212);
nand (n2224,n2214,n2212);
nand (n2225,n2208,n2214);
xor (n2226,n2227,n2236);
xor (n2227,n2228,n2232);
xor (n2228,n2229,n46);
or (n2229,n2230,n2231);
and (n2230,n540,n40);
and (n2231,n653,n44);
xor (n2232,n2233,n42);
or (n2233,n2234,n2235);
and (n2234,n277,n298);
and (n2235,n455,n302);
xor (n2236,n2237,n56);
or (n2237,n2238,n2239);
and (n2238,n657,n50);
and (n2239,n659,n54);
nand (n2240,n2241,n2255,n2260);
nand (n2241,n2242,n2246);
xor (n2242,n2243,n42);
or (n2243,n2244,n2245);
and (n2244,n455,n298);
and (n2245,n540,n302);
and (n2246,n2247,n2251);
xnor (n2247,n2248,n558);
nor (n2248,n2249,n2250);
and (n2249,n203,n668);
and (n2250,n162,n670);
xor (n2251,n2252,n300);
or (n2252,n2253,n2254);
and (n2253,n277,n556);
and (n2254,n455,n560);
nand (n2255,n2256,n2246);
xor (n2256,n2257,n56);
or (n2257,n2258,n2259);
and (n2258,n659,n50);
and (n2259,n682,n54);
nand (n2260,n2242,n2256);
nand (n2261,n2175,n2220);
xor (n2262,n2263,n2277);
xor (n2263,n2264,n2273);
xor (n2264,n2265,n2271);
xor (n2265,n2266,n2270);
xor (n2266,n2267,n64);
or (n2267,n2268,n2269);
and (n2268,n659,n80);
and (n2269,n682,n84);
xor (n2270,n1424,n69);
xor (n2271,n2272,n1467);
xor (n2272,n1460,n1464);
nand (n2273,n2274,n2275,n2276);
nand (n2274,n2222,n2226);
nand (n2275,n2240,n2226);
nand (n2276,n2222,n2240);
xor (n2277,n2278,n2287);
xor (n2278,n2279,n2283);
nand (n2279,n2280,n2281,n2282);
nand (n2280,n2177,n2178);
nand (n2281,n2182,n2178);
nand (n2282,n2177,n2182);
nand (n2283,n2284,n2285,n2286);
nand (n2284,n2228,n2232);
nand (n2285,n2236,n2232);
nand (n2286,n2228,n2236);
xor (n2287,n2288,n1489);
xor (n2288,n1475,n1479);
nor (n2289,n2290,n2294);
nand (n2290,n2291,n2292,n2293);
nand (n2291,n2264,n2273);
nand (n2292,n2277,n2273);
nand (n2293,n2264,n2277);
xor (n2294,n2295,n2302);
xor (n2295,n2296,n2298);
xor (n2296,n2297,n1473);
xor (n2297,n1454,n1458);
nand (n2298,n2299,n2300,n2301);
nand (n2299,n2279,n2283);
nand (n2300,n2287,n2283);
nand (n2301,n2279,n2287);
xor (n2302,n2303,n2308);
xor (n2303,n2304,n2306);
xor (n2304,n2305,n1423);
xor (n2305,n1414,n1418);
xor (n2306,n2307,n1438);
xor (n2307,n1432,n1436);
nand (n2308,n2309,n2310,n2311);
nand (n2309,n2266,n2270);
nand (n2310,n2271,n2270);
nand (n2311,n2266,n2271);
nor (n2312,n2313,n2328);
nor (n2313,n2314,n2318);
nand (n2314,n2315,n2316,n2317);
nand (n2315,n2296,n2298);
nand (n2316,n2302,n2298);
nand (n2317,n2296,n2302);
xor (n2318,n2319,n2326);
xor (n2319,n2320,n2322);
xor (n2320,n2321,n1430);
xor (n2321,n1410,n1412);
nand (n2322,n2323,n2324,n2325);
nand (n2323,n2304,n2306);
nand (n2324,n2308,n2306);
nand (n2325,n2304,n2308);
xor (n2326,n2327,n1452);
xor (n2327,n1447,n1449);
nor (n2328,n2329,n2333);
nand (n2329,n2330,n2331,n2332);
nand (n2330,n2320,n2322);
nand (n2331,n2326,n2322);
nand (n2332,n2320,n2326);
xor (n2333,n2334,n1445);
xor (n2334,n1320,n1371);
nor (n2335,n2336,n2458);
nor (n2336,n2337,n2434);
nor (n2337,n2338,n2431);
nor (n2338,n2339,n2407);
nand (n2339,n2340,n2379);
or (n2340,n2341,n2365,n2378);
and (n2341,n2342,n2351);
xor (n2342,n2343,n2347);
xnor (n2343,n2344,n558);
nor (n2344,n2345,n2346);
and (n2345,n455,n668);
and (n2346,n277,n670);
xnor (n2347,n2348,n300);
nor (n2348,n2349,n2350);
and (n2349,n653,n560);
and (n2350,n540,n556);
or (n2351,n2352,n2359,n2364);
and (n2352,n2353,n2355);
not (n2353,n2354);
nand (n2354,n696,n40);
xnor (n2355,n2356,n558);
nor (n2356,n2357,n2358);
and (n2357,n540,n668);
and (n2358,n455,n670);
and (n2359,n2355,n2360);
xnor (n2360,n2361,n300);
nor (n2361,n2362,n2363);
and (n2362,n657,n560);
and (n2363,n653,n556);
and (n2364,n2353,n2360);
and (n2365,n2351,n2366);
xor (n2366,n2367,n2374);
xor (n2367,n2368,n2370);
and (n2368,n46,n2369);
xnor (n2369,n2354,n46);
xnor (n2370,n2371,n42);
nor (n2371,n2372,n2373);
and (n2372,n659,n302);
and (n2373,n657,n298);
xnor (n2374,n2375,n46);
nor (n2375,n2376,n2377);
and (n2376,n696,n44);
and (n2377,n682,n40);
and (n2378,n2342,n2366);
xor (n2379,n2380,n2396);
xor (n2380,n2381,n2385);
or (n2381,n2382,n2383,n2384);
and (n2382,n2368,n2370);
and (n2383,n2370,n2374);
and (n2384,n2368,n2374);
xor (n2385,n2386,n2392);
xor (n2386,n2387,n2388);
and (n2387,n2343,n2347);
xnor (n2388,n2389,n42);
nor (n2389,n2390,n2391);
and (n2390,n657,n302);
and (n2391,n653,n298);
xnor (n2392,n2393,n46);
nor (n2393,n2394,n2395);
and (n2394,n682,n44);
and (n2395,n659,n40);
xor (n2396,n2397,n2403);
xor (n2397,n2398,n2399);
not (n2398,n2203);
xnor (n2399,n2400,n558);
nor (n2400,n2401,n2402);
and (n2401,n277,n668);
and (n2402,n203,n670);
xnor (n2403,n2404,n300);
nor (n2404,n2405,n2406);
and (n2405,n540,n560);
and (n2406,n455,n556);
nor (n2407,n2408,n2412);
or (n2408,n2409,n2410,n2411);
and (n2409,n2381,n2385);
and (n2410,n2385,n2396);
and (n2411,n2381,n2396);
xor (n2412,n2413,n2420);
xor (n2413,n2414,n2418);
or (n2414,n2415,n2416,n2417);
and (n2415,n2387,n2388);
and (n2416,n2388,n2392);
and (n2417,n2387,n2392);
xor (n2418,n2419,n2201);
xor (n2419,n2192,n2196);
xor (n2420,n2421,n2427);
xor (n2421,n2422,n2426);
xor (n2422,n2423,n56);
or (n2423,n2424,n2425);
and (n2424,n682,n50);
and (n2425,n696,n54);
xor (n2426,n2247,n2251);
or (n2427,n2428,n2429,n2430);
and (n2428,n2398,n2399);
and (n2429,n2399,n2403);
and (n2430,n2398,n2403);
not (n2431,n2432);
not (n2432,n2433);
and (n2433,n2408,n2412);
not (n2434,n2435);
nor (n2435,n2436,n2451);
nor (n2436,n2437,n2441);
nand (n2437,n2438,n2439,n2440);
nand (n2438,n2414,n2418);
nand (n2439,n2420,n2418);
nand (n2440,n2414,n2420);
xor (n2441,n2442,n2449);
xor (n2442,n2443,n2445);
xor (n2443,n2444,n2256);
xor (n2444,n2242,n2246);
nand (n2445,n2446,n2447,n2448);
nand (n2446,n2422,n2426);
nand (n2447,n2427,n2426);
nand (n2448,n2422,n2427);
xor (n2449,n2450,n2206);
xor (n2450,n2189,n2190);
nor (n2451,n2452,n2456);
nand (n2452,n2453,n2454,n2455);
nand (n2453,n2443,n2445);
nand (n2454,n2449,n2445);
nand (n2455,n2443,n2449);
xor (n2456,n2457,n2220);
xor (n2457,n2175,n2187);
not (n2458,n2459);
nor (n2459,n2460,n2462);
nor (n2460,n2461,n2451);
nand (n2461,n2437,n2441);
not (n2462,n2463);
nand (n2463,n2452,n2456);
not (n2464,n2465);
nor (n2465,n2466,n2473);
nor (n2466,n2467,n2472);
nor (n2467,n2468,n2470);
nor (n2468,n2469,n2289);
nand (n2469,n2173,n2262);
not (n2470,n2471);
nand (n2471,n2290,n2294);
not (n2472,n2312);
not (n2473,n2474);
nor (n2474,n2475,n2477);
nor (n2475,n2476,n2328);
nand (n2476,n2314,n2318);
not (n2477,n2478);
nand (n2478,n2329,n2333);
nand (n2479,n2480,n2484);
nor (n2480,n2481,n2170);
nand (n2481,n2482,n2435);
nor (n2482,n2483,n2407);
nor (n2483,n2340,n2379);
or (n2484,n2485,n2507);
and (n2485,n2486,n2488);
xor (n2486,n2487,n2366);
xor (n2487,n2342,n2351);
or (n2488,n2489,n2503,n2506);
and (n2489,n2490,n2499);
and (n2490,n2491,n2495);
xnor (n2491,n2492,n558);
nor (n2492,n2493,n2494);
and (n2493,n653,n668);
and (n2494,n540,n670);
xnor (n2495,n2496,n300);
nor (n2496,n2497,n2498);
and (n2497,n659,n560);
and (n2498,n657,n556);
xnor (n2499,n2500,n42);
nor (n2500,n2501,n2502);
and (n2501,n682,n302);
and (n2502,n659,n298);
and (n2503,n2499,n2504);
xor (n2504,n2505,n2360);
xor (n2505,n2353,n2355);
and (n2506,n2490,n2504);
and (n2507,n2508,n2509);
xor (n2508,n2486,n2488);
or (n2509,n2510,n2525);
and (n2510,n2511,n2523);
or (n2511,n2512,n2517,n2522);
and (n2512,n2513,n2514);
xor (n2513,n2491,n2495);
and (n2514,n42,n2515);
xnor (n2515,n2516,n42);
nand (n2516,n696,n298);
and (n2517,n2514,n2518);
xnor (n2518,n2519,n42);
nor (n2519,n2520,n2521);
and (n2520,n696,n302);
and (n2521,n682,n298);
and (n2522,n2513,n2518);
xor (n2523,n2524,n2504);
xor (n2524,n2490,n2499);
and (n2525,n2526,n2527);
xor (n2526,n2511,n2523);
or (n2527,n2528,n2544);
and (n2528,n2529,n2531);
xor (n2529,n2530,n2518);
xor (n2530,n2513,n2514);
or (n2531,n2532,n2538,n2543);
and (n2532,n2533,n2534);
not (n2533,n2516);
xnor (n2534,n2535,n558);
nor (n2535,n2536,n2537);
and (n2536,n657,n668);
and (n2537,n653,n670);
and (n2538,n2534,n2539);
xnor (n2539,n2540,n300);
nor (n2540,n2541,n2542);
and (n2541,n682,n560);
and (n2542,n659,n556);
and (n2543,n2533,n2539);
and (n2544,n2545,n2546);
xor (n2545,n2529,n2531);
or (n2546,n2547,n2558);
and (n2547,n2548,n2550);
xor (n2548,n2549,n2539);
xor (n2549,n2533,n2534);
and (n2550,n2551,n2554);
and (n2551,n300,n2552);
xnor (n2552,n2553,n300);
nand (n2553,n696,n556);
xnor (n2554,n2555,n558);
nor (n2555,n2556,n2557);
and (n2556,n659,n668);
and (n2557,n657,n670);
and (n2558,n2559,n2560);
xor (n2559,n2548,n2550);
or (n2560,n2561,n2567);
and (n2561,n2562,n2566);
xnor (n2562,n2563,n300);
nor (n2563,n2564,n2565);
and (n2564,n696,n560);
and (n2565,n682,n556);
xor (n2566,n2551,n2554);
and (n2567,n2568,n2569);
xor (n2568,n2562,n2566);
or (n2569,n2570,n2576);
and (n2570,n2571,n2575);
xnor (n2571,n2572,n558);
nor (n2572,n2573,n2574);
and (n2573,n682,n668);
and (n2574,n659,n670);
not (n2575,n2553);
and (n2576,n2577,n2578);
xor (n2577,n2571,n2575);
and (n2578,n2579,n2583);
xnor (n2579,n2580,n558);
nor (n2580,n2581,n2582);
and (n2581,n696,n668);
and (n2582,n682,n670);
and (n2583,n2584,n558);
xnor (n2584,n2585,n558);
nand (n2585,n696,n670);
not (n2586,n2587);
nand (n2587,n2588,n1608);
nor (n2588,n2589,n640);
nand (n2589,n2590,n1563);
nor (n2590,n2591,n1535);
nor (n2591,n1318,n1497);
not (n2592,n2593);
nor (n2593,n3,n322);
nand (n2594,n2595,n2664);
not (n2595,n2596);
nor (n2596,n2597,n2601);
nand (n2597,n2598,n2599,n2600);
nand (n2598,n324,n352);
nand (n2599,n386,n352);
nand (n2600,n324,n386);
xor (n2601,n2602,n2660);
xor (n2602,n2603,n2607);
nand (n2603,n2604,n2605,n2606);
nand (n2604,n326,n340);
nand (n2605,n348,n340);
nand (n2606,n326,n348);
xor (n2607,n2608,n2633);
xor (n2608,n2609,n2613);
nand (n2609,n2610,n2611,n2612);
nand (n2610,n356,n370);
nand (n2611,n374,n370);
nand (n2612,n356,n374);
xor (n2613,n2614,n2629);
xor (n2614,n2615,n2625);
xor (n2615,n2616,n2621);
xor (n2616,n328,n2617);
xor (n2617,n2618,n69);
or (n2618,n2619,n2620);
and (n2619,n39,n62);
and (n2620,n53,n67);
xor (n2621,n2622,n15);
or (n2622,n2623,n2624);
and (n2623,n61,n118);
and (n2624,n66,n121);
nand (n2625,n2626,n2627,n2628);
nand (n2626,n358,n362);
nand (n2627,n366,n362);
nand (n2628,n358,n366);
nand (n2629,n2630,n2631,n2632);
nand (n2630,n328,n332);
nand (n2631,n336,n332);
nand (n2632,n328,n336);
xor (n2633,n2634,n2655);
xor (n2634,n2635,n2645);
xor (n2635,n2636,n74);
xor (n2636,n2637,n2641);
xor (n2637,n2638,n31);
or (n2638,n2639,n2640);
and (n2639,n117,n25);
and (n2640,n12,n29);
xor (n2641,n2642,n74);
or (n2642,n2643,n2644);
and (n2643,n17,n159);
and (n2644,n24,n163);
xor (n2645,n2646,n2651);
xor (n2646,n2647,n329);
xor (n2647,n2648,n100);
or (n2648,n2649,n2650);
and (n2649,n83,n94);
and (n2650,n89,n98);
xor (n2651,n2652,n20);
or (n2652,n2653,n2654);
and (n2653,n97,n13);
and (n2654,n112,n18);
nand (n2655,n2656,n2658,n2659);
nand (n2656,n2657,n74);
xor (n2657,n341,n74);
nand (n2658,n344,n74);
nand (n2659,n2657,n344);
nand (n2660,n2661,n2662,n2663);
nand (n2661,n354,n378);
nand (n2662,n382,n378);
nand (n2663,n354,n382);
nand (n2664,n2597,n2601);
xor (n2665,n2666,n2840);
xor (n2666,n2667,n2763);
xor (n2667,n2668,n2729);
xor (n2668,n2669,n2702);
or (n2669,n2670,n2684,n2701);
and (n2670,n2671,n2674);
xor (n2671,n2672,n344);
xor (n2672,n2657,n2673);
not (n2673,n326);
or (n2674,n2675,n2677,n2683);
and (n2675,n2676,n127);
not (n2676,n8);
and (n2677,n127,n2678);
xor (n2678,n2679,n167);
or (n2679,n2680,n2681,n2682);
and (n2680,n130,n151);
not (n2681,n150);
and (n2682,n130,n155);
and (n2683,n2676,n2678);
and (n2684,n2674,n2685);
or (n2685,n2686,n2697,n2700);
and (n2686,n2687,n2692);
or (n2687,n2688,n2690,n2691);
and (n2688,n75,n2689);
not (n2689,n209);
and (n2690,n2689,n207);
and (n2691,n75,n207);
or (n2692,n2693,n2695,n2696);
and (n2693,n102,n2694);
not (n2694,n194);
and (n2695,n2694,n33);
and (n2696,n102,n33);
and (n2697,n2692,n2698);
xor (n2698,n2699,n141);
xor (n2699,n183,n187);
and (n2700,n2687,n2698);
and (n2701,n2671,n2685);
xor (n2702,n2703,n2720);
xor (n2703,n2704,n2711);
xor (n2704,n2705,n2710);
xor (n2705,n2625,n2706);
or (n2706,n2707,n2708,n2709);
and (n2707,n329,n332);
not (n2708,n2631);
and (n2709,n329,n336);
xor (n2710,n2616,n2647);
or (n2711,n2712,n2714,n2719);
and (n2712,n355,n2713);
and (n2713,n2679,n167);
and (n2714,n2713,n2715);
or (n2715,n2716,n2717,n2718);
not (n2716,n376);
and (n2717,n187,n141);
and (n2718,n183,n141);
and (n2719,n355,n2715);
xor (n2720,n2721,n2727);
xor (n2721,n2722,n2723);
not (n2722,n2610);
or (n2723,n2724,n2725,n2726);
and (n2724,n2657,n2673);
and (n2725,n2673,n344);
not (n2726,n2659);
xor (n2727,n2728,n2636);
xor (n2728,n2621,n2651);
or (n2729,n2730,n2759,n2762);
and (n2730,n2731,n2733);
xor (n2731,n2732,n2715);
xor (n2732,n355,n2713);
or (n2733,n2734,n2755,n2758);
and (n2734,n2735,n2753);
or (n2735,n2736,n2749,n2752);
and (n2736,n2737,n2741);
or (n2737,n2738,n2739,n2740);
and (n2738,n216,n245);
and (n2739,n245,n285);
and (n2740,n216,n285);
or (n2741,n2742,n2743,n2748);
and (n2742,n221,n248);
and (n2743,n248,n2744);
or (n2744,n2745,n2746,n2747);
and (n2745,n36,n279);
not (n2746,n283);
and (n2747,n36,n273);
and (n2748,n221,n2744);
and (n2749,n2741,n2750);
xor (n2750,n2751,n207);
xor (n2751,n75,n2689);
and (n2752,n2737,n2750);
xor (n2753,n2754,n2678);
xor (n2754,n2676,n127);
and (n2755,n2753,n2756);
xor (n2756,n2757,n2698);
xor (n2757,n2687,n2692);
and (n2758,n2735,n2756);
and (n2759,n2733,n2760);
xor (n2760,n2761,n2685);
xor (n2761,n2671,n2674);
and (n2762,n2731,n2760);
or (n2763,n2764,n2766);
xor (n2764,n2765,n2760);
xor (n2765,n2731,n2733);
or (n2766,n2767,n2790,n2839);
and (n2767,n2768,n2788);
or (n2768,n2769,n2784,n2787);
and (n2769,n2770,n2772);
xor (n2770,n2771,n33);
xor (n2771,n102,n2694);
or (n2772,n2773,n2780,n2783);
and (n2773,n243,n2774);
or (n2774,n2775,n2777,n2779);
and (n2775,n311,n2776);
not (n2776,n458);
and (n2777,n2776,n2778);
not (n2778,n446);
and (n2779,n311,n2778);
and (n2780,n2774,n2781);
xor (n2781,n2782,n285);
xor (n2782,n216,n245);
and (n2783,n243,n2781);
and (n2784,n2772,n2785);
xor (n2785,n2786,n2750);
xor (n2786,n2737,n2741);
and (n2787,n2770,n2785);
xor (n2788,n2789,n2756);
xor (n2789,n2735,n2753);
and (n2790,n2788,n2791);
or (n2791,n2792,n2803,n2838);
and (n2792,n2793,n2801);
or (n2793,n2794,n2797,n2800);
and (n2794,n2795,n401);
xor (n2795,n2796,n2744);
xor (n2796,n221,n248);
and (n2797,n401,n2798);
xor (n2798,n2799,n2781);
xor (n2799,n243,n2774);
and (n2800,n2795,n2798);
xor (n2801,n2802,n2785);
xor (n2802,n2770,n2772);
and (n2803,n2801,n2804);
or (n2804,n2805,n2834,n2837);
and (n2805,n2806,n2819);
or (n2806,n2807,n2817,n2818);
and (n2807,n2808,n488);
or (n2808,n2809,n2814,n2816);
and (n2809,n2810,n482);
or (n2810,n2811,n2812,n2813);
and (n2811,n294,n472);
not (n2812,n476);
and (n2813,n294,n477);
and (n2814,n482,n2815);
not (n2815,n485);
and (n2816,n2810,n2815);
not (n2817,n523);
and (n2818,n2808,n524);
or (n2819,n2820,n2827,n2833);
and (n2820,n2821,n2825);
or (n2821,n2822,n2823,n2824);
and (n2822,n295,n291);
not (n2823,n309);
and (n2824,n295,n305);
xor (n2825,n2826,n2778);
xor (n2826,n311,n2776);
and (n2827,n2825,n2828);
or (n2828,n2829,n2830,n2832);
and (n2829,n294,n565);
and (n2830,n565,n2831);
not (n2831,n2088);
and (n2832,n294,n2831);
and (n2833,n2821,n2828);
and (n2834,n2819,n2835);
xor (n2835,n2836,n2798);
xor (n2836,n2795,n401);
and (n2837,n2806,n2835);
and (n2838,n2793,n2804);
and (n2839,n2768,n2791);
and (n2840,n2841,n2842);
xnor (n2841,n2764,n2766);
or (n2842,n2843,n2928);
and (n2843,n2844,n2846);
xor (n2844,n2845,n2791);
xor (n2845,n2768,n2788);
or (n2846,n2847,n2849);
xor (n2847,n2848,n2804);
xor (n2848,n2793,n2801);
or (n2849,n2850,n2872,n2927);
and (n2850,n2851,n2870);
or (n2851,n2852,n2866,n2869);
and (n2852,n2853,n2855);
xor (n2853,n2854,n524);
xor (n2854,n2808,n488);
or (n2855,n2856,n2859,n2865);
and (n2856,n2857,n2091);
xor (n2857,n2858,n2815);
xor (n2858,n2810,n482);
and (n2859,n2091,n2860);
or (n2860,n2861,n2862,n2864);
not (n2861,n604);
and (n2862,n588,n2863);
not (n2863,n585);
and (n2864,n569,n2863);
and (n2865,n2857,n2860);
and (n2866,n2855,n2867);
xor (n2867,n2868,n2828);
xor (n2868,n2821,n2825);
and (n2869,n2853,n2867);
xor (n2870,n2871,n2835);
xor (n2871,n2806,n2819);
and (n2872,n2870,n2873);
or (n2873,n2874,n2889,n2926);
and (n2874,n2875,n2887);
or (n2875,n2876,n2883,n2886);
and (n2876,n2877,n2881);
or (n2877,n2878,n2879,n2880);
and (n2878,n536,n2061);
and (n2879,n2061,n2042);
and (n2880,n536,n2042);
xor (n2881,n2882,n2831);
xor (n2882,n294,n565);
and (n2883,n2881,n2884);
and (n2884,n2037,n2885);
not (n2885,n2035);
and (n2886,n2877,n2884);
xor (n2887,n2888,n2867);
xor (n2888,n2853,n2855);
and (n2889,n2887,n2890);
or (n2890,n2891,n2911,n2925);
and (n2891,n2892,n2909);
or (n2892,n2893,n2898,n2908);
and (n2893,n2894,n2064);
or (n2894,n2895,n2896,n2897);
and (n2895,n553,n544);
not (n2896,n543);
and (n2897,n553,n547);
and (n2898,n2064,n2899);
or (n2899,n2900,n2905,n2907);
and (n2900,n552,n2901);
or (n2901,n2902,n2903,n2904);
and (n2902,n552,n1865);
not (n2903,n1979);
and (n2904,n552,n1869);
and (n2905,n2901,n2906);
not (n2906,n1974);
and (n2907,n552,n2906);
and (n2908,n2894,n2899);
xor (n2909,n2910,n2860);
xor (n2910,n2857,n2091);
and (n2911,n2909,n2912);
or (n2912,n2913,n2917,n2924);
and (n2913,n2914,n2916);
xor (n2914,n2915,n2042);
xor (n2915,n536,n2061);
not (n2916,n2034);
and (n2917,n2916,n2918);
or (n2918,n2919,n2922,n2923);
and (n2919,n2920,n1980);
and (n2920,n1849,n2921);
not (n2921,n1863);
and (n2922,n1980,n2002);
and (n2923,n2920,n2002);
and (n2924,n2914,n2918);
and (n2925,n2892,n2912);
and (n2926,n2875,n2890);
and (n2927,n2851,n2873);
and (n2928,n2929,n2930);
xor (n2929,n2844,n2846);
and (n2930,n2931,n2932);
xnor (n2931,n2847,n2849);
or (n2932,n2933,n3137);
and (n2933,n2934,n2936);
xor (n2934,n2935,n2873);
xor (n2935,n2851,n2870);
or (n2936,n2937,n3012,n3136);
and (n2937,n2938,n3010);
or (n2938,n2939,n3006,n3009);
and (n2939,n2940,n2942);
xor (n2940,n2941,n2884);
xor (n2941,n2877,n2881);
or (n2942,n2943,n2977,n3005);
and (n2943,n2944,n2975);
or (n2944,n2945,n2963,n2974);
and (n2945,n2946,n2955);
and (n2946,n2947,n1889);
or (n2947,n2948,n2953,n2954);
and (n2948,n2949,n1759);
or (n2949,n2950,n2951,n2952);
and (n2950,n1828,n1624);
not (n2951,n1768);
and (n2952,n1828,n1628);
not (n2953,n1901);
and (n2954,n2949,n1763);
or (n2955,n2956,n2961,n2962);
and (n2956,n1929,n2957);
or (n2957,n2958,n2959,n2960);
and (n2958,n1828,n1748);
not (n2959,n1876);
and (n2960,n1828,n1753);
and (n2961,n2957,n1910);
and (n2962,n1929,n1910);
and (n2963,n2955,n2964);
or (n2964,n2965,n2971,n2973);
and (n2965,n2966,n2967);
not (n2966,n1848);
or (n2967,n2968,n2969,n2970);
and (n2968,n1632,n1824);
not (n2969,n1928);
and (n2970,n1632,n1829);
and (n2971,n2967,n2972);
not (n2972,n1905);
and (n2973,n2966,n2972);
and (n2974,n2946,n2964);
xor (n2975,n2976,n2899);
xor (n2976,n2894,n2064);
and (n2977,n2975,n2978);
or (n2978,n2979,n3001,n3004);
and (n2979,n2980,n2982);
xor (n2980,n2981,n2906);
xor (n2981,n552,n2901);
or (n2982,n2983,n2992,n3000);
and (n2983,n2984,n2991);
or (n2984,n2985,n2987,n2990);
and (n2985,n1808,n2986);
not (n2986,n1805);
and (n2987,n2986,n2988);
xor (n2988,n2989,n1753);
xor (n2989,n1828,n1748);
and (n2990,n1808,n2988);
xor (n2991,n2947,n1889);
and (n2992,n2991,n2993);
or (n2993,n2994,n2998,n2999);
and (n2994,n2995,n2996);
not (n2995,n1822);
xor (n2996,n2997,n1763);
xor (n2997,n2949,n1759);
and (n2998,n2996,n1782);
and (n2999,n2995,n1782);
and (n3000,n2984,n2993);
and (n3001,n2982,n3002);
xor (n3002,n3003,n2002);
xor (n3003,n2920,n1980);
and (n3004,n2980,n3002);
and (n3005,n2944,n2978);
and (n3006,n2942,n3007);
xor (n3007,n3008,n2912);
xor (n3008,n2892,n2909);
and (n3009,n2940,n3007);
xor (n3010,n3011,n2890);
xor (n3011,n2875,n2887);
and (n3012,n3010,n3013);
or (n3013,n3014,n3047,n3135);
and (n3014,n3015,n3045);
or (n3015,n3016,n3041,n3044);
and (n3016,n3017,n3019);
xor (n3017,n3018,n2918);
xor (n3018,n2914,n2916);
or (n3019,n3020,n3037,n3040);
and (n3020,n3021,n3023);
xor (n3021,n3022,n2964);
xor (n3022,n2946,n2955);
or (n3023,n3024,n3029,n3036);
and (n3024,n3025,n3027);
xor (n3025,n3026,n1910);
xor (n3026,n1929,n2957);
xor (n3027,n3028,n2972);
xor (n3028,n2966,n2967);
and (n3029,n3027,n3030);
and (n3030,n1773,n3031);
or (n3031,n3032,n3033,n3035);
not (n3032,n1779);
and (n3033,n1639,n3034);
not (n3034,n1622);
and (n3035,n1635,n3034);
and (n3036,n3025,n3030);
and (n3037,n3023,n3038);
xor (n3038,n3039,n3002);
xor (n3039,n2980,n2982);
and (n3040,n3021,n3038);
and (n3041,n3019,n3042);
xor (n3042,n3043,n2978);
xor (n3043,n2944,n2975);
and (n3044,n3017,n3042);
xor (n3045,n3046,n3007);
xor (n3046,n2940,n2942);
and (n3047,n3045,n3048);
or (n3048,n3049,n3106,n3134);
and (n3049,n3050,n3052);
xor (n3050,n3051,n3042);
xor (n3051,n3017,n3019);
or (n3052,n3053,n3085,n3105);
and (n3053,n3054,n3083);
or (n3054,n3055,n3068,n3082);
and (n3055,n3056,n3066);
or (n3056,n3057,n3064,n3065);
and (n3057,n3058,n3062);
or (n3058,n3059,n3060,n3061);
and (n3059,n1687,n1672);
and (n3060,n1672,n1655);
and (n3061,n1687,n1655);
xor (n3062,n3063,n2988);
xor (n3063,n1808,n2986);
and (n3064,n3062,n1833);
and (n3065,n3058,n1833);
xor (n3066,n3067,n2993);
xor (n3067,n2984,n2991);
and (n3068,n3066,n3069);
or (n3069,n3070,n3079,n3081);
and (n3070,n3071,n3077);
or (n3071,n3072,n3073,n3076);
and (n3072,n1677,n1671);
and (n3073,n1671,n3074);
xor (n3074,n3075,n1655);
xor (n3075,n1687,n1672);
and (n3076,n1677,n3074);
xor (n3077,n3078,n1782);
xor (n3078,n2995,n2996);
and (n3079,n3077,n3080);
xor (n3080,n1773,n3031);
and (n3081,n3071,n3080);
and (n3082,n3056,n3069);
xor (n3083,n3084,n3038);
xor (n3084,n3021,n3023);
and (n3085,n3083,n3086);
or (n3086,n3087,n3101,n3104);
and (n3087,n3088,n3090);
xor (n3088,n3089,n3030);
xor (n3089,n3025,n3027);
or (n3090,n3091,n3099,n3100);
and (n3091,n3092,n3094);
xor (n3092,n3093,n1833);
xor (n3093,n3058,n3062);
or (n3094,n3095,n3096,n3098);
not (n3095,n1732);
and (n3096,n1647,n3097);
not (n3097,n1620);
and (n3098,n1643,n3097);
and (n3099,n3094,n1734);
and (n3100,n3092,n1734);
and (n3101,n3090,n3102);
xor (n3102,n3103,n3069);
xor (n3103,n3056,n3066);
and (n3104,n3088,n3102);
and (n3105,n3054,n3086);
and (n3106,n3052,n3107);
or (n3107,n3108,n3110);
xor (n3108,n3109,n3086);
xor (n3109,n3054,n3083);
or (n3110,n3111,n3127,n3133);
and (n3111,n3112,n3125);
or (n3112,n3113,n3121,n3124);
and (n3113,n3114,n3116);
xor (n3114,n3115,n3080);
xor (n3115,n3071,n3077);
or (n3116,n3117,n3119,n3120);
and (n3117,n3118,n1719);
not (n3118,n1618);
not (n3119,n1726);
and (n3120,n3118,n1651);
and (n3121,n3116,n3122);
xor (n3122,n3123,n1734);
xor (n3123,n3092,n3094);
and (n3124,n3114,n3122);
xor (n3125,n3126,n3102);
xor (n3126,n3088,n3090);
and (n3127,n3125,n3128);
or (n3128,n3129,n3131);
or (n3129,n1612,n3130);
not (n3130,n1616);
xor (n3131,n3132,n3122);
xor (n3132,n3114,n3116);
and (n3133,n3112,n3128);
and (n3134,n3050,n3107);
and (n3135,n3015,n3048);
and (n3136,n2938,n3013);
and (n3137,n3138,n3139);
xor (n3138,n2934,n2936);
and (n3139,n3140,n3142);
xor (n3140,n3141,n3013);
xor (n3141,n2938,n3010);
or (n3142,n3143,n3145);
xor (n3143,n3144,n3048);
xor (n3144,n3015,n3045);
and (n3145,n3146,n3147);
not (n3146,n3143);
and (n3147,n3148,n3150);
xor (n3148,n3149,n3107);
xor (n3149,n3050,n3052);
and (n3150,n3151,n3152);
xnor (n3151,n3108,n3110);
and (n3152,n3153,n3155);
xor (n3153,n3154,n3128);
xor (n3154,n3112,n3125);
and (n3155,n3156,n3157);
xnor (n3156,n3129,n3131);
and (n3157,n3158,n3161);
not (n3158,n3159);
nand (n3159,n3160,n2141);
not (n3160,n1611);
nand (n3161,n638,n3162);
nand (n3162,n2588,n2167);
endmodule
