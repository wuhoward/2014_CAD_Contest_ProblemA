module top (out,n15,n19,n21,n23,n28,n29,n34,n39,n52
        ,n53,n60,n61,n71,n78,n79,n82,n88,n89,n98
        ,n107,n118,n123,n135,n143,n166,n172,n177,n188,n196
        ,n204,n228,n244,n273,n509,n540,n599,n623,n724,n728
        ,n790,n794,n826,n923,n927,n934);
output out;
input n15;
input n19;
input n21;
input n23;
input n28;
input n29;
input n34;
input n39;
input n52;
input n53;
input n60;
input n61;
input n71;
input n78;
input n79;
input n82;
input n88;
input n89;
input n98;
input n107;
input n118;
input n123;
input n135;
input n143;
input n166;
input n172;
input n177;
input n188;
input n196;
input n204;
input n228;
input n244;
input n273;
input n509;
input n540;
input n599;
input n623;
input n724;
input n728;
input n790;
input n794;
input n826;
input n923;
input n927;
input n934;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n16;
wire n17;
wire n18;
wire n20;
wire n22;
wire n24;
wire n25;
wire n26;
wire n27;
wire n30;
wire n31;
wire n32;
wire n33;
wire n35;
wire n36;
wire n37;
wire n38;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n80;
wire n81;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n119;
wire n120;
wire n121;
wire n122;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n173;
wire n174;
wire n175;
wire n176;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n725;
wire n726;
wire n727;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n791;
wire n792;
wire n793;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n924;
wire n925;
wire n926;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
xor (out,n0,n946);
nand (n0,n1,n945);
or (n1,n2,n849);
nand (n2,n3,n843);
or (n3,n4,n486);
not (n4,n5);
and (n5,n6,n443);
nand (n6,n7,n393);
not (n7,n8);
xor (n8,n9,n294);
xor (n9,n10,n156);
xor (n10,n11,n110);
xor (n11,n12,n43);
or (n12,n13,n42);
and (n13,n14,n24);
xor (n14,n15,n16);
and (n16,n17,n23);
nand (n17,n18,n22);
or (n18,n19,n20);
not (n20,n21);
nand (n22,n20,n19);
nand (n24,n25,n36);
or (n25,n26,n30);
nand (n26,n27,n29);
not (n27,n28);
not (n30,n31);
nand (n31,n32,n35);
or (n32,n33,n29);
not (n33,n34);
nand (n35,n29,n33);
nand (n36,n37,n28);
nand (n37,n38,n41);
or (n38,n39,n40);
not (n40,n29);
nand (n41,n40,n39);
and (n42,n15,n16);
or (n43,n44,n109);
and (n44,n45,n83);
xor (n45,n46,n73);
nand (n46,n47,n64);
or (n47,n48,n55);
not (n48,n49);
nand (n49,n50,n54);
or (n50,n51,n53);
not (n51,n52);
nand (n54,n53,n51);
not (n55,n56);
nand (n56,n57,n62);
nand (n57,n58,n61);
nor (n58,n59,n53);
not (n59,n60);
nand (n62,n63,n53,n59);
not (n63,n61);
nand (n64,n65,n68);
nor (n65,n66,n67);
and (n66,n59,n63);
and (n67,n60,n61);
nand (n68,n69,n72);
or (n69,n70,n53);
not (n70,n71);
nand (n72,n70,n53);
nor (n73,n74,n81);
nand (n74,n75,n21);
or (n75,n76,n80);
nor (n76,n77,n79);
and (n77,n23,n78);
nor (n80,n23,n78);
not (n81,n82);
nand (n83,n84,n100);
or (n84,n85,n93);
not (n85,n86);
nor (n86,n87,n90);
and (n87,n88,n89);
and (n90,n91,n92);
not (n91,n88);
not (n92,n89);
not (n93,n94);
nand (n94,n95,n99);
nand (n95,n96,n97,n89);
not (n96,n53);
not (n97,n98);
nand (n99,n92,n98,n53);
nand (n100,n101,n104);
nand (n101,n102,n103);
or (n102,n98,n96);
nand (n103,n96,n98);
nand (n104,n105,n108);
or (n105,n106,n89);
not (n106,n107);
nand (n108,n89,n106);
and (n109,n46,n73);
xor (n110,n111,n137);
xor (n111,n112,n120);
nand (n112,n113,n115);
or (n113,n26,n114);
not (n114,n37);
nand (n115,n116,n28);
nand (n116,n117,n119);
or (n117,n118,n40);
nand (n119,n40,n118);
nand (n120,n121,n136);
or (n121,n122,n124);
not (n122,n123);
not (n124,n125);
nand (n125,n126,n135);
or (n126,n127,n131);
not (n127,n128);
nand (n128,n129,n130);
not (n129,n23);
not (n130,n19);
not (n131,n132);
nand (n132,n133,n20);
not (n133,n134);
and (n134,n23,n19);
nand (n136,n124,n122);
nand (n137,n138,n146);
or (n138,n139,n145);
not (n139,n140);
nand (n140,n141,n144);
or (n141,n135,n142);
not (n142,n143);
nand (n144,n142,n135);
not (n145,n17);
nand (n146,n147,n153);
nand (n147,n148,n152);
or (n148,n149,n151);
not (n149,n150);
nor (n150,n21,n19);
not (n151,n135);
nand (n152,n151,n19,n21);
nand (n153,n154,n155);
or (n154,n151,n23);
nand (n155,n23,n151);
or (n156,n157,n293);
and (n157,n158,n231);
xor (n158,n159,n230);
xor (n159,n160,n207);
xor (n160,n161,n182);
nand (n161,n162,n174);
or (n162,n163,n168);
not (n163,n164);
nand (n164,n165,n167);
or (n165,n166,n63);
nand (n167,n63,n166);
not (n168,n169);
nand (n169,n170,n173);
nand (n170,n61,n40,n171);
not (n171,n172);
nand (n173,n63,n29,n172);
nand (n174,n175,n179);
nand (n175,n176,n178);
or (n176,n177,n63);
nand (n178,n63,n177);
nand (n179,n180,n181);
or (n180,n40,n172);
nand (n181,n40,n172);
nand (n182,n183,n198);
or (n183,n184,n190);
not (n184,n185);
nand (n185,n186,n189);
or (n186,n79,n187);
not (n187,n188);
nand (n189,n187,n79);
not (n190,n191);
nand (n191,n192,n197);
or (n192,n193,n92);
not (n193,n194);
nor (n194,n79,n195);
not (n195,n196);
nand (n197,n92,n79,n195);
nand (n198,n199,n202);
nand (n199,n200,n201);
or (n200,n195,n89);
nand (n201,n89,n195);
nand (n202,n203,n206);
or (n203,n204,n205);
not (n205,n79);
nand (n206,n205,n204);
nand (n207,n208,n224);
or (n208,n209,n213);
not (n209,n210);
nor (n210,n211,n212);
and (n211,n20,n142);
and (n212,n143,n21);
nand (n213,n214,n220);
or (n214,n215,n217);
not (n215,n216);
nand (n216,n20,n78);
not (n217,n218);
nand (n218,n21,n219);
not (n219,n78);
not (n220,n221);
nand (n221,n222,n223);
or (n222,n78,n205);
nand (n223,n205,n78);
nand (n224,n225,n221);
nor (n225,n226,n229);
and (n226,n20,n227);
not (n227,n228);
and (n229,n228,n21);
xor (n230,n45,n83);
or (n231,n232,n292);
and (n232,n233,n258);
xor (n233,n234,n241);
nand (n234,n235,n240);
or (n235,n236,n213);
not (n236,n237);
nand (n237,n238,n239);
or (n238,n23,n20);
or (n239,n129,n21);
nand (n240,n210,n221);
or (n241,n242,n257);
and (n242,n243,n246);
xor (n243,n244,n245);
and (n245,n221,n23);
nand (n246,n247,n252);
or (n247,n26,n248);
not (n248,n249);
nand (n249,n250,n251);
or (n250,n166,n40);
nand (n251,n40,n166);
nand (n252,n253,n28);
nand (n253,n254,n256);
or (n254,n255,n29);
not (n255,n177);
nand (n256,n29,n255);
and (n257,n244,n245);
or (n258,n259,n291);
and (n259,n260,n280);
xor (n260,n261,n272);
nand (n261,n262,n268);
or (n262,n263,n267);
not (n263,n264);
nand (n264,n265,n266);
or (n265,n106,n53);
nand (n266,n53,n106);
not (n267,n65);
nand (n268,n269,n56);
nand (n269,n270,n271);
or (n270,n91,n53);
nand (n271,n53,n91);
and (n272,n273,n274);
nor (n274,n275,n205);
and (n275,n276,n279);
nand (n276,n277,n92);
not (n277,n278);
and (n278,n23,n196);
nand (n279,n129,n195);
nand (n280,n281,n286);
or (n281,n93,n282);
not (n282,n283);
nor (n283,n284,n285);
and (n284,n187,n92);
and (n285,n188,n89);
nand (n286,n101,n287);
nor (n287,n288,n290);
and (n288,n289,n92);
not (n289,n204);
and (n290,n204,n89);
and (n291,n261,n272);
and (n292,n234,n241);
and (n293,n159,n230);
xor (n294,n295,n374);
xor (n295,n296,n327);
xor (n296,n297,n320);
xor (n297,n298,n313);
nand (n298,n299,n306,n309,n311);
nand (n299,n300,n302);
not (n300,n301);
nand (n301,n63,n60);
nand (n302,n303,n305);
or (n303,n304,n53);
not (n304,n166);
nand (n305,n304,n53);
nand (n306,n307,n302);
not (n307,n308);
nand (n308,n59,n61);
nand (n309,n310,n68);
not (n310,n57);
nand (n311,n312,n68);
not (n312,n62);
nand (n313,n314,n316);
or (n314,n315,n93);
not (n315,n104);
nand (n316,n317,n101);
nand (n317,n318,n319);
or (n318,n51,n89);
nand (n319,n89,n51);
nand (n320,n321,n323);
or (n321,n322,n168);
not (n322,n175);
nand (n323,n179,n324);
nand (n324,n325,n326);
or (n325,n33,n61);
nand (n326,n61,n33);
or (n327,n328,n373);
and (n328,n329,n359);
xor (n329,n330,n358);
or (n330,n331,n357);
and (n331,n332,n350);
xor (n332,n333,n338);
nand (n333,n334,n335,n336);
nand (n334,n101,n86);
nand (n335,n53,n92,n204,n98);
nand (n336,n337,n96,n89);
nor (n337,n204,n98);
nand (n338,n339,n344,n346,n348);
nand (n339,n340,n341);
not (n340,n173);
nand (n341,n342,n343);
or (n342,n71,n63);
nand (n343,n63,n71);
nand (n344,n341,n345);
not (n345,n170);
nand (n346,n164,n347);
not (n347,n181);
nand (n348,n164,n349);
not (n349,n180);
nand (n350,n351,n356);
or (n351,n352,n190);
not (n352,n353);
nand (n353,n354,n355);
or (n354,n79,n227);
nand (n355,n227,n79);
nand (n356,n199,n185);
and (n357,n333,n338);
xor (n358,n14,n24);
or (n359,n360,n372);
and (n360,n361,n369);
xor (n361,n362,n366);
nand (n362,n363,n365);
or (n363,n26,n364);
not (n364,n253);
nand (n365,n31,n28);
nand (n366,n367,n368);
or (n367,n82,n74);
nand (n368,n74,n82);
nand (n369,n370,n371);
or (n370,n263,n55);
nand (n371,n65,n49);
and (n372,n362,n366);
and (n373,n330,n358);
xor (n374,n375,n390);
xor (n375,n376,n383);
nand (n376,n377,n379);
or (n377,n378,n190);
not (n378,n202);
nand (n379,n199,n380);
nand (n380,n381,n382);
or (n381,n91,n79);
nand (n382,n79,n91);
nand (n383,n384,n386);
or (n384,n385,n213);
not (n385,n225);
nand (n386,n387,n221);
nor (n387,n388,n389);
and (n388,n20,n187);
and (n389,n188,n21);
or (n390,n391,n392);
and (n391,n160,n207);
and (n392,n161,n182);
not (n393,n394);
or (n394,n395,n442);
and (n395,n396,n399);
xor (n396,n397,n398);
xor (n397,n329,n359);
xor (n398,n158,n231);
or (n399,n400,n441);
and (n400,n401,n404);
xor (n401,n402,n403);
xor (n402,n332,n350);
xor (n403,n361,n369);
or (n404,n405,n440);
and (n405,n406,n421);
xor (n406,n407,n414);
nand (n407,n408,n413);
or (n408,n409,n190);
not (n409,n410);
nand (n410,n411,n412);
or (n411,n143,n205);
nand (n412,n143,n205);
nand (n413,n199,n353);
nand (n414,n415,n420);
or (n415,n168,n416);
not (n416,n417);
nand (n417,n418,n419);
or (n418,n51,n61);
nand (n419,n61,n51);
nand (n420,n179,n341);
or (n421,n422,n439);
and (n422,n423,n432);
xor (n423,n424,n431);
nand (n424,n425,n430);
or (n425,n26,n426);
not (n426,n427);
nand (n427,n428,n429);
or (n428,n70,n29);
nand (n429,n29,n70);
nand (n430,n249,n28);
xor (n431,n273,n274);
nand (n432,n433,n438);
or (n433,n434,n55);
not (n434,n435);
nand (n435,n436,n437);
or (n436,n204,n96);
nand (n437,n96,n204);
nand (n438,n65,n269);
and (n439,n424,n431);
and (n440,n407,n414);
and (n441,n402,n403);
and (n442,n397,n398);
nand (n443,n444,n446);
not (n444,n445);
xor (n445,n396,n399);
not (n446,n447);
or (n447,n448,n485);
and (n448,n449,n484);
xor (n449,n450,n483);
or (n450,n451,n482);
and (n451,n452,n481);
xor (n452,n453,n480);
or (n453,n454,n479);
and (n454,n455,n472);
xor (n455,n456,n463);
nand (n456,n457,n462);
or (n457,n458,n93);
not (n458,n459);
nand (n459,n460,n461);
or (n460,n227,n89);
nand (n461,n89,n227);
nand (n462,n101,n283);
nand (n463,n464,n466);
or (n464,n465,n409);
not (n465,n199);
nand (n466,n465,n467,n470);
nand (n467,n468,n469);
or (n468,n205,n23);
nand (n469,n23,n205);
nand (n470,n193,n471);
nand (n471,n79,n195);
nand (n472,n473,n478);
or (n473,n474,n168);
not (n474,n475);
nand (n475,n476,n477);
or (n476,n106,n61);
nand (n477,n61,n106);
nand (n478,n417,n179);
and (n479,n456,n463);
xor (n480,n243,n246);
xor (n481,n260,n280);
and (n482,n453,n480);
xor (n483,n233,n258);
xor (n484,n401,n404);
and (n485,n450,n483);
not (n486,n487);
nand (n487,n488,n672);
or (n488,n489,n668);
nor (n489,n490,n661);
and (n490,n491,n648);
and (n491,n492,n612);
nand (n492,n493,n574);
not (n493,n494);
xor (n494,n495,n551);
xor (n495,n496,n497);
xor (n496,n455,n472);
or (n497,n498,n550);
and (n498,n499,n518);
xor (n499,n500,n507);
nand (n500,n501,n506);
or (n501,n502,n168);
not (n502,n503);
nor (n503,n504,n505);
and (n504,n88,n61);
and (n505,n91,n63);
nand (n506,n179,n475);
xor (n507,n508,n511);
xor (n508,n509,n510);
and (n510,n199,n23);
nand (n511,n512,n517);
or (n512,n26,n513);
not (n513,n514);
nand (n514,n515,n516);
or (n515,n52,n40);
nand (n516,n40,n52);
nand (n517,n427,n28);
or (n518,n519,n549);
and (n519,n520,n538);
xor (n520,n521,n528);
nand (n521,n522,n527);
or (n522,n26,n523);
not (n523,n524);
nand (n524,n525,n526);
or (n525,n106,n29);
nand (n526,n29,n106);
nand (n527,n514,n28);
nand (n528,n529,n534);
or (n529,n530,n55);
not (n530,n531);
nand (n531,n532,n533);
or (n532,n227,n53);
nand (n533,n53,n227);
nand (n534,n65,n535);
nand (n535,n536,n537);
or (n536,n53,n187);
nand (n537,n53,n187);
nand (n538,n539,n548);
or (n539,n540,n541);
not (n541,n542);
nor (n542,n543,n92);
and (n543,n544,n547);
nand (n544,n545,n96);
not (n545,n546);
and (n546,n23,n98);
nand (n547,n129,n97);
nand (n548,n541,n540);
and (n549,n521,n528);
and (n550,n500,n507);
xor (n551,n552,n573);
xor (n552,n553,n556);
or (n553,n554,n555);
and (n554,n508,n511);
and (n555,n509,n510);
or (n556,n557,n572);
and (n557,n558,n570);
xor (n558,n559,n563);
nand (n559,n560,n562);
or (n560,n561,n55);
not (n561,n535);
nand (n562,n65,n435);
nand (n563,n564,n569);
or (n564,n565,n93);
not (n565,n566);
nand (n566,n567,n568);
or (n567,n89,n142);
nand (n568,n89,n142);
nand (n569,n101,n459);
nor (n570,n541,n571);
not (n571,n540);
and (n572,n559,n563);
xor (n573,n423,n432);
not (n574,n575);
or (n575,n576,n611);
and (n576,n577,n610);
xor (n577,n578,n579);
xor (n578,n558,n570);
or (n579,n580,n609);
and (n580,n581,n596);
xor (n581,n582,n589);
nand (n582,n583,n588);
or (n583,n584,n93);
not (n584,n585);
nand (n585,n586,n587);
or (n586,n92,n23);
or (n587,n129,n89);
nand (n588,n101,n566);
nand (n589,n590,n595);
or (n590,n591,n168);
not (n591,n592);
nor (n592,n593,n594);
and (n593,n204,n61);
and (n594,n289,n63);
nand (n595,n179,n503);
or (n596,n597,n608);
and (n597,n598,n601);
xor (n598,n599,n600);
and (n600,n101,n23);
nand (n601,n602,n607);
or (n602,n603,n55);
not (n603,n604);
nand (n604,n605,n606);
or (n605,n142,n53);
nand (n606,n53,n142);
nand (n607,n65,n531);
and (n608,n599,n600);
and (n609,n582,n589);
xor (n610,n499,n518);
and (n611,n578,n579);
nand (n612,n613,n614);
nand (n613,n494,n575);
nand (n614,n615,n616);
xor (n615,n577,n610);
or (n616,n617,n647);
and (n617,n618,n646);
xor (n618,n619,n645);
or (n619,n620,n644);
and (n620,n621,n637);
xor (n621,n622,n630);
and (n622,n623,n624);
nor (n624,n625,n96);
and (n625,n626,n629);
nand (n626,n627,n63);
not (n627,n628);
and (n628,n23,n60);
nand (n629,n59,n129);
nand (n630,n631,n636);
or (n631,n26,n632);
not (n632,n633);
nand (n633,n634,n635);
or (n634,n88,n40);
nand (n635,n40,n88);
nand (n636,n524,n28);
nand (n637,n638,n643);
or (n638,n639,n168);
not (n639,n640);
nor (n640,n641,n642);
and (n641,n188,n61);
and (n642,n187,n63);
nand (n643,n179,n592);
and (n644,n622,n630);
xor (n645,n520,n538);
xor (n646,n581,n596);
and (n647,n619,n645);
nand (n648,n649,n657);
not (n649,n650);
xor (n650,n651,n654);
xor (n651,n652,n653);
xor (n652,n406,n421);
xor (n653,n452,n481);
or (n654,n655,n656);
and (n655,n552,n573);
and (n656,n553,n556);
not (n657,n658);
or (n658,n659,n660);
and (n659,n495,n551);
and (n660,n496,n497);
nand (n661,n662,n667);
nand (n662,n663,n664);
xor (n663,n449,n484);
or (n664,n665,n666);
and (n665,n651,n654);
and (n666,n652,n653);
nand (n667,n650,n658);
not (n668,n669);
nand (n669,n670,n671);
not (n670,n663);
not (n671,n664);
nand (n672,n673,n839,n669,n648);
nand (n673,n674,n838);
or (n674,n675,n703);
not (n675,n676);
or (n676,n677,n678);
xor (n677,n618,n646);
or (n678,n679,n702);
and (n679,n680,n701);
xor (n680,n681,n682);
xor (n681,n598,n601);
or (n682,n683,n700);
and (n683,n684,n693);
xor (n684,n685,n692);
nand (n685,n686,n691);
or (n686,n687,n55);
not (n687,n688);
nand (n688,n689,n690);
or (n689,n53,n129);
nand (n690,n129,n53);
nand (n691,n604,n65);
xor (n692,n623,n624);
nand (n693,n694,n699);
or (n694,n26,n695);
not (n695,n696);
nand (n696,n697,n698);
or (n697,n204,n40);
nand (n698,n40,n204);
nand (n699,n633,n28);
and (n700,n685,n692);
xor (n701,n621,n637);
and (n702,n681,n682);
not (n703,n704);
nand (n704,n705,n837);
or (n705,n706,n737);
not (n706,n707);
nand (n707,n708,n710);
not (n708,n709);
xor (n709,n680,n701);
not (n710,n711);
or (n711,n712,n736);
and (n712,n713,n735);
xor (n713,n714,n721);
nand (n714,n715,n720);
or (n715,n716,n168);
not (n716,n717);
nand (n717,n718,n719);
or (n718,n228,n63);
nand (n719,n63,n228);
nand (n720,n179,n640);
or (n721,n722,n734);
and (n722,n723,n726);
xor (n723,n724,n725);
and (n725,n65,n23);
nor (n726,n727,n729);
not (n727,n728);
nand (n729,n730,n61);
or (n730,n731,n733);
nor (n731,n732,n29);
and (n732,n23,n172);
nor (n733,n23,n172);
and (n734,n724,n725);
xor (n735,n684,n693);
and (n736,n714,n721);
not (n737,n738);
or (n738,n739,n836);
and (n739,n740,n760);
xor (n740,n741,n759);
or (n741,n742,n758);
and (n742,n743,n757);
xor (n743,n744,n751);
nand (n744,n745,n746);
or (n745,n27,n695);
nand (n746,n747,n748);
not (n747,n26);
nand (n748,n749,n750);
or (n749,n188,n40);
nand (n750,n40,n188);
nand (n751,n752,n756);
nand (n752,n169,n753);
nand (n753,n754,n755);
or (n754,n143,n63);
nand (n755,n63,n143);
nand (n756,n717,n179);
xor (n757,n723,n726);
and (n758,n744,n751);
xor (n759,n713,n735);
nand (n760,n761,n835);
or (n761,n762,n830);
nor (n762,n763,n829);
and (n763,n764,n799);
nand (n764,n765,n786);
not (n765,n766);
xor (n766,n767,n779);
xor (n767,n768,n775);
nand (n768,n769,n771);
or (n769,n27,n770);
not (n770,n748);
nand (n771,n772,n747);
nand (n772,n773,n774);
or (n773,n228,n40);
nand (n774,n40,n228);
nand (n775,n776,n778);
or (n776,n727,n777);
not (n777,n729);
nand (n778,n727,n777);
nand (n779,n780,n785);
or (n780,n781,n168);
not (n781,n782);
nand (n782,n783,n784);
or (n783,n63,n23);
nand (n784,n23,n63);
nand (n785,n179,n753);
not (n786,n787);
or (n787,n788,n798);
and (n788,n789,n792);
xor (n789,n790,n791);
and (n791,n179,n23);
nor (n792,n793,n795);
not (n793,n794);
nand (n795,n796,n29);
not (n796,n797);
and (n797,n23,n28);
and (n798,n790,n791);
nand (n799,n800,n828);
or (n800,n801,n811);
nor (n801,n802,n803);
xor (n802,n789,n792);
nand (n803,n804,n809);
or (n804,n805,n26);
not (n805,n806);
nor (n806,n807,n808);
and (n807,n142,n40);
and (n808,n143,n29);
or (n809,n810,n27);
not (n810,n772);
nor (n811,n812,n827);
and (n812,n813,n825);
nand (n813,n814,n818);
nor (n814,n815,n817);
and (n815,n816,n793);
not (n816,n795);
and (n817,n795,n794);
not (n818,n819);
nand (n819,n820,n821);
or (n820,n27,n805);
nand (n821,n822,n747);
nand (n822,n823,n824);
or (n823,n23,n40);
nand (n824,n40,n23);
and (n825,n797,n826);
nor (n827,n814,n818);
nand (n828,n802,n803);
nor (n829,n765,n786);
nor (n830,n831,n832);
xor (n831,n743,n757);
or (n832,n833,n834);
and (n833,n767,n779);
and (n834,n768,n775);
nand (n835,n831,n832);
and (n836,n741,n759);
nand (n837,n709,n711);
nand (n838,n677,n678);
and (n839,n492,n840);
nand (n840,n841,n842);
not (n841,n615);
not (n842,n616);
nand (n843,n844,n6);
or (n844,n845,n847);
not (n845,n846);
nand (n846,n445,n447);
not (n847,n848);
nand (n848,n8,n394);
nand (n849,n850,n944);
not (n850,n851);
nor (n851,n852,n940);
not (n852,n853);
xor (n853,n854,n904);
xor (n854,n855,n901);
xor (n855,n856,n878);
xor (n856,n857,n860);
or (n857,n858,n859);
and (n858,n111,n137);
and (n859,n112,n120);
xor (n860,n861,n871);
xor (n861,n862,n863);
nor (n862,n125,n122);
nand (n863,n864,n866);
or (n864,n865,n168);
not (n865,n324);
nand (n866,n867,n179);
nand (n867,n868,n870);
or (n868,n869,n61);
not (n869,n39);
nand (n870,n61,n869);
nand (n871,n872,n874);
or (n872,n873,n190);
not (n873,n380);
nand (n874,n875,n199);
nand (n875,n876,n877);
or (n876,n106,n79);
nand (n877,n79,n106);
xor (n878,n879,n894);
xor (n879,n880,n887);
nand (n880,n881,n883);
or (n881,n882,n139);
not (n882,n147);
nand (n883,n17,n884);
nand (n884,n885,n886);
or (n885,n135,n227);
nand (n886,n227,n135);
nand (n887,n888,n890);
or (n888,n55,n889);
not (n889,n302);
nand (n890,n65,n891);
nand (n891,n892,n893);
or (n892,n177,n96);
or (n893,n53,n255);
nand (n894,n895,n897);
or (n895,n896,n93);
not (n896,n317);
nand (n897,n101,n898);
nand (n898,n899,n900);
or (n899,n70,n89);
or (n900,n92,n71);
or (n901,n902,n903);
and (n902,n295,n374);
and (n903,n296,n327);
xor (n904,n905,n937);
xor (n905,n906,n909);
or (n906,n907,n908);
and (n907,n375,n390);
and (n908,n376,n383);
xor (n909,n910,n921);
xor (n910,n911,n918);
nand (n911,n912,n914);
or (n912,n913,n213);
not (n913,n387);
nand (n914,n915,n221);
nand (n915,n916,n917);
or (n916,n20,n204);
or (n917,n289,n21);
or (n918,n919,n920);
and (n919,n297,n320);
and (n920,n298,n313);
xor (n921,n922,n928);
xor (n922,n923,n924);
nor (n924,n129,n925);
not (n925,n926);
xor (n926,n135,n927);
nand (n928,n929,n936);
or (n929,n27,n930);
not (n930,n931);
nand (n931,n932,n935);
or (n932,n933,n29);
not (n933,n934);
nand (n935,n29,n933);
nand (n936,n747,n116);
or (n937,n938,n939);
and (n938,n11,n110);
and (n939,n12,n43);
not (n940,n941);
or (n941,n942,n943);
and (n942,n9,n294);
and (n943,n10,n156);
nand (n944,n852,n940);
nand (n945,n2,n849);
xor (n946,n947,n1481);
xor (n947,n948,n923);
xor (n948,n949,n1480);
xor (n949,n950,n1477);
xor (n950,n951,n1476);
xor (n951,n952,n1468);
xor (n952,n953,n1467);
xor (n953,n954,n1454);
xor (n954,n955,n389);
xor (n955,n956,n1434);
xor (n956,n957,n1433);
xor (n957,n958,n1406);
xor (n958,n959,n1405);
xor (n959,n960,n1373);
xor (n960,n961,n1372);
xor (n961,n962,n1336);
xor (n962,n963,n1335);
xor (n963,n964,n1291);
xor (n964,n965,n1290);
xor (n965,n966,n1239);
xor (n966,n967,n1238);
xor (n967,n968,n1182);
xor (n968,n969,n1181);
xor (n969,n970,n1121);
xor (n970,n971,n1120);
xor (n971,n972,n1052);
xor (n972,n973,n1051);
xor (n973,n974,n977);
xor (n974,n975,n976);
and (n975,n934,n28);
and (n976,n118,n29);
or (n977,n978,n981);
and (n978,n979,n980);
and (n979,n118,n28);
and (n980,n39,n29);
and (n981,n982,n983);
xor (n982,n979,n980);
or (n983,n984,n987);
and (n984,n985,n986);
and (n985,n39,n28);
and (n986,n34,n29);
and (n987,n988,n989);
xor (n988,n985,n986);
or (n989,n990,n993);
and (n990,n991,n992);
and (n991,n34,n28);
and (n992,n177,n29);
and (n993,n994,n995);
xor (n994,n991,n992);
or (n995,n996,n999);
and (n996,n997,n998);
and (n997,n177,n28);
and (n998,n166,n29);
and (n999,n1000,n1001);
xor (n1000,n997,n998);
or (n1001,n1002,n1005);
and (n1002,n1003,n1004);
and (n1003,n166,n28);
and (n1004,n71,n29);
and (n1005,n1006,n1007);
xor (n1006,n1003,n1004);
or (n1007,n1008,n1011);
and (n1008,n1009,n1010);
and (n1009,n71,n28);
and (n1010,n52,n29);
and (n1011,n1012,n1013);
xor (n1012,n1009,n1010);
or (n1013,n1014,n1017);
and (n1014,n1015,n1016);
and (n1015,n52,n28);
and (n1016,n107,n29);
and (n1017,n1018,n1019);
xor (n1018,n1015,n1016);
or (n1019,n1020,n1023);
and (n1020,n1021,n1022);
and (n1021,n107,n28);
and (n1022,n88,n29);
and (n1023,n1024,n1025);
xor (n1024,n1021,n1022);
or (n1025,n1026,n1029);
and (n1026,n1027,n1028);
and (n1027,n88,n28);
and (n1028,n204,n29);
and (n1029,n1030,n1031);
xor (n1030,n1027,n1028);
or (n1031,n1032,n1035);
and (n1032,n1033,n1034);
and (n1033,n204,n28);
and (n1034,n188,n29);
and (n1035,n1036,n1037);
xor (n1036,n1033,n1034);
or (n1037,n1038,n1041);
and (n1038,n1039,n1040);
and (n1039,n188,n28);
and (n1040,n228,n29);
and (n1041,n1042,n1043);
xor (n1042,n1039,n1040);
or (n1043,n1044,n1046);
and (n1044,n1045,n808);
and (n1045,n228,n28);
and (n1046,n1047,n1048);
xor (n1047,n1045,n808);
and (n1048,n1049,n1050);
and (n1049,n143,n28);
and (n1050,n23,n29);
and (n1051,n39,n172);
or (n1052,n1053,n1056);
and (n1053,n1054,n1055);
xor (n1054,n982,n983);
and (n1055,n34,n172);
and (n1056,n1057,n1058);
xor (n1057,n1054,n1055);
or (n1058,n1059,n1062);
and (n1059,n1060,n1061);
xor (n1060,n988,n989);
and (n1061,n177,n172);
and (n1062,n1063,n1064);
xor (n1063,n1060,n1061);
or (n1064,n1065,n1068);
and (n1065,n1066,n1067);
xor (n1066,n994,n995);
and (n1067,n166,n172);
and (n1068,n1069,n1070);
xor (n1069,n1066,n1067);
or (n1070,n1071,n1074);
and (n1071,n1072,n1073);
xor (n1072,n1000,n1001);
and (n1073,n71,n172);
and (n1074,n1075,n1076);
xor (n1075,n1072,n1073);
or (n1076,n1077,n1080);
and (n1077,n1078,n1079);
xor (n1078,n1006,n1007);
and (n1079,n52,n172);
and (n1080,n1081,n1082);
xor (n1081,n1078,n1079);
or (n1082,n1083,n1086);
and (n1083,n1084,n1085);
xor (n1084,n1012,n1013);
and (n1085,n107,n172);
and (n1086,n1087,n1088);
xor (n1087,n1084,n1085);
or (n1088,n1089,n1092);
and (n1089,n1090,n1091);
xor (n1090,n1018,n1019);
and (n1091,n88,n172);
and (n1092,n1093,n1094);
xor (n1093,n1090,n1091);
or (n1094,n1095,n1098);
and (n1095,n1096,n1097);
xor (n1096,n1024,n1025);
and (n1097,n204,n172);
and (n1098,n1099,n1100);
xor (n1099,n1096,n1097);
or (n1100,n1101,n1104);
and (n1101,n1102,n1103);
xor (n1102,n1030,n1031);
and (n1103,n188,n172);
and (n1104,n1105,n1106);
xor (n1105,n1102,n1103);
or (n1106,n1107,n1110);
and (n1107,n1108,n1109);
xor (n1108,n1036,n1037);
and (n1109,n228,n172);
and (n1110,n1111,n1112);
xor (n1111,n1108,n1109);
or (n1112,n1113,n1116);
and (n1113,n1114,n1115);
xor (n1114,n1042,n1043);
and (n1115,n143,n172);
and (n1116,n1117,n1118);
xor (n1117,n1114,n1115);
and (n1118,n1119,n732);
xor (n1119,n1047,n1048);
and (n1120,n34,n61);
or (n1121,n1122,n1125);
and (n1122,n1123,n1124);
xor (n1123,n1057,n1058);
and (n1124,n177,n61);
and (n1125,n1126,n1127);
xor (n1126,n1123,n1124);
or (n1127,n1128,n1131);
and (n1128,n1129,n1130);
xor (n1129,n1063,n1064);
and (n1130,n166,n61);
and (n1131,n1132,n1133);
xor (n1132,n1129,n1130);
or (n1133,n1134,n1137);
and (n1134,n1135,n1136);
xor (n1135,n1069,n1070);
and (n1136,n71,n61);
and (n1137,n1138,n1139);
xor (n1138,n1135,n1136);
or (n1139,n1140,n1143);
and (n1140,n1141,n1142);
xor (n1141,n1075,n1076);
and (n1142,n52,n61);
and (n1143,n1144,n1145);
xor (n1144,n1141,n1142);
or (n1145,n1146,n1149);
and (n1146,n1147,n1148);
xor (n1147,n1081,n1082);
and (n1148,n107,n61);
and (n1149,n1150,n1151);
xor (n1150,n1147,n1148);
or (n1151,n1152,n1154);
and (n1152,n1153,n504);
xor (n1153,n1087,n1088);
and (n1154,n1155,n1156);
xor (n1155,n1153,n504);
or (n1156,n1157,n1159);
and (n1157,n1158,n593);
xor (n1158,n1093,n1094);
and (n1159,n1160,n1161);
xor (n1160,n1158,n593);
or (n1161,n1162,n1164);
and (n1162,n1163,n641);
xor (n1163,n1099,n1100);
and (n1164,n1165,n1166);
xor (n1165,n1163,n641);
or (n1166,n1167,n1170);
and (n1167,n1168,n1169);
xor (n1168,n1105,n1106);
and (n1169,n228,n61);
and (n1170,n1171,n1172);
xor (n1171,n1168,n1169);
or (n1172,n1173,n1176);
and (n1173,n1174,n1175);
xor (n1174,n1111,n1112);
and (n1175,n143,n61);
and (n1176,n1177,n1178);
xor (n1177,n1174,n1175);
and (n1178,n1179,n1180);
xor (n1179,n1117,n1118);
and (n1180,n23,n61);
and (n1181,n177,n60);
or (n1182,n1183,n1186);
and (n1183,n1184,n1185);
xor (n1184,n1126,n1127);
and (n1185,n166,n60);
and (n1186,n1187,n1188);
xor (n1187,n1184,n1185);
or (n1188,n1189,n1192);
and (n1189,n1190,n1191);
xor (n1190,n1132,n1133);
and (n1191,n71,n60);
and (n1192,n1193,n1194);
xor (n1193,n1190,n1191);
or (n1194,n1195,n1198);
and (n1195,n1196,n1197);
xor (n1196,n1138,n1139);
and (n1197,n52,n60);
and (n1198,n1199,n1200);
xor (n1199,n1196,n1197);
or (n1200,n1201,n1204);
and (n1201,n1202,n1203);
xor (n1202,n1144,n1145);
and (n1203,n107,n60);
and (n1204,n1205,n1206);
xor (n1205,n1202,n1203);
or (n1206,n1207,n1210);
and (n1207,n1208,n1209);
xor (n1208,n1150,n1151);
and (n1209,n88,n60);
and (n1210,n1211,n1212);
xor (n1211,n1208,n1209);
or (n1212,n1213,n1216);
and (n1213,n1214,n1215);
xor (n1214,n1155,n1156);
and (n1215,n204,n60);
and (n1216,n1217,n1218);
xor (n1217,n1214,n1215);
or (n1218,n1219,n1222);
and (n1219,n1220,n1221);
xor (n1220,n1160,n1161);
and (n1221,n188,n60);
and (n1222,n1223,n1224);
xor (n1223,n1220,n1221);
or (n1224,n1225,n1228);
and (n1225,n1226,n1227);
xor (n1226,n1165,n1166);
and (n1227,n228,n60);
and (n1228,n1229,n1230);
xor (n1229,n1226,n1227);
or (n1230,n1231,n1234);
and (n1231,n1232,n1233);
xor (n1232,n1171,n1172);
and (n1233,n143,n60);
and (n1234,n1235,n1236);
xor (n1235,n1232,n1233);
and (n1236,n1237,n628);
xor (n1237,n1177,n1178);
and (n1238,n166,n53);
or (n1239,n1240,n1243);
and (n1240,n1241,n1242);
xor (n1241,n1187,n1188);
and (n1242,n71,n53);
and (n1243,n1244,n1245);
xor (n1244,n1241,n1242);
or (n1245,n1246,n1249);
and (n1246,n1247,n1248);
xor (n1247,n1193,n1194);
and (n1248,n52,n53);
and (n1249,n1250,n1251);
xor (n1250,n1247,n1248);
or (n1251,n1252,n1255);
and (n1252,n1253,n1254);
xor (n1253,n1199,n1200);
and (n1254,n107,n53);
and (n1255,n1256,n1257);
xor (n1256,n1253,n1254);
or (n1257,n1258,n1261);
and (n1258,n1259,n1260);
xor (n1259,n1205,n1206);
and (n1260,n88,n53);
and (n1261,n1262,n1263);
xor (n1262,n1259,n1260);
or (n1263,n1264,n1267);
and (n1264,n1265,n1266);
xor (n1265,n1211,n1212);
and (n1266,n204,n53);
and (n1267,n1268,n1269);
xor (n1268,n1265,n1266);
or (n1269,n1270,n1273);
and (n1270,n1271,n1272);
xor (n1271,n1217,n1218);
and (n1272,n188,n53);
and (n1273,n1274,n1275);
xor (n1274,n1271,n1272);
or (n1275,n1276,n1279);
and (n1276,n1277,n1278);
xor (n1277,n1223,n1224);
and (n1278,n228,n53);
and (n1279,n1280,n1281);
xor (n1280,n1277,n1278);
or (n1281,n1282,n1285);
and (n1282,n1283,n1284);
xor (n1283,n1229,n1230);
and (n1284,n143,n53);
and (n1285,n1286,n1287);
xor (n1286,n1283,n1284);
and (n1287,n1288,n1289);
xor (n1288,n1235,n1236);
and (n1289,n23,n53);
and (n1290,n71,n98);
or (n1291,n1292,n1295);
and (n1292,n1293,n1294);
xor (n1293,n1244,n1245);
and (n1294,n52,n98);
and (n1295,n1296,n1297);
xor (n1296,n1293,n1294);
or (n1297,n1298,n1301);
and (n1298,n1299,n1300);
xor (n1299,n1250,n1251);
and (n1300,n107,n98);
and (n1301,n1302,n1303);
xor (n1302,n1299,n1300);
or (n1303,n1304,n1307);
and (n1304,n1305,n1306);
xor (n1305,n1256,n1257);
and (n1306,n88,n98);
and (n1307,n1308,n1309);
xor (n1308,n1305,n1306);
or (n1309,n1310,n1313);
and (n1310,n1311,n1312);
xor (n1311,n1262,n1263);
and (n1312,n204,n98);
and (n1313,n1314,n1315);
xor (n1314,n1311,n1312);
or (n1315,n1316,n1319);
and (n1316,n1317,n1318);
xor (n1317,n1268,n1269);
and (n1318,n188,n98);
and (n1319,n1320,n1321);
xor (n1320,n1317,n1318);
or (n1321,n1322,n1325);
and (n1322,n1323,n1324);
xor (n1323,n1274,n1275);
and (n1324,n228,n98);
and (n1325,n1326,n1327);
xor (n1326,n1323,n1324);
or (n1327,n1328,n1331);
and (n1328,n1329,n1330);
xor (n1329,n1280,n1281);
and (n1330,n143,n98);
and (n1331,n1332,n1333);
xor (n1332,n1329,n1330);
and (n1333,n1334,n546);
xor (n1334,n1286,n1287);
and (n1335,n52,n89);
or (n1336,n1337,n1340);
and (n1337,n1338,n1339);
xor (n1338,n1296,n1297);
and (n1339,n107,n89);
and (n1340,n1341,n1342);
xor (n1341,n1338,n1339);
or (n1342,n1343,n1345);
and (n1343,n1344,n87);
xor (n1344,n1302,n1303);
and (n1345,n1346,n1347);
xor (n1346,n1344,n87);
or (n1347,n1348,n1350);
and (n1348,n1349,n290);
xor (n1349,n1308,n1309);
and (n1350,n1351,n1352);
xor (n1351,n1349,n290);
or (n1352,n1353,n1355);
and (n1353,n1354,n285);
xor (n1354,n1314,n1315);
and (n1355,n1356,n1357);
xor (n1356,n1354,n285);
or (n1357,n1358,n1361);
and (n1358,n1359,n1360);
xor (n1359,n1320,n1321);
and (n1360,n228,n89);
and (n1361,n1362,n1363);
xor (n1362,n1359,n1360);
or (n1363,n1364,n1367);
and (n1364,n1365,n1366);
xor (n1365,n1326,n1327);
and (n1366,n143,n89);
and (n1367,n1368,n1369);
xor (n1368,n1365,n1366);
and (n1369,n1370,n1371);
xor (n1370,n1332,n1333);
and (n1371,n23,n89);
and (n1372,n107,n196);
or (n1373,n1374,n1377);
and (n1374,n1375,n1376);
xor (n1375,n1341,n1342);
and (n1376,n88,n196);
and (n1377,n1378,n1379);
xor (n1378,n1375,n1376);
or (n1379,n1380,n1383);
and (n1380,n1381,n1382);
xor (n1381,n1346,n1347);
and (n1382,n204,n196);
and (n1383,n1384,n1385);
xor (n1384,n1381,n1382);
or (n1385,n1386,n1389);
and (n1386,n1387,n1388);
xor (n1387,n1351,n1352);
and (n1388,n188,n196);
and (n1389,n1390,n1391);
xor (n1390,n1387,n1388);
or (n1391,n1392,n1395);
and (n1392,n1393,n1394);
xor (n1393,n1356,n1357);
and (n1394,n228,n196);
and (n1395,n1396,n1397);
xor (n1396,n1393,n1394);
or (n1397,n1398,n1401);
and (n1398,n1399,n1400);
xor (n1399,n1362,n1363);
and (n1400,n143,n196);
and (n1401,n1402,n1403);
xor (n1402,n1399,n1400);
and (n1403,n1404,n278);
xor (n1404,n1368,n1369);
and (n1405,n88,n79);
or (n1406,n1407,n1410);
and (n1407,n1408,n1409);
xor (n1408,n1378,n1379);
and (n1409,n204,n79);
and (n1410,n1411,n1412);
xor (n1411,n1408,n1409);
or (n1412,n1413,n1416);
and (n1413,n1414,n1415);
xor (n1414,n1384,n1385);
and (n1415,n188,n79);
and (n1416,n1417,n1418);
xor (n1417,n1414,n1415);
or (n1418,n1419,n1422);
and (n1419,n1420,n1421);
xor (n1420,n1390,n1391);
and (n1421,n228,n79);
and (n1422,n1423,n1424);
xor (n1423,n1420,n1421);
or (n1424,n1425,n1428);
and (n1425,n1426,n1427);
xor (n1426,n1396,n1397);
and (n1427,n143,n79);
and (n1428,n1429,n1430);
xor (n1429,n1426,n1427);
and (n1430,n1431,n1432);
xor (n1431,n1402,n1403);
and (n1432,n23,n79);
and (n1433,n204,n78);
or (n1434,n1435,n1438);
and (n1435,n1436,n1437);
xor (n1436,n1411,n1412);
and (n1437,n188,n78);
and (n1438,n1439,n1440);
xor (n1439,n1436,n1437);
or (n1440,n1441,n1444);
and (n1441,n1442,n1443);
xor (n1442,n1417,n1418);
and (n1443,n228,n78);
and (n1444,n1445,n1446);
xor (n1445,n1442,n1443);
or (n1446,n1447,n1450);
and (n1447,n1448,n1449);
xor (n1448,n1423,n1424);
and (n1449,n143,n78);
and (n1450,n1451,n1452);
xor (n1451,n1448,n1449);
and (n1452,n1453,n77);
xor (n1453,n1429,n1430);
or (n1454,n1455,n1457);
and (n1455,n1456,n229);
xor (n1456,n1439,n1440);
and (n1457,n1458,n1459);
xor (n1458,n1456,n229);
or (n1459,n1460,n1462);
and (n1460,n1461,n212);
xor (n1461,n1445,n1446);
and (n1462,n1463,n1464);
xor (n1463,n1461,n212);
and (n1464,n1465,n1466);
xor (n1465,n1451,n1452);
and (n1466,n23,n21);
and (n1467,n228,n19);
or (n1468,n1469,n1472);
and (n1469,n1470,n1471);
xor (n1470,n1458,n1459);
and (n1471,n143,n19);
and (n1472,n1473,n1474);
xor (n1473,n1470,n1471);
and (n1474,n1475,n134);
xor (n1475,n1463,n1464);
and (n1476,n143,n135);
and (n1477,n1478,n1479);
xor (n1478,n1473,n1474);
and (n1479,n23,n135);
and (n1480,n23,n927);
or (n1481,n1482,n1484,n1545);
and (n1482,n1483,n123);
xor (n1483,n1478,n1479);
and (n1484,n123,n1485);
or (n1485,n1486,n1488,n1544);
and (n1486,n1487,n15);
xor (n1487,n1475,n134);
and (n1488,n15,n1489);
or (n1489,n1490,n1492,n1543);
and (n1490,n1491,n82);
xor (n1491,n1465,n1466);
and (n1492,n82,n1493);
or (n1493,n1494,n1496,n1542);
and (n1494,n1495,n244);
xor (n1495,n1453,n77);
and (n1496,n244,n1497);
or (n1497,n1498,n1500,n1541);
and (n1498,n1499,n273);
xor (n1499,n1431,n1432);
and (n1500,n273,n1501);
or (n1501,n1502,n1504,n1540);
and (n1502,n1503,n509);
xor (n1503,n1404,n278);
and (n1504,n509,n1505);
or (n1505,n1506,n1508,n1539);
and (n1506,n1507,n540);
xor (n1507,n1370,n1371);
and (n1508,n540,n1509);
or (n1509,n1510,n1512,n1538);
and (n1510,n1511,n599);
xor (n1511,n1334,n546);
and (n1512,n599,n1513);
or (n1513,n1514,n1516,n1537);
and (n1514,n1515,n623);
xor (n1515,n1288,n1289);
and (n1516,n623,n1517);
or (n1517,n1518,n1520,n1536);
and (n1518,n1519,n724);
xor (n1519,n1237,n628);
and (n1520,n724,n1521);
or (n1521,n1522,n1524,n1535);
and (n1522,n1523,n728);
xor (n1523,n1179,n1180);
and (n1524,n728,n1525);
or (n1525,n1526,n1528,n1534);
and (n1526,n1527,n790);
xor (n1527,n1119,n732);
and (n1528,n790,n1529);
or (n1529,n1530,n1532,n1533);
and (n1530,n1531,n794);
xor (n1531,n1049,n1050);
and (n1532,n794,n825);
and (n1533,n1531,n825);
and (n1534,n1527,n1529);
and (n1535,n1523,n1525);
and (n1536,n1519,n1521);
and (n1537,n1515,n1517);
and (n1538,n1511,n1513);
and (n1539,n1507,n1509);
and (n1540,n1503,n1505);
and (n1541,n1499,n1501);
and (n1542,n1495,n1497);
and (n1543,n1491,n1493);
and (n1544,n1487,n1489);
and (n1545,n1483,n1485);
endmodule
