module top (out,n3,n4,n5,n26,n28,n35,n36,n46,n55
        ,n56,n61,n66,n72,n76,n88,n95,n96,n105,n114
        ,n116,n121,n131,n140,n147,n153,n197,n201,n206,n215
        ,n230,n819);
output out;
input n3;
input n4;
input n5;
input n26;
input n28;
input n35;
input n36;
input n46;
input n55;
input n56;
input n61;
input n66;
input n72;
input n76;
input n88;
input n95;
input n96;
input n105;
input n114;
input n116;
input n121;
input n131;
input n140;
input n147;
input n153;
input n197;
input n201;
input n206;
input n215;
input n230;
input n819;
wire n0;
wire n1;
wire n2;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n24;
wire n25;
wire n27;
wire n29;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n57;
wire n58;
wire n59;
wire n60;
wire n62;
wire n63;
wire n64;
wire n65;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n73;
wire n74;
wire n75;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n115;
wire n117;
wire n118;
wire n119;
wire n120;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n198;
wire n199;
wire n200;
wire n202;
wire n203;
wire n204;
wire n205;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
xnor (out,n0,n845);
nor (n0,n1,n6);
and (n1,n2,n5);
nor (n2,n3,n4);
and (n6,n7,n842);
nand (n7,n8,n841);
or (n8,n9,n768);
nand (n9,n10,n767);
or (n10,n11,n360);
not (n11,n12);
nand (n12,n13,n327);
not (n13,n14);
xor (n14,n15,n271);
xor (n15,n16,n158);
nand (n16,n17,n157);
or (n17,n18,n78);
or (n18,n19,n77);
and (n19,n20,n75);
xor (n20,n21,n49);
nand (n21,n22,n42);
or (n22,n23,n31);
not (n23,n24);
nand (n24,n25,n29);
or (n25,n26,n27);
not (n27,n28);
or (n29,n30,n28);
not (n30,n26);
nand (n31,n32,n39);
nor (n32,n33,n37);
and (n33,n34,n36);
not (n34,n35);
and (n37,n35,n38);
not (n38,n36);
nand (n39,n40,n41);
or (n40,n36,n30);
nand (n41,n30,n36);
nand (n42,n43,n48);
nor (n43,n44,n47);
and (n44,n45,n30);
not (n45,n46);
and (n47,n26,n46);
not (n48,n32);
nand (n49,n50,n69);
or (n50,n51,n63);
nand (n51,n52,n59);
nor (n52,n53,n57);
and (n53,n54,n56);
not (n54,n55);
and (n57,n55,n58);
not (n58,n56);
nand (n59,n60,n62);
or (n60,n58,n61);
nand (n62,n58,n61);
nor (n63,n64,n67);
and (n64,n65,n66);
not (n65,n61);
and (n67,n68,n61);
not (n68,n66);
or (n69,n52,n70);
nor (n70,n71,n73);
and (n71,n65,n72);
and (n73,n61,n74);
not (n74,n72);
and (n75,n61,n76);
and (n77,n21,n49);
not (n78,n79);
or (n79,n80,n156);
and (n80,n81,n133);
xor (n81,n82,n108);
nand (n82,n83,n102);
or (n83,n84,n90);
not (n84,n85);
nor (n85,n86,n89);
and (n86,n87,n34);
not (n87,n88);
and (n89,n35,n88);
not (n90,n91);
nor (n91,n92,n98);
nand (n92,n93,n97);
or (n93,n94,n96);
not (n94,n95);
nand (n97,n94,n96);
nor (n98,n99,n100);
and (n99,n34,n96);
and (n100,n35,n101);
not (n101,n96);
nand (n102,n92,n103);
nor (n103,n104,n106);
and (n104,n35,n105);
and (n106,n107,n34);
not (n107,n105);
nand (n108,n109,n127);
or (n109,n110,n118);
not (n110,n111);
nor (n111,n112,n117);
and (n112,n113,n115);
not (n113,n114);
not (n115,n116);
and (n117,n116,n114);
nand (n118,n119,n123);
nand (n119,n120,n122);
or (n120,n121,n115);
nand (n122,n115,n121);
not (n123,n124);
nand (n124,n125,n126);
or (n125,n30,n121);
nand (n126,n30,n121);
nand (n127,n124,n128);
nor (n128,n129,n132);
and (n129,n130,n115);
not (n130,n131);
and (n132,n116,n131);
nand (n133,n134,n150);
or (n134,n135,n145);
not (n135,n136);
and (n136,n137,n142);
not (n137,n138);
nand (n138,n139,n141);
or (n139,n140,n115);
nand (n141,n140,n115);
nand (n142,n143,n144);
or (n143,n140,n54);
nand (n144,n54,n140);
nor (n145,n146,n148);
and (n146,n54,n147);
and (n148,n55,n149);
not (n149,n147);
or (n150,n137,n151);
nor (n151,n152,n154);
and (n152,n54,n153);
and (n154,n55,n155);
not (n155,n153);
and (n156,n82,n108);
nand (n157,n78,n18);
xor (n158,n159,n217);
xor (n159,n160,n182);
xor (n160,n161,n175);
xor (n161,n162,n169);
nand (n162,n163,n165);
or (n163,n164,n118);
not (n164,n128);
nand (n165,n166,n124);
nor (n166,n167,n168);
and (n167,n27,n115);
and (n168,n116,n28);
nand (n169,n170,n171);
or (n170,n135,n151);
nand (n171,n138,n172);
nand (n172,n173,n174);
or (n173,n55,n113);
or (n174,n54,n114);
nand (n175,n176,n178);
or (n176,n177,n31);
not (n177,n43);
or (n178,n32,n179);
nor (n179,n180,n181);
and (n180,n30,n88);
and (n181,n26,n87);
xor (n182,n183,n191);
xor (n183,n184,n190);
nand (n184,n185,n186);
or (n185,n70,n51);
or (n186,n52,n187);
nor (n187,n188,n189);
and (n188,n147,n65);
and (n189,n149,n61);
and (n190,n61,n66);
xor (n191,n192,n208);
nand (n192,n193,n202);
or (n193,n194,n199);
nor (n194,n195,n198);
and (n195,n196,n95);
not (n196,n197);
and (n198,n197,n94);
nand (n199,n95,n200);
not (n200,n201);
or (n202,n203,n200);
not (n203,n204);
nand (n204,n205,n207);
or (n205,n206,n94);
nand (n207,n94,n206);
nand (n208,n209,n211);
or (n209,n210,n90);
not (n210,n103);
nand (n211,n92,n212);
nand (n212,n213,n216);
or (n213,n35,n214);
not (n214,n215);
or (n216,n34,n215);
or (n217,n218,n270);
and (n218,n219,n245);
xor (n219,n220,n226);
nand (n220,n221,n225);
or (n221,n222,n199);
nor (n222,n223,n224);
and (n223,n214,n95);
and (n224,n215,n94);
or (n225,n194,n200);
or (n226,n227,n244);
and (n227,n228,n238);
xor (n228,n229,n231);
and (n229,n61,n230);
nand (n231,n232,n237);
or (n232,n233,n90);
not (n233,n234);
nand (n234,n235,n236);
or (n235,n35,n45);
or (n236,n34,n46);
nand (n237,n85,n92);
nand (n238,n239,n240);
or (n239,n110,n123);
or (n240,n118,n241);
nor (n241,n242,n243);
and (n242,n115,n153);
and (n243,n116,n155);
and (n244,n229,n231);
or (n245,n246,n269);
and (n246,n247,n260);
xor (n247,n248,n254);
nand (n248,n249,n253);
or (n249,n135,n250);
nor (n250,n251,n252);
and (n251,n54,n72);
and (n252,n55,n74);
or (n253,n137,n145);
nand (n254,n255,n259);
or (n255,n256,n199);
nor (n256,n257,n258);
and (n257,n107,n95);
and (n258,n105,n94);
or (n259,n222,n200);
nand (n260,n261,n266);
or (n261,n262,n51);
nor (n262,n263,n264);
and (n263,n76,n65);
and (n264,n265,n61);
not (n265,n76);
nand (n266,n267,n268);
not (n267,n63);
not (n268,n52);
and (n269,n248,n254);
and (n270,n220,n226);
or (n271,n272,n326);
and (n272,n273,n276);
xor (n273,n274,n275);
xor (n274,n20,n75);
xor (n275,n81,n133);
or (n276,n277,n325);
and (n277,n278,n300);
xor (n278,n279,n285);
nand (n279,n280,n284);
or (n280,n31,n281);
nor (n281,n282,n283);
and (n282,n30,n131);
and (n283,n26,n130);
or (n284,n32,n23);
nor (n285,n286,n294);
not (n286,n287);
nand (n287,n288,n293);
or (n288,n289,n90);
not (n289,n290);
nor (n290,n291,n292);
and (n291,n27,n34);
and (n292,n35,n28);
nand (n293,n92,n234);
nand (n294,n295,n61);
nand (n295,n296,n297);
or (n296,n55,n56);
nand (n297,n298,n299);
or (n298,n58,n54);
not (n299,n230);
or (n300,n301,n324);
and (n301,n302,n318);
xor (n302,n303,n311);
nand (n303,n304,n309);
or (n304,n305,n118);
not (n305,n306);
nand (n306,n307,n308);
or (n307,n116,n149);
or (n308,n115,n147);
nand (n309,n310,n124);
not (n310,n241);
nand (n311,n312,n317);
or (n312,n313,n135);
not (n313,n314);
nand (n314,n315,n316);
or (n315,n55,n68);
or (n316,n54,n66);
or (n317,n137,n250);
nand (n318,n319,n323);
or (n319,n320,n199);
nor (n320,n321,n322);
and (n321,n94,n88);
and (n322,n95,n87);
or (n323,n256,n200);
and (n324,n303,n311);
and (n325,n279,n285);
and (n326,n274,n275);
not (n327,n328);
or (n328,n329,n359);
and (n329,n330,n358);
xor (n330,n331,n332);
xor (n331,n219,n245);
or (n332,n333,n357);
and (n333,n334,n337);
xor (n334,n335,n336);
xor (n335,n247,n260);
xor (n336,n228,n238);
or (n337,n338,n356);
and (n338,n339,n352);
xor (n339,n340,n346);
nand (n340,n341,n345);
or (n341,n51,n342);
nor (n342,n343,n344);
and (n343,n65,n230);
and (n344,n299,n61);
or (n345,n52,n262);
nand (n346,n347,n351);
or (n347,n31,n348);
nor (n348,n349,n350);
and (n349,n30,n114);
and (n350,n26,n113);
or (n351,n32,n281);
nand (n352,n353,n355);
or (n353,n354,n286);
not (n354,n294);
or (n355,n287,n294);
and (n356,n340,n346);
and (n357,n335,n336);
xor (n358,n273,n276);
and (n359,n331,n332);
not (n360,n361);
nand (n361,n362,n761);
or (n362,n363,n472);
not (n363,n364);
and (n364,n365,n422);
nand (n365,n366,n368);
not (n366,n367);
xor (n367,n330,n358);
not (n368,n369);
or (n369,n370,n421);
and (n370,n371,n420);
xor (n371,n372,n373);
xor (n372,n278,n300);
or (n373,n374,n419);
and (n374,n375,n418);
xor (n375,n376,n395);
or (n376,n377,n394);
and (n377,n378,n387);
xor (n378,n379,n380);
and (n379,n268,n230);
nand (n380,n381,n386);
or (n381,n382,n90);
not (n382,n383);
nand (n383,n384,n385);
or (n384,n35,n130);
or (n385,n34,n131);
nand (n386,n92,n290);
nand (n387,n388,n393);
or (n388,n389,n118);
not (n389,n390);
nor (n390,n391,n392);
and (n391,n74,n115);
and (n392,n116,n72);
nand (n393,n124,n306);
and (n394,n379,n380);
or (n395,n396,n417);
and (n396,n397,n411);
xor (n397,n398,n405);
nand (n398,n399,n404);
or (n399,n400,n135);
not (n400,n401);
nand (n401,n402,n403);
or (n402,n55,n265);
or (n403,n54,n76);
nand (n404,n138,n314);
nand (n405,n406,n410);
or (n406,n407,n199);
nor (n407,n408,n409);
and (n408,n94,n46);
and (n409,n95,n45);
or (n410,n320,n200);
nand (n411,n412,n416);
or (n412,n31,n413);
nor (n413,n414,n415);
and (n414,n30,n153);
and (n415,n26,n155);
or (n416,n348,n32);
and (n417,n398,n405);
xor (n418,n302,n318);
and (n419,n376,n395);
xor (n420,n334,n337);
and (n421,n372,n373);
or (n422,n423,n424);
xor (n423,n371,n420);
or (n424,n425,n471);
and (n425,n426,n429);
xor (n426,n427,n428);
xor (n427,n339,n352);
xor (n428,n375,n418);
or (n429,n430,n470);
and (n430,n431,n469);
xor (n431,n432,n447);
and (n432,n433,n439);
and (n433,n434,n55);
nand (n434,n435,n436);
or (n435,n116,n140);
nand (n436,n437,n299);
or (n437,n438,n115);
not (n438,n140);
nand (n439,n440,n442);
or (n440,n441,n382);
not (n441,n92);
nand (n442,n443,n91);
not (n443,n444);
nor (n444,n445,n446);
and (n445,n34,n114);
and (n446,n35,n113);
or (n447,n448,n468);
and (n448,n449,n462);
xor (n449,n450,n456);
nand (n450,n451,n455);
or (n451,n118,n452);
nor (n452,n453,n454);
and (n453,n68,n116);
and (n454,n66,n115);
nand (n455,n390,n124);
nand (n456,n457,n458);
or (n457,n137,n400);
nand (n458,n136,n459);
nand (n459,n460,n461);
or (n460,n55,n299);
or (n461,n54,n230);
nand (n462,n463,n467);
or (n463,n199,n464);
nor (n464,n465,n466);
and (n465,n94,n28);
and (n466,n95,n27);
or (n467,n407,n200);
and (n468,n450,n456);
xor (n469,n378,n387);
and (n470,n432,n447);
and (n471,n427,n428);
not (n472,n473);
nand (n473,n474,n751,n760);
nand (n474,n475,n610,n617);
nor (n475,n476,n549);
not (n476,n477);
nand (n477,n478,n512);
not (n478,n479);
xor (n479,n480,n511);
xor (n480,n481,n482);
xor (n481,n397,n411);
or (n482,n483,n510);
and (n483,n484,n492);
xor (n484,n485,n491);
nand (n485,n486,n490);
or (n486,n31,n487);
nor (n487,n488,n489);
and (n488,n147,n30);
and (n489,n26,n149);
or (n490,n413,n32);
xor (n491,n433,n439);
or (n492,n493,n509);
and (n493,n494,n502);
xor (n494,n495,n496);
and (n495,n138,n230);
nand (n496,n497,n501);
or (n497,n498,n199);
nor (n498,n499,n500);
and (n499,n130,n95);
and (n500,n131,n94);
or (n501,n464,n200);
nand (n502,n503,n508);
or (n503,n118,n504);
not (n504,n505);
nor (n505,n506,n507);
and (n506,n265,n115);
and (n507,n116,n76);
or (n508,n123,n452);
and (n509,n495,n496);
and (n510,n485,n491);
xor (n511,n431,n469);
not (n512,n513);
or (n513,n514,n548);
and (n514,n515,n547);
xor (n515,n516,n517);
xor (n516,n449,n462);
or (n517,n518,n546);
and (n518,n519,n532);
xor (n519,n520,n526);
nand (n520,n521,n525);
or (n521,n90,n522);
nor (n522,n523,n524);
and (n523,n155,n35);
and (n524,n153,n34);
or (n525,n441,n444);
nand (n526,n527,n531);
or (n527,n31,n528);
nor (n528,n529,n530);
and (n529,n72,n30);
and (n530,n26,n74);
or (n531,n32,n487);
and (n532,n533,n539);
nor (n533,n534,n115);
nor (n534,n535,n537);
and (n535,n536,n299);
nand (n536,n26,n121);
and (n537,n30,n538);
not (n538,n121);
nand (n539,n540,n545);
or (n540,n199,n541);
not (n541,n542);
nor (n542,n543,n544);
and (n543,n95,n114);
and (n544,n113,n94);
or (n545,n498,n200);
and (n546,n520,n526);
xor (n547,n484,n492);
and (n548,n516,n517);
nand (n549,n550,n584);
not (n550,n551);
nor (n551,n552,n553);
xor (n552,n515,n547);
or (n553,n554,n583);
and (n554,n555,n582);
xor (n555,n556,n581);
or (n556,n557,n580);
and (n557,n558,n574);
xor (n558,n559,n566);
nand (n559,n560,n565);
or (n560,n561,n118);
not (n561,n562);
nand (n562,n563,n564);
or (n563,n116,n299);
or (n564,n115,n230);
nand (n565,n505,n124);
nand (n566,n567,n572);
or (n567,n568,n90);
not (n568,n569);
nand (n569,n570,n571);
or (n570,n35,n149);
or (n571,n34,n147);
nand (n572,n573,n92);
not (n573,n522);
nand (n574,n575,n579);
or (n575,n31,n576);
nor (n576,n577,n578);
and (n577,n30,n66);
and (n578,n26,n68);
or (n579,n32,n528);
and (n580,n559,n566);
xor (n581,n494,n502);
xor (n582,n519,n532);
and (n583,n556,n581);
or (n584,n585,n586);
xor (n585,n555,n582);
or (n586,n587,n609);
and (n587,n588,n608);
xor (n588,n589,n590);
xor (n589,n533,n539);
or (n590,n591,n607);
and (n591,n592,n600);
xor (n592,n593,n594);
and (n593,n124,n230);
nand (n594,n595,n596);
or (n595,n200,n541);
or (n596,n199,n597);
nor (n597,n598,n599);
and (n598,n94,n153);
and (n599,n95,n155);
nand (n600,n601,n606);
or (n601,n602,n90);
not (n602,n603);
nor (n603,n604,n605);
and (n604,n35,n72);
and (n605,n74,n34);
nand (n606,n92,n569);
and (n607,n593,n594);
xor (n608,n558,n574);
and (n609,n589,n590);
nand (n610,n611,n613);
not (n611,n612);
xor (n612,n426,n429);
not (n613,n614);
or (n614,n615,n616);
and (n615,n480,n511);
and (n616,n481,n482);
or (n617,n618,n750);
and (n618,n619,n644);
xor (n619,n620,n643);
or (n620,n621,n642);
and (n621,n622,n641);
xor (n622,n623,n629);
nand (n623,n624,n628);
or (n624,n31,n625);
nor (n625,n626,n627);
and (n626,n30,n76);
and (n627,n26,n265);
or (n628,n32,n576);
and (n629,n630,n635);
and (n630,n631,n26);
nand (n631,n632,n633);
or (n632,n35,n36);
nand (n633,n634,n299);
or (n634,n38,n34);
nand (n635,n636,n640);
or (n636,n637,n199);
nor (n637,n638,n639);
and (n638,n94,n147);
and (n639,n95,n149);
or (n640,n597,n200);
xor (n641,n592,n600);
and (n642,n623,n629);
xor (n643,n588,n608);
or (n644,n645,n749);
and (n645,n646,n667);
xor (n646,n647,n666);
or (n647,n648,n665);
and (n648,n649,n664);
xor (n649,n650,n657);
nand (n650,n651,n656);
or (n651,n652,n90);
not (n652,n653);
nor (n653,n654,n655);
and (n654,n68,n34);
and (n655,n35,n66);
nand (n656,n92,n603);
nand (n657,n658,n663);
or (n658,n659,n31);
not (n659,n660);
nand (n660,n661,n662);
or (n661,n299,n26);
or (n662,n30,n230);
or (n663,n32,n625);
xor (n664,n630,n635);
and (n665,n650,n657);
xor (n666,n622,n641);
or (n667,n668,n748);
and (n668,n669,n689);
xor (n669,n670,n688);
or (n670,n671,n687);
and (n671,n672,n680);
xor (n672,n673,n674);
nor (n673,n32,n299);
nand (n674,n675,n679);
or (n675,n676,n90);
nor (n676,n677,n678);
and (n677,n76,n34);
and (n678,n265,n35);
nand (n679,n653,n92);
nand (n680,n681,n686);
or (n681,n199,n682);
not (n682,n683);
nand (n683,n684,n685);
or (n684,n72,n94);
nand (n685,n94,n72);
or (n686,n637,n200);
and (n687,n673,n674);
xor (n688,n649,n664);
or (n689,n690,n747);
and (n690,n691,n746);
xor (n691,n692,n707);
nor (n692,n693,n701);
not (n693,n694);
nand (n694,n695,n700);
or (n695,n199,n696);
not (n696,n697);
nand (n697,n698,n699);
or (n698,n66,n94);
nand (n699,n94,n66);
nand (n700,n683,n201);
nand (n701,n702,n35);
nand (n702,n703,n706);
nand (n703,n704,n299);
not (n704,n705);
and (n705,n95,n96);
or (n706,n96,n95);
nand (n707,n708,n745);
nand (n708,n709,n722);
or (n709,n710,n717);
not (n710,n711);
nor (n711,n712,n716);
and (n712,n91,n713);
nand (n713,n714,n715);
or (n714,n35,n299);
or (n715,n34,n230);
nor (n716,n441,n676);
not (n717,n718);
nor (n718,n719,n720);
and (n719,n701,n694);
and (n720,n721,n693);
not (n721,n701);
nand (n722,n723,n744);
or (n723,n724,n734);
nor (n724,n725,n727);
not (n725,n726);
nand (n726,n92,n230);
nand (n727,n728,n729);
or (n728,n200,n696);
nand (n729,n730,n733);
nand (n730,n731,n732);
or (n731,n265,n95);
nand (n732,n95,n265);
not (n733,n199);
nand (n734,n735,n742);
nand (n735,n736,n740);
or (n736,n737,n199);
nor (n737,n738,n739);
and (n738,n299,n95);
and (n739,n230,n94);
or (n740,n741,n200);
not (n741,n730);
nor (n742,n743,n94);
and (n743,n230,n201);
nand (n744,n725,n727);
or (n745,n718,n711);
xor (n746,n672,n680);
and (n747,n692,n707);
and (n748,n670,n688);
and (n749,n647,n666);
and (n750,n620,n643);
nand (n751,n752,n610);
nand (n752,n753,n759);
or (n753,n754,n476);
not (n754,n755);
nand (n755,n756,n758);
or (n756,n551,n757);
nand (n757,n585,n586);
nand (n758,n552,n553);
nand (n759,n479,n513);
nand (n760,n612,n614);
nand (n761,n762,n365);
or (n762,n763,n765);
not (n763,n764);
nand (n764,n423,n424);
not (n765,n766);
nand (n766,n367,n369);
nand (n767,n14,n328);
nand (n768,n769,n840);
nand (n769,n770,n836);
not (n770,n771);
xor (n771,n772,n833);
xor (n772,n773,n801);
xor (n773,n774,n779);
xor (n774,n775,n776);
and (n775,n192,n208);
or (n776,n777,n778);
and (n777,n161,n175);
and (n778,n162,n169);
xor (n779,n780,n795);
xor (n780,n781,n788);
nand (n781,n782,n784);
or (n782,n783,n118);
not (n783,n166);
nand (n784,n785,n124);
nor (n785,n786,n787);
and (n786,n116,n46);
and (n787,n45,n115);
nand (n788,n789,n791);
or (n789,n790,n135);
not (n790,n172);
nand (n791,n138,n792);
nand (n792,n793,n794);
or (n793,n55,n130);
or (n794,n54,n131);
nand (n795,n796,n797);
or (n796,n31,n179);
or (n797,n798,n32);
nor (n798,n799,n800);
and (n799,n30,n105);
and (n800,n26,n107);
xor (n801,n802,n832);
xor (n802,n803,n829);
xor (n803,n804,n812);
xor (n804,n805,n811);
nand (n805,n806,n807);
or (n806,n51,n187);
or (n807,n52,n808);
nor (n808,n809,n810);
and (n809,n153,n65);
and (n810,n155,n61);
and (n811,n61,n72);
xor (n812,n813,n822);
nand (n813,n814,n821);
or (n814,n200,n815);
not (n815,n816);
nor (n816,n817,n820);
and (n817,n818,n94);
not (n818,n819);
and (n820,n95,n819);
nand (n821,n204,n733);
nand (n822,n823,n825);
or (n823,n824,n90);
not (n824,n212);
nand (n825,n92,n826);
nor (n826,n827,n828);
and (n827,n35,n197);
and (n828,n196,n34);
or (n829,n830,n831);
and (n830,n183,n191);
and (n831,n184,n190);
and (n832,n79,n18);
or (n833,n834,n835);
and (n834,n159,n217);
and (n835,n160,n182);
not (n836,n837);
or (n837,n838,n839);
and (n838,n15,n271);
and (n839,n16,n158);
nand (n840,n771,n837);
nand (n841,n9,n768);
not (n842,n843);
nand (n843,n844,n3);
not (n844,n4);
wire s0n845,s1n845,notn845;
or (n845,s0n845,s1n845);
not(notn845,n4);
and (s0n845,notn845,n846);
and (s1n845,n4,1'b0);
wire s0n846,s1n846,notn846;
or (n846,s0n846,s1n846);
not(notn846,n3);
and (s0n846,notn846,n5);
and (s1n846,n3,n847);
xor (n847,n848,n1429);
xor (n848,n849,n1426);
xor (n849,n850,n1425);
xor (n850,n851,n1416);
xor (n851,n852,n1415);
xor (n852,n853,n1400);
xor (n853,n854,n1399);
xor (n854,n855,n1379);
xor (n855,n856,n1378);
xor (n856,n857,n1352);
xor (n857,n858,n1351);
xor (n858,n859,n1319);
xor (n859,n860,n1318);
xor (n860,n861,n1280);
xor (n861,n862,n168);
xor (n862,n863,n1236);
xor (n863,n864,n1235);
xor (n864,n865,n1186);
xor (n865,n866,n1185);
xor (n866,n867,n1128);
xor (n867,n868,n1127);
xor (n868,n869,n1064);
xor (n869,n870,n1063);
or (n870,n871,n1000);
and (n871,n872,n811);
or (n872,n873,n936);
and (n873,n874,n190);
and (n874,n75,n875);
or (n875,n876,n878);
and (n876,n229,n877);
and (n877,n56,n76);
and (n878,n879,n880);
xor (n879,n229,n877);
or (n880,n881,n884);
and (n881,n882,n883);
and (n882,n56,n230);
and (n883,n55,n76);
and (n884,n885,n886);
xor (n885,n882,n883);
or (n886,n887,n890);
and (n887,n888,n889);
and (n888,n55,n230);
and (n889,n140,n76);
and (n890,n891,n892);
xor (n891,n888,n889);
or (n892,n893,n895);
and (n893,n894,n507);
and (n894,n140,n230);
and (n895,n896,n897);
xor (n896,n894,n507);
or (n897,n898,n901);
and (n898,n899,n900);
and (n899,n116,n230);
and (n900,n121,n76);
and (n901,n902,n903);
xor (n902,n899,n900);
or (n903,n904,n907);
and (n904,n905,n906);
and (n905,n121,n230);
and (n906,n26,n76);
and (n907,n908,n909);
xor (n908,n905,n906);
or (n909,n910,n913);
and (n910,n911,n912);
and (n911,n26,n230);
and (n912,n36,n76);
and (n913,n914,n915);
xor (n914,n911,n912);
or (n915,n916,n919);
and (n916,n917,n918);
and (n917,n36,n230);
and (n918,n35,n76);
and (n919,n920,n921);
xor (n920,n917,n918);
or (n921,n922,n925);
and (n922,n923,n924);
and (n923,n35,n230);
and (n924,n96,n76);
and (n925,n926,n927);
xor (n926,n923,n924);
or (n927,n928,n931);
and (n928,n929,n930);
and (n929,n96,n230);
and (n930,n95,n76);
and (n931,n932,n933);
xor (n932,n929,n930);
and (n933,n934,n935);
and (n934,n95,n230);
and (n935,n201,n76);
and (n936,n937,n938);
xor (n937,n874,n190);
or (n938,n939,n942);
and (n939,n940,n941);
xor (n940,n75,n875);
and (n941,n56,n66);
and (n942,n943,n944);
xor (n943,n940,n941);
or (n944,n945,n948);
and (n945,n946,n947);
xor (n946,n879,n880);
and (n947,n55,n66);
and (n948,n949,n950);
xor (n949,n946,n947);
or (n950,n951,n954);
and (n951,n952,n953);
xor (n952,n885,n886);
and (n953,n140,n66);
and (n954,n955,n956);
xor (n955,n952,n953);
or (n956,n957,n960);
and (n957,n958,n959);
xor (n958,n891,n892);
and (n959,n116,n66);
and (n960,n961,n962);
xor (n961,n958,n959);
or (n962,n963,n966);
and (n963,n964,n965);
xor (n964,n896,n897);
and (n965,n121,n66);
and (n966,n967,n968);
xor (n967,n964,n965);
or (n968,n969,n972);
and (n969,n970,n971);
xor (n970,n902,n903);
and (n971,n26,n66);
and (n972,n973,n974);
xor (n973,n970,n971);
or (n974,n975,n978);
and (n975,n976,n977);
xor (n976,n908,n909);
and (n977,n36,n66);
and (n978,n979,n980);
xor (n979,n976,n977);
or (n980,n981,n983);
and (n981,n982,n655);
xor (n982,n914,n915);
and (n983,n984,n985);
xor (n984,n982,n655);
or (n985,n986,n989);
and (n986,n987,n988);
xor (n987,n920,n921);
and (n988,n96,n66);
and (n989,n990,n991);
xor (n990,n987,n988);
or (n991,n992,n995);
and (n992,n993,n994);
xor (n993,n926,n927);
and (n994,n95,n66);
and (n995,n996,n997);
xor (n996,n993,n994);
and (n997,n998,n999);
xor (n998,n932,n933);
and (n999,n201,n66);
and (n1000,n1001,n1002);
xor (n1001,n872,n811);
or (n1002,n1003,n1006);
and (n1003,n1004,n1005);
xor (n1004,n937,n938);
and (n1005,n56,n72);
and (n1006,n1007,n1008);
xor (n1007,n1004,n1005);
or (n1008,n1009,n1012);
and (n1009,n1010,n1011);
xor (n1010,n943,n944);
and (n1011,n55,n72);
and (n1012,n1013,n1014);
xor (n1013,n1010,n1011);
or (n1014,n1015,n1018);
and (n1015,n1016,n1017);
xor (n1016,n949,n950);
and (n1017,n140,n72);
and (n1018,n1019,n1020);
xor (n1019,n1016,n1017);
or (n1020,n1021,n1023);
and (n1021,n1022,n392);
xor (n1022,n955,n956);
and (n1023,n1024,n1025);
xor (n1024,n1022,n392);
or (n1025,n1026,n1029);
and (n1026,n1027,n1028);
xor (n1027,n961,n962);
and (n1028,n121,n72);
and (n1029,n1030,n1031);
xor (n1030,n1027,n1028);
or (n1031,n1032,n1035);
and (n1032,n1033,n1034);
xor (n1033,n967,n968);
and (n1034,n26,n72);
and (n1035,n1036,n1037);
xor (n1036,n1033,n1034);
or (n1037,n1038,n1041);
and (n1038,n1039,n1040);
xor (n1039,n973,n974);
and (n1040,n36,n72);
and (n1041,n1042,n1043);
xor (n1042,n1039,n1040);
or (n1043,n1044,n1046);
and (n1044,n1045,n604);
xor (n1045,n979,n980);
and (n1046,n1047,n1048);
xor (n1047,n1045,n604);
or (n1048,n1049,n1052);
and (n1049,n1050,n1051);
xor (n1050,n984,n985);
and (n1051,n96,n72);
and (n1052,n1053,n1054);
xor (n1053,n1050,n1051);
or (n1054,n1055,n1058);
and (n1055,n1056,n1057);
xor (n1056,n990,n991);
and (n1057,n95,n72);
and (n1058,n1059,n1060);
xor (n1059,n1056,n1057);
and (n1060,n1061,n1062);
xor (n1061,n996,n997);
and (n1062,n201,n72);
and (n1063,n61,n147);
or (n1064,n1065,n1068);
and (n1065,n1066,n1067);
xor (n1066,n1001,n1002);
and (n1067,n56,n147);
and (n1068,n1069,n1070);
xor (n1069,n1066,n1067);
or (n1070,n1071,n1074);
and (n1071,n1072,n1073);
xor (n1072,n1007,n1008);
and (n1073,n55,n147);
and (n1074,n1075,n1076);
xor (n1075,n1072,n1073);
or (n1076,n1077,n1080);
and (n1077,n1078,n1079);
xor (n1078,n1013,n1014);
and (n1079,n140,n147);
and (n1080,n1081,n1082);
xor (n1081,n1078,n1079);
or (n1082,n1083,n1086);
and (n1083,n1084,n1085);
xor (n1084,n1019,n1020);
and (n1085,n116,n147);
and (n1086,n1087,n1088);
xor (n1087,n1084,n1085);
or (n1088,n1089,n1092);
and (n1089,n1090,n1091);
xor (n1090,n1024,n1025);
and (n1091,n121,n147);
and (n1092,n1093,n1094);
xor (n1093,n1090,n1091);
or (n1094,n1095,n1098);
and (n1095,n1096,n1097);
xor (n1096,n1030,n1031);
and (n1097,n26,n147);
and (n1098,n1099,n1100);
xor (n1099,n1096,n1097);
or (n1100,n1101,n1104);
and (n1101,n1102,n1103);
xor (n1102,n1036,n1037);
and (n1103,n36,n147);
and (n1104,n1105,n1106);
xor (n1105,n1102,n1103);
or (n1106,n1107,n1110);
and (n1107,n1108,n1109);
xor (n1108,n1042,n1043);
and (n1109,n35,n147);
and (n1110,n1111,n1112);
xor (n1111,n1108,n1109);
or (n1112,n1113,n1116);
and (n1113,n1114,n1115);
xor (n1114,n1047,n1048);
and (n1115,n96,n147);
and (n1116,n1117,n1118);
xor (n1117,n1114,n1115);
or (n1118,n1119,n1122);
and (n1119,n1120,n1121);
xor (n1120,n1053,n1054);
and (n1121,n95,n147);
and (n1122,n1123,n1124);
xor (n1123,n1120,n1121);
and (n1124,n1125,n1126);
xor (n1125,n1059,n1060);
and (n1126,n201,n147);
and (n1127,n56,n153);
or (n1128,n1129,n1132);
and (n1129,n1130,n1131);
xor (n1130,n1069,n1070);
and (n1131,n55,n153);
and (n1132,n1133,n1134);
xor (n1133,n1130,n1131);
or (n1134,n1135,n1138);
and (n1135,n1136,n1137);
xor (n1136,n1075,n1076);
and (n1137,n140,n153);
and (n1138,n1139,n1140);
xor (n1139,n1136,n1137);
or (n1140,n1141,n1144);
and (n1141,n1142,n1143);
xor (n1142,n1081,n1082);
and (n1143,n116,n153);
and (n1144,n1145,n1146);
xor (n1145,n1142,n1143);
or (n1146,n1147,n1150);
and (n1147,n1148,n1149);
xor (n1148,n1087,n1088);
and (n1149,n121,n153);
and (n1150,n1151,n1152);
xor (n1151,n1148,n1149);
or (n1152,n1153,n1156);
and (n1153,n1154,n1155);
xor (n1154,n1093,n1094);
and (n1155,n26,n153);
and (n1156,n1157,n1158);
xor (n1157,n1154,n1155);
or (n1158,n1159,n1162);
and (n1159,n1160,n1161);
xor (n1160,n1099,n1100);
and (n1161,n36,n153);
and (n1162,n1163,n1164);
xor (n1163,n1160,n1161);
or (n1164,n1165,n1168);
and (n1165,n1166,n1167);
xor (n1166,n1105,n1106);
and (n1167,n35,n153);
and (n1168,n1169,n1170);
xor (n1169,n1166,n1167);
or (n1170,n1171,n1174);
and (n1171,n1172,n1173);
xor (n1172,n1111,n1112);
and (n1173,n96,n153);
and (n1174,n1175,n1176);
xor (n1175,n1172,n1173);
or (n1176,n1177,n1180);
and (n1177,n1178,n1179);
xor (n1178,n1117,n1118);
and (n1179,n95,n153);
and (n1180,n1181,n1182);
xor (n1181,n1178,n1179);
and (n1182,n1183,n1184);
xor (n1183,n1123,n1124);
and (n1184,n201,n153);
and (n1185,n55,n114);
or (n1186,n1187,n1190);
and (n1187,n1188,n1189);
xor (n1188,n1133,n1134);
and (n1189,n140,n114);
and (n1190,n1191,n1192);
xor (n1191,n1188,n1189);
or (n1192,n1193,n1195);
and (n1193,n1194,n117);
xor (n1194,n1139,n1140);
and (n1195,n1196,n1197);
xor (n1196,n1194,n117);
or (n1197,n1198,n1201);
and (n1198,n1199,n1200);
xor (n1199,n1145,n1146);
and (n1200,n121,n114);
and (n1201,n1202,n1203);
xor (n1202,n1199,n1200);
or (n1203,n1204,n1207);
and (n1204,n1205,n1206);
xor (n1205,n1151,n1152);
and (n1206,n26,n114);
and (n1207,n1208,n1209);
xor (n1208,n1205,n1206);
or (n1209,n1210,n1213);
and (n1210,n1211,n1212);
xor (n1211,n1157,n1158);
and (n1212,n36,n114);
and (n1213,n1214,n1215);
xor (n1214,n1211,n1212);
or (n1215,n1216,n1219);
and (n1216,n1217,n1218);
xor (n1217,n1163,n1164);
and (n1218,n35,n114);
and (n1219,n1220,n1221);
xor (n1220,n1217,n1218);
or (n1221,n1222,n1225);
and (n1222,n1223,n1224);
xor (n1223,n1169,n1170);
and (n1224,n96,n114);
and (n1225,n1226,n1227);
xor (n1226,n1223,n1224);
or (n1227,n1228,n1230);
and (n1228,n1229,n543);
xor (n1229,n1175,n1176);
and (n1230,n1231,n1232);
xor (n1231,n1229,n543);
and (n1232,n1233,n1234);
xor (n1233,n1181,n1182);
and (n1234,n201,n114);
and (n1235,n140,n131);
or (n1236,n1237,n1239);
and (n1237,n1238,n132);
xor (n1238,n1191,n1192);
and (n1239,n1240,n1241);
xor (n1240,n1238,n132);
or (n1241,n1242,n1245);
and (n1242,n1243,n1244);
xor (n1243,n1196,n1197);
and (n1244,n121,n131);
and (n1245,n1246,n1247);
xor (n1246,n1243,n1244);
or (n1247,n1248,n1251);
and (n1248,n1249,n1250);
xor (n1249,n1202,n1203);
and (n1250,n26,n131);
and (n1251,n1252,n1253);
xor (n1252,n1249,n1250);
or (n1253,n1254,n1257);
and (n1254,n1255,n1256);
xor (n1255,n1208,n1209);
and (n1256,n36,n131);
and (n1257,n1258,n1259);
xor (n1258,n1255,n1256);
or (n1259,n1260,n1263);
and (n1260,n1261,n1262);
xor (n1261,n1214,n1215);
and (n1262,n35,n131);
and (n1263,n1264,n1265);
xor (n1264,n1261,n1262);
or (n1265,n1266,n1269);
and (n1266,n1267,n1268);
xor (n1267,n1220,n1221);
and (n1268,n96,n131);
and (n1269,n1270,n1271);
xor (n1270,n1267,n1268);
or (n1271,n1272,n1275);
and (n1272,n1273,n1274);
xor (n1273,n1226,n1227);
and (n1274,n95,n131);
and (n1275,n1276,n1277);
xor (n1276,n1273,n1274);
and (n1277,n1278,n1279);
xor (n1278,n1231,n1232);
and (n1279,n201,n131);
or (n1280,n1281,n1284);
and (n1281,n1282,n1283);
xor (n1282,n1240,n1241);
and (n1283,n121,n28);
and (n1284,n1285,n1286);
xor (n1285,n1282,n1283);
or (n1286,n1287,n1290);
and (n1287,n1288,n1289);
xor (n1288,n1246,n1247);
and (n1289,n26,n28);
and (n1290,n1291,n1292);
xor (n1291,n1288,n1289);
or (n1292,n1293,n1296);
and (n1293,n1294,n1295);
xor (n1294,n1252,n1253);
and (n1295,n36,n28);
and (n1296,n1297,n1298);
xor (n1297,n1294,n1295);
or (n1298,n1299,n1301);
and (n1299,n1300,n292);
xor (n1300,n1258,n1259);
and (n1301,n1302,n1303);
xor (n1302,n1300,n292);
or (n1303,n1304,n1307);
and (n1304,n1305,n1306);
xor (n1305,n1264,n1265);
and (n1306,n96,n28);
and (n1307,n1308,n1309);
xor (n1308,n1305,n1306);
or (n1309,n1310,n1313);
and (n1310,n1311,n1312);
xor (n1311,n1270,n1271);
and (n1312,n95,n28);
and (n1313,n1314,n1315);
xor (n1314,n1311,n1312);
and (n1315,n1316,n1317);
xor (n1316,n1276,n1277);
and (n1317,n201,n28);
and (n1318,n121,n46);
or (n1319,n1320,n1322);
and (n1320,n1321,n47);
xor (n1321,n1285,n1286);
and (n1322,n1323,n1324);
xor (n1323,n1321,n47);
or (n1324,n1325,n1328);
and (n1325,n1326,n1327);
xor (n1326,n1291,n1292);
and (n1327,n36,n46);
and (n1328,n1329,n1330);
xor (n1329,n1326,n1327);
or (n1330,n1331,n1334);
and (n1331,n1332,n1333);
xor (n1332,n1297,n1298);
and (n1333,n35,n46);
and (n1334,n1335,n1336);
xor (n1335,n1332,n1333);
or (n1336,n1337,n1340);
and (n1337,n1338,n1339);
xor (n1338,n1302,n1303);
and (n1339,n96,n46);
and (n1340,n1341,n1342);
xor (n1341,n1338,n1339);
or (n1342,n1343,n1346);
and (n1343,n1344,n1345);
xor (n1344,n1308,n1309);
and (n1345,n95,n46);
and (n1346,n1347,n1348);
xor (n1347,n1344,n1345);
and (n1348,n1349,n1350);
xor (n1349,n1314,n1315);
and (n1350,n201,n46);
and (n1351,n26,n88);
or (n1352,n1353,n1356);
and (n1353,n1354,n1355);
xor (n1354,n1323,n1324);
and (n1355,n36,n88);
and (n1356,n1357,n1358);
xor (n1357,n1354,n1355);
or (n1358,n1359,n1361);
and (n1359,n1360,n89);
xor (n1360,n1329,n1330);
and (n1361,n1362,n1363);
xor (n1362,n1360,n89);
or (n1363,n1364,n1367);
and (n1364,n1365,n1366);
xor (n1365,n1335,n1336);
and (n1366,n96,n88);
and (n1367,n1368,n1369);
xor (n1368,n1365,n1366);
or (n1369,n1370,n1373);
and (n1370,n1371,n1372);
xor (n1371,n1341,n1342);
and (n1372,n95,n88);
and (n1373,n1374,n1375);
xor (n1374,n1371,n1372);
and (n1375,n1376,n1377);
xor (n1376,n1347,n1348);
and (n1377,n201,n88);
and (n1378,n36,n105);
or (n1379,n1380,n1382);
and (n1380,n1381,n104);
xor (n1381,n1357,n1358);
and (n1382,n1383,n1384);
xor (n1383,n1381,n104);
or (n1384,n1385,n1388);
and (n1385,n1386,n1387);
xor (n1386,n1362,n1363);
and (n1387,n96,n105);
and (n1388,n1389,n1390);
xor (n1389,n1386,n1387);
or (n1390,n1391,n1394);
and (n1391,n1392,n1393);
xor (n1392,n1368,n1369);
and (n1393,n95,n105);
and (n1394,n1395,n1396);
xor (n1395,n1392,n1393);
and (n1396,n1397,n1398);
xor (n1397,n1374,n1375);
and (n1398,n201,n105);
and (n1399,n35,n215);
or (n1400,n1401,n1404);
and (n1401,n1402,n1403);
xor (n1402,n1383,n1384);
and (n1403,n96,n215);
and (n1404,n1405,n1406);
xor (n1405,n1402,n1403);
or (n1406,n1407,n1410);
and (n1407,n1408,n1409);
xor (n1408,n1389,n1390);
and (n1409,n95,n215);
and (n1410,n1411,n1412);
xor (n1411,n1408,n1409);
and (n1412,n1413,n1414);
xor (n1413,n1395,n1396);
and (n1414,n201,n215);
and (n1415,n96,n197);
or (n1416,n1417,n1420);
and (n1417,n1418,n1419);
xor (n1418,n1405,n1406);
and (n1419,n95,n197);
and (n1420,n1421,n1422);
xor (n1421,n1418,n1419);
and (n1422,n1423,n1424);
xor (n1423,n1411,n1412);
and (n1424,n201,n197);
and (n1425,n95,n206);
and (n1426,n1427,n1428);
xor (n1427,n1421,n1422);
and (n1428,n201,n206);
and (n1429,n201,n819);
endmodule
