module top (out,n7,n10,n11,n15,n18,n19,n23,n29,n38
        ,n39,n76,n80,n94,n95,n148,n151,n190,n198,n199
        ,n245,n303,n304,n356,n361,n407,n408,n445,n514,n578
        ,n672,n745,n830);
output out;
input n7;
input n10;
input n11;
input n15;
input n18;
input n19;
input n23;
input n29;
input n38;
input n39;
input n76;
input n80;
input n94;
input n95;
input n148;
input n151;
input n190;
input n198;
input n199;
input n245;
input n303;
input n304;
input n356;
input n361;
input n407;
input n408;
input n445;
input n514;
input n578;
input n672;
input n745;
input n830;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n8;
wire n9;
wire n12;
wire n13;
wire n14;
wire n16;
wire n17;
wire n20;
wire n21;
wire n22;
wire n24;
wire n25;
wire n26;
wire n27;
wire n28;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n77;
wire n78;
wire n79;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n149;
wire n150;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n357;
wire n358;
wire n359;
wire n360;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
xor (out,n0,n1487);
xor (n0,n1,n123);
xor (n1,n2,n62);
xor (n2,n3,n55);
xor (n3,n4,n31);
or (n4,n5,n27,n30);
and (n5,n6,n12);
and (n6,n7,n8);
not (n8,n9);
and (n9,n10,n11);
xnor (n12,n13,n24);
nor (n13,n14,n22);
and (n14,n15,n16);
and (n16,n17,n20);
xor (n17,n18,n19);
not (n20,n21);
xor (n21,n19,n7);
and (n22,n23,n21);
and (n24,n18,n25);
not (n25,n26);
and (n26,n19,n7);
and (n27,n12,n28);
and (n28,n29,n18);
and (n30,n6,n28);
or (n31,n32,n53);
or (n32,n33,n47,n52);
and (n33,n34,n40);
not (n34,n35);
and (n35,n11,n36);
not (n36,n37);
and (n37,n38,n39);
xnor (n40,n41,n6);
not (n41,n42);
and (n42,n23,n43);
and (n43,n44,n45);
xor (n44,n7,n10);
not (n45,n46);
xor (n46,n10,n11);
and (n47,n40,n48);
xnor (n48,n49,n24);
nor (n49,n50,n51);
and (n50,n29,n16);
and (n51,n15,n21);
and (n52,n34,n48);
xor (n53,n54,n28);
xor (n54,n6,n12);
xor (n55,n56,n61);
xor (n56,n57,n58);
not (n57,n6);
xnor (n58,n59,n24);
not (n59,n60);
and (n60,n23,n16);
and (n61,n15,n18);
or (n62,n63,n120,n122);
and (n63,n64,n84);
or (n64,n65,n81,n83);
and (n65,n66,n79);
or (n66,n67,n72,n78);
and (n67,n35,n68);
xnor (n68,n69,n6);
nor (n69,n70,n71);
and (n70,n15,n43);
and (n71,n23,n46);
and (n72,n68,n73);
xnor (n73,n74,n24);
nor (n74,n75,n77);
and (n75,n76,n16);
and (n77,n29,n21);
and (n78,n35,n73);
and (n79,n80,n18);
and (n81,n79,n82);
and (n82,n76,n18);
and (n83,n66,n82);
or (n84,n85,n116,n119);
and (n85,n86,n114);
or (n86,n87,n111,n113);
and (n87,n88,n109);
or (n88,n89,n103,n108);
and (n89,n90,n96);
not (n90,n91);
and (n91,n39,n92);
not (n92,n93);
and (n93,n94,n95);
xnor (n96,n97,n35);
not (n97,n98);
and (n98,n23,n99);
and (n99,n100,n101);
xor (n100,n11,n38);
not (n101,n102);
xor (n102,n38,n39);
and (n103,n96,n104);
xnor (n104,n105,n6);
nor (n105,n106,n107);
and (n106,n29,n43);
and (n107,n15,n46);
and (n108,n90,n104);
xor (n109,n110,n73);
xor (n110,n35,n68);
and (n111,n109,n112);
not (n112,n79);
and (n113,n88,n112);
xor (n114,n115,n48);
xor (n115,n34,n40);
and (n116,n114,n117);
xor (n117,n118,n82);
xor (n118,n66,n79);
and (n119,n86,n117);
and (n120,n84,n121);
xnor (n121,n32,n53);
and (n122,n64,n121);
or (n123,n124,n168);
and (n124,n125,n127);
xor (n125,n126,n121);
xor (n126,n64,n84);
and (n127,n128,n166);
or (n128,n129,n162,n165);
and (n129,n130,n158);
or (n130,n131,n152,n157);
and (n131,n132,n144);
or (n132,n133,n138,n143);
and (n133,n91,n134);
xnor (n134,n135,n35);
nor (n135,n136,n137);
and (n136,n15,n99);
and (n137,n23,n102);
and (n138,n134,n139);
xnor (n139,n140,n6);
nor (n140,n141,n142);
and (n141,n76,n43);
and (n142,n29,n46);
and (n143,n91,n139);
or (n144,n145,n150);
xnor (n145,n146,n24);
nor (n146,n147,n149);
and (n147,n148,n16);
and (n149,n80,n21);
and (n150,n151,n18);
and (n152,n144,n153);
xnor (n153,n154,n24);
nor (n154,n155,n156);
and (n155,n80,n16);
and (n156,n76,n21);
and (n157,n132,n153);
and (n158,n159,n160);
and (n159,n148,n18);
xor (n160,n161,n104);
xor (n161,n90,n96);
and (n162,n158,n163);
xor (n163,n164,n112);
xor (n164,n88,n109);
and (n165,n130,n163);
xor (n166,n167,n117);
xor (n167,n86,n114);
and (n168,n169,n170);
xor (n169,n125,n127);
or (n170,n171,n223);
and (n171,n172,n173);
xor (n172,n128,n166);
and (n173,n174,n221);
or (n174,n175,n218,n220);
and (n175,n176,n216);
or (n176,n177,n213,n215);
and (n177,n178,n192);
or (n178,n179,n188,n191);
and (n179,n180,n184);
xnor (n180,n181,n6);
nor (n181,n182,n183);
and (n182,n80,n43);
and (n183,n76,n46);
xnor (n184,n185,n24);
nor (n185,n186,n187);
and (n186,n151,n16);
and (n187,n148,n21);
and (n188,n184,n189);
and (n189,n190,n18);
and (n191,n180,n189);
or (n192,n193,n207,n212);
and (n193,n194,n200);
not (n194,n195);
and (n195,n95,n196);
not (n196,n197);
and (n197,n198,n199);
xnor (n200,n201,n91);
not (n201,n202);
and (n202,n23,n203);
and (n203,n204,n205);
xor (n204,n39,n94);
not (n205,n206);
xor (n206,n94,n95);
and (n207,n200,n208);
xnor (n208,n209,n35);
nor (n209,n210,n211);
and (n210,n29,n99);
and (n211,n15,n102);
and (n212,n194,n208);
and (n213,n192,n214);
xnor (n214,n145,n150);
and (n215,n178,n214);
xor (n216,n217,n153);
xor (n217,n132,n144);
and (n218,n216,n219);
xor (n219,n159,n160);
and (n220,n176,n219);
xor (n221,n222,n163);
xor (n222,n130,n158);
and (n223,n224,n225);
xor (n224,n172,n173);
or (n225,n226,n271);
and (n226,n227,n228);
xor (n227,n174,n221);
and (n228,n229,n269);
or (n229,n230,n265,n268);
and (n230,n231,n263);
or (n231,n232,n259,n262);
and (n232,n233,n247);
or (n233,n234,n243,n246);
and (n234,n235,n239);
xnor (n235,n236,n6);
nor (n236,n237,n238);
and (n237,n148,n43);
and (n238,n80,n46);
xnor (n239,n240,n24);
nor (n240,n241,n242);
and (n241,n190,n16);
and (n242,n151,n21);
and (n243,n239,n244);
and (n244,n245,n18);
and (n246,n235,n244);
or (n247,n248,n253,n258);
and (n248,n195,n249);
xnor (n249,n250,n91);
nor (n250,n251,n252);
and (n251,n15,n203);
and (n252,n23,n206);
and (n253,n249,n254);
xnor (n254,n255,n35);
nor (n255,n256,n257);
and (n256,n76,n99);
and (n257,n29,n102);
and (n258,n195,n254);
and (n259,n247,n260);
xor (n260,n261,n189);
xor (n261,n180,n184);
and (n262,n233,n260);
xor (n263,n264,n139);
xor (n264,n91,n134);
and (n265,n263,n266);
xor (n266,n267,n214);
xor (n267,n178,n192);
and (n268,n231,n266);
xor (n269,n270,n219);
xor (n270,n176,n216);
and (n271,n272,n273);
xor (n272,n227,n228);
or (n273,n274,n388);
and (n274,n275,n276);
xor (n275,n229,n269);
or (n276,n277,n384,n387);
and (n277,n278,n324);
or (n278,n279,n320,n323);
and (n279,n280,n318);
or (n280,n281,n297);
or (n281,n282,n291,n296);
and (n282,n283,n287);
xnor (n283,n284,n35);
nor (n284,n285,n286);
and (n285,n80,n99);
and (n286,n76,n102);
xnor (n287,n288,n6);
nor (n288,n289,n290);
and (n289,n151,n43);
and (n290,n148,n46);
and (n291,n287,n292);
xnor (n292,n293,n24);
nor (n293,n294,n295);
and (n294,n245,n16);
and (n295,n190,n21);
and (n296,n283,n292);
or (n297,n298,n312,n317);
and (n298,n299,n305);
not (n299,n300);
and (n300,n199,n301);
not (n301,n302);
and (n302,n303,n304);
xnor (n305,n306,n195);
not (n306,n307);
and (n307,n23,n308);
and (n308,n309,n310);
xor (n309,n95,n198);
not (n310,n311);
xor (n311,n198,n199);
and (n312,n305,n313);
xnor (n313,n314,n91);
nor (n314,n315,n316);
and (n315,n29,n203);
and (n316,n15,n206);
and (n317,n299,n313);
xor (n318,n319,n208);
xor (n319,n194,n200);
and (n320,n318,n321);
xor (n321,n322,n260);
xor (n322,n233,n247);
and (n323,n280,n321);
or (n324,n325,n380,n383);
and (n325,n326,n376);
or (n326,n327,n372,n375);
and (n327,n328,n363);
or (n328,n329,n359,n362);
and (n329,n330,n342);
or (n330,n331,n336,n341);
and (n331,n300,n332);
xnor (n332,n333,n195);
nor (n333,n334,n335);
and (n334,n15,n308);
and (n335,n23,n311);
and (n336,n332,n337);
xnor (n337,n338,n91);
nor (n338,n339,n340);
and (n339,n76,n203);
and (n340,n29,n206);
and (n341,n300,n337);
or (n342,n343,n352,n358);
and (n343,n344,n348);
xnor (n344,n345,n35);
nor (n345,n346,n347);
and (n346,n148,n99);
and (n347,n80,n102);
xnor (n348,n349,n6);
nor (n349,n350,n351);
and (n350,n190,n43);
and (n351,n151,n46);
and (n352,n348,n353);
xnor (n353,n354,n24);
nor (n354,n355,n357);
and (n355,n356,n16);
and (n357,n245,n21);
and (n358,n344,n353);
and (n359,n342,n360);
and (n360,n361,n18);
and (n362,n330,n360);
or (n363,n364,n368,n371);
and (n364,n365,n366);
and (n365,n356,n18);
xor (n366,n367,n292);
xor (n367,n283,n287);
and (n368,n366,n369);
xor (n369,n370,n313);
xor (n370,n299,n305);
and (n371,n365,n369);
and (n372,n363,n373);
xor (n373,n374,n244);
xor (n374,n235,n239);
and (n375,n328,n373);
and (n376,n377,n379);
xor (n377,n378,n254);
xor (n378,n195,n249);
xnor (n379,n281,n297);
and (n380,n376,n381);
xor (n381,n382,n321);
xor (n382,n280,n318);
and (n383,n326,n381);
and (n384,n324,n385);
xor (n385,n386,n266);
xor (n386,n231,n263);
and (n387,n278,n385);
and (n388,n389,n390);
xor (n389,n275,n276);
or (n390,n391,n467);
and (n391,n392,n394);
xor (n392,n393,n385);
xor (n393,n278,n324);
and (n394,n395,n465);
or (n395,n396,n462,n464);
and (n396,n397,n460);
or (n397,n398,n456,n459);
and (n398,n399,n447);
or (n399,n400,n438,n446);
and (n400,n401,n422);
or (n401,n402,n416,n421);
and (n402,n403,n409);
not (n403,n404);
and (n404,n304,n405);
not (n405,n406);
and (n406,n407,n408);
xnor (n409,n410,n300);
not (n410,n411);
and (n411,n23,n412);
and (n412,n413,n414);
xor (n413,n199,n303);
not (n414,n415);
xor (n415,n303,n304);
and (n416,n409,n417);
xnor (n417,n418,n195);
nor (n418,n419,n420);
and (n419,n29,n308);
and (n420,n15,n311);
and (n421,n403,n417);
or (n422,n423,n432,n437);
and (n423,n424,n428);
xnor (n424,n425,n91);
nor (n425,n426,n427);
and (n426,n80,n203);
and (n427,n76,n206);
xnor (n428,n429,n35);
nor (n429,n430,n431);
and (n430,n151,n99);
and (n431,n148,n102);
and (n432,n428,n433);
xnor (n433,n434,n6);
nor (n434,n435,n436);
and (n435,n245,n43);
and (n436,n190,n46);
and (n437,n424,n433);
and (n438,n422,n439);
and (n439,n440,n444);
xnor (n440,n441,n24);
nor (n441,n442,n443);
and (n442,n361,n16);
and (n443,n356,n21);
and (n444,n445,n18);
and (n446,n401,n439);
or (n447,n448,n453,n455);
and (n448,n449,n451);
xor (n449,n450,n337);
xor (n450,n300,n332);
xor (n451,n452,n353);
xor (n452,n344,n348);
and (n453,n451,n454);
not (n454,n360);
and (n455,n449,n454);
and (n456,n447,n457);
xor (n457,n458,n369);
xor (n458,n365,n366);
and (n459,n399,n457);
xor (n460,n461,n373);
xor (n461,n328,n363);
and (n462,n460,n463);
xor (n463,n377,n379);
and (n464,n397,n463);
xor (n465,n466,n381);
xor (n466,n326,n376);
and (n467,n468,n469);
xor (n468,n392,n394);
or (n469,n470,n538);
and (n470,n471,n472);
xor (n471,n395,n465);
and (n472,n473,n536);
or (n473,n474,n532,n535);
and (n474,n475,n530);
or (n475,n476,n525,n529);
and (n476,n477,n516);
or (n477,n478,n507,n515);
and (n478,n479,n491);
or (n479,n480,n485,n490);
and (n480,n404,n481);
xnor (n481,n482,n300);
nor (n482,n483,n484);
and (n483,n15,n412);
and (n484,n23,n415);
and (n485,n481,n486);
xnor (n486,n487,n195);
nor (n487,n488,n489);
and (n488,n76,n308);
and (n489,n29,n311);
and (n490,n404,n486);
or (n491,n492,n501,n506);
and (n492,n493,n497);
xnor (n493,n494,n91);
nor (n494,n495,n496);
and (n495,n148,n203);
and (n496,n80,n206);
xnor (n497,n498,n35);
nor (n498,n499,n500);
and (n499,n190,n99);
and (n500,n151,n102);
and (n501,n497,n502);
xnor (n502,n503,n6);
nor (n503,n504,n505);
and (n504,n356,n43);
and (n505,n245,n46);
and (n506,n493,n502);
and (n507,n491,n508);
or (n508,n509,n513);
xnor (n509,n510,n24);
nor (n510,n511,n512);
and (n511,n445,n16);
and (n512,n361,n21);
and (n513,n514,n18);
and (n515,n479,n508);
or (n516,n517,n522,n524);
and (n517,n518,n520);
xor (n518,n519,n417);
xor (n519,n403,n409);
xor (n520,n521,n433);
xor (n521,n424,n428);
and (n522,n520,n523);
xor (n523,n440,n444);
and (n524,n518,n523);
and (n525,n516,n526);
xor (n526,n527,n451);
xor (n527,n360,n528);
not (n528,n449);
and (n529,n477,n526);
xor (n530,n531,n360);
xor (n531,n330,n342);
and (n532,n530,n533);
xor (n533,n534,n457);
xor (n534,n399,n447);
and (n535,n475,n533);
xor (n536,n537,n463);
xor (n537,n397,n460);
and (n538,n539,n540);
xor (n539,n471,n472);
or (n540,n541,n619);
and (n541,n542,n543);
xor (n542,n473,n536);
and (n543,n544,n617);
or (n544,n545,n613,n616);
and (n545,n546,n611);
or (n546,n547,n607,n610);
and (n547,n548,n598);
or (n548,n549,n580,n597);
and (n549,n550,n566);
or (n550,n551,n560,n565);
and (n551,n552,n553);
not (n552,n408);
xnor (n553,n554,n404);
not (n554,n555);
and (n555,n23,n556);
and (n556,n557,n558);
xor (n557,n304,n407);
not (n558,n559);
xor (n559,n407,n408);
and (n560,n553,n561);
xnor (n561,n562,n300);
nor (n562,n563,n564);
and (n563,n29,n412);
and (n564,n15,n415);
and (n565,n552,n561);
or (n566,n567,n576,n579);
and (n567,n568,n572);
xnor (n568,n569,n6);
nor (n569,n570,n571);
and (n570,n361,n43);
and (n571,n356,n46);
xnor (n572,n573,n24);
nor (n573,n574,n575);
and (n574,n514,n16);
and (n575,n445,n21);
and (n576,n572,n577);
and (n577,n578,n18);
and (n579,n568,n577);
and (n580,n566,n581);
or (n581,n582,n591,n596);
and (n582,n583,n587);
xnor (n583,n584,n195);
nor (n584,n585,n586);
and (n585,n80,n308);
and (n586,n76,n311);
xnor (n587,n588,n91);
nor (n588,n589,n590);
and (n589,n151,n203);
and (n590,n148,n206);
and (n591,n587,n592);
xnor (n592,n593,n35);
nor (n593,n594,n595);
and (n594,n245,n99);
and (n595,n190,n102);
and (n596,n583,n592);
and (n597,n550,n581);
or (n598,n599,n604,n606);
and (n599,n600,n602);
xor (n600,n601,n486);
xor (n601,n404,n481);
xor (n602,n603,n502);
xor (n603,n493,n497);
and (n604,n602,n605);
xnor (n605,n509,n513);
and (n606,n600,n605);
and (n607,n598,n608);
xor (n608,n609,n523);
xor (n609,n518,n520);
and (n610,n548,n608);
xor (n611,n612,n439);
xor (n612,n401,n422);
and (n613,n611,n614);
xor (n614,n615,n526);
xor (n615,n477,n516);
and (n616,n546,n614);
xor (n617,n618,n533);
xor (n618,n475,n530);
and (n619,n620,n621);
xor (n620,n542,n543);
or (n621,n622,n694);
and (n622,n623,n624);
xor (n623,n544,n617);
and (n624,n625,n692);
or (n625,n626,n688,n691);
and (n626,n627,n686);
or (n627,n628,n680,n685);
and (n628,n629,n675);
or (n629,n630,n659,n674);
and (n630,n631,n647);
or (n631,n632,n641,n646);
and (n632,n633,n637);
xnor (n633,n634,n195);
nor (n634,n635,n636);
and (n635,n148,n308);
and (n636,n80,n311);
xnor (n637,n638,n91);
nor (n638,n639,n640);
and (n639,n190,n203);
and (n640,n151,n206);
and (n641,n637,n642);
xnor (n642,n643,n35);
nor (n643,n644,n645);
and (n644,n356,n99);
and (n645,n245,n102);
and (n646,n633,n642);
or (n647,n648,n653,n658);
and (n648,n408,n649);
xnor (n649,n650,n404);
nor (n650,n651,n652);
and (n651,n15,n556);
and (n652,n23,n559);
and (n653,n649,n654);
xnor (n654,n655,n300);
nor (n655,n656,n657);
and (n656,n76,n412);
and (n657,n29,n415);
and (n658,n408,n654);
and (n659,n647,n660);
or (n660,n661,n670,n673);
and (n661,n662,n666);
xnor (n662,n663,n6);
nor (n663,n664,n665);
and (n664,n445,n43);
and (n665,n361,n46);
xnor (n666,n667,n24);
nor (n667,n668,n669);
and (n668,n578,n16);
and (n669,n514,n21);
and (n670,n666,n671);
and (n671,n672,n18);
and (n673,n662,n671);
and (n674,n631,n660);
or (n675,n676,n678);
xor (n676,n677,n577);
xor (n677,n568,n572);
xor (n678,n679,n592);
xor (n679,n583,n587);
and (n680,n675,n681);
xor (n681,n682,n684);
xor (n682,n683,n602);
not (n683,n600);
not (n684,n605);
and (n685,n629,n681);
xor (n686,n687,n508);
xor (n687,n479,n491);
and (n688,n686,n689);
xor (n689,n690,n608);
xor (n690,n548,n598);
and (n691,n627,n689);
xor (n692,n693,n614);
xor (n693,n546,n611);
and (n694,n695,n696);
xor (n695,n623,n624);
or (n696,n697,n776);
and (n697,n698,n699);
xor (n698,n625,n692);
and (n699,n700,n774);
or (n700,n701,n770,n773);
and (n701,n702,n766);
or (n702,n703,n762,n765);
and (n703,n704,n752);
or (n704,n705,n738,n751);
and (n705,n706,n722);
or (n706,n707,n716,n721);
and (n707,n708,n712);
xnor (n708,n709,n300);
nor (n709,n710,n711);
and (n710,n80,n412);
and (n711,n76,n415);
xnor (n712,n713,n195);
nor (n713,n714,n715);
and (n714,n151,n308);
and (n715,n148,n311);
and (n716,n712,n717);
xnor (n717,n718,n91);
nor (n718,n719,n720);
and (n719,n245,n203);
and (n720,n190,n206);
and (n721,n708,n717);
or (n722,n723,n732,n737);
and (n723,n724,n728);
xnor (n724,n725,n35);
nor (n725,n726,n727);
and (n726,n361,n99);
and (n727,n356,n102);
xnor (n728,n729,n6);
nor (n729,n730,n731);
and (n730,n514,n43);
and (n731,n445,n46);
and (n732,n728,n733);
xnor (n733,n734,n24);
nor (n734,n735,n736);
and (n735,n672,n16);
and (n736,n578,n21);
and (n737,n724,n733);
and (n738,n722,n739);
and (n739,n740,n747);
xnor (n740,n741,n408);
not (n741,n742);
and (n742,n23,n743);
and (n743,n744,n746);
xor (n744,n408,n745);
not (n746,n745);
xnor (n747,n748,n404);
nor (n748,n749,n750);
and (n749,n29,n556);
and (n750,n15,n559);
and (n751,n706,n739);
or (n752,n753,n758,n761);
and (n753,n754,n756);
xor (n754,n755,n642);
xor (n755,n633,n637);
xor (n756,n757,n654);
xor (n757,n408,n649);
and (n758,n756,n759);
xor (n759,n760,n671);
xor (n760,n662,n666);
and (n761,n754,n759);
and (n762,n752,n763);
xor (n763,n764,n561);
xor (n764,n552,n553);
and (n765,n704,n763);
and (n766,n767,n769);
xor (n767,n768,n660);
xor (n768,n631,n647);
xnor (n769,n676,n678);
and (n770,n766,n771);
xor (n771,n772,n581);
xor (n772,n550,n566);
and (n773,n702,n771);
xor (n774,n775,n689);
xor (n775,n627,n686);
and (n776,n777,n778);
xor (n777,n698,n699);
or (n778,n779,n858);
and (n779,n780,n781);
xor (n780,n700,n774);
or (n781,n782,n854,n857);
and (n782,n783,n852);
or (n783,n784,n849,n851);
and (n784,n785,n847);
or (n785,n786,n843,n846);
and (n786,n787,n833);
or (n787,n788,n821,n832);
and (n788,n789,n805);
or (n789,n790,n799,n804);
and (n790,n791,n795);
xnor (n791,n792,n408);
nor (n792,n793,n794);
and (n793,n15,n743);
and (n794,n23,n745);
xnor (n795,n796,n404);
nor (n796,n797,n798);
and (n797,n76,n556);
and (n798,n29,n559);
and (n799,n795,n800);
xnor (n800,n801,n300);
nor (n801,n802,n803);
and (n802,n148,n412);
and (n803,n80,n415);
and (n804,n791,n800);
or (n805,n806,n815,n820);
and (n806,n807,n811);
xnor (n807,n808,n195);
nor (n808,n809,n810);
and (n809,n190,n308);
and (n810,n151,n311);
xnor (n811,n812,n91);
nor (n812,n813,n814);
and (n813,n356,n203);
and (n814,n245,n206);
and (n815,n811,n816);
xnor (n816,n817,n35);
nor (n817,n818,n819);
and (n818,n445,n99);
and (n819,n361,n102);
and (n820,n807,n816);
and (n821,n805,n822);
and (n822,n823,n827);
xnor (n823,n824,n6);
nor (n824,n825,n826);
and (n825,n578,n43);
and (n826,n514,n46);
xnor (n827,n828,n24);
nor (n828,n829,n831);
and (n829,n830,n16);
and (n831,n672,n21);
and (n832,n789,n822);
or (n833,n834,n839,n842);
and (n834,n835,n837);
not (n835,n836);
nand (n836,n830,n18);
xor (n837,n838,n717);
xor (n838,n708,n712);
and (n839,n837,n840);
xor (n840,n841,n733);
xor (n841,n724,n728);
and (n842,n835,n840);
and (n843,n833,n844);
xor (n844,n845,n759);
xor (n845,n754,n756);
and (n846,n787,n844);
xor (n847,n848,n763);
xor (n848,n704,n752);
and (n849,n847,n850);
xor (n850,n767,n769);
and (n851,n785,n850);
xor (n852,n853,n771);
xor (n853,n702,n766);
and (n854,n852,n855);
xor (n855,n856,n681);
xor (n856,n629,n675);
and (n857,n783,n855);
and (n858,n859,n860);
xor (n859,n780,n781);
or (n860,n861,n938);
and (n861,n862,n864);
xor (n862,n863,n855);
xor (n863,n783,n852);
and (n864,n865,n936);
or (n865,n866,n932,n935);
and (n866,n867,n927);
or (n867,n868,n924,n926);
and (n868,n869,n915);
or (n869,n870,n897,n914);
and (n870,n871,n885);
or (n871,n872,n881,n884);
and (n872,n873,n877);
xnor (n873,n874,n35);
nor (n874,n875,n876);
and (n875,n514,n99);
and (n876,n445,n102);
xnor (n877,n878,n6);
nor (n878,n879,n880);
and (n879,n672,n43);
and (n880,n578,n46);
and (n881,n877,n882);
xnor (n882,n883,n24);
nand (n883,n830,n21);
and (n884,n873,n882);
or (n885,n886,n895,n896);
and (n886,n887,n891);
xnor (n887,n888,n408);
nor (n888,n889,n890);
and (n889,n29,n743);
and (n890,n15,n745);
xnor (n891,n892,n404);
nor (n892,n893,n894);
and (n893,n80,n556);
and (n894,n76,n559);
and (n895,n891,n24);
and (n896,n887,n24);
and (n897,n885,n898);
or (n898,n899,n908,n913);
and (n899,n900,n904);
xnor (n900,n901,n300);
nor (n901,n902,n903);
and (n902,n151,n412);
and (n903,n148,n415);
xnor (n904,n905,n195);
nor (n905,n906,n907);
and (n906,n245,n308);
and (n907,n190,n311);
and (n908,n904,n909);
xnor (n909,n910,n91);
nor (n910,n911,n912);
and (n911,n361,n203);
and (n912,n356,n206);
and (n913,n900,n909);
and (n914,n871,n898);
or (n915,n916,n921,n923);
and (n916,n917,n919);
xor (n917,n918,n800);
xor (n918,n791,n795);
xor (n919,n920,n816);
xor (n920,n807,n811);
and (n921,n919,n922);
xor (n922,n823,n827);
and (n923,n917,n922);
and (n924,n915,n925);
xor (n925,n740,n747);
and (n926,n869,n925);
and (n927,n928,n930);
xor (n928,n929,n822);
xor (n929,n789,n805);
xor (n930,n931,n840);
xor (n931,n835,n837);
and (n932,n927,n933);
xor (n933,n934,n739);
xor (n934,n706,n722);
and (n935,n867,n933);
xor (n936,n937,n850);
xor (n937,n785,n847);
and (n938,n939,n940);
xor (n939,n862,n864);
or (n940,n941,n948);
and (n941,n942,n943);
xor (n942,n865,n936);
and (n943,n944,n946);
xor (n944,n945,n933);
xor (n945,n867,n927);
xor (n946,n947,n844);
xor (n947,n787,n833);
and (n948,n949,n950);
xor (n949,n942,n943);
or (n950,n951,n1014);
and (n951,n952,n958);
xor (n952,n953,n956);
xor (n953,n933,n954);
xor (n954,n947,n955);
not (n955,n756);
xor (n956,n945,n957);
xnor (n957,n754,n759);
or (n958,n959,n1011,n1013);
and (n959,n960,n1009);
or (n960,n961,n1005,n1008);
and (n961,n962,n1000);
or (n962,n963,n996,n999);
and (n963,n964,n980);
or (n964,n965,n974,n979);
and (n965,n966,n970);
xnor (n966,n967,n408);
nor (n967,n968,n969);
and (n968,n76,n743);
and (n969,n29,n745);
xnor (n970,n971,n404);
nor (n971,n972,n973);
and (n972,n148,n556);
and (n973,n80,n559);
and (n974,n970,n975);
xnor (n975,n976,n300);
nor (n976,n977,n978);
and (n977,n190,n412);
and (n978,n151,n415);
and (n979,n966,n975);
or (n980,n981,n990,n995);
and (n981,n982,n986);
xnor (n982,n983,n195);
nor (n983,n984,n985);
and (n984,n356,n308);
and (n985,n245,n311);
xnor (n986,n987,n91);
nor (n987,n988,n989);
and (n988,n445,n203);
and (n989,n361,n206);
and (n990,n986,n991);
xnor (n991,n992,n35);
nor (n992,n993,n994);
and (n993,n578,n99);
and (n994,n514,n102);
and (n995,n982,n991);
and (n996,n980,n997);
xor (n997,n998,n882);
xor (n998,n873,n877);
and (n999,n964,n997);
and (n1000,n1001,n1003);
xor (n1001,n1002,n24);
xor (n1002,n887,n891);
xor (n1003,n1004,n909);
xor (n1004,n900,n904);
and (n1005,n1000,n1006);
xor (n1006,n1007,n922);
xor (n1007,n917,n919);
and (n1008,n962,n1006);
xor (n1009,n1010,n925);
xor (n1010,n869,n915);
and (n1011,n1009,n1012);
xor (n1012,n928,n930);
and (n1013,n960,n1012);
and (n1014,n1015,n1016);
xor (n1015,n952,n958);
or (n1016,n1017,n1071);
and (n1017,n1018,n1020);
xor (n1018,n1019,n1012);
xor (n1019,n960,n1009);
or (n1020,n1021,n1067,n1070);
and (n1021,n1022,n1065);
or (n1022,n1023,n1062,n1064);
and (n1023,n1024,n1060);
or (n1024,n1025,n1054,n1059);
and (n1025,n1026,n1038);
or (n1026,n1027,n1036,n1037);
and (n1027,n1028,n1032);
xnor (n1028,n1029,n408);
nor (n1029,n1030,n1031);
and (n1030,n80,n743);
and (n1031,n76,n745);
xnor (n1032,n1033,n404);
nor (n1033,n1034,n1035);
and (n1034,n151,n556);
and (n1035,n148,n559);
and (n1036,n1032,n6);
and (n1037,n1028,n6);
or (n1038,n1039,n1048,n1053);
and (n1039,n1040,n1044);
xnor (n1040,n1041,n300);
nor (n1041,n1042,n1043);
and (n1042,n245,n412);
and (n1043,n190,n415);
xnor (n1044,n1045,n195);
nor (n1045,n1046,n1047);
and (n1046,n361,n308);
and (n1047,n356,n311);
and (n1048,n1044,n1049);
xnor (n1049,n1050,n91);
nor (n1050,n1051,n1052);
and (n1051,n514,n203);
and (n1052,n445,n206);
and (n1053,n1040,n1049);
and (n1054,n1038,n1055);
xnor (n1055,n1056,n6);
nor (n1056,n1057,n1058);
and (n1057,n830,n43);
and (n1058,n672,n46);
and (n1059,n1026,n1055);
xor (n1060,n1061,n997);
xor (n1061,n964,n980);
and (n1062,n1060,n1063);
xor (n1063,n1001,n1003);
and (n1064,n1024,n1063);
xor (n1065,n1066,n898);
xor (n1066,n871,n885);
and (n1067,n1065,n1068);
xor (n1068,n1069,n1006);
xor (n1069,n962,n1000);
and (n1070,n1022,n1068);
and (n1071,n1072,n1073);
xor (n1072,n1018,n1020);
or (n1073,n1074,n1144);
and (n1074,n1075,n1077);
xor (n1075,n1076,n1068);
xor (n1076,n1022,n1065);
or (n1077,n1078,n1140,n1143);
and (n1078,n1079,n1135);
or (n1079,n1080,n1131,n1134);
and (n1080,n1081,n1121);
or (n1081,n1082,n1115,n1120);
and (n1082,n1083,n1099);
or (n1083,n1084,n1093,n1098);
and (n1084,n1085,n1089);
xnor (n1085,n1086,n195);
nor (n1086,n1087,n1088);
and (n1087,n445,n308);
and (n1088,n361,n311);
xnor (n1089,n1090,n91);
nor (n1090,n1091,n1092);
and (n1091,n578,n203);
and (n1092,n514,n206);
and (n1093,n1089,n1094);
xnor (n1094,n1095,n35);
nor (n1095,n1096,n1097);
and (n1096,n830,n99);
and (n1097,n672,n102);
and (n1098,n1085,n1094);
or (n1099,n1100,n1109,n1114);
and (n1100,n1101,n1105);
xnor (n1101,n1102,n408);
nor (n1102,n1103,n1104);
and (n1103,n148,n743);
and (n1104,n80,n745);
xnor (n1105,n1106,n404);
nor (n1106,n1107,n1108);
and (n1107,n190,n556);
and (n1108,n151,n559);
and (n1109,n1105,n1110);
xnor (n1110,n1111,n300);
nor (n1111,n1112,n1113);
and (n1112,n356,n412);
and (n1113,n245,n415);
and (n1114,n1101,n1110);
and (n1115,n1099,n1116);
xnor (n1116,n1117,n35);
nor (n1117,n1118,n1119);
and (n1118,n672,n99);
and (n1119,n578,n102);
and (n1120,n1083,n1116);
or (n1121,n1122,n1127,n1130);
and (n1122,n1123,n1125);
xnor (n1123,n1124,n6);
nand (n1124,n830,n46);
xor (n1125,n1126,n6);
xor (n1126,n1028,n1032);
and (n1127,n1125,n1128);
xor (n1128,n1129,n1049);
xor (n1129,n1040,n1044);
and (n1130,n1123,n1128);
and (n1131,n1121,n1132);
xor (n1132,n1133,n991);
xor (n1133,n982,n986);
and (n1134,n1081,n1132);
and (n1135,n1136,n1138);
xor (n1136,n1137,n975);
xor (n1137,n966,n970);
xor (n1138,n1139,n1055);
xor (n1139,n1026,n1038);
and (n1140,n1135,n1141);
xor (n1141,n1142,n1063);
xor (n1142,n1024,n1060);
and (n1143,n1079,n1141);
and (n1144,n1145,n1146);
xor (n1145,n1075,n1077);
or (n1146,n1147,n1199);
and (n1147,n1148,n1150);
xor (n1148,n1149,n1141);
xor (n1149,n1079,n1135);
or (n1150,n1151,n1196,n1198);
and (n1151,n1152,n1194);
or (n1152,n1153,n1190,n1193);
and (n1153,n1154,n1188);
or (n1154,n1155,n1184,n1187);
and (n1155,n1156,n1172);
or (n1156,n1157,n1166,n1171);
and (n1157,n1158,n1162);
xnor (n1158,n1159,n300);
nor (n1159,n1160,n1161);
and (n1160,n361,n412);
and (n1161,n356,n415);
xnor (n1162,n1163,n195);
nor (n1163,n1164,n1165);
and (n1164,n514,n308);
and (n1165,n445,n311);
and (n1166,n1162,n1167);
xnor (n1167,n1168,n91);
nor (n1168,n1169,n1170);
and (n1169,n672,n203);
and (n1170,n578,n206);
and (n1171,n1158,n1167);
or (n1172,n1173,n1182,n1183);
and (n1173,n1174,n1178);
xnor (n1174,n1175,n408);
nor (n1175,n1176,n1177);
and (n1176,n151,n743);
and (n1177,n148,n745);
xnor (n1178,n1179,n404);
nor (n1179,n1180,n1181);
and (n1180,n245,n556);
and (n1181,n190,n559);
and (n1182,n1178,n35);
and (n1183,n1174,n35);
and (n1184,n1172,n1185);
xor (n1185,n1186,n1094);
xor (n1186,n1085,n1089);
and (n1187,n1156,n1185);
xor (n1188,n1189,n1116);
xor (n1189,n1083,n1099);
and (n1190,n1188,n1191);
xor (n1191,n1192,n1128);
xor (n1192,n1123,n1125);
and (n1193,n1154,n1191);
xor (n1194,n1195,n1132);
xor (n1195,n1081,n1121);
and (n1196,n1194,n1197);
xor (n1197,n1136,n1138);
and (n1198,n1152,n1197);
and (n1199,n1200,n1201);
xor (n1200,n1148,n1150);
or (n1201,n1202,n1240);
and (n1202,n1203,n1205);
xor (n1203,n1204,n1197);
xor (n1204,n1152,n1194);
and (n1205,n1206,n1238);
or (n1206,n1207,n1234,n1237);
and (n1207,n1208,n1232);
or (n1208,n1209,n1228,n1231);
and (n1209,n1210,n1226);
or (n1210,n1211,n1220,n1225);
and (n1211,n1212,n1216);
xnor (n1212,n1213,n408);
nor (n1213,n1214,n1215);
and (n1214,n190,n743);
and (n1215,n151,n745);
xnor (n1216,n1217,n404);
nor (n1217,n1218,n1219);
and (n1218,n356,n556);
and (n1219,n245,n559);
and (n1220,n1216,n1221);
xnor (n1221,n1222,n300);
nor (n1222,n1223,n1224);
and (n1223,n445,n412);
and (n1224,n361,n415);
and (n1225,n1212,n1221);
xnor (n1226,n1227,n35);
nand (n1227,n830,n102);
and (n1228,n1226,n1229);
xor (n1229,n1230,n1167);
xor (n1230,n1158,n1162);
and (n1231,n1210,n1229);
xor (n1232,n1233,n1110);
xor (n1233,n1101,n1105);
and (n1234,n1232,n1235);
xor (n1235,n1236,n1185);
xor (n1236,n1156,n1172);
and (n1237,n1208,n1235);
xor (n1238,n1239,n1191);
xor (n1239,n1154,n1188);
and (n1240,n1241,n1242);
xor (n1241,n1203,n1205);
or (n1242,n1243,n1295);
and (n1243,n1244,n1245);
xor (n1244,n1206,n1238);
and (n1245,n1246,n1293);
or (n1246,n1247,n1289,n1292);
and (n1247,n1248,n1282);
or (n1248,n1249,n1276,n1281);
and (n1249,n1250,n1264);
or (n1250,n1251,n1260,n1263);
and (n1251,n1252,n1256);
xnor (n1252,n1253,n300);
nor (n1253,n1254,n1255);
and (n1254,n514,n412);
and (n1255,n445,n415);
xnor (n1256,n1257,n195);
nor (n1257,n1258,n1259);
and (n1258,n672,n308);
and (n1259,n578,n311);
and (n1260,n1256,n1261);
xnor (n1261,n1262,n91);
nand (n1262,n830,n206);
and (n1263,n1252,n1261);
or (n1264,n1265,n1274,n1275);
and (n1265,n1266,n1270);
xnor (n1266,n1267,n408);
nor (n1267,n1268,n1269);
and (n1268,n245,n743);
and (n1269,n190,n745);
xnor (n1270,n1271,n404);
nor (n1271,n1272,n1273);
and (n1272,n361,n556);
and (n1273,n356,n559);
and (n1274,n1270,n91);
and (n1275,n1266,n91);
and (n1276,n1264,n1277);
xnor (n1277,n1278,n195);
nor (n1278,n1279,n1280);
and (n1279,n578,n308);
and (n1280,n514,n311);
and (n1281,n1250,n1277);
and (n1282,n1283,n1287);
xnor (n1283,n1284,n91);
nor (n1284,n1285,n1286);
and (n1285,n830,n203);
and (n1286,n672,n206);
xor (n1287,n1288,n1221);
xor (n1288,n1212,n1216);
and (n1289,n1282,n1290);
xor (n1290,n1291,n35);
xor (n1291,n1174,n1178);
and (n1292,n1248,n1290);
xor (n1293,n1294,n1235);
xor (n1294,n1208,n1232);
and (n1295,n1296,n1297);
xor (n1296,n1244,n1245);
or (n1297,n1298,n1305);
and (n1298,n1299,n1300);
xor (n1299,n1246,n1293);
and (n1300,n1301,n1303);
xor (n1301,n1302,n1229);
xor (n1302,n1210,n1226);
xor (n1303,n1304,n1290);
xor (n1304,n1248,n1282);
and (n1305,n1306,n1307);
xor (n1306,n1299,n1300);
or (n1307,n1308,n1341);
and (n1308,n1309,n1310);
xor (n1309,n1301,n1303);
or (n1310,n1311,n1338,n1340);
and (n1311,n1312,n1336);
or (n1312,n1313,n1332,n1335);
and (n1313,n1314,n1330);
or (n1314,n1315,n1324,n1329);
and (n1315,n1316,n1320);
xnor (n1316,n1317,n408);
nor (n1317,n1318,n1319);
and (n1318,n356,n743);
and (n1319,n245,n745);
xnor (n1320,n1321,n404);
nor (n1321,n1322,n1323);
and (n1322,n445,n556);
and (n1323,n361,n559);
and (n1324,n1320,n1325);
xnor (n1325,n1326,n300);
nor (n1326,n1327,n1328);
and (n1327,n578,n412);
and (n1328,n514,n415);
and (n1329,n1316,n1325);
xor (n1330,n1331,n1261);
xor (n1331,n1252,n1256);
and (n1332,n1330,n1333);
xor (n1333,n1334,n91);
xor (n1334,n1266,n1270);
and (n1335,n1314,n1333);
xor (n1336,n1337,n1277);
xor (n1337,n1250,n1264);
and (n1338,n1336,n1339);
xor (n1339,n1283,n1287);
and (n1340,n1312,n1339);
and (n1341,n1342,n1343);
xor (n1342,n1309,n1310);
or (n1343,n1344,n1377);
and (n1344,n1345,n1347);
xor (n1345,n1346,n1339);
xor (n1346,n1312,n1336);
and (n1347,n1348,n1375);
or (n1348,n1349,n1369,n1374);
and (n1349,n1350,n1362);
or (n1350,n1351,n1360,n1361);
and (n1351,n1352,n1356);
xnor (n1352,n1353,n408);
nor (n1353,n1354,n1355);
and (n1354,n361,n743);
and (n1355,n356,n745);
xnor (n1356,n1357,n404);
nor (n1357,n1358,n1359);
and (n1358,n514,n556);
and (n1359,n445,n559);
and (n1360,n1356,n195);
and (n1361,n1352,n195);
and (n1362,n1363,n1367);
xnor (n1363,n1364,n300);
nor (n1364,n1365,n1366);
and (n1365,n672,n412);
and (n1366,n578,n415);
xnor (n1367,n1368,n195);
nand (n1368,n830,n311);
and (n1369,n1362,n1370);
xnor (n1370,n1371,n195);
nor (n1371,n1372,n1373);
and (n1372,n830,n308);
and (n1373,n672,n311);
and (n1374,n1350,n1370);
xor (n1375,n1376,n1333);
xor (n1376,n1314,n1330);
and (n1377,n1378,n1379);
xor (n1378,n1345,n1347);
or (n1379,n1380,n1387);
and (n1380,n1381,n1382);
xor (n1381,n1348,n1375);
and (n1382,n1383,n1385);
xor (n1383,n1384,n1325);
xor (n1384,n1316,n1320);
xor (n1385,n1386,n1370);
xor (n1386,n1350,n1362);
and (n1387,n1388,n1389);
xor (n1388,n1381,n1382);
or (n1389,n1390,n1415);
and (n1390,n1391,n1392);
xor (n1391,n1383,n1385);
or (n1392,n1393,n1412,n1414);
and (n1393,n1394,n1410);
or (n1394,n1395,n1404,n1409);
and (n1395,n1396,n1400);
xnor (n1396,n1397,n408);
nor (n1397,n1398,n1399);
and (n1398,n445,n743);
and (n1399,n361,n745);
xnor (n1400,n1401,n404);
nor (n1401,n1402,n1403);
and (n1402,n578,n556);
and (n1403,n514,n559);
and (n1404,n1400,n1405);
xnor (n1405,n1406,n300);
nor (n1406,n1407,n1408);
and (n1407,n830,n412);
and (n1408,n672,n415);
and (n1409,n1396,n1405);
xor (n1410,n1411,n195);
xor (n1411,n1352,n1356);
and (n1412,n1410,n1413);
xor (n1413,n1363,n1367);
and (n1414,n1394,n1413);
and (n1415,n1416,n1417);
xor (n1416,n1391,n1392);
or (n1417,n1418,n1436);
and (n1418,n1419,n1421);
xor (n1419,n1420,n1413);
xor (n1420,n1394,n1410);
and (n1421,n1422,n1434);
or (n1422,n1423,n1432,n1433);
and (n1423,n1424,n1428);
xnor (n1424,n1425,n408);
nor (n1425,n1426,n1427);
and (n1426,n514,n743);
and (n1427,n445,n745);
xnor (n1428,n1429,n404);
nor (n1429,n1430,n1431);
and (n1430,n672,n556);
and (n1431,n578,n559);
and (n1432,n1428,n300);
and (n1433,n1424,n300);
xor (n1434,n1435,n1405);
xor (n1435,n1396,n1400);
and (n1436,n1437,n1438);
xor (n1437,n1419,n1421);
or (n1438,n1439,n1446);
and (n1439,n1440,n1441);
xor (n1440,n1422,n1434);
and (n1441,n1442,n1444);
xnor (n1442,n1443,n300);
nand (n1443,n830,n415);
xor (n1444,n1445,n300);
xor (n1445,n1424,n1428);
and (n1446,n1447,n1448);
xor (n1447,n1440,n1441);
or (n1448,n1449,n1460);
and (n1449,n1450,n1451);
xor (n1450,n1442,n1444);
and (n1451,n1452,n1456);
xnor (n1452,n1453,n408);
nor (n1453,n1454,n1455);
and (n1454,n578,n743);
and (n1455,n514,n745);
xnor (n1456,n1457,n404);
nor (n1457,n1458,n1459);
and (n1458,n830,n556);
and (n1459,n672,n559);
and (n1460,n1461,n1462);
xor (n1461,n1450,n1451);
or (n1462,n1463,n1470);
and (n1463,n1464,n1465);
xor (n1464,n1452,n1456);
and (n1465,n1466,n404);
xnor (n1466,n1467,n408);
nor (n1467,n1468,n1469);
and (n1468,n672,n743);
and (n1469,n578,n745);
and (n1470,n1471,n1472);
xor (n1471,n1464,n1465);
or (n1472,n1473,n1477);
and (n1473,n1474,n1476);
xnor (n1474,n1475,n404);
nand (n1475,n830,n559);
xor (n1476,n1466,n404);
and (n1477,n1478,n1479);
xor (n1478,n1474,n1476);
and (n1479,n1480,n1484);
xnor (n1480,n1481,n408);
nor (n1481,n1482,n1483);
and (n1482,n830,n743);
and (n1483,n672,n745);
and (n1484,n1485,n408);
xnor (n1485,n1486,n408);
nand (n1486,n830,n745);
xor (n1487,n1488,n1508);
xor (n1488,n1489,n1494);
xor (n1489,n1490,n1493);
or (n1490,n1491,n27,n1492);
and (n1491,n57,n12);
and (n1492,n57,n28);
xnor (n1493,n58,n61);
or (n1494,n1495,n1505,n1507);
and (n1495,n1496,n1499);
or (n1496,n47,n1497,n1498);
and (n1497,n48,n82);
and (n1498,n40,n82);
or (n1499,n1500,n1503);
or (n1500,n1501,n72,n1502);
and (n1501,n34,n68);
and (n1502,n34,n73);
xor (n1503,n1504,n82);
xor (n1504,n40,n48);
and (n1505,n1499,n1506);
not (n1506,n53);
and (n1507,n1496,n1506);
or (n1508,n1509,n1541);
and (n1509,n1510,n1512);
xor (n1510,n1511,n1506);
xor (n1511,n1496,n1499);
or (n1512,n1513,n1538,n1540);
and (n1513,n1514,n1521);
or (n1514,n1515,n1519,n1520);
and (n1515,n1516,n159);
or (n1516,n103,n1517,n1518);
and (n1517,n104,n153);
and (n1518,n96,n153);
and (n1519,n159,n79);
and (n1520,n1516,n79);
or (n1521,n1522,n1534,n1537);
and (n1522,n1523,n1533);
or (n1523,n1524,n1530,n1532);
and (n1524,n1525,n1528);
or (n1525,n1526,n138,n1527);
and (n1526,n90,n134);
and (n1527,n90,n139);
xor (n1528,n1529,n153);
xor (n1529,n96,n104);
and (n1530,n1528,n1531);
not (n1531,n159);
and (n1532,n1525,n1531);
not (n1533,n109);
and (n1534,n1533,n1535);
xor (n1535,n1536,n79);
xor (n1536,n1516,n159);
and (n1537,n1523,n1535);
and (n1538,n1521,n1539);
xnor (n1539,n1500,n1503);
and (n1540,n1514,n1539);
and (n1541,n1542,n1543);
xor (n1542,n1510,n1512);
or (n1543,n1544,n1566);
and (n1544,n1545,n1547);
xor (n1545,n1546,n1539);
xor (n1546,n1514,n1521);
and (n1547,n1548,n1564);
or (n1548,n1549,n1560,n1563);
and (n1549,n1550,n1558);
or (n1550,n1551,n1556,n1557);
and (n1551,n1552,n1555);
or (n1552,n207,n1553,n1554);
and (n1553,n208,n180);
and (n1554,n200,n180);
or (n1555,n184,n189);
and (n1556,n1555,n145);
and (n1557,n1552,n145);
and (n1558,n150,n1559);
not (n1559,n263);
and (n1560,n1558,n1561);
xor (n1561,n1562,n1531);
xor (n1562,n1525,n1528);
and (n1563,n1550,n1561);
xor (n1564,n1565,n1535);
xor (n1565,n1523,n1533);
and (n1566,n1567,n1568);
xor (n1567,n1545,n1547);
or (n1568,n1569,n1589);
and (n1569,n1570,n1571);
xor (n1570,n1548,n1564);
and (n1571,n1572,n1587);
or (n1572,n1573,n1584,n1586);
and (n1573,n1574,n1582);
or (n1574,n1575,n1579,n1581);
and (n1575,n233,n1576);
or (n1576,n1577,n253,n1578);
and (n1577,n194,n249);
and (n1578,n194,n254);
and (n1579,n1576,n1580);
xnor (n1580,n184,n189);
and (n1581,n233,n1580);
xor (n1582,n1583,n145);
xor (n1583,n1552,n1555);
and (n1584,n1582,n1585);
xor (n1585,n150,n1559);
and (n1586,n1574,n1585);
xor (n1587,n1588,n1561);
xor (n1588,n1550,n1558);
and (n1589,n1590,n1591);
xor (n1590,n1570,n1571);
or (n1591,n1592,n1615);
and (n1592,n1593,n1594);
xor (n1593,n1572,n1587);
and (n1594,n1595,n1613);
or (n1595,n1596,n1609,n1612);
and (n1596,n1597,n1607);
or (n1597,n1598,n1605,n1606);
and (n1598,n1599,n1602);
or (n1599,n291,n1600,n1601);
and (n1600,n292,n365);
and (n1601,n287,n365);
or (n1602,n312,n1603,n1604);
and (n1603,n313,n283);
and (n1604,n305,n283);
and (n1605,n1602,n373);
and (n1606,n1599,n373);
xor (n1607,n1608,n180);
xor (n1608,n200,n208);
and (n1609,n1607,n1610);
xor (n1610,n1611,n1580);
xor (n1611,n233,n1576);
and (n1612,n1597,n1610);
xor (n1613,n1614,n1585);
xor (n1614,n1574,n1582);
and (n1615,n1616,n1617);
xor (n1616,n1593,n1594);
or (n1617,n1618,n1667);
and (n1618,n1619,n1620);
xor (n1619,n1595,n1613);
or (n1620,n1621,n1663,n1666);
and (n1621,n1622,n1633);
or (n1622,n1623,n1629,n1632);
and (n1623,n1624,n1628);
or (n1624,n1625,n342);
or (n1625,n1626,n336,n1627);
and (n1626,n299,n332);
and (n1627,n299,n337);
not (n1628,n377);
and (n1629,n1628,n1630);
xor (n1630,n1631,n373);
xor (n1631,n1599,n1602);
and (n1632,n1624,n1630);
or (n1633,n1634,n1659,n1662);
and (n1634,n1635,n1655);
or (n1635,n1636,n1651,n1654);
and (n1636,n1637,n1647);
or (n1637,n1638,n1645,n1646);
and (n1638,n1639,n1642);
or (n1639,n416,n1640,n1641);
and (n1640,n417,n424);
and (n1641,n409,n424);
or (n1642,n432,n1643,n1644);
and (n1643,n433,n440);
and (n1644,n428,n440);
and (n1645,n1642,n444);
and (n1646,n1639,n444);
or (n1647,n1648,n1649,n1650);
and (n1648,n360,n528);
and (n1649,n528,n451);
and (n1650,n360,n451);
and (n1651,n1647,n1652);
xor (n1652,n1653,n365);
xor (n1653,n287,n292);
and (n1654,n1637,n1652);
and (n1655,n1656,n1658);
xor (n1656,n1657,n283);
xor (n1657,n305,n313);
xnor (n1658,n1625,n342);
and (n1659,n1655,n1660);
xor (n1660,n1661,n1630);
xor (n1661,n1624,n1628);
and (n1662,n1635,n1660);
and (n1663,n1633,n1664);
xor (n1664,n1665,n1610);
xor (n1665,n1597,n1607);
and (n1666,n1622,n1664);
and (n1667,n1668,n1669);
xor (n1668,n1619,n1620);
or (n1669,n1670,n1704);
and (n1670,n1671,n1673);
xor (n1671,n1672,n1664);
xor (n1672,n1622,n1633);
and (n1673,n1674,n1702);
or (n1674,n1675,n1699,n1701);
and (n1675,n1676,n1697);
or (n1676,n1677,n1695,n1696);
and (n1677,n1678,n1686);
or (n1678,n1679,n1683,n1685);
and (n1679,n1680,n491);
or (n1680,n1681,n485,n1682);
and (n1681,n403,n481);
and (n1682,n403,n486);
and (n1683,n491,n1684);
and (n1684,n509,n513);
and (n1685,n1680,n1684);
or (n1686,n1687,n1692,n1694);
and (n1687,n1688,n1690);
xor (n1688,n1689,n424);
xor (n1689,n409,n417);
xor (n1690,n1691,n440);
xor (n1691,n428,n433);
and (n1692,n1690,n1693);
not (n1693,n444);
and (n1694,n1688,n1693);
and (n1695,n1686,n526);
and (n1696,n1678,n526);
xor (n1697,n1698,n1652);
xor (n1698,n1637,n1647);
and (n1699,n1697,n1700);
xor (n1700,n1656,n1658);
and (n1701,n1676,n1700);
xor (n1702,n1703,n1660);
xor (n1703,n1635,n1655);
and (n1704,n1705,n1706);
xor (n1705,n1671,n1673);
or (n1706,n1707,n1741);
and (n1707,n1708,n1709);
xor (n1708,n1674,n1702);
and (n1709,n1710,n1739);
or (n1710,n1711,n1735,n1738);
and (n1711,n1712,n1733);
or (n1712,n1713,n1729,n1732);
and (n1713,n1714,n1725);
or (n1714,n1715,n1722,n1724);
and (n1715,n1716,n1719);
or (n1716,n560,n1717,n1718);
and (n1717,n561,n583);
and (n1718,n553,n583);
or (n1719,n591,n1720,n1721);
and (n1720,n592,n568);
and (n1721,n587,n568);
and (n1722,n1719,n1723);
or (n1723,n572,n577);
and (n1724,n1716,n1723);
or (n1725,n1726,n1727,n1728);
and (n1726,n683,n602);
and (n1727,n602,n684);
and (n1728,n683,n684);
and (n1729,n1725,n1730);
xor (n1730,n1731,n1693);
xor (n1731,n1688,n1690);
and (n1732,n1714,n1730);
xor (n1733,n1734,n444);
xor (n1734,n1639,n1642);
and (n1735,n1733,n1736);
xor (n1736,n1737,n526);
xor (n1737,n1678,n1686);
and (n1738,n1712,n1736);
xor (n1739,n1740,n1700);
xor (n1740,n1676,n1697);
and (n1741,n1742,n1743);
xor (n1742,n1708,n1709);
or (n1743,n1744,n1776);
and (n1744,n1745,n1746);
xor (n1745,n1710,n1739);
and (n1746,n1747,n1774);
or (n1747,n1748,n1770,n1773);
and (n1748,n1749,n1768);
or (n1749,n1750,n1766,n1767);
and (n1750,n1751,n1757);
or (n1751,n1752,n1756,n674);
and (n1752,n631,n1753);
or (n1753,n1754,n653,n1755);
and (n1754,n552,n649);
and (n1755,n552,n654);
and (n1756,n1753,n660);
or (n1757,n1758,n1763,n1765);
and (n1758,n1759,n1761);
xor (n1759,n1760,n583);
xor (n1760,n553,n561);
xor (n1761,n1762,n568);
xor (n1762,n587,n592);
and (n1763,n1761,n1764);
xnor (n1764,n572,n577);
and (n1765,n1759,n1764);
and (n1766,n1757,n681);
and (n1767,n1751,n681);
xor (n1768,n1769,n1684);
xor (n1769,n1680,n491);
and (n1770,n1768,n1771);
xor (n1771,n1772,n1730);
xor (n1772,n1714,n1725);
and (n1773,n1749,n1771);
xor (n1774,n1775,n1736);
xor (n1775,n1712,n1733);
and (n1776,n1777,n1778);
xor (n1777,n1745,n1746);
or (n1778,n1779,n1799);
and (n1779,n1780,n1781);
xor (n1780,n1747,n1774);
and (n1781,n1782,n1797);
or (n1782,n1783,n1793,n1796);
and (n1783,n1784,n1791);
or (n1784,n1785,n1787,n1790);
and (n1785,n704,n1786);
or (n1786,n754,n759);
and (n1787,n1786,n1788);
xor (n1788,n1789,n1764);
xor (n1789,n1759,n1761);
and (n1790,n704,n1788);
xor (n1791,n1792,n1723);
xor (n1792,n1716,n1719);
and (n1793,n1791,n1794);
xor (n1794,n1795,n681);
xor (n1795,n1751,n1757);
and (n1796,n1784,n1794);
xor (n1797,n1798,n1771);
xor (n1798,n1749,n1768);
and (n1799,n1800,n1801);
xor (n1800,n1780,n1781);
or (n1801,n1802,n1818);
and (n1802,n1803,n1804);
xor (n1803,n1782,n1797);
and (n1804,n1805,n1816);
or (n1805,n1806,n1812,n1815);
and (n1806,n1807,n1810);
or (n1807,n786,n1808,n1809);
and (n1808,n833,n955);
and (n1809,n787,n955);
xor (n1810,n1811,n660);
xor (n1811,n631,n1753);
and (n1812,n1810,n1813);
xor (n1813,n1814,n1788);
xor (n1814,n704,n1786);
and (n1815,n1807,n1813);
xor (n1816,n1817,n1794);
xor (n1817,n1784,n1791);
and (n1818,n1819,n1820);
xor (n1819,n1803,n1804);
or (n1820,n1821,n1829);
and (n1821,n1822,n1823);
xor (n1822,n1805,n1816);
and (n1823,n1824,n1827);
or (n1824,n866,n1825,n1826);
and (n1825,n927,n957);
and (n1826,n867,n957);
xor (n1827,n1828,n1813);
xor (n1828,n1807,n1810);
and (n1829,n1830,n1831);
xor (n1830,n1822,n1823);
or (n1831,n1832,n948);
and (n1832,n1833,n1834);
xor (n1833,n1824,n1827);
or (n1834,n1835,n1836,n1837);
and (n1835,n933,n954);
and (n1836,n954,n956);
and (n1837,n933,n956);
endmodule
