module top (out,n7,n10,n11,n15,n18,n19,n27,n41,n50
        ,n51,n89,n93,n107,n108,n163,n166,n205,n213,n214
        ,n260,n318,n319,n371,n376,n422,n423,n460,n529,n593
        ,n687,n760,n845);
output out;
input n7;
input n10;
input n11;
input n15;
input n18;
input n19;
input n27;
input n41;
input n50;
input n51;
input n89;
input n93;
input n107;
input n108;
input n163;
input n166;
input n205;
input n213;
input n214;
input n260;
input n318;
input n319;
input n371;
input n376;
input n422;
input n423;
input n460;
input n529;
input n593;
input n687;
input n760;
input n845;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n8;
wire n9;
wire n12;
wire n13;
wire n14;
wire n16;
wire n17;
wire n20;
wire n21;
wire n22;
wire n23;
wire n24;
wire n25;
wire n26;
wire n28;
wire n29;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n90;
wire n91;
wire n92;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n164;
wire n165;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n372;
wire n373;
wire n374;
wire n375;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
xor (out,n0,n1502);
xor (n0,n1,n71);
xor (n1,n2,n31);
xor (n2,n3,n29);
or (n3,n4,n25,n28);
and (n4,n5,n12);
not (n5,n6);
and (n6,n7,n8);
not (n8,n9);
and (n9,n10,n11);
xnor (n12,n13,n22);
not (n13,n14);
and (n14,n15,n16);
and (n16,n17,n20);
xor (n17,n18,n19);
not (n20,n21);
xor (n21,n19,n7);
and (n22,n18,n23);
not (n23,n24);
and (n24,n19,n7);
and (n25,n12,n26);
and (n26,n27,n18);
and (n28,n5,n26);
xnor (n29,n22,n30);
and (n30,n15,n18);
or (n31,n32,n67,n70);
and (n32,n33,n43);
or (n33,n34,n39,n42);
and (n34,n6,n35);
xnor (n35,n36,n22);
nor (n36,n37,n38);
and (n37,n27,n16);
and (n38,n15,n21);
and (n39,n35,n40);
and (n40,n41,n18);
and (n42,n6,n40);
or (n43,n44,n65);
or (n44,n45,n59,n64);
and (n45,n46,n52);
not (n46,n47);
and (n47,n11,n48);
not (n48,n49);
and (n49,n50,n51);
xnor (n52,n53,n6);
not (n53,n54);
and (n54,n15,n55);
and (n55,n56,n57);
xor (n56,n7,n10);
not (n57,n58);
xor (n58,n10,n11);
and (n59,n52,n60);
xnor (n60,n61,n22);
nor (n61,n62,n63);
and (n62,n41,n16);
and (n63,n27,n21);
and (n64,n46,n60);
xor (n65,n66,n40);
xor (n66,n6,n35);
and (n67,n43,n68);
xor (n68,n69,n26);
xor (n69,n5,n12);
and (n70,n33,n68);
or (n71,n72,n136);
and (n72,n73,n75);
xor (n73,n74,n68);
xor (n74,n33,n43);
or (n75,n76,n133,n135);
and (n76,n77,n97);
or (n77,n78,n94,n96);
and (n78,n79,n92);
or (n79,n80,n85,n91);
and (n80,n47,n81);
xnor (n81,n82,n6);
nor (n82,n83,n84);
and (n83,n27,n55);
and (n84,n15,n58);
and (n85,n81,n86);
xnor (n86,n87,n22);
nor (n87,n88,n90);
and (n88,n89,n16);
and (n90,n41,n21);
and (n91,n47,n86);
and (n92,n93,n18);
and (n94,n92,n95);
and (n95,n89,n18);
and (n96,n79,n95);
or (n97,n98,n129,n132);
and (n98,n99,n127);
or (n99,n100,n124,n126);
and (n100,n101,n122);
or (n101,n102,n116,n121);
and (n102,n103,n109);
not (n103,n104);
and (n104,n51,n105);
not (n105,n106);
and (n106,n107,n108);
xnor (n109,n110,n47);
not (n110,n111);
and (n111,n15,n112);
and (n112,n113,n114);
xor (n113,n11,n50);
not (n114,n115);
xor (n115,n50,n51);
and (n116,n109,n117);
xnor (n117,n118,n6);
nor (n118,n119,n120);
and (n119,n41,n55);
and (n120,n27,n58);
and (n121,n103,n117);
xor (n122,n123,n86);
xor (n123,n47,n81);
and (n124,n122,n125);
not (n125,n92);
and (n126,n101,n125);
xor (n127,n128,n60);
xor (n128,n46,n52);
and (n129,n127,n130);
xor (n130,n131,n95);
xor (n131,n79,n92);
and (n132,n99,n130);
and (n133,n97,n134);
xnor (n134,n44,n65);
and (n135,n77,n134);
and (n136,n137,n138);
xor (n137,n73,n75);
or (n138,n139,n183);
and (n139,n140,n142);
xor (n140,n141,n134);
xor (n141,n77,n97);
and (n142,n143,n181);
or (n143,n144,n177,n180);
and (n144,n145,n173);
or (n145,n146,n167,n172);
and (n146,n147,n159);
or (n147,n148,n153,n158);
and (n148,n104,n149);
xnor (n149,n150,n47);
nor (n150,n151,n152);
and (n151,n27,n112);
and (n152,n15,n115);
and (n153,n149,n154);
xnor (n154,n155,n6);
nor (n155,n156,n157);
and (n156,n89,n55);
and (n157,n41,n58);
and (n158,n104,n154);
or (n159,n160,n165);
xnor (n160,n161,n22);
nor (n161,n162,n164);
and (n162,n163,n16);
and (n164,n93,n21);
and (n165,n166,n18);
and (n167,n159,n168);
xnor (n168,n169,n22);
nor (n169,n170,n171);
and (n170,n93,n16);
and (n171,n89,n21);
and (n172,n147,n168);
and (n173,n174,n175);
and (n174,n163,n18);
xor (n175,n176,n117);
xor (n176,n103,n109);
and (n177,n173,n178);
xor (n178,n179,n125);
xor (n179,n101,n122);
and (n180,n145,n178);
xor (n181,n182,n130);
xor (n182,n99,n127);
and (n183,n184,n185);
xor (n184,n140,n142);
or (n185,n186,n238);
and (n186,n187,n188);
xor (n187,n143,n181);
and (n188,n189,n236);
or (n189,n190,n233,n235);
and (n190,n191,n231);
or (n191,n192,n228,n230);
and (n192,n193,n207);
or (n193,n194,n203,n206);
and (n194,n195,n199);
xnor (n195,n196,n6);
nor (n196,n197,n198);
and (n197,n93,n55);
and (n198,n89,n58);
xnor (n199,n200,n22);
nor (n200,n201,n202);
and (n201,n166,n16);
and (n202,n163,n21);
and (n203,n199,n204);
and (n204,n205,n18);
and (n206,n195,n204);
or (n207,n208,n222,n227);
and (n208,n209,n215);
not (n209,n210);
and (n210,n108,n211);
not (n211,n212);
and (n212,n213,n214);
xnor (n215,n216,n104);
not (n216,n217);
and (n217,n15,n218);
and (n218,n219,n220);
xor (n219,n51,n107);
not (n220,n221);
xor (n221,n107,n108);
and (n222,n215,n223);
xnor (n223,n224,n47);
nor (n224,n225,n226);
and (n225,n41,n112);
and (n226,n27,n115);
and (n227,n209,n223);
and (n228,n207,n229);
xnor (n229,n160,n165);
and (n230,n193,n229);
xor (n231,n232,n168);
xor (n232,n147,n159);
and (n233,n231,n234);
xor (n234,n174,n175);
and (n235,n191,n234);
xor (n236,n237,n178);
xor (n237,n145,n173);
and (n238,n239,n240);
xor (n239,n187,n188);
or (n240,n241,n286);
and (n241,n242,n243);
xor (n242,n189,n236);
and (n243,n244,n284);
or (n244,n245,n280,n283);
and (n245,n246,n278);
or (n246,n247,n274,n277);
and (n247,n248,n262);
or (n248,n249,n258,n261);
and (n249,n250,n254);
xnor (n250,n251,n6);
nor (n251,n252,n253);
and (n252,n163,n55);
and (n253,n93,n58);
xnor (n254,n255,n22);
nor (n255,n256,n257);
and (n256,n205,n16);
and (n257,n166,n21);
and (n258,n254,n259);
and (n259,n260,n18);
and (n261,n250,n259);
or (n262,n263,n268,n273);
and (n263,n210,n264);
xnor (n264,n265,n104);
nor (n265,n266,n267);
and (n266,n27,n218);
and (n267,n15,n221);
and (n268,n264,n269);
xnor (n269,n270,n47);
nor (n270,n271,n272);
and (n271,n89,n112);
and (n272,n41,n115);
and (n273,n210,n269);
and (n274,n262,n275);
xor (n275,n276,n204);
xor (n276,n195,n199);
and (n277,n248,n275);
xor (n278,n279,n154);
xor (n279,n104,n149);
and (n280,n278,n281);
xor (n281,n282,n229);
xor (n282,n193,n207);
and (n283,n246,n281);
xor (n284,n285,n234);
xor (n285,n191,n231);
and (n286,n287,n288);
xor (n287,n242,n243);
or (n288,n289,n403);
and (n289,n290,n291);
xor (n290,n244,n284);
or (n291,n292,n399,n402);
and (n292,n293,n339);
or (n293,n294,n335,n338);
and (n294,n295,n333);
or (n295,n296,n312);
or (n296,n297,n306,n311);
and (n297,n298,n302);
xnor (n298,n299,n47);
nor (n299,n300,n301);
and (n300,n93,n112);
and (n301,n89,n115);
xnor (n302,n303,n6);
nor (n303,n304,n305);
and (n304,n166,n55);
and (n305,n163,n58);
and (n306,n302,n307);
xnor (n307,n308,n22);
nor (n308,n309,n310);
and (n309,n260,n16);
and (n310,n205,n21);
and (n311,n298,n307);
or (n312,n313,n327,n332);
and (n313,n314,n320);
not (n314,n315);
and (n315,n214,n316);
not (n316,n317);
and (n317,n318,n319);
xnor (n320,n321,n210);
not (n321,n322);
and (n322,n15,n323);
and (n323,n324,n325);
xor (n324,n108,n213);
not (n325,n326);
xor (n326,n213,n214);
and (n327,n320,n328);
xnor (n328,n329,n104);
nor (n329,n330,n331);
and (n330,n41,n218);
and (n331,n27,n221);
and (n332,n314,n328);
xor (n333,n334,n223);
xor (n334,n209,n215);
and (n335,n333,n336);
xor (n336,n337,n275);
xor (n337,n248,n262);
and (n338,n295,n336);
or (n339,n340,n395,n398);
and (n340,n341,n391);
or (n341,n342,n387,n390);
and (n342,n343,n378);
or (n343,n344,n374,n377);
and (n344,n345,n357);
or (n345,n346,n351,n356);
and (n346,n315,n347);
xnor (n347,n348,n210);
nor (n348,n349,n350);
and (n349,n27,n323);
and (n350,n15,n326);
and (n351,n347,n352);
xnor (n352,n353,n104);
nor (n353,n354,n355);
and (n354,n89,n218);
and (n355,n41,n221);
and (n356,n315,n352);
or (n357,n358,n367,n373);
and (n358,n359,n363);
xnor (n359,n360,n47);
nor (n360,n361,n362);
and (n361,n163,n112);
and (n362,n93,n115);
xnor (n363,n364,n6);
nor (n364,n365,n366);
and (n365,n205,n55);
and (n366,n166,n58);
and (n367,n363,n368);
xnor (n368,n369,n22);
nor (n369,n370,n372);
and (n370,n371,n16);
and (n372,n260,n21);
and (n373,n359,n368);
and (n374,n357,n375);
and (n375,n376,n18);
and (n377,n345,n375);
or (n378,n379,n383,n386);
and (n379,n380,n381);
and (n380,n371,n18);
xor (n381,n382,n307);
xor (n382,n298,n302);
and (n383,n381,n384);
xor (n384,n385,n328);
xor (n385,n314,n320);
and (n386,n380,n384);
and (n387,n378,n388);
xor (n388,n389,n259);
xor (n389,n250,n254);
and (n390,n343,n388);
and (n391,n392,n394);
xor (n392,n393,n269);
xor (n393,n210,n264);
xnor (n394,n296,n312);
and (n395,n391,n396);
xor (n396,n397,n336);
xor (n397,n295,n333);
and (n398,n341,n396);
and (n399,n339,n400);
xor (n400,n401,n281);
xor (n401,n246,n278);
and (n402,n293,n400);
and (n403,n404,n405);
xor (n404,n290,n291);
or (n405,n406,n482);
and (n406,n407,n409);
xor (n407,n408,n400);
xor (n408,n293,n339);
and (n409,n410,n480);
or (n410,n411,n477,n479);
and (n411,n412,n475);
or (n412,n413,n471,n474);
and (n413,n414,n462);
or (n414,n415,n453,n461);
and (n415,n416,n437);
or (n416,n417,n431,n436);
and (n417,n418,n424);
not (n418,n419);
and (n419,n319,n420);
not (n420,n421);
and (n421,n422,n423);
xnor (n424,n425,n315);
not (n425,n426);
and (n426,n15,n427);
and (n427,n428,n429);
xor (n428,n214,n318);
not (n429,n430);
xor (n430,n318,n319);
and (n431,n424,n432);
xnor (n432,n433,n210);
nor (n433,n434,n435);
and (n434,n41,n323);
and (n435,n27,n326);
and (n436,n418,n432);
or (n437,n438,n447,n452);
and (n438,n439,n443);
xnor (n439,n440,n104);
nor (n440,n441,n442);
and (n441,n93,n218);
and (n442,n89,n221);
xnor (n443,n444,n47);
nor (n444,n445,n446);
and (n445,n166,n112);
and (n446,n163,n115);
and (n447,n443,n448);
xnor (n448,n449,n6);
nor (n449,n450,n451);
and (n450,n260,n55);
and (n451,n205,n58);
and (n452,n439,n448);
and (n453,n437,n454);
and (n454,n455,n459);
xnor (n455,n456,n22);
nor (n456,n457,n458);
and (n457,n376,n16);
and (n458,n371,n21);
and (n459,n460,n18);
and (n461,n416,n454);
or (n462,n463,n468,n470);
and (n463,n464,n466);
xor (n464,n465,n352);
xor (n465,n315,n347);
xor (n466,n467,n368);
xor (n467,n359,n363);
and (n468,n466,n469);
not (n469,n375);
and (n470,n464,n469);
and (n471,n462,n472);
xor (n472,n473,n384);
xor (n473,n380,n381);
and (n474,n414,n472);
xor (n475,n476,n388);
xor (n476,n343,n378);
and (n477,n475,n478);
xor (n478,n392,n394);
and (n479,n412,n478);
xor (n480,n481,n396);
xor (n481,n341,n391);
and (n482,n483,n484);
xor (n483,n407,n409);
or (n484,n485,n553);
and (n485,n486,n487);
xor (n486,n410,n480);
and (n487,n488,n551);
or (n488,n489,n547,n550);
and (n489,n490,n545);
or (n490,n491,n540,n544);
and (n491,n492,n531);
or (n492,n493,n522,n530);
and (n493,n494,n506);
or (n494,n495,n500,n505);
and (n495,n419,n496);
xnor (n496,n497,n315);
nor (n497,n498,n499);
and (n498,n27,n427);
and (n499,n15,n430);
and (n500,n496,n501);
xnor (n501,n502,n210);
nor (n502,n503,n504);
and (n503,n89,n323);
and (n504,n41,n326);
and (n505,n419,n501);
or (n506,n507,n516,n521);
and (n507,n508,n512);
xnor (n508,n509,n104);
nor (n509,n510,n511);
and (n510,n163,n218);
and (n511,n93,n221);
xnor (n512,n513,n47);
nor (n513,n514,n515);
and (n514,n205,n112);
and (n515,n166,n115);
and (n516,n512,n517);
xnor (n517,n518,n6);
nor (n518,n519,n520);
and (n519,n371,n55);
and (n520,n260,n58);
and (n521,n508,n517);
and (n522,n506,n523);
or (n523,n524,n528);
xnor (n524,n525,n22);
nor (n525,n526,n527);
and (n526,n460,n16);
and (n527,n376,n21);
and (n528,n529,n18);
and (n530,n494,n523);
or (n531,n532,n537,n539);
and (n532,n533,n535);
xor (n533,n534,n432);
xor (n534,n418,n424);
xor (n535,n536,n448);
xor (n536,n439,n443);
and (n537,n535,n538);
xor (n538,n455,n459);
and (n539,n533,n538);
and (n540,n531,n541);
xor (n541,n542,n466);
xor (n542,n375,n543);
not (n543,n464);
and (n544,n492,n541);
xor (n545,n546,n375);
xor (n546,n345,n357);
and (n547,n545,n548);
xor (n548,n549,n472);
xor (n549,n414,n462);
and (n550,n490,n548);
xor (n551,n552,n478);
xor (n552,n412,n475);
and (n553,n554,n555);
xor (n554,n486,n487);
or (n555,n556,n634);
and (n556,n557,n558);
xor (n557,n488,n551);
and (n558,n559,n632);
or (n559,n560,n628,n631);
and (n560,n561,n626);
or (n561,n562,n622,n625);
and (n562,n563,n613);
or (n563,n564,n595,n612);
and (n564,n565,n581);
or (n565,n566,n575,n580);
and (n566,n567,n568);
not (n567,n423);
xnor (n568,n569,n419);
not (n569,n570);
and (n570,n15,n571);
and (n571,n572,n573);
xor (n572,n319,n422);
not (n573,n574);
xor (n574,n422,n423);
and (n575,n568,n576);
xnor (n576,n577,n315);
nor (n577,n578,n579);
and (n578,n41,n427);
and (n579,n27,n430);
and (n580,n567,n576);
or (n581,n582,n591,n594);
and (n582,n583,n587);
xnor (n583,n584,n6);
nor (n584,n585,n586);
and (n585,n376,n55);
and (n586,n371,n58);
xnor (n587,n588,n22);
nor (n588,n589,n590);
and (n589,n529,n16);
and (n590,n460,n21);
and (n591,n587,n592);
and (n592,n593,n18);
and (n594,n583,n592);
and (n595,n581,n596);
or (n596,n597,n606,n611);
and (n597,n598,n602);
xnor (n598,n599,n210);
nor (n599,n600,n601);
and (n600,n93,n323);
and (n601,n89,n326);
xnor (n602,n603,n104);
nor (n603,n604,n605);
and (n604,n166,n218);
and (n605,n163,n221);
and (n606,n602,n607);
xnor (n607,n608,n47);
nor (n608,n609,n610);
and (n609,n260,n112);
and (n610,n205,n115);
and (n611,n598,n607);
and (n612,n565,n596);
or (n613,n614,n619,n621);
and (n614,n615,n617);
xor (n615,n616,n501);
xor (n616,n419,n496);
xor (n617,n618,n517);
xor (n618,n508,n512);
and (n619,n617,n620);
xnor (n620,n524,n528);
and (n621,n615,n620);
and (n622,n613,n623);
xor (n623,n624,n538);
xor (n624,n533,n535);
and (n625,n563,n623);
xor (n626,n627,n454);
xor (n627,n416,n437);
and (n628,n626,n629);
xor (n629,n630,n541);
xor (n630,n492,n531);
and (n631,n561,n629);
xor (n632,n633,n548);
xor (n633,n490,n545);
and (n634,n635,n636);
xor (n635,n557,n558);
or (n636,n637,n709);
and (n637,n638,n639);
xor (n638,n559,n632);
and (n639,n640,n707);
or (n640,n641,n703,n706);
and (n641,n642,n701);
or (n642,n643,n695,n700);
and (n643,n644,n690);
or (n644,n645,n674,n689);
and (n645,n646,n662);
or (n646,n647,n656,n661);
and (n647,n648,n652);
xnor (n648,n649,n210);
nor (n649,n650,n651);
and (n650,n163,n323);
and (n651,n93,n326);
xnor (n652,n653,n104);
nor (n653,n654,n655);
and (n654,n205,n218);
and (n655,n166,n221);
and (n656,n652,n657);
xnor (n657,n658,n47);
nor (n658,n659,n660);
and (n659,n371,n112);
and (n660,n260,n115);
and (n661,n648,n657);
or (n662,n663,n668,n673);
and (n663,n423,n664);
xnor (n664,n665,n419);
nor (n665,n666,n667);
and (n666,n27,n571);
and (n667,n15,n574);
and (n668,n664,n669);
xnor (n669,n670,n315);
nor (n670,n671,n672);
and (n671,n89,n427);
and (n672,n41,n430);
and (n673,n423,n669);
and (n674,n662,n675);
or (n675,n676,n685,n688);
and (n676,n677,n681);
xnor (n677,n678,n6);
nor (n678,n679,n680);
and (n679,n460,n55);
and (n680,n376,n58);
xnor (n681,n682,n22);
nor (n682,n683,n684);
and (n683,n593,n16);
and (n684,n529,n21);
and (n685,n681,n686);
and (n686,n687,n18);
and (n688,n677,n686);
and (n689,n646,n675);
or (n690,n691,n693);
xor (n691,n692,n592);
xor (n692,n583,n587);
xor (n693,n694,n607);
xor (n694,n598,n602);
and (n695,n690,n696);
xor (n696,n697,n699);
xor (n697,n698,n617);
not (n698,n615);
not (n699,n620);
and (n700,n644,n696);
xor (n701,n702,n523);
xor (n702,n494,n506);
and (n703,n701,n704);
xor (n704,n705,n623);
xor (n705,n563,n613);
and (n706,n642,n704);
xor (n707,n708,n629);
xor (n708,n561,n626);
and (n709,n710,n711);
xor (n710,n638,n639);
or (n711,n712,n791);
and (n712,n713,n714);
xor (n713,n640,n707);
and (n714,n715,n789);
or (n715,n716,n785,n788);
and (n716,n717,n781);
or (n717,n718,n777,n780);
and (n718,n719,n767);
or (n719,n720,n753,n766);
and (n720,n721,n737);
or (n721,n722,n731,n736);
and (n722,n723,n727);
xnor (n723,n724,n315);
nor (n724,n725,n726);
and (n725,n93,n427);
and (n726,n89,n430);
xnor (n727,n728,n210);
nor (n728,n729,n730);
and (n729,n166,n323);
and (n730,n163,n326);
and (n731,n727,n732);
xnor (n732,n733,n104);
nor (n733,n734,n735);
and (n734,n260,n218);
and (n735,n205,n221);
and (n736,n723,n732);
or (n737,n738,n747,n752);
and (n738,n739,n743);
xnor (n739,n740,n47);
nor (n740,n741,n742);
and (n741,n376,n112);
and (n742,n371,n115);
xnor (n743,n744,n6);
nor (n744,n745,n746);
and (n745,n529,n55);
and (n746,n460,n58);
and (n747,n743,n748);
xnor (n748,n749,n22);
nor (n749,n750,n751);
and (n750,n687,n16);
and (n751,n593,n21);
and (n752,n739,n748);
and (n753,n737,n754);
and (n754,n755,n762);
xnor (n755,n756,n423);
not (n756,n757);
and (n757,n15,n758);
and (n758,n759,n761);
xor (n759,n423,n760);
not (n761,n760);
xnor (n762,n763,n419);
nor (n763,n764,n765);
and (n764,n41,n571);
and (n765,n27,n574);
and (n766,n721,n754);
or (n767,n768,n773,n776);
and (n768,n769,n771);
xor (n769,n770,n657);
xor (n770,n648,n652);
xor (n771,n772,n669);
xor (n772,n423,n664);
and (n773,n771,n774);
xor (n774,n775,n686);
xor (n775,n677,n681);
and (n776,n769,n774);
and (n777,n767,n778);
xor (n778,n779,n576);
xor (n779,n567,n568);
and (n780,n719,n778);
and (n781,n782,n784);
xor (n782,n783,n675);
xor (n783,n646,n662);
xnor (n784,n691,n693);
and (n785,n781,n786);
xor (n786,n787,n596);
xor (n787,n565,n581);
and (n788,n717,n786);
xor (n789,n790,n704);
xor (n790,n642,n701);
and (n791,n792,n793);
xor (n792,n713,n714);
or (n793,n794,n873);
and (n794,n795,n796);
xor (n795,n715,n789);
or (n796,n797,n869,n872);
and (n797,n798,n867);
or (n798,n799,n864,n866);
and (n799,n800,n862);
or (n800,n801,n858,n861);
and (n801,n802,n848);
or (n802,n803,n836,n847);
and (n803,n804,n820);
or (n804,n805,n814,n819);
and (n805,n806,n810);
xnor (n806,n807,n423);
nor (n807,n808,n809);
and (n808,n27,n758);
and (n809,n15,n760);
xnor (n810,n811,n419);
nor (n811,n812,n813);
and (n812,n89,n571);
and (n813,n41,n574);
and (n814,n810,n815);
xnor (n815,n816,n315);
nor (n816,n817,n818);
and (n817,n163,n427);
and (n818,n93,n430);
and (n819,n806,n815);
or (n820,n821,n830,n835);
and (n821,n822,n826);
xnor (n822,n823,n210);
nor (n823,n824,n825);
and (n824,n205,n323);
and (n825,n166,n326);
xnor (n826,n827,n104);
nor (n827,n828,n829);
and (n828,n371,n218);
and (n829,n260,n221);
and (n830,n826,n831);
xnor (n831,n832,n47);
nor (n832,n833,n834);
and (n833,n460,n112);
and (n834,n376,n115);
and (n835,n822,n831);
and (n836,n820,n837);
and (n837,n838,n842);
xnor (n838,n839,n6);
nor (n839,n840,n841);
and (n840,n593,n55);
and (n841,n529,n58);
xnor (n842,n843,n22);
nor (n843,n844,n846);
and (n844,n845,n16);
and (n846,n687,n21);
and (n847,n804,n837);
or (n848,n849,n854,n857);
and (n849,n850,n852);
not (n850,n851);
nand (n851,n845,n18);
xor (n852,n853,n732);
xor (n853,n723,n727);
and (n854,n852,n855);
xor (n855,n856,n748);
xor (n856,n739,n743);
and (n857,n850,n855);
and (n858,n848,n859);
xor (n859,n860,n774);
xor (n860,n769,n771);
and (n861,n802,n859);
xor (n862,n863,n778);
xor (n863,n719,n767);
and (n864,n862,n865);
xor (n865,n782,n784);
and (n866,n800,n865);
xor (n867,n868,n786);
xor (n868,n717,n781);
and (n869,n867,n870);
xor (n870,n871,n696);
xor (n871,n644,n690);
and (n872,n798,n870);
and (n873,n874,n875);
xor (n874,n795,n796);
or (n875,n876,n953);
and (n876,n877,n879);
xor (n877,n878,n870);
xor (n878,n798,n867);
and (n879,n880,n951);
or (n880,n881,n947,n950);
and (n881,n882,n942);
or (n882,n883,n939,n941);
and (n883,n884,n930);
or (n884,n885,n912,n929);
and (n885,n886,n900);
or (n886,n887,n896,n899);
and (n887,n888,n892);
xnor (n888,n889,n47);
nor (n889,n890,n891);
and (n890,n529,n112);
and (n891,n460,n115);
xnor (n892,n893,n6);
nor (n893,n894,n895);
and (n894,n687,n55);
and (n895,n593,n58);
and (n896,n892,n897);
xnor (n897,n898,n22);
nand (n898,n845,n21);
and (n899,n888,n897);
or (n900,n901,n910,n911);
and (n901,n902,n906);
xnor (n902,n903,n423);
nor (n903,n904,n905);
and (n904,n41,n758);
and (n905,n27,n760);
xnor (n906,n907,n419);
nor (n907,n908,n909);
and (n908,n93,n571);
and (n909,n89,n574);
and (n910,n906,n22);
and (n911,n902,n22);
and (n912,n900,n913);
or (n913,n914,n923,n928);
and (n914,n915,n919);
xnor (n915,n916,n315);
nor (n916,n917,n918);
and (n917,n166,n427);
and (n918,n163,n430);
xnor (n919,n920,n210);
nor (n920,n921,n922);
and (n921,n260,n323);
and (n922,n205,n326);
and (n923,n919,n924);
xnor (n924,n925,n104);
nor (n925,n926,n927);
and (n926,n376,n218);
and (n927,n371,n221);
and (n928,n915,n924);
and (n929,n886,n913);
or (n930,n931,n936,n938);
and (n931,n932,n934);
xor (n932,n933,n815);
xor (n933,n806,n810);
xor (n934,n935,n831);
xor (n935,n822,n826);
and (n936,n934,n937);
xor (n937,n838,n842);
and (n938,n932,n937);
and (n939,n930,n940);
xor (n940,n755,n762);
and (n941,n884,n940);
and (n942,n943,n945);
xor (n943,n944,n837);
xor (n944,n804,n820);
xor (n945,n946,n855);
xor (n946,n850,n852);
and (n947,n942,n948);
xor (n948,n949,n754);
xor (n949,n721,n737);
and (n950,n882,n948);
xor (n951,n952,n865);
xor (n952,n800,n862);
and (n953,n954,n955);
xor (n954,n877,n879);
or (n955,n956,n963);
and (n956,n957,n958);
xor (n957,n880,n951);
and (n958,n959,n961);
xor (n959,n960,n948);
xor (n960,n882,n942);
xor (n961,n962,n859);
xor (n962,n802,n848);
and (n963,n964,n965);
xor (n964,n957,n958);
or (n965,n966,n1029);
and (n966,n967,n973);
xor (n967,n968,n971);
xor (n968,n948,n969);
xor (n969,n962,n970);
not (n970,n771);
xor (n971,n960,n972);
xnor (n972,n769,n774);
or (n973,n974,n1026,n1028);
and (n974,n975,n1024);
or (n975,n976,n1020,n1023);
and (n976,n977,n1015);
or (n977,n978,n1011,n1014);
and (n978,n979,n995);
or (n979,n980,n989,n994);
and (n980,n981,n985);
xnor (n981,n982,n423);
nor (n982,n983,n984);
and (n983,n89,n758);
and (n984,n41,n760);
xnor (n985,n986,n419);
nor (n986,n987,n988);
and (n987,n163,n571);
and (n988,n93,n574);
and (n989,n985,n990);
xnor (n990,n991,n315);
nor (n991,n992,n993);
and (n992,n205,n427);
and (n993,n166,n430);
and (n994,n981,n990);
or (n995,n996,n1005,n1010);
and (n996,n997,n1001);
xnor (n997,n998,n210);
nor (n998,n999,n1000);
and (n999,n371,n323);
and (n1000,n260,n326);
xnor (n1001,n1002,n104);
nor (n1002,n1003,n1004);
and (n1003,n460,n218);
and (n1004,n376,n221);
and (n1005,n1001,n1006);
xnor (n1006,n1007,n47);
nor (n1007,n1008,n1009);
and (n1008,n593,n112);
and (n1009,n529,n115);
and (n1010,n997,n1006);
and (n1011,n995,n1012);
xor (n1012,n1013,n897);
xor (n1013,n888,n892);
and (n1014,n979,n1012);
and (n1015,n1016,n1018);
xor (n1016,n1017,n22);
xor (n1017,n902,n906);
xor (n1018,n1019,n924);
xor (n1019,n915,n919);
and (n1020,n1015,n1021);
xor (n1021,n1022,n937);
xor (n1022,n932,n934);
and (n1023,n977,n1021);
xor (n1024,n1025,n940);
xor (n1025,n884,n930);
and (n1026,n1024,n1027);
xor (n1027,n943,n945);
and (n1028,n975,n1027);
and (n1029,n1030,n1031);
xor (n1030,n967,n973);
or (n1031,n1032,n1086);
and (n1032,n1033,n1035);
xor (n1033,n1034,n1027);
xor (n1034,n975,n1024);
or (n1035,n1036,n1082,n1085);
and (n1036,n1037,n1080);
or (n1037,n1038,n1077,n1079);
and (n1038,n1039,n1075);
or (n1039,n1040,n1069,n1074);
and (n1040,n1041,n1053);
or (n1041,n1042,n1051,n1052);
and (n1042,n1043,n1047);
xnor (n1043,n1044,n423);
nor (n1044,n1045,n1046);
and (n1045,n93,n758);
and (n1046,n89,n760);
xnor (n1047,n1048,n419);
nor (n1048,n1049,n1050);
and (n1049,n166,n571);
and (n1050,n163,n574);
and (n1051,n1047,n6);
and (n1052,n1043,n6);
or (n1053,n1054,n1063,n1068);
and (n1054,n1055,n1059);
xnor (n1055,n1056,n315);
nor (n1056,n1057,n1058);
and (n1057,n260,n427);
and (n1058,n205,n430);
xnor (n1059,n1060,n210);
nor (n1060,n1061,n1062);
and (n1061,n376,n323);
and (n1062,n371,n326);
and (n1063,n1059,n1064);
xnor (n1064,n1065,n104);
nor (n1065,n1066,n1067);
and (n1066,n529,n218);
and (n1067,n460,n221);
and (n1068,n1055,n1064);
and (n1069,n1053,n1070);
xnor (n1070,n1071,n6);
nor (n1071,n1072,n1073);
and (n1072,n845,n55);
and (n1073,n687,n58);
and (n1074,n1041,n1070);
xor (n1075,n1076,n1012);
xor (n1076,n979,n995);
and (n1077,n1075,n1078);
xor (n1078,n1016,n1018);
and (n1079,n1039,n1078);
xor (n1080,n1081,n913);
xor (n1081,n886,n900);
and (n1082,n1080,n1083);
xor (n1083,n1084,n1021);
xor (n1084,n977,n1015);
and (n1085,n1037,n1083);
and (n1086,n1087,n1088);
xor (n1087,n1033,n1035);
or (n1088,n1089,n1159);
and (n1089,n1090,n1092);
xor (n1090,n1091,n1083);
xor (n1091,n1037,n1080);
or (n1092,n1093,n1155,n1158);
and (n1093,n1094,n1150);
or (n1094,n1095,n1146,n1149);
and (n1095,n1096,n1136);
or (n1096,n1097,n1130,n1135);
and (n1097,n1098,n1114);
or (n1098,n1099,n1108,n1113);
and (n1099,n1100,n1104);
xnor (n1100,n1101,n210);
nor (n1101,n1102,n1103);
and (n1102,n460,n323);
and (n1103,n376,n326);
xnor (n1104,n1105,n104);
nor (n1105,n1106,n1107);
and (n1106,n593,n218);
and (n1107,n529,n221);
and (n1108,n1104,n1109);
xnor (n1109,n1110,n47);
nor (n1110,n1111,n1112);
and (n1111,n845,n112);
and (n1112,n687,n115);
and (n1113,n1100,n1109);
or (n1114,n1115,n1124,n1129);
and (n1115,n1116,n1120);
xnor (n1116,n1117,n423);
nor (n1117,n1118,n1119);
and (n1118,n163,n758);
and (n1119,n93,n760);
xnor (n1120,n1121,n419);
nor (n1121,n1122,n1123);
and (n1122,n205,n571);
and (n1123,n166,n574);
and (n1124,n1120,n1125);
xnor (n1125,n1126,n315);
nor (n1126,n1127,n1128);
and (n1127,n371,n427);
and (n1128,n260,n430);
and (n1129,n1116,n1125);
and (n1130,n1114,n1131);
xnor (n1131,n1132,n47);
nor (n1132,n1133,n1134);
and (n1133,n687,n112);
and (n1134,n593,n115);
and (n1135,n1098,n1131);
or (n1136,n1137,n1142,n1145);
and (n1137,n1138,n1140);
xnor (n1138,n1139,n6);
nand (n1139,n845,n58);
xor (n1140,n1141,n6);
xor (n1141,n1043,n1047);
and (n1142,n1140,n1143);
xor (n1143,n1144,n1064);
xor (n1144,n1055,n1059);
and (n1145,n1138,n1143);
and (n1146,n1136,n1147);
xor (n1147,n1148,n1006);
xor (n1148,n997,n1001);
and (n1149,n1096,n1147);
and (n1150,n1151,n1153);
xor (n1151,n1152,n990);
xor (n1152,n981,n985);
xor (n1153,n1154,n1070);
xor (n1154,n1041,n1053);
and (n1155,n1150,n1156);
xor (n1156,n1157,n1078);
xor (n1157,n1039,n1075);
and (n1158,n1094,n1156);
and (n1159,n1160,n1161);
xor (n1160,n1090,n1092);
or (n1161,n1162,n1214);
and (n1162,n1163,n1165);
xor (n1163,n1164,n1156);
xor (n1164,n1094,n1150);
or (n1165,n1166,n1211,n1213);
and (n1166,n1167,n1209);
or (n1167,n1168,n1205,n1208);
and (n1168,n1169,n1203);
or (n1169,n1170,n1199,n1202);
and (n1170,n1171,n1187);
or (n1171,n1172,n1181,n1186);
and (n1172,n1173,n1177);
xnor (n1173,n1174,n315);
nor (n1174,n1175,n1176);
and (n1175,n376,n427);
and (n1176,n371,n430);
xnor (n1177,n1178,n210);
nor (n1178,n1179,n1180);
and (n1179,n529,n323);
and (n1180,n460,n326);
and (n1181,n1177,n1182);
xnor (n1182,n1183,n104);
nor (n1183,n1184,n1185);
and (n1184,n687,n218);
and (n1185,n593,n221);
and (n1186,n1173,n1182);
or (n1187,n1188,n1197,n1198);
and (n1188,n1189,n1193);
xnor (n1189,n1190,n423);
nor (n1190,n1191,n1192);
and (n1191,n166,n758);
and (n1192,n163,n760);
xnor (n1193,n1194,n419);
nor (n1194,n1195,n1196);
and (n1195,n260,n571);
and (n1196,n205,n574);
and (n1197,n1193,n47);
and (n1198,n1189,n47);
and (n1199,n1187,n1200);
xor (n1200,n1201,n1109);
xor (n1201,n1100,n1104);
and (n1202,n1171,n1200);
xor (n1203,n1204,n1131);
xor (n1204,n1098,n1114);
and (n1205,n1203,n1206);
xor (n1206,n1207,n1143);
xor (n1207,n1138,n1140);
and (n1208,n1169,n1206);
xor (n1209,n1210,n1147);
xor (n1210,n1096,n1136);
and (n1211,n1209,n1212);
xor (n1212,n1151,n1153);
and (n1213,n1167,n1212);
and (n1214,n1215,n1216);
xor (n1215,n1163,n1165);
or (n1216,n1217,n1255);
and (n1217,n1218,n1220);
xor (n1218,n1219,n1212);
xor (n1219,n1167,n1209);
and (n1220,n1221,n1253);
or (n1221,n1222,n1249,n1252);
and (n1222,n1223,n1247);
or (n1223,n1224,n1243,n1246);
and (n1224,n1225,n1241);
or (n1225,n1226,n1235,n1240);
and (n1226,n1227,n1231);
xnor (n1227,n1228,n423);
nor (n1228,n1229,n1230);
and (n1229,n205,n758);
and (n1230,n166,n760);
xnor (n1231,n1232,n419);
nor (n1232,n1233,n1234);
and (n1233,n371,n571);
and (n1234,n260,n574);
and (n1235,n1231,n1236);
xnor (n1236,n1237,n315);
nor (n1237,n1238,n1239);
and (n1238,n460,n427);
and (n1239,n376,n430);
and (n1240,n1227,n1236);
xnor (n1241,n1242,n47);
nand (n1242,n845,n115);
and (n1243,n1241,n1244);
xor (n1244,n1245,n1182);
xor (n1245,n1173,n1177);
and (n1246,n1225,n1244);
xor (n1247,n1248,n1125);
xor (n1248,n1116,n1120);
and (n1249,n1247,n1250);
xor (n1250,n1251,n1200);
xor (n1251,n1171,n1187);
and (n1252,n1223,n1250);
xor (n1253,n1254,n1206);
xor (n1254,n1169,n1203);
and (n1255,n1256,n1257);
xor (n1256,n1218,n1220);
or (n1257,n1258,n1310);
and (n1258,n1259,n1260);
xor (n1259,n1221,n1253);
and (n1260,n1261,n1308);
or (n1261,n1262,n1304,n1307);
and (n1262,n1263,n1297);
or (n1263,n1264,n1291,n1296);
and (n1264,n1265,n1279);
or (n1265,n1266,n1275,n1278);
and (n1266,n1267,n1271);
xnor (n1267,n1268,n315);
nor (n1268,n1269,n1270);
and (n1269,n529,n427);
and (n1270,n460,n430);
xnor (n1271,n1272,n210);
nor (n1272,n1273,n1274);
and (n1273,n687,n323);
and (n1274,n593,n326);
and (n1275,n1271,n1276);
xnor (n1276,n1277,n104);
nand (n1277,n845,n221);
and (n1278,n1267,n1276);
or (n1279,n1280,n1289,n1290);
and (n1280,n1281,n1285);
xnor (n1281,n1282,n423);
nor (n1282,n1283,n1284);
and (n1283,n260,n758);
and (n1284,n205,n760);
xnor (n1285,n1286,n419);
nor (n1286,n1287,n1288);
and (n1287,n376,n571);
and (n1288,n371,n574);
and (n1289,n1285,n104);
and (n1290,n1281,n104);
and (n1291,n1279,n1292);
xnor (n1292,n1293,n210);
nor (n1293,n1294,n1295);
and (n1294,n593,n323);
and (n1295,n529,n326);
and (n1296,n1265,n1292);
and (n1297,n1298,n1302);
xnor (n1298,n1299,n104);
nor (n1299,n1300,n1301);
and (n1300,n845,n218);
and (n1301,n687,n221);
xor (n1302,n1303,n1236);
xor (n1303,n1227,n1231);
and (n1304,n1297,n1305);
xor (n1305,n1306,n47);
xor (n1306,n1189,n1193);
and (n1307,n1263,n1305);
xor (n1308,n1309,n1250);
xor (n1309,n1223,n1247);
and (n1310,n1311,n1312);
xor (n1311,n1259,n1260);
or (n1312,n1313,n1320);
and (n1313,n1314,n1315);
xor (n1314,n1261,n1308);
and (n1315,n1316,n1318);
xor (n1316,n1317,n1244);
xor (n1317,n1225,n1241);
xor (n1318,n1319,n1305);
xor (n1319,n1263,n1297);
and (n1320,n1321,n1322);
xor (n1321,n1314,n1315);
or (n1322,n1323,n1356);
and (n1323,n1324,n1325);
xor (n1324,n1316,n1318);
or (n1325,n1326,n1353,n1355);
and (n1326,n1327,n1351);
or (n1327,n1328,n1347,n1350);
and (n1328,n1329,n1345);
or (n1329,n1330,n1339,n1344);
and (n1330,n1331,n1335);
xnor (n1331,n1332,n423);
nor (n1332,n1333,n1334);
and (n1333,n371,n758);
and (n1334,n260,n760);
xnor (n1335,n1336,n419);
nor (n1336,n1337,n1338);
and (n1337,n460,n571);
and (n1338,n376,n574);
and (n1339,n1335,n1340);
xnor (n1340,n1341,n315);
nor (n1341,n1342,n1343);
and (n1342,n593,n427);
and (n1343,n529,n430);
and (n1344,n1331,n1340);
xor (n1345,n1346,n1276);
xor (n1346,n1267,n1271);
and (n1347,n1345,n1348);
xor (n1348,n1349,n104);
xor (n1349,n1281,n1285);
and (n1350,n1329,n1348);
xor (n1351,n1352,n1292);
xor (n1352,n1265,n1279);
and (n1353,n1351,n1354);
xor (n1354,n1298,n1302);
and (n1355,n1327,n1354);
and (n1356,n1357,n1358);
xor (n1357,n1324,n1325);
or (n1358,n1359,n1392);
and (n1359,n1360,n1362);
xor (n1360,n1361,n1354);
xor (n1361,n1327,n1351);
and (n1362,n1363,n1390);
or (n1363,n1364,n1384,n1389);
and (n1364,n1365,n1377);
or (n1365,n1366,n1375,n1376);
and (n1366,n1367,n1371);
xnor (n1367,n1368,n423);
nor (n1368,n1369,n1370);
and (n1369,n376,n758);
and (n1370,n371,n760);
xnor (n1371,n1372,n419);
nor (n1372,n1373,n1374);
and (n1373,n529,n571);
and (n1374,n460,n574);
and (n1375,n1371,n210);
and (n1376,n1367,n210);
and (n1377,n1378,n1382);
xnor (n1378,n1379,n315);
nor (n1379,n1380,n1381);
and (n1380,n687,n427);
and (n1381,n593,n430);
xnor (n1382,n1383,n210);
nand (n1383,n845,n326);
and (n1384,n1377,n1385);
xnor (n1385,n1386,n210);
nor (n1386,n1387,n1388);
and (n1387,n845,n323);
and (n1388,n687,n326);
and (n1389,n1365,n1385);
xor (n1390,n1391,n1348);
xor (n1391,n1329,n1345);
and (n1392,n1393,n1394);
xor (n1393,n1360,n1362);
or (n1394,n1395,n1402);
and (n1395,n1396,n1397);
xor (n1396,n1363,n1390);
and (n1397,n1398,n1400);
xor (n1398,n1399,n1340);
xor (n1399,n1331,n1335);
xor (n1400,n1401,n1385);
xor (n1401,n1365,n1377);
and (n1402,n1403,n1404);
xor (n1403,n1396,n1397);
or (n1404,n1405,n1430);
and (n1405,n1406,n1407);
xor (n1406,n1398,n1400);
or (n1407,n1408,n1427,n1429);
and (n1408,n1409,n1425);
or (n1409,n1410,n1419,n1424);
and (n1410,n1411,n1415);
xnor (n1411,n1412,n423);
nor (n1412,n1413,n1414);
and (n1413,n460,n758);
and (n1414,n376,n760);
xnor (n1415,n1416,n419);
nor (n1416,n1417,n1418);
and (n1417,n593,n571);
and (n1418,n529,n574);
and (n1419,n1415,n1420);
xnor (n1420,n1421,n315);
nor (n1421,n1422,n1423);
and (n1422,n845,n427);
and (n1423,n687,n430);
and (n1424,n1411,n1420);
xor (n1425,n1426,n210);
xor (n1426,n1367,n1371);
and (n1427,n1425,n1428);
xor (n1428,n1378,n1382);
and (n1429,n1409,n1428);
and (n1430,n1431,n1432);
xor (n1431,n1406,n1407);
or (n1432,n1433,n1451);
and (n1433,n1434,n1436);
xor (n1434,n1435,n1428);
xor (n1435,n1409,n1425);
and (n1436,n1437,n1449);
or (n1437,n1438,n1447,n1448);
and (n1438,n1439,n1443);
xnor (n1439,n1440,n423);
nor (n1440,n1441,n1442);
and (n1441,n529,n758);
and (n1442,n460,n760);
xnor (n1443,n1444,n419);
nor (n1444,n1445,n1446);
and (n1445,n687,n571);
and (n1446,n593,n574);
and (n1447,n1443,n315);
and (n1448,n1439,n315);
xor (n1449,n1450,n1420);
xor (n1450,n1411,n1415);
and (n1451,n1452,n1453);
xor (n1452,n1434,n1436);
or (n1453,n1454,n1461);
and (n1454,n1455,n1456);
xor (n1455,n1437,n1449);
and (n1456,n1457,n1459);
xnor (n1457,n1458,n315);
nand (n1458,n845,n430);
xor (n1459,n1460,n315);
xor (n1460,n1439,n1443);
and (n1461,n1462,n1463);
xor (n1462,n1455,n1456);
or (n1463,n1464,n1475);
and (n1464,n1465,n1466);
xor (n1465,n1457,n1459);
and (n1466,n1467,n1471);
xnor (n1467,n1468,n423);
nor (n1468,n1469,n1470);
and (n1469,n593,n758);
and (n1470,n529,n760);
xnor (n1471,n1472,n419);
nor (n1472,n1473,n1474);
and (n1473,n845,n571);
and (n1474,n687,n574);
and (n1475,n1476,n1477);
xor (n1476,n1465,n1466);
or (n1477,n1478,n1485);
and (n1478,n1479,n1480);
xor (n1479,n1467,n1471);
and (n1480,n1481,n419);
xnor (n1481,n1482,n423);
nor (n1482,n1483,n1484);
and (n1483,n687,n758);
and (n1484,n593,n760);
and (n1485,n1486,n1487);
xor (n1486,n1479,n1480);
or (n1487,n1488,n1492);
and (n1488,n1489,n1491);
xnor (n1489,n1490,n419);
nand (n1490,n845,n574);
xor (n1491,n1481,n419);
and (n1492,n1493,n1494);
xor (n1493,n1489,n1491);
and (n1494,n1495,n1499);
xnor (n1495,n1496,n423);
nor (n1496,n1497,n1498);
and (n1497,n845,n758);
and (n1498,n687,n760);
and (n1499,n1500,n423);
xnor (n1500,n1501,n423);
nand (n1501,n845,n760);
xor (n1502,n1503,n1513);
xor (n1503,n1504,n1508);
xor (n1504,n1505,n30);
xor (n1505,n1506,n1507);
or (n1506,n12,n26);
not (n1507,n22);
and (n1508,n1509,n1512);
or (n1509,n1510,n39,n1511);
and (n1510,n5,n35);
and (n1511,n5,n40);
xnor (n1512,n12,n26);
or (n1513,n1514,n1530);
and (n1514,n1515,n1516);
xor (n1515,n1509,n1512);
or (n1516,n1517,n1527,n1529);
and (n1517,n1518,n1521);
or (n1518,n59,n1519,n1520);
and (n1519,n60,n95);
and (n1520,n52,n95);
or (n1521,n1522,n1525);
or (n1522,n1523,n85,n1524);
and (n1523,n46,n81);
and (n1524,n46,n86);
xor (n1525,n1526,n95);
xor (n1526,n52,n60);
and (n1527,n1521,n1528);
not (n1528,n65);
and (n1529,n1518,n1528);
and (n1530,n1531,n1532);
xor (n1531,n1515,n1516);
or (n1532,n1533,n1565);
and (n1533,n1534,n1536);
xor (n1534,n1535,n1528);
xor (n1535,n1518,n1521);
or (n1536,n1537,n1562,n1564);
and (n1537,n1538,n1545);
or (n1538,n1539,n1543,n1544);
and (n1539,n1540,n174);
or (n1540,n116,n1541,n1542);
and (n1541,n117,n168);
and (n1542,n109,n168);
and (n1543,n174,n92);
and (n1544,n1540,n92);
or (n1545,n1546,n1558,n1561);
and (n1546,n1547,n1557);
or (n1547,n1548,n1554,n1556);
and (n1548,n1549,n1552);
or (n1549,n1550,n153,n1551);
and (n1550,n103,n149);
and (n1551,n103,n154);
xor (n1552,n1553,n168);
xor (n1553,n109,n117);
and (n1554,n1552,n1555);
not (n1555,n174);
and (n1556,n1549,n1555);
not (n1557,n122);
and (n1558,n1557,n1559);
xor (n1559,n1560,n92);
xor (n1560,n1540,n174);
and (n1561,n1547,n1559);
and (n1562,n1545,n1563);
xnor (n1563,n1522,n1525);
and (n1564,n1538,n1563);
and (n1565,n1566,n1567);
xor (n1566,n1534,n1536);
or (n1567,n1568,n1590);
and (n1568,n1569,n1571);
xor (n1569,n1570,n1563);
xor (n1570,n1538,n1545);
and (n1571,n1572,n1588);
or (n1572,n1573,n1584,n1587);
and (n1573,n1574,n1582);
or (n1574,n1575,n1580,n1581);
and (n1575,n1576,n1579);
or (n1576,n222,n1577,n1578);
and (n1577,n223,n195);
and (n1578,n215,n195);
or (n1579,n199,n204);
and (n1580,n1579,n160);
and (n1581,n1576,n160);
and (n1582,n165,n1583);
not (n1583,n278);
and (n1584,n1582,n1585);
xor (n1585,n1586,n1555);
xor (n1586,n1549,n1552);
and (n1587,n1574,n1585);
xor (n1588,n1589,n1559);
xor (n1589,n1547,n1557);
and (n1590,n1591,n1592);
xor (n1591,n1569,n1571);
or (n1592,n1593,n1613);
and (n1593,n1594,n1595);
xor (n1594,n1572,n1588);
and (n1595,n1596,n1611);
or (n1596,n1597,n1608,n1610);
and (n1597,n1598,n1606);
or (n1598,n1599,n1603,n1605);
and (n1599,n248,n1600);
or (n1600,n1601,n268,n1602);
and (n1601,n209,n264);
and (n1602,n209,n269);
and (n1603,n1600,n1604);
xnor (n1604,n199,n204);
and (n1605,n248,n1604);
xor (n1606,n1607,n160);
xor (n1607,n1576,n1579);
and (n1608,n1606,n1609);
xor (n1609,n165,n1583);
and (n1610,n1598,n1609);
xor (n1611,n1612,n1585);
xor (n1612,n1574,n1582);
and (n1613,n1614,n1615);
xor (n1614,n1594,n1595);
or (n1615,n1616,n1639);
and (n1616,n1617,n1618);
xor (n1617,n1596,n1611);
and (n1618,n1619,n1637);
or (n1619,n1620,n1633,n1636);
and (n1620,n1621,n1631);
or (n1621,n1622,n1629,n1630);
and (n1622,n1623,n1626);
or (n1623,n306,n1624,n1625);
and (n1624,n307,n380);
and (n1625,n302,n380);
or (n1626,n327,n1627,n1628);
and (n1627,n328,n298);
and (n1628,n320,n298);
and (n1629,n1626,n388);
and (n1630,n1623,n388);
xor (n1631,n1632,n195);
xor (n1632,n215,n223);
and (n1633,n1631,n1634);
xor (n1634,n1635,n1604);
xor (n1635,n248,n1600);
and (n1636,n1621,n1634);
xor (n1637,n1638,n1609);
xor (n1638,n1598,n1606);
and (n1639,n1640,n1641);
xor (n1640,n1617,n1618);
or (n1641,n1642,n1691);
and (n1642,n1643,n1644);
xor (n1643,n1619,n1637);
or (n1644,n1645,n1687,n1690);
and (n1645,n1646,n1657);
or (n1646,n1647,n1653,n1656);
and (n1647,n1648,n1652);
or (n1648,n1649,n357);
or (n1649,n1650,n351,n1651);
and (n1650,n314,n347);
and (n1651,n314,n352);
not (n1652,n392);
and (n1653,n1652,n1654);
xor (n1654,n1655,n388);
xor (n1655,n1623,n1626);
and (n1656,n1648,n1654);
or (n1657,n1658,n1683,n1686);
and (n1658,n1659,n1679);
or (n1659,n1660,n1675,n1678);
and (n1660,n1661,n1671);
or (n1661,n1662,n1669,n1670);
and (n1662,n1663,n1666);
or (n1663,n431,n1664,n1665);
and (n1664,n432,n439);
and (n1665,n424,n439);
or (n1666,n447,n1667,n1668);
and (n1667,n448,n455);
and (n1668,n443,n455);
and (n1669,n1666,n459);
and (n1670,n1663,n459);
or (n1671,n1672,n1673,n1674);
and (n1672,n375,n543);
and (n1673,n543,n466);
and (n1674,n375,n466);
and (n1675,n1671,n1676);
xor (n1676,n1677,n380);
xor (n1677,n302,n307);
and (n1678,n1661,n1676);
and (n1679,n1680,n1682);
xor (n1680,n1681,n298);
xor (n1681,n320,n328);
xnor (n1682,n1649,n357);
and (n1683,n1679,n1684);
xor (n1684,n1685,n1654);
xor (n1685,n1648,n1652);
and (n1686,n1659,n1684);
and (n1687,n1657,n1688);
xor (n1688,n1689,n1634);
xor (n1689,n1621,n1631);
and (n1690,n1646,n1688);
and (n1691,n1692,n1693);
xor (n1692,n1643,n1644);
or (n1693,n1694,n1728);
and (n1694,n1695,n1697);
xor (n1695,n1696,n1688);
xor (n1696,n1646,n1657);
and (n1697,n1698,n1726);
or (n1698,n1699,n1723,n1725);
and (n1699,n1700,n1721);
or (n1700,n1701,n1719,n1720);
and (n1701,n1702,n1710);
or (n1702,n1703,n1707,n1709);
and (n1703,n1704,n506);
or (n1704,n1705,n500,n1706);
and (n1705,n418,n496);
and (n1706,n418,n501);
and (n1707,n506,n1708);
and (n1708,n524,n528);
and (n1709,n1704,n1708);
or (n1710,n1711,n1716,n1718);
and (n1711,n1712,n1714);
xor (n1712,n1713,n439);
xor (n1713,n424,n432);
xor (n1714,n1715,n455);
xor (n1715,n443,n448);
and (n1716,n1714,n1717);
not (n1717,n459);
and (n1718,n1712,n1717);
and (n1719,n1710,n541);
and (n1720,n1702,n541);
xor (n1721,n1722,n1676);
xor (n1722,n1661,n1671);
and (n1723,n1721,n1724);
xor (n1724,n1680,n1682);
and (n1725,n1700,n1724);
xor (n1726,n1727,n1684);
xor (n1727,n1659,n1679);
and (n1728,n1729,n1730);
xor (n1729,n1695,n1697);
or (n1730,n1731,n1765);
and (n1731,n1732,n1733);
xor (n1732,n1698,n1726);
and (n1733,n1734,n1763);
or (n1734,n1735,n1759,n1762);
and (n1735,n1736,n1757);
or (n1736,n1737,n1753,n1756);
and (n1737,n1738,n1749);
or (n1738,n1739,n1746,n1748);
and (n1739,n1740,n1743);
or (n1740,n575,n1741,n1742);
and (n1741,n576,n598);
and (n1742,n568,n598);
or (n1743,n606,n1744,n1745);
and (n1744,n607,n583);
and (n1745,n602,n583);
and (n1746,n1743,n1747);
or (n1747,n587,n592);
and (n1748,n1740,n1747);
or (n1749,n1750,n1751,n1752);
and (n1750,n698,n617);
and (n1751,n617,n699);
and (n1752,n698,n699);
and (n1753,n1749,n1754);
xor (n1754,n1755,n1717);
xor (n1755,n1712,n1714);
and (n1756,n1738,n1754);
xor (n1757,n1758,n459);
xor (n1758,n1663,n1666);
and (n1759,n1757,n1760);
xor (n1760,n1761,n541);
xor (n1761,n1702,n1710);
and (n1762,n1736,n1760);
xor (n1763,n1764,n1724);
xor (n1764,n1700,n1721);
and (n1765,n1766,n1767);
xor (n1766,n1732,n1733);
or (n1767,n1768,n1800);
and (n1768,n1769,n1770);
xor (n1769,n1734,n1763);
and (n1770,n1771,n1798);
or (n1771,n1772,n1794,n1797);
and (n1772,n1773,n1792);
or (n1773,n1774,n1790,n1791);
and (n1774,n1775,n1781);
or (n1775,n1776,n1780,n689);
and (n1776,n646,n1777);
or (n1777,n1778,n668,n1779);
and (n1778,n567,n664);
and (n1779,n567,n669);
and (n1780,n1777,n675);
or (n1781,n1782,n1787,n1789);
and (n1782,n1783,n1785);
xor (n1783,n1784,n598);
xor (n1784,n568,n576);
xor (n1785,n1786,n583);
xor (n1786,n602,n607);
and (n1787,n1785,n1788);
xnor (n1788,n587,n592);
and (n1789,n1783,n1788);
and (n1790,n1781,n696);
and (n1791,n1775,n696);
xor (n1792,n1793,n1708);
xor (n1793,n1704,n506);
and (n1794,n1792,n1795);
xor (n1795,n1796,n1754);
xor (n1796,n1738,n1749);
and (n1797,n1773,n1795);
xor (n1798,n1799,n1760);
xor (n1799,n1736,n1757);
and (n1800,n1801,n1802);
xor (n1801,n1769,n1770);
or (n1802,n1803,n1823);
and (n1803,n1804,n1805);
xor (n1804,n1771,n1798);
and (n1805,n1806,n1821);
or (n1806,n1807,n1817,n1820);
and (n1807,n1808,n1815);
or (n1808,n1809,n1811,n1814);
and (n1809,n719,n1810);
or (n1810,n769,n774);
and (n1811,n1810,n1812);
xor (n1812,n1813,n1788);
xor (n1813,n1783,n1785);
and (n1814,n719,n1812);
xor (n1815,n1816,n1747);
xor (n1816,n1740,n1743);
and (n1817,n1815,n1818);
xor (n1818,n1819,n696);
xor (n1819,n1775,n1781);
and (n1820,n1808,n1818);
xor (n1821,n1822,n1795);
xor (n1822,n1773,n1792);
and (n1823,n1824,n1825);
xor (n1824,n1804,n1805);
or (n1825,n1826,n1842);
and (n1826,n1827,n1828);
xor (n1827,n1806,n1821);
and (n1828,n1829,n1840);
or (n1829,n1830,n1836,n1839);
and (n1830,n1831,n1834);
or (n1831,n801,n1832,n1833);
and (n1832,n848,n970);
and (n1833,n802,n970);
xor (n1834,n1835,n675);
xor (n1835,n646,n1777);
and (n1836,n1834,n1837);
xor (n1837,n1838,n1812);
xor (n1838,n719,n1810);
and (n1839,n1831,n1837);
xor (n1840,n1841,n1818);
xor (n1841,n1808,n1815);
and (n1842,n1843,n1844);
xor (n1843,n1827,n1828);
or (n1844,n1845,n1853);
and (n1845,n1846,n1847);
xor (n1846,n1829,n1840);
and (n1847,n1848,n1851);
or (n1848,n881,n1849,n1850);
and (n1849,n942,n972);
and (n1850,n882,n972);
xor (n1851,n1852,n1837);
xor (n1852,n1831,n1834);
and (n1853,n1854,n1855);
xor (n1854,n1846,n1847);
or (n1855,n1856,n963);
and (n1856,n1857,n1858);
xor (n1857,n1848,n1851);
or (n1858,n1859,n1860,n1861);
and (n1859,n948,n969);
and (n1860,n969,n971);
and (n1861,n948,n971);
endmodule
