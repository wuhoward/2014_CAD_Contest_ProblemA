module top (out,n13,n16,n17,n20,n22,n29,n32,n33,n37
        ,n45,n48,n49,n53,n62,n65,n66,n70,n73,n74
        ,n84,n87,n91,n178,n183,n254,n255,n292,n360,n423
        ,n519,n590,n676);
output out;
input n13;
input n16;
input n17;
input n20;
input n22;
input n29;
input n32;
input n33;
input n37;
input n45;
input n48;
input n49;
input n53;
input n62;
input n65;
input n66;
input n70;
input n73;
input n74;
input n84;
input n87;
input n91;
input n178;
input n183;
input n254;
input n255;
input n292;
input n360;
input n423;
input n519;
input n590;
input n676;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n14;
wire n15;
wire n18;
wire n19;
wire n21;
wire n23;
wire n24;
wire n25;
wire n26;
wire n27;
wire n28;
wire n30;
wire n31;
wire n34;
wire n35;
wire n36;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n46;
wire n47;
wire n50;
wire n51;
wire n52;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n63;
wire n64;
wire n67;
wire n68;
wire n69;
wire n71;
wire n72;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n85;
wire n86;
wire n88;
wire n89;
wire n90;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n179;
wire n180;
wire n181;
wire n182;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
xor (out,n0,n1360);
buf (n0,n1);
xor (n1,n2,n315);
xor (n2,n3,n241);
xor (n3,n4,n207);
xor (n4,n5,n146);
or (n5,n6,n106,n145);
nand (n6,n7,n96);
or (n7,n8,n58);
or (n8,n9,n41,n57);
and (n9,n10,n26);
xnor (n10,n11,n23);
nor (n11,n12,n21);
and (n12,n13,n14);
and (n14,n15,n18);
xor (n15,n16,n17);
not (n18,n19);
xor (n19,n17,n20);
and (n21,n22,n19);
and (n23,n16,n24);
not (n24,n25);
and (n25,n17,n20);
xnor (n26,n27,n38);
nor (n27,n28,n36);
and (n28,n29,n30);
and (n30,n31,n34);
xor (n31,n32,n33);
not (n34,n35);
xor (n35,n33,n16);
and (n36,n37,n35);
and (n38,n32,n39);
not (n39,n40);
and (n40,n33,n16);
and (n41,n26,n42);
xnor (n42,n43,n54);
nor (n43,n44,n52);
and (n44,n45,n46);
and (n46,n47,n50);
xor (n47,n48,n49);
not (n50,n51);
xor (n51,n49,n32);
and (n52,n53,n51);
and (n54,n48,n55);
not (n55,n56);
and (n56,n49,n32);
and (n57,n10,n42);
or (n58,n59,n80,n95);
and (n59,n60,n67);
not (n60,n61);
and (n61,n62,n63);
not (n63,n64);
and (n64,n65,n66);
xnor (n67,n68,n77);
not (n68,n69);
and (n69,n70,n71);
and (n71,n72,n75);
xor (n72,n73,n74);
not (n75,n76);
xor (n76,n74,n62);
and (n77,n73,n78);
not (n78,n79);
and (n79,n74,n62);
and (n80,n67,n81);
xnor (n81,n82,n92);
nor (n82,n83,n90);
and (n83,n84,n85);
and (n85,n86,n88);
xor (n86,n20,n87);
not (n88,n89);
xor (n89,n87,n73);
and (n90,n91,n89);
and (n92,n20,n93);
not (n93,n94);
and (n94,n87,n73);
and (n95,n60,n81);
xor (n96,n97,n102);
xor (n97,n98,n99);
not (n98,n77);
xnor (n99,n100,n92);
not (n100,n101);
and (n101,n70,n85);
xnor (n102,n103,n23);
nor (n103,n104,n105);
and (n104,n84,n14);
and (n105,n91,n19);
and (n106,n96,n107);
xor (n107,n108,n134);
xor (n108,n109,n122);
or (n109,n110,n119,n121);
and (n110,n111,n115);
xnor (n111,n112,n38);
nor (n112,n113,n114);
and (n113,n37,n30);
and (n114,n13,n35);
xnor (n115,n116,n54);
nor (n116,n117,n118);
and (n117,n53,n46);
and (n118,n29,n51);
and (n119,n115,n120);
and (n120,n45,n48);
and (n121,n111,n120);
or (n122,n123,n128,n133);
and (n123,n77,n124);
xnor (n124,n125,n92);
nor (n125,n126,n127);
and (n126,n91,n85);
and (n127,n70,n89);
and (n128,n124,n129);
xnor (n129,n130,n23);
nor (n130,n131,n132);
and (n131,n22,n14);
and (n132,n84,n19);
and (n133,n77,n129);
xor (n134,n135,n144);
xor (n135,n136,n140);
xnor (n136,n137,n38);
nor (n137,n138,n139);
and (n138,n13,n30);
and (n139,n22,n35);
xnor (n140,n141,n54);
nor (n141,n142,n143);
and (n142,n29,n46);
and (n143,n37,n51);
and (n144,n53,n48);
and (n145,n7,n107);
or (n146,n147,n203,n206);
and (n147,n148,n198);
or (n148,n149,n194,n197);
and (n149,n150,n185);
or (n150,n151,n181,n184);
and (n151,n152,n164);
or (n152,n153,n158,n163);
and (n153,n61,n154);
xnor (n154,n155,n77);
nor (n155,n156,n157);
and (n156,n91,n71);
and (n157,n70,n76);
and (n158,n154,n159);
xnor (n159,n160,n92);
nor (n160,n161,n162);
and (n161,n22,n85);
and (n162,n84,n89);
and (n163,n61,n159);
or (n164,n165,n174,n180);
and (n165,n166,n170);
xnor (n166,n167,n23);
nor (n167,n168,n169);
and (n168,n37,n14);
and (n169,n13,n19);
xnor (n170,n171,n38);
nor (n171,n172,n173);
and (n172,n53,n30);
and (n173,n29,n35);
and (n174,n170,n175);
xnor (n175,n176,n54);
nor (n176,n177,n179);
and (n177,n178,n46);
and (n179,n45,n51);
and (n180,n166,n175);
and (n181,n164,n182);
and (n182,n183,n48);
and (n184,n152,n182);
or (n185,n186,n190,n193);
and (n186,n187,n188);
and (n187,n178,n48);
xor (n188,n189,n42);
xor (n189,n10,n26);
and (n190,n188,n191);
xor (n191,n192,n81);
xor (n192,n60,n67);
and (n193,n187,n191);
and (n194,n185,n195);
xor (n195,n196,n120);
xor (n196,n111,n115);
and (n197,n150,n195);
and (n198,n199,n202);
not (n199,n200);
xor (n200,n201,n129);
xor (n201,n98,n124);
xnor (n202,n8,n58);
and (n203,n198,n204);
xor (n204,n205,n107);
xor (n205,n7,n96);
and (n206,n148,n204);
xor (n207,n208,n225);
xor (n208,n209,n213);
or (n209,n210,n211,n212);
and (n210,n109,n122);
and (n211,n122,n134);
and (n212,n109,n134);
not (n213,n214);
xor (n214,n215,n221);
xor (n215,n216,n217);
not (n216,n92);
xnor (n217,n218,n23);
nor (n218,n219,n220);
and (n219,n91,n14);
and (n220,n70,n19);
xnor (n221,n222,n38);
nor (n222,n223,n224);
and (n223,n22,n30);
and (n224,n84,n35);
xor (n225,n226,n235);
xor (n226,n227,n231);
or (n227,n228,n229,n230);
and (n228,n136,n140);
and (n229,n140,n144);
and (n230,n136,n144);
or (n231,n232,n233,n234);
and (n232,n98,n99);
and (n233,n99,n102);
and (n234,n98,n102);
xnor (n235,n236,n240);
xnor (n236,n237,n54);
nor (n237,n238,n239);
and (n238,n37,n46);
and (n239,n13,n51);
and (n240,n29,n48);
and (n241,n242,n313);
or (n242,n243,n310,n312);
and (n243,n244,n308);
or (n244,n245,n304,n307);
and (n245,n246,n294);
or (n246,n247,n285,n293);
and (n247,n248,n269);
or (n248,n249,n263,n268);
and (n249,n250,n256);
not (n250,n251);
and (n251,n66,n252);
not (n252,n253);
and (n253,n254,n255);
xnor (n256,n257,n61);
not (n257,n258);
and (n258,n70,n259);
and (n259,n260,n261);
xor (n260,n62,n65);
not (n261,n262);
xor (n262,n65,n66);
and (n263,n256,n264);
xnor (n264,n265,n77);
nor (n265,n266,n267);
and (n266,n84,n71);
and (n267,n91,n76);
and (n268,n250,n264);
or (n269,n270,n279,n284);
and (n270,n271,n275);
xnor (n271,n272,n92);
nor (n272,n273,n274);
and (n273,n13,n85);
and (n274,n22,n89);
xnor (n275,n276,n23);
nor (n276,n277,n278);
and (n277,n29,n14);
and (n278,n37,n19);
and (n279,n275,n280);
xnor (n280,n281,n38);
nor (n281,n282,n283);
and (n282,n45,n30);
and (n283,n53,n35);
and (n284,n271,n280);
and (n285,n269,n286);
and (n286,n287,n291);
xnor (n287,n288,n54);
nor (n288,n289,n290);
and (n289,n183,n46);
and (n290,n178,n51);
and (n291,n292,n48);
and (n293,n248,n286);
or (n294,n295,n301,n303);
and (n295,n296,n299);
not (n296,n297);
xor (n297,n298,n159);
xor (n298,n60,n154);
xor (n299,n300,n175);
xor (n300,n166,n170);
and (n301,n299,n302);
not (n302,n182);
and (n303,n296,n302);
and (n304,n294,n305);
xor (n305,n306,n191);
xor (n306,n187,n188);
and (n307,n246,n305);
xor (n308,n309,n195);
xor (n309,n150,n185);
and (n310,n308,n311);
xor (n311,n199,n202);
and (n312,n244,n311);
xor (n313,n314,n204);
xor (n314,n148,n198);
or (n315,n316,n383);
and (n316,n317,n318);
xor (n317,n242,n313);
and (n318,n319,n381);
or (n319,n320,n377,n380);
and (n320,n321,n375);
or (n321,n322,n371,n374);
and (n322,n323,n362);
or (n323,n324,n353,n361);
and (n324,n325,n337);
or (n325,n326,n331,n336);
and (n326,n251,n327);
xnor (n327,n328,n61);
nor (n328,n329,n330);
and (n329,n91,n259);
and (n330,n70,n262);
and (n331,n327,n332);
xnor (n332,n333,n77);
nor (n333,n334,n335);
and (n334,n22,n71);
and (n335,n84,n76);
and (n336,n251,n332);
or (n337,n338,n347,n352);
and (n338,n339,n343);
xnor (n339,n340,n92);
nor (n340,n341,n342);
and (n341,n37,n85);
and (n342,n13,n89);
xnor (n343,n344,n23);
nor (n344,n345,n346);
and (n345,n53,n14);
and (n346,n29,n19);
and (n347,n343,n348);
xnor (n348,n349,n38);
nor (n349,n350,n351);
and (n350,n178,n30);
and (n351,n45,n35);
and (n352,n339,n348);
and (n353,n337,n354);
or (n354,n355,n359);
xnor (n355,n356,n54);
nor (n356,n357,n358);
and (n357,n292,n46);
and (n358,n183,n51);
and (n359,n360,n48);
and (n361,n325,n354);
or (n362,n363,n368,n370);
and (n363,n364,n366);
xor (n364,n365,n264);
xor (n365,n250,n256);
xor (n366,n367,n280);
xor (n367,n271,n275);
and (n368,n366,n369);
xor (n369,n287,n291);
and (n370,n364,n369);
and (n371,n362,n372);
xor (n372,n373,n299);
xor (n373,n182,n297);
and (n374,n323,n372);
xor (n375,n376,n182);
xor (n376,n152,n164);
and (n377,n375,n378);
xor (n378,n379,n305);
xor (n379,n246,n294);
and (n380,n321,n378);
xor (n381,n382,n311);
xor (n382,n244,n308);
and (n383,n384,n385);
xor (n384,n317,n318);
or (n385,n386,n466);
and (n386,n387,n388);
xor (n387,n319,n381);
and (n388,n389,n464);
or (n389,n390,n460,n463);
and (n390,n391,n458);
or (n391,n392,n454,n457);
and (n392,n393,n443);
or (n393,n394,n425,n442);
and (n394,n395,n411);
or (n395,n396,n405,n410);
and (n396,n397,n398);
not (n397,n255);
xnor (n398,n399,n251);
not (n399,n400);
and (n400,n70,n401);
and (n401,n402,n403);
xor (n402,n66,n254);
not (n403,n404);
xor (n404,n254,n255);
and (n405,n398,n406);
xnor (n406,n407,n61);
nor (n407,n408,n409);
and (n408,n84,n259);
and (n409,n91,n262);
and (n410,n397,n406);
or (n411,n412,n421,n424);
and (n412,n413,n417);
xnor (n413,n414,n38);
nor (n414,n415,n416);
and (n415,n183,n30);
and (n416,n178,n35);
xnor (n417,n418,n54);
nor (n418,n419,n420);
and (n419,n360,n46);
and (n420,n292,n51);
and (n421,n417,n422);
and (n422,n423,n48);
and (n424,n413,n422);
and (n425,n411,n426);
or (n426,n427,n436,n441);
and (n427,n428,n432);
xnor (n428,n429,n77);
nor (n429,n430,n431);
and (n430,n13,n71);
and (n431,n22,n76);
xnor (n432,n433,n92);
nor (n433,n434,n435);
and (n434,n29,n85);
and (n435,n37,n89);
and (n436,n432,n437);
xnor (n437,n438,n23);
nor (n438,n439,n440);
and (n439,n45,n14);
and (n440,n53,n19);
and (n441,n428,n437);
and (n442,n395,n426);
or (n443,n444,n450,n453);
and (n444,n445,n448);
not (n445,n446);
xor (n446,n447,n332);
xor (n447,n250,n327);
xor (n448,n449,n348);
xor (n449,n339,n343);
and (n450,n448,n451);
not (n451,n452);
xor (n452,n355,n359);
and (n453,n445,n451);
and (n454,n443,n455);
xor (n455,n456,n369);
xor (n456,n364,n366);
and (n457,n393,n455);
xor (n458,n459,n286);
xor (n459,n248,n269);
and (n460,n458,n461);
xor (n461,n462,n372);
xor (n462,n323,n362);
and (n463,n391,n461);
xor (n464,n465,n378);
xor (n465,n321,n375);
and (n466,n467,n468);
xor (n467,n387,n388);
or (n468,n469,n539);
and (n469,n470,n471);
xor (n470,n389,n464);
and (n471,n472,n537);
or (n472,n473,n533,n536);
and (n473,n474,n531);
or (n474,n475,n527,n530);
and (n475,n476,n522);
or (n476,n477,n506,n521);
and (n477,n478,n494);
or (n478,n479,n488,n493);
and (n479,n480,n484);
xnor (n480,n481,n77);
nor (n481,n482,n483);
and (n482,n37,n71);
and (n483,n13,n76);
xnor (n484,n485,n92);
nor (n485,n486,n487);
and (n486,n53,n85);
and (n487,n29,n89);
and (n488,n484,n489);
xnor (n489,n490,n23);
nor (n490,n491,n492);
and (n491,n178,n14);
and (n492,n45,n19);
and (n493,n480,n489);
or (n494,n495,n500,n505);
and (n495,n255,n496);
xnor (n496,n497,n251);
nor (n497,n498,n499);
and (n498,n91,n401);
and (n499,n70,n404);
and (n500,n496,n501);
xnor (n501,n502,n61);
nor (n502,n503,n504);
and (n503,n22,n259);
and (n504,n84,n262);
and (n505,n255,n501);
and (n506,n494,n507);
or (n507,n508,n517,n520);
and (n508,n509,n513);
xnor (n509,n510,n38);
nor (n510,n511,n512);
and (n511,n292,n30);
and (n512,n183,n35);
xnor (n513,n514,n54);
nor (n514,n515,n516);
and (n515,n423,n46);
and (n516,n360,n51);
and (n517,n513,n518);
and (n518,n519,n48);
and (n520,n509,n518);
and (n521,n478,n507);
or (n522,n523,n525);
xor (n523,n524,n422);
xor (n524,n413,n417);
xor (n525,n526,n437);
xor (n526,n428,n432);
and (n527,n522,n528);
xor (n528,n529,n452);
xor (n529,n446,n448);
and (n530,n476,n528);
xor (n531,n532,n354);
xor (n532,n325,n337);
and (n533,n531,n534);
xor (n534,n535,n455);
xor (n535,n393,n443);
and (n536,n474,n534);
xor (n537,n538,n461);
xor (n538,n391,n458);
and (n539,n540,n541);
xor (n540,n470,n471);
or (n541,n542,n622);
and (n542,n543,n544);
xor (n543,n472,n537);
and (n544,n545,n620);
or (n545,n546,n616,n619);
and (n546,n547,n612);
or (n547,n548,n608,n611);
and (n548,n549,n597);
or (n549,n550,n583,n596);
and (n550,n551,n567);
or (n551,n552,n561,n566);
and (n552,n553,n557);
xnor (n553,n554,n61);
nor (n554,n555,n556);
and (n555,n13,n259);
and (n556,n22,n262);
xnor (n557,n558,n77);
nor (n558,n559,n560);
and (n559,n29,n71);
and (n560,n37,n76);
and (n561,n557,n562);
xnor (n562,n563,n92);
nor (n563,n564,n565);
and (n564,n45,n85);
and (n565,n53,n89);
and (n566,n553,n562);
or (n567,n568,n577,n582);
and (n568,n569,n573);
xnor (n569,n570,n23);
nor (n570,n571,n572);
and (n571,n183,n14);
and (n572,n178,n19);
xnor (n573,n574,n38);
nor (n574,n575,n576);
and (n575,n360,n30);
and (n576,n292,n35);
and (n577,n573,n578);
xnor (n578,n579,n54);
nor (n579,n580,n581);
and (n580,n519,n46);
and (n581,n423,n51);
and (n582,n569,n578);
and (n583,n567,n584);
and (n584,n585,n592);
xnor (n585,n586,n255);
not (n586,n587);
and (n587,n70,n588);
and (n588,n589,n591);
xor (n589,n255,n590);
not (n591,n590);
xnor (n592,n593,n251);
nor (n593,n594,n595);
and (n594,n84,n401);
and (n595,n91,n404);
and (n596,n551,n584);
or (n597,n598,n604,n607);
and (n598,n599,n601);
xor (n599,n600,n489);
xor (n600,n480,n484);
not (n601,n602);
xor (n602,n603,n501);
xor (n603,n397,n496);
and (n604,n601,n605);
xor (n605,n606,n518);
xor (n606,n509,n513);
and (n607,n599,n605);
and (n608,n597,n609);
xor (n609,n610,n406);
xor (n610,n397,n398);
and (n611,n549,n609);
and (n612,n613,n615);
xor (n613,n614,n507);
xor (n614,n478,n494);
xnor (n615,n523,n525);
and (n616,n612,n617);
xor (n617,n618,n426);
xor (n618,n395,n411);
and (n619,n547,n617);
xor (n620,n621,n534);
xor (n621,n474,n531);
and (n622,n623,n624);
xor (n623,n543,n544);
or (n624,n625,n704);
and (n625,n626,n627);
xor (n626,n545,n620);
or (n627,n628,n700,n703);
and (n628,n629,n698);
or (n629,n630,n695,n697);
and (n630,n631,n693);
or (n631,n632,n689,n692);
and (n632,n633,n679);
or (n633,n634,n667,n678);
and (n634,n635,n651);
or (n635,n636,n645,n650);
and (n636,n637,n641);
xnor (n637,n638,n255);
nor (n638,n639,n640);
and (n639,n91,n588);
and (n640,n70,n590);
xnor (n641,n642,n251);
nor (n642,n643,n644);
and (n643,n22,n401);
and (n644,n84,n404);
and (n645,n641,n646);
xnor (n646,n647,n61);
nor (n647,n648,n649);
and (n648,n37,n259);
and (n649,n13,n262);
and (n650,n637,n646);
or (n651,n652,n661,n666);
and (n652,n653,n657);
xnor (n653,n654,n77);
nor (n654,n655,n656);
and (n655,n53,n71);
and (n656,n29,n76);
xnor (n657,n658,n92);
nor (n658,n659,n660);
and (n659,n178,n85);
and (n660,n45,n89);
and (n661,n657,n662);
xnor (n662,n663,n23);
nor (n663,n664,n665);
and (n664,n292,n14);
and (n665,n183,n19);
and (n666,n653,n662);
and (n667,n651,n668);
and (n668,n669,n673);
xnor (n669,n670,n38);
nor (n670,n671,n672);
and (n671,n423,n30);
and (n672,n360,n35);
xnor (n673,n674,n54);
nor (n674,n675,n677);
and (n675,n676,n46);
and (n677,n519,n51);
and (n678,n635,n668);
or (n679,n680,n685,n688);
and (n680,n681,n683);
not (n681,n682);
nand (n682,n676,n48);
xor (n683,n684,n562);
xor (n684,n553,n557);
and (n685,n683,n686);
xor (n686,n687,n578);
xor (n687,n569,n573);
and (n688,n681,n686);
and (n689,n679,n690);
xor (n690,n691,n605);
xor (n691,n599,n601);
and (n692,n633,n690);
xor (n693,n694,n609);
xor (n694,n549,n597);
and (n695,n693,n696);
xor (n696,n613,n615);
and (n697,n631,n696);
xor (n698,n699,n617);
xor (n699,n547,n612);
and (n700,n698,n701);
xor (n701,n702,n528);
xor (n702,n476,n522);
and (n703,n629,n701);
and (n704,n705,n706);
xor (n705,n626,n627);
or (n706,n707,n784);
and (n707,n708,n710);
xor (n708,n709,n701);
xor (n709,n629,n698);
and (n710,n711,n782);
or (n711,n712,n778,n781);
and (n712,n713,n773);
or (n713,n714,n770,n772);
and (n714,n715,n761);
or (n715,n716,n743,n760);
and (n716,n717,n731);
or (n717,n718,n727,n730);
and (n718,n719,n723);
xnor (n719,n720,n23);
nor (n720,n721,n722);
and (n721,n360,n14);
and (n722,n292,n19);
xnor (n723,n724,n38);
nor (n724,n725,n726);
and (n725,n519,n30);
and (n726,n423,n35);
and (n727,n723,n728);
xnor (n728,n729,n54);
nand (n729,n676,n51);
and (n730,n719,n728);
or (n731,n732,n741,n742);
and (n732,n733,n737);
xnor (n733,n734,n255);
nor (n734,n735,n736);
and (n735,n84,n588);
and (n736,n91,n590);
xnor (n737,n738,n251);
nor (n738,n739,n740);
and (n739,n13,n401);
and (n740,n22,n404);
and (n741,n737,n54);
and (n742,n733,n54);
and (n743,n731,n744);
or (n744,n745,n754,n759);
and (n745,n746,n750);
xnor (n746,n747,n61);
nor (n747,n748,n749);
and (n748,n29,n259);
and (n749,n37,n262);
xnor (n750,n751,n77);
nor (n751,n752,n753);
and (n752,n45,n71);
and (n753,n53,n76);
and (n754,n750,n755);
xnor (n755,n756,n92);
nor (n756,n757,n758);
and (n757,n183,n85);
and (n758,n178,n89);
and (n759,n746,n755);
and (n760,n717,n744);
or (n761,n762,n767,n769);
and (n762,n763,n765);
xor (n763,n764,n646);
xor (n764,n637,n641);
xor (n765,n766,n662);
xor (n766,n653,n657);
and (n767,n765,n768);
xor (n768,n669,n673);
and (n769,n763,n768);
and (n770,n761,n771);
xor (n771,n585,n592);
and (n772,n715,n771);
and (n773,n774,n776);
xor (n774,n775,n668);
xor (n775,n635,n651);
xor (n776,n777,n686);
xor (n777,n681,n683);
and (n778,n773,n779);
xor (n779,n780,n584);
xor (n780,n551,n567);
and (n781,n713,n779);
xor (n782,n783,n696);
xor (n783,n631,n693);
and (n784,n785,n786);
xor (n785,n708,n710);
or (n786,n787,n794);
and (n787,n788,n789);
xor (n788,n711,n782);
and (n789,n790,n792);
xor (n790,n791,n779);
xor (n791,n713,n773);
xor (n792,n793,n690);
xor (n793,n633,n679);
and (n794,n795,n827);
xor (n795,n796,n821);
xor (n796,n797,n801);
or (n797,n712,n798,n800);
and (n798,n773,n799);
xnor (n799,n599,n605);
and (n800,n713,n799);
xor (n801,n802,n811);
xor (n802,n803,n806);
or (n803,n632,n804,n805);
and (n804,n679,n602);
and (n805,n633,n602);
xor (n806,n807,n507);
xor (n807,n478,n808);
or (n808,n809,n500,n810);
and (n809,n397,n496);
and (n810,n397,n501);
xor (n811,n812,n814);
xor (n812,n549,n813);
or (n813,n599,n605);
xor (n814,n815,n820);
xor (n815,n816,n818);
xor (n816,n817,n428);
xor (n817,n398,n406);
xor (n818,n819,n413);
xor (n819,n432,n437);
xnor (n820,n417,n422);
or (n821,n822,n824,n826);
and (n822,n779,n823);
xor (n823,n793,n602);
and (n824,n823,n825);
xor (n825,n791,n799);
and (n826,n779,n825);
or (n827,n828,n887);
and (n828,n829,n831);
xor (n829,n830,n825);
xor (n830,n779,n823);
or (n831,n832,n884,n886);
and (n832,n833,n882);
or (n833,n834,n878,n881);
and (n834,n835,n873);
or (n835,n836,n869,n872);
and (n836,n837,n853);
or (n837,n838,n847,n852);
and (n838,n839,n843);
xnor (n839,n840,n255);
nor (n840,n841,n842);
and (n841,n22,n588);
and (n842,n84,n590);
xnor (n843,n844,n251);
nor (n844,n845,n846);
and (n845,n37,n401);
and (n846,n13,n404);
and (n847,n843,n848);
xnor (n848,n849,n61);
nor (n849,n850,n851);
and (n850,n53,n259);
and (n851,n29,n262);
and (n852,n839,n848);
or (n853,n854,n863,n868);
and (n854,n855,n859);
xnor (n855,n856,n77);
nor (n856,n857,n858);
and (n857,n178,n71);
and (n858,n45,n76);
xnor (n859,n860,n92);
nor (n860,n861,n862);
and (n861,n292,n85);
and (n862,n183,n89);
and (n863,n859,n864);
xnor (n864,n865,n23);
nor (n865,n866,n867);
and (n866,n423,n14);
and (n867,n360,n19);
and (n868,n855,n864);
and (n869,n853,n870);
xor (n870,n871,n728);
xor (n871,n719,n723);
and (n872,n837,n870);
and (n873,n874,n876);
xor (n874,n875,n54);
xor (n875,n733,n737);
xor (n876,n877,n755);
xor (n877,n746,n750);
and (n878,n873,n879);
xor (n879,n880,n768);
xor (n880,n763,n765);
and (n881,n835,n879);
xor (n882,n883,n771);
xor (n883,n715,n761);
and (n884,n882,n885);
xor (n885,n774,n776);
and (n886,n833,n885);
and (n887,n888,n889);
xor (n888,n829,n831);
or (n889,n890,n944);
and (n890,n891,n893);
xor (n891,n892,n885);
xor (n892,n833,n882);
or (n893,n894,n940,n943);
and (n894,n895,n938);
or (n895,n896,n935,n937);
and (n896,n897,n933);
or (n897,n898,n927,n932);
and (n898,n899,n911);
or (n899,n900,n909,n910);
and (n900,n901,n905);
xnor (n901,n902,n255);
nor (n902,n903,n904);
and (n903,n13,n588);
and (n904,n22,n590);
xnor (n905,n906,n251);
nor (n906,n907,n908);
and (n907,n29,n401);
and (n908,n37,n404);
and (n909,n905,n38);
and (n910,n901,n38);
or (n911,n912,n921,n926);
and (n912,n913,n917);
xnor (n913,n914,n61);
nor (n914,n915,n916);
and (n915,n45,n259);
and (n916,n53,n262);
xnor (n917,n918,n77);
nor (n918,n919,n920);
and (n919,n183,n71);
and (n920,n178,n76);
and (n921,n917,n922);
xnor (n922,n923,n92);
nor (n923,n924,n925);
and (n924,n360,n85);
and (n925,n292,n89);
and (n926,n913,n922);
and (n927,n911,n928);
xnor (n928,n929,n38);
nor (n929,n930,n931);
and (n930,n676,n30);
and (n931,n519,n35);
and (n932,n899,n928);
xor (n933,n934,n870);
xor (n934,n837,n853);
and (n935,n933,n936);
xor (n936,n874,n876);
and (n937,n897,n936);
xor (n938,n939,n744);
xor (n939,n717,n731);
and (n940,n938,n941);
xor (n941,n942,n879);
xor (n942,n835,n873);
and (n943,n895,n941);
and (n944,n945,n946);
xor (n945,n891,n893);
or (n946,n947,n1017);
and (n947,n948,n950);
xor (n948,n949,n941);
xor (n949,n895,n938);
or (n950,n951,n1013,n1016);
and (n951,n952,n1008);
or (n952,n953,n1004,n1007);
and (n953,n954,n994);
or (n954,n955,n988,n993);
and (n955,n956,n972);
or (n956,n957,n966,n971);
and (n957,n958,n962);
xnor (n958,n959,n77);
nor (n959,n960,n961);
and (n960,n292,n71);
and (n961,n183,n76);
xnor (n962,n963,n92);
nor (n963,n964,n965);
and (n964,n423,n85);
and (n965,n360,n89);
and (n966,n962,n967);
xnor (n967,n968,n23);
nor (n968,n969,n970);
and (n969,n676,n14);
and (n970,n519,n19);
and (n971,n958,n967);
or (n972,n973,n982,n987);
and (n973,n974,n978);
xnor (n974,n975,n255);
nor (n975,n976,n977);
and (n976,n37,n588);
and (n977,n13,n590);
xnor (n978,n979,n251);
nor (n979,n980,n981);
and (n980,n53,n401);
and (n981,n29,n404);
and (n982,n978,n983);
xnor (n983,n984,n61);
nor (n984,n985,n986);
and (n985,n178,n259);
and (n986,n45,n262);
and (n987,n974,n983);
and (n988,n972,n989);
xnor (n989,n990,n23);
nor (n990,n991,n992);
and (n991,n519,n14);
and (n992,n423,n19);
and (n993,n956,n989);
or (n994,n995,n1000,n1003);
and (n995,n996,n998);
xnor (n996,n997,n38);
nand (n997,n676,n35);
xor (n998,n999,n38);
xor (n999,n901,n905);
and (n1000,n998,n1001);
xor (n1001,n1002,n922);
xor (n1002,n913,n917);
and (n1003,n996,n1001);
and (n1004,n994,n1005);
xor (n1005,n1006,n864);
xor (n1006,n855,n859);
and (n1007,n954,n1005);
and (n1008,n1009,n1011);
xor (n1009,n1010,n848);
xor (n1010,n839,n843);
xor (n1011,n1012,n928);
xor (n1012,n899,n911);
and (n1013,n1008,n1014);
xor (n1014,n1015,n936);
xor (n1015,n897,n933);
and (n1016,n952,n1014);
and (n1017,n1018,n1019);
xor (n1018,n948,n950);
or (n1019,n1020,n1072);
and (n1020,n1021,n1023);
xor (n1021,n1022,n1014);
xor (n1022,n952,n1008);
or (n1023,n1024,n1069,n1071);
and (n1024,n1025,n1067);
or (n1025,n1026,n1063,n1066);
and (n1026,n1027,n1061);
or (n1027,n1028,n1057,n1060);
and (n1028,n1029,n1045);
or (n1029,n1030,n1039,n1044);
and (n1030,n1031,n1035);
xnor (n1031,n1032,n61);
nor (n1032,n1033,n1034);
and (n1033,n183,n259);
and (n1034,n178,n262);
xnor (n1035,n1036,n77);
nor (n1036,n1037,n1038);
and (n1037,n360,n71);
and (n1038,n292,n76);
and (n1039,n1035,n1040);
xnor (n1040,n1041,n92);
nor (n1041,n1042,n1043);
and (n1042,n519,n85);
and (n1043,n423,n89);
and (n1044,n1031,n1040);
or (n1045,n1046,n1055,n1056);
and (n1046,n1047,n1051);
xnor (n1047,n1048,n255);
nor (n1048,n1049,n1050);
and (n1049,n29,n588);
and (n1050,n37,n590);
xnor (n1051,n1052,n251);
nor (n1052,n1053,n1054);
and (n1053,n45,n401);
and (n1054,n53,n404);
and (n1055,n1051,n23);
and (n1056,n1047,n23);
and (n1057,n1045,n1058);
xor (n1058,n1059,n967);
xor (n1059,n958,n962);
and (n1060,n1029,n1058);
xor (n1061,n1062,n989);
xor (n1062,n956,n972);
and (n1063,n1061,n1064);
xor (n1064,n1065,n1001);
xor (n1065,n996,n998);
and (n1066,n1027,n1064);
xor (n1067,n1068,n1005);
xor (n1068,n954,n994);
and (n1069,n1067,n1070);
xor (n1070,n1009,n1011);
and (n1071,n1025,n1070);
and (n1072,n1073,n1074);
xor (n1073,n1021,n1023);
or (n1074,n1075,n1113);
and (n1075,n1076,n1078);
xor (n1076,n1077,n1070);
xor (n1077,n1025,n1067);
and (n1078,n1079,n1111);
or (n1079,n1080,n1107,n1110);
and (n1080,n1081,n1105);
or (n1081,n1082,n1101,n1104);
and (n1082,n1083,n1099);
or (n1083,n1084,n1093,n1098);
and (n1084,n1085,n1089);
xnor (n1085,n1086,n255);
nor (n1086,n1087,n1088);
and (n1087,n53,n588);
and (n1088,n29,n590);
xnor (n1089,n1090,n251);
nor (n1090,n1091,n1092);
and (n1091,n178,n401);
and (n1092,n45,n404);
and (n1093,n1089,n1094);
xnor (n1094,n1095,n61);
nor (n1095,n1096,n1097);
and (n1096,n292,n259);
and (n1097,n183,n262);
and (n1098,n1085,n1094);
xnor (n1099,n1100,n23);
nand (n1100,n676,n19);
and (n1101,n1099,n1102);
xor (n1102,n1103,n1040);
xor (n1103,n1031,n1035);
and (n1104,n1083,n1102);
xor (n1105,n1106,n983);
xor (n1106,n974,n978);
and (n1107,n1105,n1108);
xor (n1108,n1109,n1058);
xor (n1109,n1029,n1045);
and (n1110,n1081,n1108);
xor (n1111,n1112,n1064);
xor (n1112,n1027,n1061);
and (n1113,n1114,n1115);
xor (n1114,n1076,n1078);
or (n1115,n1116,n1168);
and (n1116,n1117,n1118);
xor (n1117,n1079,n1111);
and (n1118,n1119,n1166);
or (n1119,n1120,n1162,n1165);
and (n1120,n1121,n1155);
or (n1121,n1122,n1149,n1154);
and (n1122,n1123,n1137);
or (n1123,n1124,n1133,n1136);
and (n1124,n1125,n1129);
xnor (n1125,n1126,n61);
nor (n1126,n1127,n1128);
and (n1127,n360,n259);
and (n1128,n292,n262);
xnor (n1129,n1130,n77);
nor (n1130,n1131,n1132);
and (n1131,n519,n71);
and (n1132,n423,n76);
and (n1133,n1129,n1134);
xnor (n1134,n1135,n92);
nand (n1135,n676,n89);
and (n1136,n1125,n1134);
or (n1137,n1138,n1147,n1148);
and (n1138,n1139,n1143);
xnor (n1139,n1140,n255);
nor (n1140,n1141,n1142);
and (n1141,n45,n588);
and (n1142,n53,n590);
xnor (n1143,n1144,n251);
nor (n1144,n1145,n1146);
and (n1145,n183,n401);
and (n1146,n178,n404);
and (n1147,n1143,n92);
and (n1148,n1139,n92);
and (n1149,n1137,n1150);
xnor (n1150,n1151,n77);
nor (n1151,n1152,n1153);
and (n1152,n423,n71);
and (n1153,n360,n76);
and (n1154,n1123,n1150);
and (n1155,n1156,n1160);
xnor (n1156,n1157,n92);
nor (n1157,n1158,n1159);
and (n1158,n676,n85);
and (n1159,n519,n89);
xor (n1160,n1161,n1094);
xor (n1161,n1085,n1089);
and (n1162,n1155,n1163);
xor (n1163,n1164,n23);
xor (n1164,n1047,n1051);
and (n1165,n1121,n1163);
xor (n1166,n1167,n1108);
xor (n1167,n1081,n1105);
and (n1168,n1169,n1170);
xor (n1169,n1117,n1118);
or (n1170,n1171,n1178);
and (n1171,n1172,n1173);
xor (n1172,n1119,n1166);
and (n1173,n1174,n1176);
xor (n1174,n1175,n1102);
xor (n1175,n1083,n1099);
xor (n1176,n1177,n1163);
xor (n1177,n1121,n1155);
and (n1178,n1179,n1180);
xor (n1179,n1172,n1173);
or (n1180,n1181,n1214);
and (n1181,n1182,n1183);
xor (n1182,n1174,n1176);
or (n1183,n1184,n1211,n1213);
and (n1184,n1185,n1209);
or (n1185,n1186,n1205,n1208);
and (n1186,n1187,n1203);
or (n1187,n1188,n1197,n1202);
and (n1188,n1189,n1193);
xnor (n1189,n1190,n255);
nor (n1190,n1191,n1192);
and (n1191,n178,n588);
and (n1192,n45,n590);
xnor (n1193,n1194,n251);
nor (n1194,n1195,n1196);
and (n1195,n292,n401);
and (n1196,n183,n404);
and (n1197,n1193,n1198);
xnor (n1198,n1199,n61);
nor (n1199,n1200,n1201);
and (n1200,n423,n259);
and (n1201,n360,n262);
and (n1202,n1189,n1198);
xor (n1203,n1204,n1134);
xor (n1204,n1125,n1129);
and (n1205,n1203,n1206);
xor (n1206,n1207,n92);
xor (n1207,n1139,n1143);
and (n1208,n1187,n1206);
xor (n1209,n1210,n1150);
xor (n1210,n1123,n1137);
and (n1211,n1209,n1212);
xor (n1212,n1156,n1160);
and (n1213,n1185,n1212);
and (n1214,n1215,n1216);
xor (n1215,n1182,n1183);
or (n1216,n1217,n1250);
and (n1217,n1218,n1220);
xor (n1218,n1219,n1212);
xor (n1219,n1185,n1209);
and (n1220,n1221,n1248);
or (n1221,n1222,n1242,n1247);
and (n1222,n1223,n1235);
or (n1223,n1224,n1233,n1234);
and (n1224,n1225,n1229);
xnor (n1225,n1226,n255);
nor (n1226,n1227,n1228);
and (n1227,n183,n588);
and (n1228,n178,n590);
xnor (n1229,n1230,n251);
nor (n1230,n1231,n1232);
and (n1231,n360,n401);
and (n1232,n292,n404);
and (n1233,n1229,n77);
and (n1234,n1225,n77);
and (n1235,n1236,n1240);
xnor (n1236,n1237,n61);
nor (n1237,n1238,n1239);
and (n1238,n519,n259);
and (n1239,n423,n262);
xnor (n1240,n1241,n77);
nand (n1241,n676,n76);
and (n1242,n1235,n1243);
xnor (n1243,n1244,n77);
nor (n1244,n1245,n1246);
and (n1245,n676,n71);
and (n1246,n519,n76);
and (n1247,n1223,n1243);
xor (n1248,n1249,n1206);
xor (n1249,n1187,n1203);
and (n1250,n1251,n1252);
xor (n1251,n1218,n1220);
or (n1252,n1253,n1260);
and (n1253,n1254,n1255);
xor (n1254,n1221,n1248);
and (n1255,n1256,n1258);
xor (n1256,n1257,n1198);
xor (n1257,n1189,n1193);
xor (n1258,n1259,n1243);
xor (n1259,n1223,n1235);
and (n1260,n1261,n1262);
xor (n1261,n1254,n1255);
or (n1262,n1263,n1288);
and (n1263,n1264,n1265);
xor (n1264,n1256,n1258);
or (n1265,n1266,n1285,n1287);
and (n1266,n1267,n1283);
or (n1267,n1268,n1277,n1282);
and (n1268,n1269,n1273);
xnor (n1269,n1270,n255);
nor (n1270,n1271,n1272);
and (n1271,n292,n588);
and (n1272,n183,n590);
xnor (n1273,n1274,n251);
nor (n1274,n1275,n1276);
and (n1275,n423,n401);
and (n1276,n360,n404);
and (n1277,n1273,n1278);
xnor (n1278,n1279,n61);
nor (n1279,n1280,n1281);
and (n1280,n676,n259);
and (n1281,n519,n262);
and (n1282,n1269,n1278);
xor (n1283,n1284,n77);
xor (n1284,n1225,n1229);
and (n1285,n1283,n1286);
xor (n1286,n1236,n1240);
and (n1287,n1267,n1286);
and (n1288,n1289,n1290);
xor (n1289,n1264,n1265);
or (n1290,n1291,n1309);
and (n1291,n1292,n1294);
xor (n1292,n1293,n1286);
xor (n1293,n1267,n1283);
and (n1294,n1295,n1307);
or (n1295,n1296,n1305,n1306);
and (n1296,n1297,n1301);
xnor (n1297,n1298,n255);
nor (n1298,n1299,n1300);
and (n1299,n360,n588);
and (n1300,n292,n590);
xnor (n1301,n1302,n251);
nor (n1302,n1303,n1304);
and (n1303,n519,n401);
and (n1304,n423,n404);
and (n1305,n1301,n61);
and (n1306,n1297,n61);
xor (n1307,n1308,n1278);
xor (n1308,n1269,n1273);
and (n1309,n1310,n1311);
xor (n1310,n1292,n1294);
or (n1311,n1312,n1319);
and (n1312,n1313,n1314);
xor (n1313,n1295,n1307);
and (n1314,n1315,n1317);
xnor (n1315,n1316,n61);
nand (n1316,n676,n262);
xor (n1317,n1318,n61);
xor (n1318,n1297,n1301);
and (n1319,n1320,n1321);
xor (n1320,n1313,n1314);
or (n1321,n1322,n1333);
and (n1322,n1323,n1324);
xor (n1323,n1315,n1317);
and (n1324,n1325,n1329);
xnor (n1325,n1326,n255);
nor (n1326,n1327,n1328);
and (n1327,n423,n588);
and (n1328,n360,n590);
xnor (n1329,n1330,n251);
nor (n1330,n1331,n1332);
and (n1331,n676,n401);
and (n1332,n519,n404);
and (n1333,n1334,n1335);
xor (n1334,n1323,n1324);
or (n1335,n1336,n1343);
and (n1336,n1337,n1338);
xor (n1337,n1325,n1329);
and (n1338,n1339,n251);
xnor (n1339,n1340,n255);
nor (n1340,n1341,n1342);
and (n1341,n519,n588);
and (n1342,n423,n590);
and (n1343,n1344,n1345);
xor (n1344,n1337,n1338);
or (n1345,n1346,n1350);
and (n1346,n1347,n1349);
xnor (n1347,n1348,n251);
nand (n1348,n676,n404);
xor (n1349,n1339,n251);
and (n1350,n1351,n1352);
xor (n1351,n1347,n1349);
and (n1352,n1353,n1357);
xnor (n1353,n1354,n255);
nor (n1354,n1355,n1356);
and (n1355,n676,n588);
and (n1356,n519,n590);
and (n1357,n1358,n255);
xnor (n1358,n1359,n255);
nand (n1359,n676,n590);
buf (n1360,n1361);
xor (n1361,n1362,n1446);
xor (n1362,n1363,n1399);
xor (n1363,n1364,n1386);
or (n1364,n1365,n1378,n1385);
and (n1365,n1366,n1376);
or (n1366,n1367,n1374,n1375);
and (n1367,n1368,n1371);
or (n1368,n41,n1369,n1370);
and (n1369,n42,n187);
and (n1370,n26,n187);
or (n1371,n80,n1372,n1373);
and (n1372,n81,n10);
and (n1373,n67,n10);
and (n1374,n1371,n195);
and (n1375,n1368,n195);
xor (n1376,n1377,n136);
xor (n1377,n99,n102);
and (n1378,n1376,n1379);
xor (n1379,n1380,n1384);
xor (n1380,n109,n1381);
or (n1381,n1382,n128,n1383);
and (n1382,n98,n124);
and (n1383,n98,n129);
xnor (n1384,n140,n144);
and (n1385,n1366,n1379);
xor (n1386,n1387,n1398);
xor (n1387,n1388,n1392);
or (n1388,n1389,n1390,n1391);
and (n1389,n109,n1381);
and (n1390,n1381,n1384);
and (n1391,n109,n1384);
xor (n1392,n1393,n236);
xor (n1393,n1394,n1397);
or (n1394,n233,n1395,n1396);
and (n1395,n102,n136);
and (n1396,n99,n136);
or (n1397,n140,n144);
xor (n1398,n240,n214);
or (n1399,n1400,n1442,n1445);
and (n1400,n1401,n1411);
or (n1401,n1402,n1407,n1410);
and (n1402,n1403,n200);
or (n1403,n1404,n164);
or (n1404,n1405,n158,n1406);
and (n1405,n60,n154);
and (n1406,n60,n159);
and (n1407,n200,n1408);
xor (n1408,n1409,n195);
xor (n1409,n1368,n1371);
and (n1410,n1403,n1408);
or (n1411,n1412,n1438,n1441);
and (n1412,n1413,n1434);
or (n1413,n1414,n1430,n1433);
and (n1414,n1415,n1426);
or (n1415,n1416,n1423,n1425);
and (n1416,n1417,n1420);
or (n1417,n263,n1418,n1419);
and (n1418,n264,n271);
and (n1419,n256,n271);
or (n1420,n279,n1421,n1422);
and (n1421,n280,n287);
and (n1422,n275,n287);
and (n1423,n1420,n1424);
buf (n1424,n291);
and (n1425,n1417,n1424);
or (n1426,n1427,n1428,n1429);
and (n1427,n182,n297);
and (n1428,n297,n299);
and (n1429,n182,n299);
and (n1430,n1426,n1431);
xor (n1431,n1432,n187);
xor (n1432,n26,n42);
and (n1433,n1415,n1431);
and (n1434,n1435,n1437);
xor (n1435,n1436,n10);
xor (n1436,n67,n81);
xnor (n1437,n1404,n164);
and (n1438,n1434,n1439);
xor (n1439,n1440,n1408);
xor (n1440,n1403,n200);
and (n1441,n1413,n1439);
and (n1442,n1411,n1443);
xor (n1443,n1444,n1379);
xor (n1444,n1366,n1376);
and (n1445,n1401,n1443);
or (n1446,n1447,n1481);
and (n1447,n1448,n1450);
xor (n1448,n1449,n1443);
xor (n1449,n1401,n1411);
and (n1450,n1451,n1479);
or (n1451,n1452,n1476,n1478);
and (n1452,n1453,n1474);
or (n1453,n1454,n1472,n1473);
and (n1454,n1455,n1463);
or (n1455,n1456,n1460,n1462);
and (n1456,n1457,n337);
or (n1457,n1458,n331,n1459);
and (n1458,n250,n327);
and (n1459,n250,n332);
and (n1460,n337,n1461);
and (n1461,n355,n359);
and (n1462,n1457,n1461);
or (n1463,n1464,n1469,n1471);
and (n1464,n1465,n1467);
xor (n1465,n1466,n271);
xor (n1466,n256,n264);
xor (n1467,n1468,n287);
xor (n1468,n275,n280);
and (n1469,n1467,n1470);
not (n1470,n291);
and (n1471,n1465,n1470);
and (n1472,n1463,n372);
and (n1473,n1455,n372);
xor (n1474,n1475,n1431);
xor (n1475,n1415,n1426);
and (n1476,n1474,n1477);
xor (n1477,n1435,n1437);
and (n1478,n1453,n1477);
xor (n1479,n1480,n1439);
xor (n1480,n1413,n1434);
and (n1481,n1482,n1483);
xor (n1482,n1448,n1450);
or (n1483,n1484,n1518);
and (n1484,n1485,n1486);
xor (n1485,n1451,n1479);
and (n1486,n1487,n1516);
or (n1487,n1488,n1512,n1515);
and (n1488,n1489,n1510);
or (n1489,n1490,n1506,n1509);
and (n1490,n1491,n1502);
or (n1491,n1492,n1499,n1501);
and (n1492,n1493,n1496);
or (n1493,n405,n1494,n1495);
and (n1494,n406,n428);
and (n1495,n398,n428);
or (n1496,n436,n1497,n1498);
and (n1497,n437,n413);
and (n1498,n432,n413);
and (n1499,n1496,n1500);
or (n1500,n417,n422);
and (n1501,n1493,n1500);
or (n1502,n1503,n1504,n1505);
and (n1503,n446,n448);
and (n1504,n448,n452);
and (n1505,n446,n452);
and (n1506,n1502,n1507);
xor (n1507,n1508,n1470);
xor (n1508,n1465,n1467);
and (n1509,n1491,n1507);
xor (n1510,n1511,n1424);
xor (n1511,n1417,n1420);
and (n1512,n1510,n1513);
xor (n1513,n1514,n372);
xor (n1514,n1455,n1463);
and (n1515,n1489,n1513);
xor (n1516,n1517,n1477);
xor (n1517,n1453,n1474);
and (n1518,n1519,n1520);
xor (n1519,n1485,n1486);
or (n1520,n1521,n1545);
and (n1521,n1522,n1523);
xor (n1522,n1487,n1516);
and (n1523,n1524,n1543);
or (n1524,n1525,n1539,n1542);
and (n1525,n1526,n1537);
or (n1526,n1527,n1535,n1536);
and (n1527,n1528,n1531);
or (n1528,n1529,n1530,n521);
and (n1529,n478,n808);
and (n1530,n808,n507);
or (n1531,n1532,n1533,n1534);
and (n1532,n816,n818);
and (n1533,n818,n820);
and (n1534,n816,n820);
and (n1535,n1531,n528);
and (n1536,n1528,n528);
xor (n1537,n1538,n1461);
xor (n1538,n1457,n337);
and (n1539,n1537,n1540);
xor (n1540,n1541,n1507);
xor (n1541,n1491,n1502);
and (n1542,n1526,n1540);
xor (n1543,n1544,n1513);
xor (n1544,n1489,n1510);
and (n1545,n1546,n1547);
xor (n1546,n1522,n1523);
or (n1547,n1548,n1565);
and (n1548,n1549,n1550);
xor (n1549,n1524,n1543);
and (n1550,n1551,n1563);
or (n1551,n1552,n1559,n1562);
and (n1552,n1553,n1557);
or (n1553,n1554,n1555,n1556);
and (n1554,n549,n813);
and (n1555,n813,n814);
and (n1556,n549,n814);
xor (n1557,n1558,n1500);
xor (n1558,n1493,n1496);
and (n1559,n1557,n1560);
xor (n1560,n1561,n528);
xor (n1561,n1528,n1531);
and (n1562,n1553,n1560);
xor (n1563,n1564,n1540);
xor (n1564,n1526,n1537);
and (n1565,n1566,n1567);
xor (n1566,n1549,n1550);
or (n1567,n1568,n1577);
and (n1568,n1569,n1570);
xor (n1569,n1551,n1563);
and (n1570,n1571,n1575);
or (n1571,n1572,n1573,n1574);
and (n1572,n803,n806);
and (n1573,n806,n811);
and (n1574,n803,n811);
xor (n1575,n1576,n1560);
xor (n1576,n1553,n1557);
and (n1577,n1578,n1579);
xor (n1578,n1569,n1570);
or (n1579,n1580,n1583);
and (n1580,n1581,n1582);
xor (n1581,n1571,n1575);
and (n1582,n797,n801);
and (n1583,n1584,n1585);
xor (n1584,n1581,n1582);
or (n1585,n1586,n794);
and (n1586,n796,n821);
endmodule
