module top (out,n16,n18,n19,n21,n24,n25,n31,n33,n34
        ,n36,n39,n43,n45,n46,n48,n51,n56,n58,n60
        ,n72,n81,n83,n85,n88,n100,n107,n109,n111,n114
        ,n122,n123,n135,n147,n185,n189,n191,n193,n221,n222
        ,n329,n346,n347,n727,n731,n733,n744,n756,n770);
output out;
input n16;
input n18;
input n19;
input n21;
input n24;
input n25;
input n31;
input n33;
input n34;
input n36;
input n39;
input n43;
input n45;
input n46;
input n48;
input n51;
input n56;
input n58;
input n60;
input n72;
input n81;
input n83;
input n85;
input n88;
input n100;
input n107;
input n109;
input n111;
input n114;
input n122;
input n123;
input n135;
input n147;
input n185;
input n189;
input n191;
input n193;
input n221;
input n222;
input n329;
input n346;
input n347;
input n727;
input n731;
input n733;
input n744;
input n756;
input n770;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n17;
wire n20;
wire n22;
wire n23;
wire n26;
wire n27;
wire n28;
wire n29;
wire n30;
wire n32;
wire n35;
wire n37;
wire n38;
wire n40;
wire n41;
wire n42;
wire n44;
wire n47;
wire n49;
wire n50;
wire n52;
wire n53;
wire n54;
wire n55;
wire n57;
wire n59;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n82;
wire n84;
wire n86;
wire n87;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n108;
wire n110;
wire n112;
wire n113;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n186;
wire n187;
wire n188;
wire n190;
wire n192;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n728;
wire n729;
wire n730;
wire n732;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2988;
wire n2989;
wire n2990;
wire n2991;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2996;
wire n2997;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3003;
wire n3004;
wire n3005;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3010;
wire n3011;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3038;
wire n3039;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
wire n3056;
wire n3057;
wire n3058;
wire n3059;
wire n3060;
wire n3061;
wire n3062;
wire n3063;
wire n3064;
wire n3065;
wire n3066;
wire n3067;
wire n3068;
wire n3069;
wire n3070;
wire n3071;
wire n3072;
wire n3073;
wire n3074;
wire n3075;
wire n3076;
wire n3077;
wire n3078;
wire n3079;
wire n3080;
wire n3081;
wire n3082;
wire n3083;
wire n3084;
wire n3085;
wire n3086;
wire n3087;
wire n3088;
wire n3089;
wire n3090;
wire n3091;
wire n3092;
wire n3093;
wire n3094;
wire n3095;
wire n3096;
wire n3097;
wire n3098;
wire n3099;
wire n3100;
wire n3101;
wire n3102;
wire n3103;
wire n3104;
wire n3105;
wire n3106;
wire n3107;
wire n3108;
wire n3109;
wire n3110;
wire n3111;
wire n3112;
wire n3113;
wire n3114;
wire n3115;
wire n3116;
wire n3117;
wire n3118;
wire n3119;
wire n3120;
wire n3121;
wire n3122;
wire n3123;
wire n3124;
wire n3125;
wire n3126;
wire n3127;
wire n3128;
wire n3129;
wire n3130;
wire n3131;
wire n3132;
wire n3133;
wire n3134;
wire n3135;
wire n3136;
wire n3137;
wire n3138;
wire n3139;
wire n3140;
wire n3141;
wire n3142;
wire n3143;
wire n3144;
wire n3145;
wire n3146;
wire n3147;
wire n3148;
wire n3149;
wire n3150;
wire n3151;
wire n3152;
wire n3153;
wire n3154;
wire n3155;
wire n3156;
wire n3157;
wire n3158;
wire n3159;
wire n3160;
wire n3161;
wire n3162;
wire n3163;
wire n3164;
wire n3165;
wire n3166;
wire n3167;
wire n3168;
wire n3169;
wire n3170;
wire n3171;
wire n3172;
wire n3173;
wire n3174;
wire n3175;
wire n3176;
wire n3177;
wire n3178;
wire n3179;
wire n3180;
wire n3181;
wire n3182;
wire n3183;
wire n3184;
wire n3185;
wire n3186;
wire n3187;
wire n3188;
wire n3189;
wire n3190;
wire n3191;
wire n3192;
wire n3193;
wire n3194;
wire n3195;
wire n3196;
wire n3197;
wire n3198;
wire n3199;
wire n3200;
wire n3201;
wire n3202;
wire n3203;
wire n3204;
wire n3205;
wire n3206;
wire n3207;
wire n3208;
wire n3209;
wire n3210;
wire n3211;
wire n3212;
wire n3213;
wire n3214;
wire n3215;
wire n3216;
wire n3217;
wire n3218;
wire n3219;
wire n3220;
wire n3221;
wire n3222;
wire n3223;
wire n3224;
wire n3225;
wire n3226;
wire n3227;
wire n3228;
wire n3229;
wire n3230;
wire n3231;
wire n3232;
wire n3233;
wire n3234;
wire n3235;
wire n3236;
wire n3237;
wire n3238;
wire n3239;
wire n3240;
wire n3241;
wire n3242;
wire n3243;
wire n3244;
wire n3245;
wire n3246;
wire n3247;
wire n3248;
wire n3249;
wire n3250;
wire n3251;
wire n3252;
wire n3253;
wire n3254;
wire n3255;
wire n3256;
wire n3257;
wire n3258;
wire n3259;
wire n3260;
wire n3261;
wire n3262;
wire n3263;
wire n3264;
wire n3265;
wire n3266;
wire n3267;
wire n3268;
wire n3269;
wire n3270;
wire n3271;
xor (out,n0,n2738);
xnor (n0,n1,n2670);
nand (n1,n2,n708);
nor (n2,n3,n702);
nor (n3,n4,n559);
nor (n4,n5,n557);
nor (n5,n6,n480);
nand (n6,n7,n400);
nand (n7,n8,n316,n399);
nand (n8,n9,n175);
xor (n9,n10,n139);
xor (n10,n11,n64);
xor (n11,n12,n26);
xor (n12,n13,n25);
xor (n13,n14,n24);
or (n14,n15,n20);
and (n15,n16,n17);
xor (n17,n18,n19);
and (n20,n21,n22);
nor (n22,n17,n23);
xnor (n23,n24,n18);
nand (n26,n27,n52,n63);
nand (n27,n28,n40);
xor (n28,n29,n39);
or (n29,n30,n35);
and (n30,n31,n32);
xor (n32,n33,n34);
and (n35,n36,n37);
nor (n37,n32,n38);
xnor (n38,n39,n33);
xor (n40,n41,n51);
or (n41,n42,n47);
and (n42,n43,n44);
xor (n44,n45,n46);
and (n47,n48,n49);
nor (n49,n44,n50);
xnor (n50,n51,n45);
nand (n52,n53,n40);
xor (n53,n54,n34);
or (n54,n55,n59);
and (n55,n56,n57);
xor (n57,n58,n51);
and (n59,n60,n61);
nor (n61,n57,n62);
xnor (n62,n34,n58);
nand (n63,n28,n53);
nand (n64,n65,n115,n138);
nand (n65,n66,n90);
nand (n66,n67,n77,n89);
nand (n67,n68,n73);
xor (n68,n69,n39);
or (n69,n70,n71);
and (n70,n36,n32);
and (n71,n72,n37);
xor (n73,n74,n51);
or (n74,n75,n76);
and (n75,n48,n44);
and (n76,n56,n49);
nand (n77,n78,n73);
xor (n78,n79,n88);
or (n79,n80,n84);
and (n80,n81,n82);
xor (n82,n83,n39);
and (n84,n85,n86);
nor (n86,n82,n87);
xnor (n87,n88,n83);
nand (n89,n68,n78);
xor (n90,n91,n104);
xor (n91,n92,n96);
xor (n92,n93,n88);
or (n93,n94,n95);
and (n94,n72,n82);
and (n95,n81,n86);
xor (n96,n97,n19);
or (n97,n98,n101);
and (n98,n85,n99);
xor (n99,n100,n88);
and (n101,n16,n102);
nor (n102,n99,n103);
xnor (n103,n19,n100);
xor (n104,n105,n114);
or (n105,n106,n110);
and (n106,n107,n108);
xor (n108,n109,n24);
and (n110,n111,n112);
nor (n112,n108,n113);
xnor (n113,n114,n109);
nand (n115,n116,n90);
nand (n116,n117,n131,n137);
nand (n117,n118,n127);
xor (n118,n119,n46);
or (n119,n120,n124);
and (n120,n43,n121);
xor (n121,n122,n123);
and (n124,n48,n125);
nor (n125,n121,n126);
xnor (n126,n46,n122);
xor (n127,n128,n19);
or (n128,n129,n130);
and (n129,n16,n99);
and (n130,n21,n102);
nand (n131,n132,n127);
xor (n132,n133,n24);
or (n133,n134,n136);
and (n134,n135,n17);
and (n136,n107,n22);
nand (n137,n118,n132);
nand (n138,n66,n116);
xor (n139,n140,n171);
xor (n140,n141,n157);
xor (n141,n142,n153);
xor (n142,n143,n149);
not (n143,n144);
xor (n144,n145,n46);
or (n145,n146,n148);
and (n146,n147,n121);
and (n148,n147,n125);
xor (n149,n150,n51);
or (n150,n151,n152);
and (n151,n147,n44);
and (n152,n43,n49);
xor (n153,n154,n39);
or (n154,n155,n156);
and (n155,n60,n32);
and (n156,n31,n37);
xor (n157,n158,n167);
xor (n158,n159,n163);
xor (n159,n160,n34);
or (n160,n161,n162);
and (n161,n48,n57);
and (n162,n56,n61);
xor (n163,n164,n88);
or (n164,n165,n166);
and (n165,n36,n82);
and (n166,n72,n86);
xor (n167,n168,n19);
or (n168,n169,n170);
and (n169,n81,n99);
and (n170,n85,n102);
nand (n171,n172,n173,n174);
nand (n172,n92,n96);
nand (n173,n104,n96);
nand (n174,n92,n104);
xor (n175,n176,n255);
xor (n176,n177,n235);
nand (n177,n178,n208,n234);
nand (n178,n179,n198);
nand (n179,n180,n196,n197);
nand (n180,n181,n186);
xor (n181,n182,n114);
or (n182,n183,n184);
and (n183,n111,n108);
and (n184,n185,n112);
xor (n186,n187,n25);
or (n187,n188,n192);
and (n188,n189,n190);
xor (n190,n191,n114);
and (n192,n193,n194);
nor (n194,n190,n195);
xnor (n195,n25,n191);
nand (n196,n25,n186);
nand (n197,n181,n25);
xor (n198,n199,n204);
xor (n199,n200,n143);
xor (n200,n201,n25);
or (n201,n202,n203);
and (n202,n185,n190);
and (n203,n189,n194);
xor (n204,n205,n24);
or (n205,n206,n207);
and (n206,n21,n17);
and (n207,n135,n22);
nand (n208,n209,n198);
xor (n209,n210,n232);
xor (n210,n25,n211);
nand (n211,n212,n226,n231);
nand (n212,n213,n216);
xor (n213,n214,n46);
or (n214,n146,n215);
and (n215,n43,n125);
not (n216,n217);
xor (n217,n218,n123);
or (n218,n219,n223);
and (n219,n147,n220);
xor (n220,n221,n222);
and (n223,n147,n224);
nor (n224,n220,n225);
xnor (n225,n123,n221);
nand (n226,n227,n216);
xor (n227,n228,n34);
or (n228,n229,n230);
and (n229,n60,n57);
and (n230,n31,n61);
nand (n231,n213,n227);
xor (n232,n233,n53);
xor (n233,n28,n40);
nand (n234,n179,n209);
xor (n235,n236,n251);
xor (n236,n237,n241);
nand (n237,n238,n239,n240);
nand (n238,n200,n143);
nand (n239,n204,n143);
nand (n240,n200,n204);
xor (n241,n242,n144);
xor (n242,n243,n247);
xor (n243,n244,n114);
or (n244,n245,n246);
and (n245,n135,n108);
and (n246,n107,n112);
xor (n247,n248,n25);
or (n248,n249,n250);
and (n249,n111,n190);
and (n250,n185,n194);
nand (n251,n252,n253,n254);
nand (n252,n25,n211);
nand (n253,n232,n211);
nand (n254,n25,n232);
nand (n255,n256,n312,n315);
nand (n256,n257,n277);
nand (n257,n258,n273,n276);
nand (n258,n259,n271);
nand (n259,n260,n265,n270);
nand (n260,n217,n261);
xor (n261,n262,n34);
or (n262,n263,n264);
and (n263,n31,n57);
and (n264,n36,n61);
nand (n265,n266,n261);
xor (n266,n267,n39);
or (n267,n268,n269);
and (n268,n72,n32);
and (n269,n81,n37);
nand (n270,n217,n266);
xor (n271,n272,n78);
xor (n272,n68,n73);
nand (n273,n274,n271);
xor (n274,n275,n227);
xor (n275,n213,n216);
nand (n276,n259,n274);
nand (n277,n278,n308,n311);
nand (n278,n279,n292);
nand (n279,n280,n286,n291);
nand (n280,n281,n285);
xor (n281,n282,n51);
or (n282,n283,n284);
and (n283,n56,n44);
and (n284,n60,n49);
not (n285,n118);
nand (n286,n287,n285);
xor (n287,n288,n88);
or (n288,n289,n290);
and (n289,n85,n82);
and (n290,n16,n86);
nand (n291,n281,n287);
nand (n292,n293,n302,n307);
nand (n293,n294,n298);
xor (n294,n295,n19);
or (n295,n296,n297);
and (n296,n21,n99);
and (n297,n135,n102);
xor (n298,n299,n24);
or (n299,n300,n301);
and (n300,n107,n17);
and (n301,n111,n22);
nand (n302,n303,n298);
xor (n303,n304,n114);
or (n304,n305,n306);
and (n305,n185,n108);
and (n306,n189,n112);
nand (n307,n294,n303);
nand (n308,n309,n292);
xor (n309,n310,n132);
xor (n310,n118,n127);
nand (n311,n279,n309);
nand (n312,n313,n277);
xor (n313,n314,n116);
xor (n314,n66,n90);
nand (n315,n257,n313);
nand (n316,n317,n175);
nand (n317,n318,n395,n398);
nand (n318,n319,n321);
xor (n319,n320,n209);
xor (n320,n179,n198);
nand (n321,n322,n355,n394);
nand (n322,n323,n353);
nand (n323,n324,n330,n352);
nand (n324,n325,n25);
xor (n325,n326,n25);
or (n326,n327,n328);
and (n327,n193,n190);
and (n328,n329,n194);
nand (n330,n331,n25);
nand (n331,n332,n340,n351);
nand (n332,n333,n336);
xor (n333,n334,n123);
or (n334,n219,n335);
and (n335,n43,n224);
xor (n336,n337,n46);
or (n337,n338,n339);
and (n338,n48,n121);
and (n339,n56,n125);
nand (n340,n341,n336);
not (n341,n342);
xor (n342,n343,n222);
or (n343,n344,n348);
and (n344,n147,n345);
xor (n345,n346,n347);
and (n348,n147,n349);
nor (n349,n345,n350);
xnor (n350,n222,n346);
nand (n351,n333,n341);
nand (n352,n325,n331);
xor (n353,n354,n25);
xor (n354,n181,n186);
nand (n355,n356,n353);
nand (n356,n357,n376,n393);
nand (n357,n358,n374);
nand (n358,n359,n368,n373);
nand (n359,n360,n364);
xor (n360,n361,n51);
or (n361,n362,n363);
and (n362,n60,n44);
and (n363,n31,n49);
xor (n364,n365,n34);
or (n365,n366,n367);
and (n366,n36,n57);
and (n367,n72,n61);
nand (n368,n369,n364);
xor (n369,n370,n39);
or (n370,n371,n372);
and (n371,n81,n32);
and (n372,n85,n37);
nand (n373,n360,n369);
xor (n374,n375,n266);
xor (n375,n217,n261);
nand (n376,n377,n374);
nand (n377,n378,n387,n392);
nand (n378,n379,n383);
xor (n379,n380,n19);
or (n380,n381,n382);
and (n381,n135,n99);
and (n382,n107,n102);
xor (n383,n384,n123);
or (n384,n385,n386);
and (n385,n43,n220);
and (n386,n48,n224);
nand (n387,n388,n383);
xor (n388,n389,n88);
or (n389,n390,n391);
and (n390,n16,n82);
and (n391,n21,n86);
nand (n392,n379,n388);
nand (n393,n358,n377);
nand (n394,n323,n356);
nand (n395,n396,n321);
xor (n396,n397,n313);
xor (n397,n257,n277);
nand (n398,n319,n396);
nand (n399,n9,n317);
xor (n400,n401,n476);
xor (n401,n402,n406);
nand (n402,n403,n404,n405);
nand (n403,n11,n64);
nand (n404,n139,n64);
nand (n405,n11,n139);
xor (n406,n407,n446);
xor (n407,n408,n412);
nand (n408,n409,n410,n411);
nand (n409,n237,n241);
nand (n410,n251,n241);
nand (n411,n237,n251);
xor (n412,n413,n432);
xor (n413,n414,n418);
nand (n414,n415,n416,n417);
nand (n415,n243,n247);
nand (n416,n144,n247);
nand (n417,n243,n144);
xor (n418,n419,n428);
xor (n419,n420,n424);
xor (n420,n421,n24);
or (n421,n422,n423);
and (n422,n85,n17);
and (n423,n16,n22);
xor (n424,n425,n114);
or (n425,n426,n427);
and (n426,n21,n108);
and (n427,n135,n112);
nand (n428,n429,n430,n431);
nand (n429,n143,n149);
nand (n430,n153,n149);
nand (n431,n143,n153);
xor (n432,n433,n442);
xor (n433,n434,n438);
xor (n434,n435,n19);
or (n435,n436,n437);
and (n436,n72,n99);
and (n437,n81,n102);
xor (n438,n439,n25);
or (n439,n440,n441);
and (n440,n107,n190);
and (n441,n111,n194);
not (n442,n443);
xor (n443,n444,n51);
or (n444,n151,n445);
and (n445,n147,n49);
xor (n446,n447,n472);
xor (n447,n448,n452);
nand (n448,n449,n450,n451);
nand (n449,n13,n25);
nand (n450,n26,n25);
nand (n451,n13,n26);
xor (n452,n453,n468);
xor (n453,n25,n454);
xor (n454,n455,n464);
xor (n455,n456,n460);
xor (n456,n457,n34);
or (n457,n458,n459);
and (n458,n43,n57);
and (n459,n48,n61);
xor (n460,n461,n39);
or (n461,n462,n463);
and (n462,n56,n32);
and (n463,n60,n37);
xor (n464,n465,n88);
or (n465,n466,n467);
and (n466,n31,n82);
and (n467,n36,n86);
nand (n468,n469,n470,n471);
nand (n469,n159,n163);
nand (n470,n167,n163);
nand (n471,n159,n167);
nand (n472,n473,n474,n475);
nand (n473,n141,n157);
nand (n474,n171,n157);
nand (n475,n141,n171);
nand (n476,n477,n478,n479);
nand (n477,n177,n235);
nand (n478,n255,n235);
nand (n479,n177,n255);
nor (n480,n481,n485);
nand (n481,n482,n483,n484);
nand (n482,n402,n406);
nand (n483,n476,n406);
nand (n484,n402,n476);
xor (n485,n486,n553);
xor (n486,n487,n513);
xor (n487,n488,n497);
xor (n488,n489,n493);
nand (n489,n490,n491,n492);
nand (n490,n420,n424);
nand (n491,n428,n424);
nand (n492,n420,n428);
nand (n493,n494,n495,n496);
nand (n494,n25,n454);
nand (n495,n468,n454);
nand (n496,n25,n468);
xor (n497,n498,n509);
xor (n498,n25,n499);
xor (n499,n500,n505);
xor (n500,n442,n501);
xor (n501,n502,n34);
or (n502,n503,n504);
and (n503,n147,n57);
and (n504,n43,n61);
xor (n505,n506,n39);
or (n506,n507,n508);
and (n507,n48,n32);
and (n508,n56,n37);
nand (n509,n510,n511,n512);
nand (n510,n456,n460);
nand (n511,n464,n460);
nand (n512,n456,n464);
xor (n513,n514,n549);
xor (n514,n515,n545);
xor (n515,n516,n535);
xor (n516,n517,n521);
nand (n517,n518,n519,n520);
nand (n518,n434,n438);
nand (n519,n442,n438);
nand (n520,n434,n442);
xor (n521,n522,n531);
xor (n522,n523,n527);
xor (n523,n524,n88);
or (n524,n525,n526);
and (n525,n60,n82);
and (n526,n31,n86);
xor (n527,n528,n19);
or (n528,n529,n530);
and (n529,n36,n99);
and (n530,n72,n102);
xor (n531,n532,n25);
or (n532,n533,n534);
and (n533,n135,n190);
and (n534,n107,n194);
xor (n535,n536,n541);
xor (n536,n443,n537);
xor (n537,n538,n24);
or (n538,n539,n540);
and (n539,n81,n17);
and (n540,n85,n22);
xor (n541,n542,n114);
or (n542,n543,n544);
and (n543,n16,n108);
and (n544,n21,n112);
nand (n545,n546,n547,n548);
nand (n546,n414,n418);
nand (n547,n432,n418);
nand (n548,n414,n432);
nand (n549,n550,n551,n552);
nand (n550,n448,n452);
nand (n551,n472,n452);
nand (n552,n448,n472);
nand (n553,n554,n555,n556);
nand (n554,n408,n412);
nand (n555,n446,n412);
nand (n556,n408,n446);
not (n557,n558);
nand (n558,n481,n485);
not (n559,n560);
nor (n560,n561,n634);
nor (n561,n562,n566);
nand (n562,n563,n564,n565);
nand (n563,n487,n513);
nand (n564,n553,n513);
nand (n565,n487,n553);
xor (n566,n567,n630);
xor (n567,n568,n596);
xor (n568,n569,n592);
xor (n569,n570,n584);
xor (n570,n571,n580);
xor (n571,n572,n576);
not (n572,n573);
xor (n573,n574,n34);
or (n574,n503,n575);
and (n575,n147,n61);
xor (n576,n577,n24);
or (n577,n578,n579);
and (n578,n72,n17);
and (n579,n81,n22);
xor (n580,n581,n114);
or (n581,n582,n583);
and (n582,n85,n108);
and (n583,n16,n112);
xor (n584,n585,n588);
or (n585,n586,n587);
and (n586,n21,n190);
and (n587,n135,n194);
nand (n588,n589,n590,n591);
nand (n589,n442,n501);
nand (n590,n505,n501);
nand (n591,n442,n505);
nand (n592,n593,n594,n595);
nand (n593,n25,n499);
nand (n594,n509,n499);
nand (n595,n25,n509);
xor (n596,n597,n626);
xor (n597,n598,n622);
xor (n598,n599,n618);
xor (n599,n600,n614);
xor (n600,n601,n610);
xor (n601,n602,n606);
xor (n602,n603,n39);
or (n603,n604,n605);
and (n604,n43,n32);
and (n605,n48,n37);
xor (n606,n607,n19);
or (n607,n608,n609);
and (n608,n31,n99);
and (n609,n36,n102);
xor (n610,n611,n88);
or (n611,n612,n613);
and (n612,n56,n82);
and (n613,n60,n86);
nand (n614,n615,n616,n617);
nand (n615,n523,n527);
nand (n616,n531,n527);
nand (n617,n523,n531);
nand (n618,n619,n620,n621);
nand (n619,n443,n537);
nand (n620,n541,n537);
nand (n621,n443,n541);
nand (n622,n623,n624,n625);
nand (n623,n517,n521);
nand (n624,n535,n521);
nand (n625,n517,n535);
nand (n626,n627,n628,n629);
nand (n627,n489,n493);
nand (n628,n497,n493);
nand (n629,n489,n497);
nand (n630,n631,n632,n633);
nand (n631,n515,n545);
nand (n632,n549,n545);
nand (n633,n515,n549);
nor (n634,n635,n639);
nand (n635,n636,n637,n638);
nand (n636,n568,n596);
nand (n637,n630,n596);
nand (n638,n568,n630);
xor (n639,n640,n698);
xor (n640,n641,n645);
nand (n641,n642,n643,n644);
nand (n642,n570,n584);
nand (n643,n592,n584);
nand (n644,n570,n592);
xor (n645,n646,n671);
xor (n646,n647,n651);
nand (n647,n648,n649,n650);
nand (n648,n600,n614);
nand (n649,n618,n614);
nand (n650,n600,n618);
xor (n651,n652,n667);
xor (n652,n653,n663);
xor (n653,n654,n659);
xor (n654,n572,n655);
xor (n655,n656,n39);
or (n656,n657,n658);
and (n657,n147,n32);
and (n658,n43,n37);
xor (n659,n660,n19);
or (n660,n661,n662);
and (n661,n60,n99);
and (n662,n31,n102);
nand (n663,n664,n665,n666);
nand (n664,n602,n606);
nand (n665,n610,n606);
nand (n666,n602,n610);
nand (n667,n668,n669,n670);
nand (n668,n572,n576);
nand (n669,n580,n576);
nand (n670,n572,n580);
xor (n671,n672,n693);
xor (n672,n673,n683);
xor (n673,n674,n25);
xor (n674,n675,n679);
xor (n675,n676,n114);
or (n676,n677,n678);
and (n677,n81,n108);
and (n678,n85,n112);
xor (n679,n680,n25);
or (n680,n681,n682);
and (n681,n16,n190);
and (n682,n21,n194);
xor (n683,n684,n689);
xor (n684,n685,n573);
xor (n685,n686,n88);
or (n686,n687,n688);
and (n687,n48,n82);
and (n688,n56,n86);
xor (n689,n690,n24);
or (n690,n691,n692);
and (n691,n36,n17);
and (n692,n72,n22);
nand (n693,n694,n696,n697);
nand (n694,n695,n25);
xor (n695,n585,n25);
nand (n696,n588,n25);
nand (n697,n695,n588);
nand (n698,n699,n700,n701);
nand (n699,n598,n622);
nand (n700,n626,n622);
nand (n701,n598,n626);
not (n702,n703);
nor (n703,n704,n706);
nor (n704,n705,n634);
nand (n705,n562,n566);
not (n706,n707);
nand (n707,n635,n639);
nand (n708,n709,n2666);
nand (n709,n710,n2240);
nor (n710,n711,n2208);
nor (n711,n712,n1681);
nor (n712,n713,n1666);
nor (n713,n714,n1387);
nand (n714,n715,n1170);
nor (n715,n716,n1069);
nor (n716,n717,n979);
nand (n717,n718,n894,n978);
nand (n718,n719,n796);
xor (n719,n720,n772);
xor (n720,n721,n746);
xor (n721,n722,n734);
xor (n722,n723,n728);
xor (n723,n724,n88);
or (n724,n725,n726);
and (n725,n329,n82);
and (n726,n727,n86);
xor (n728,n729,n19);
or (n729,n730,n732);
and (n730,n731,n99);
and (n732,n733,n102);
xor (n734,n735,n739);
xor (n735,n736,n222);
or (n736,n737,n738);
and (n737,n36,n345);
and (n738,n72,n349);
xnor (n739,n740,n347);
nor (n740,n741,n745);
and (n741,n31,n742);
and (n742,n743,n347);
not (n743,n744);
and (n745,n60,n744);
nand (n746,n747,n757,n771);
nand (n747,n748,n752);
xor (n748,n749,n88);
or (n749,n750,n751);
and (n750,n727,n82);
and (n751,n731,n86);
xor (n752,n753,n19);
or (n753,n754,n755);
and (n754,n733,n99);
and (n755,n756,n102);
nand (n757,n758,n752);
xor (n758,n759,n768);
xor (n759,n760,n764);
xor (n760,n761,n222);
or (n761,n762,n763);
and (n762,n72,n345);
and (n763,n81,n349);
xor (n764,n765,n46);
or (n765,n766,n767);
and (n766,n21,n121);
and (n767,n135,n125);
xnor (n768,n769,n24);
nand (n769,n770,n17);
nand (n771,n748,n758);
xor (n772,n773,n782);
xor (n773,n774,n778);
xor (n774,n775,n24);
or (n775,n776,n777);
and (n776,n756,n17);
and (n777,n770,n22);
nand (n778,n779,n780,n781);
nand (n779,n760,n764);
nand (n780,n768,n764);
nand (n781,n760,n768);
xor (n782,n783,n792);
xor (n783,n784,n788);
xor (n784,n785,n46);
or (n785,n786,n787);
and (n786,n16,n121);
and (n787,n21,n125);
xor (n788,n789,n123);
or (n789,n790,n791);
and (n790,n81,n220);
and (n791,n85,n224);
xor (n792,n793,n51);
or (n793,n794,n795);
and (n794,n135,n44);
and (n795,n107,n49);
nand (n796,n797,n851,n893);
nand (n797,n798,n800);
xor (n798,n799,n758);
xor (n799,n748,n752);
xor (n800,n801,n840);
xor (n801,n802,n818);
nand (n802,n803,n812,n817);
nand (n803,n804,n808);
xor (n804,n805,n46);
or (n805,n806,n807);
and (n806,n135,n121);
and (n807,n107,n125);
xor (n808,n809,n123);
or (n809,n810,n811);
and (n810,n16,n220);
and (n811,n21,n224);
nand (n812,n813,n808);
xor (n813,n814,n51);
or (n814,n815,n816);
and (n815,n111,n44);
and (n816,n185,n49);
nand (n817,n804,n813);
nand (n818,n819,n834,n839);
nand (n819,n820,n829);
xor (n820,n821,n825);
xnor (n821,n822,n347);
nor (n822,n823,n824);
and (n823,n72,n742);
and (n824,n36,n744);
xor (n825,n826,n222);
or (n826,n827,n828);
and (n827,n81,n345);
and (n828,n85,n349);
and (n829,n830,n19);
xnor (n830,n831,n347);
nor (n831,n832,n833);
and (n832,n81,n742);
and (n833,n72,n744);
nand (n834,n835,n829);
xor (n835,n836,n34);
or (n836,n837,n838);
and (n837,n189,n57);
and (n838,n193,n61);
nand (n839,n820,n835);
xor (n840,n841,n847);
xor (n841,n842,n846);
xor (n842,n843,n34);
or (n843,n844,n845);
and (n844,n185,n57);
and (n845,n189,n61);
and (n846,n821,n825);
xor (n847,n848,n39);
or (n848,n849,n850);
and (n849,n193,n32);
and (n850,n329,n37);
nand (n851,n852,n800);
nand (n852,n853,n877,n892);
nand (n853,n854,n875);
nand (n854,n855,n869,n874);
nand (n855,n856,n865);
and (n856,n857,n861);
xnor (n857,n858,n347);
nor (n858,n859,n860);
and (n859,n85,n742);
and (n860,n81,n744);
xor (n861,n862,n222);
or (n862,n863,n864);
and (n863,n16,n345);
and (n864,n21,n349);
xor (n865,n866,n34);
or (n866,n867,n868);
and (n867,n193,n57);
and (n868,n329,n61);
nand (n869,n870,n865);
xor (n870,n871,n39);
or (n871,n872,n873);
and (n872,n727,n32);
and (n873,n731,n37);
nand (n874,n856,n870);
xor (n875,n876,n835);
xor (n876,n820,n829);
nand (n877,n878,n875);
xor (n878,n879,n888);
xor (n879,n880,n884);
xor (n880,n881,n39);
or (n881,n882,n883);
and (n882,n329,n32);
and (n883,n727,n37);
xor (n884,n885,n88);
or (n885,n886,n887);
and (n886,n731,n82);
and (n887,n733,n86);
xor (n888,n889,n19);
or (n889,n890,n891);
and (n890,n756,n99);
and (n891,n770,n102);
nand (n892,n854,n878);
nand (n893,n798,n852);
nand (n894,n895,n796);
xor (n895,n896,n935);
xor (n896,n897,n901);
nand (n897,n898,n899,n900);
nand (n898,n802,n818);
nand (n899,n840,n818);
nand (n900,n802,n840);
xor (n901,n902,n924);
xor (n902,n903,n920);
nand (n903,n904,n914,n919);
nand (n904,n905,n909);
xor (n905,n906,n123);
or (n906,n907,n908);
and (n907,n85,n220);
and (n908,n16,n224);
xor (n909,n910,n24);
xnor (n910,n911,n347);
nor (n911,n912,n913);
and (n912,n36,n742);
and (n913,n31,n744);
nand (n914,n915,n909);
xor (n915,n916,n51);
or (n916,n917,n918);
and (n917,n107,n44);
and (n918,n111,n49);
nand (n919,n905,n915);
nand (n920,n921,n922,n923);
nand (n921,n842,n846);
nand (n922,n847,n846);
nand (n923,n842,n847);
xor (n924,n925,n931);
xor (n925,n926,n927);
and (n926,n910,n24);
xor (n927,n928,n34);
or (n928,n929,n930);
and (n929,n111,n57);
and (n930,n185,n61);
xor (n931,n932,n39);
or (n932,n933,n934);
and (n933,n189,n32);
and (n934,n193,n37);
nand (n935,n936,n943,n977);
nand (n936,n937,n941);
nand (n937,n938,n939,n940);
nand (n938,n880,n884);
nand (n939,n888,n884);
nand (n940,n880,n888);
xor (n941,n942,n915);
xor (n942,n905,n909);
nand (n943,n944,n941);
nand (n944,n945,n962,n976);
nand (n945,n946,n960);
nand (n946,n947,n956,n959);
nand (n947,n948,n952);
xor (n948,n949,n222);
or (n949,n950,n951);
and (n950,n85,n345);
and (n951,n16,n349);
xor (n952,n953,n46);
or (n953,n954,n955);
and (n954,n107,n121);
and (n955,n111,n125);
nand (n956,n957,n952);
xnor (n957,n958,n19);
nand (n958,n770,n99);
nand (n959,n948,n957);
xor (n960,n961,n813);
xor (n961,n804,n808);
nand (n962,n963,n960);
nand (n963,n964,n970,n975);
nand (n964,n965,n969);
xor (n965,n966,n123);
or (n966,n967,n968);
and (n967,n21,n220);
and (n968,n135,n224);
xor (n969,n830,n19);
nand (n970,n971,n969);
xor (n971,n972,n51);
or (n972,n973,n974);
and (n973,n185,n44);
and (n974,n189,n49);
nand (n975,n965,n971);
nand (n976,n946,n963);
nand (n977,n937,n944);
nand (n978,n719,n895);
xor (n979,n980,n1065);
xor (n980,n981,n1002);
xor (n981,n982,n998);
xor (n982,n983,n994);
xor (n983,n984,n990);
xor (n984,n985,n989);
xor (n985,n986,n19);
or (n986,n987,n988);
and (n987,n727,n99);
and (n988,n731,n102);
and (n989,n735,n739);
xor (n990,n991,n24);
or (n991,n992,n993);
and (n992,n733,n17);
and (n993,n756,n22);
nand (n994,n995,n996,n997);
nand (n995,n774,n778);
nand (n996,n782,n778);
nand (n997,n774,n782);
nand (n998,n999,n1000,n1001);
nand (n999,n903,n920);
nand (n1000,n924,n920);
nand (n1001,n903,n924);
xor (n1002,n1003,n1061);
xor (n1003,n1004,n1028);
xor (n1004,n1005,n1024);
xor (n1005,n1006,n1010);
nand (n1006,n1007,n1008,n1009);
nand (n1007,n926,n927);
nand (n1008,n931,n927);
nand (n1009,n926,n931);
xor (n1010,n1011,n1020);
xor (n1011,n1012,n1016);
xnor (n1012,n1013,n347);
nor (n1013,n1014,n1015);
and (n1014,n60,n742);
and (n1015,n56,n744);
xor (n1016,n1017,n46);
or (n1017,n1018,n1019);
and (n1018,n85,n121);
and (n1019,n16,n125);
xor (n1020,n1021,n123);
or (n1021,n1022,n1023);
and (n1022,n72,n220);
and (n1023,n81,n224);
nand (n1024,n1025,n1026,n1027);
nand (n1025,n784,n788);
nand (n1026,n792,n788);
nand (n1027,n784,n792);
xor (n1028,n1029,n1047);
xor (n1029,n1030,n1034);
nand (n1030,n1031,n1032,n1033);
nand (n1031,n723,n728);
nand (n1032,n734,n728);
nand (n1033,n723,n734);
xor (n1034,n1035,n1045);
xor (n1035,n1036,n1040);
xor (n1036,n1037,n51);
or (n1037,n1038,n1039);
and (n1038,n21,n44);
and (n1039,n135,n49);
xor (n1040,n114,n1041);
xor (n1041,n1042,n222);
or (n1042,n1043,n1044);
and (n1043,n31,n345);
and (n1044,n36,n349);
xnor (n1045,n1046,n114);
nand (n1046,n770,n108);
xor (n1047,n1048,n1057);
xor (n1048,n1049,n1053);
xor (n1049,n1050,n34);
or (n1050,n1051,n1052);
and (n1051,n107,n57);
and (n1052,n111,n61);
xor (n1053,n1054,n39);
or (n1054,n1055,n1056);
and (n1055,n185,n32);
and (n1056,n189,n37);
xor (n1057,n1058,n88);
or (n1058,n1059,n1060);
and (n1059,n193,n82);
and (n1060,n329,n86);
nand (n1061,n1062,n1063,n1064);
nand (n1062,n721,n746);
nand (n1063,n772,n746);
nand (n1064,n721,n772);
nand (n1065,n1066,n1067,n1068);
nand (n1066,n897,n901);
nand (n1067,n935,n901);
nand (n1068,n897,n935);
nor (n1069,n1070,n1074);
nand (n1070,n1071,n1072,n1073);
nand (n1071,n981,n1002);
nand (n1072,n1065,n1002);
nand (n1073,n981,n1065);
xor (n1074,n1075,n1084);
xor (n1075,n1076,n1080);
nand (n1076,n1077,n1078,n1079);
nand (n1077,n983,n994);
nand (n1078,n998,n994);
nand (n1079,n983,n998);
nand (n1080,n1081,n1082,n1083);
nand (n1081,n1004,n1028);
nand (n1082,n1061,n1028);
nand (n1083,n1004,n1061);
xor (n1084,n1085,n1146);
xor (n1085,n1086,n1117);
xor (n1086,n1087,n1106);
xor (n1087,n1088,n1102);
xor (n1088,n1089,n1098);
xor (n1089,n1090,n1094);
xor (n1090,n1091,n46);
or (n1091,n1092,n1093);
and (n1092,n81,n121);
and (n1093,n85,n125);
xor (n1094,n1095,n123);
or (n1095,n1096,n1097);
and (n1096,n36,n220);
and (n1097,n72,n224);
xor (n1098,n1099,n51);
or (n1099,n1100,n1101);
and (n1100,n16,n44);
and (n1101,n21,n49);
nand (n1102,n1103,n1104,n1105);
nand (n1103,n1036,n1040);
nand (n1104,n1045,n1040);
nand (n1105,n1036,n1045);
xor (n1106,n1107,n1113);
xor (n1107,n1108,n1112);
xor (n1108,n1109,n34);
or (n1109,n1110,n1111);
and (n1110,n135,n57);
and (n1111,n107,n61);
and (n1112,n114,n1041);
xor (n1113,n1114,n39);
or (n1114,n1115,n1116);
and (n1115,n111,n32);
and (n1116,n185,n37);
xor (n1117,n1118,n1142);
xor (n1118,n1119,n1123);
nand (n1119,n1120,n1121,n1122);
nand (n1120,n1049,n1053);
nand (n1121,n1057,n1053);
nand (n1122,n1049,n1057);
xor (n1123,n1124,n1133);
xor (n1124,n1125,n1129);
xor (n1125,n1126,n88);
or (n1126,n1127,n1128);
and (n1127,n189,n82);
and (n1128,n193,n86);
xor (n1129,n1130,n19);
or (n1130,n1131,n1132);
and (n1131,n329,n99);
and (n1132,n727,n102);
xor (n1133,n1134,n1138);
xnor (n1134,n1135,n347);
nor (n1135,n1136,n1137);
and (n1136,n56,n742);
and (n1137,n48,n744);
xor (n1138,n1139,n222);
or (n1139,n1140,n1141);
and (n1140,n60,n345);
and (n1141,n31,n349);
nand (n1142,n1143,n1144,n1145);
nand (n1143,n985,n989);
nand (n1144,n990,n989);
nand (n1145,n985,n990);
xor (n1146,n1147,n1166);
xor (n1147,n1148,n1162);
xor (n1148,n1149,n1158);
xor (n1149,n1150,n1154);
xor (n1150,n1151,n24);
or (n1151,n1152,n1153);
and (n1152,n731,n17);
and (n1153,n733,n22);
xor (n1154,n1155,n114);
or (n1155,n1156,n1157);
and (n1156,n756,n108);
and (n1157,n770,n112);
nand (n1158,n1159,n1160,n1161);
nand (n1159,n1012,n1016);
nand (n1160,n1020,n1016);
nand (n1161,n1012,n1020);
nand (n1162,n1163,n1164,n1165);
nand (n1163,n1006,n1010);
nand (n1164,n1024,n1010);
nand (n1165,n1006,n1024);
nand (n1166,n1167,n1168,n1169);
nand (n1167,n1030,n1034);
nand (n1168,n1047,n1034);
nand (n1169,n1030,n1047);
nor (n1170,n1171,n1276);
nor (n1171,n1172,n1176);
nand (n1172,n1173,n1174,n1175);
nand (n1173,n1076,n1080);
nand (n1174,n1084,n1080);
nand (n1175,n1076,n1084);
xor (n1176,n1177,n1272);
xor (n1177,n1178,n1212);
xor (n1178,n1179,n1208);
xor (n1179,n1180,n1184);
nand (n1180,n1181,n1182,n1183);
nand (n1181,n1088,n1102);
nand (n1182,n1106,n1102);
nand (n1183,n1088,n1106);
xor (n1184,n1185,n1194);
xor (n1185,n1186,n1190);
xor (n1186,n1187,n114);
or (n1187,n1188,n1189);
and (n1188,n733,n108);
and (n1189,n756,n112);
nand (n1190,n1191,n1192,n1193);
nand (n1191,n1108,n1112);
nand (n1192,n1113,n1112);
nand (n1193,n1108,n1113);
xor (n1194,n1195,n1204);
xor (n1195,n1196,n1200);
xor (n1196,n1197,n46);
or (n1197,n1198,n1199);
and (n1198,n72,n121);
and (n1199,n81,n125);
xnor (n1200,n1201,n347);
nor (n1201,n1202,n1203);
and (n1202,n48,n742);
and (n1203,n43,n744);
xor (n1204,n1205,n123);
or (n1205,n1206,n1207);
and (n1206,n31,n220);
and (n1207,n36,n224);
nand (n1208,n1209,n1210,n1211);
nand (n1209,n1119,n1123);
nand (n1210,n1142,n1123);
nand (n1211,n1119,n1142);
xor (n1212,n1213,n1268);
xor (n1213,n1214,n1236);
xor (n1214,n1215,n1224);
xor (n1215,n1216,n1220);
nand (n1216,n1217,n1218,n1219);
nand (n1217,n1090,n1094);
nand (n1218,n1098,n1094);
nand (n1219,n1090,n1098);
nand (n1220,n1221,n1222,n1223);
nand (n1221,n1125,n1129);
nand (n1222,n1133,n1129);
nand (n1223,n1125,n1133);
xor (n1224,n1225,n1232);
xor (n1225,n1226,n1230);
xor (n1226,n1227,n51);
or (n1227,n1228,n1229);
and (n1228,n85,n44);
and (n1229,n16,n49);
xnor (n1230,n1231,n25);
nand (n1231,n770,n190);
xor (n1232,n1233,n34);
or (n1233,n1234,n1235);
and (n1234,n21,n57);
and (n1235,n135,n61);
xor (n1236,n1237,n1256);
xor (n1237,n1238,n1242);
nand (n1238,n1239,n1240,n1241);
nand (n1239,n1150,n1154);
nand (n1240,n1158,n1154);
nand (n1241,n1150,n1158);
xor (n1242,n1243,n1252);
xor (n1243,n1244,n1248);
xor (n1244,n1245,n39);
or (n1245,n1246,n1247);
and (n1246,n107,n32);
and (n1247,n111,n37);
xor (n1248,n1249,n88);
or (n1249,n1250,n1251);
and (n1250,n185,n82);
and (n1251,n189,n86);
xor (n1252,n1253,n19);
or (n1253,n1254,n1255);
and (n1254,n193,n99);
and (n1255,n329,n102);
xor (n1256,n1257,n1264);
xor (n1257,n1258,n1263);
xor (n1258,n25,n1259);
xor (n1259,n1260,n222);
or (n1260,n1261,n1262);
and (n1261,n56,n345);
and (n1262,n60,n349);
and (n1263,n1134,n1138);
xor (n1264,n1265,n24);
or (n1265,n1266,n1267);
and (n1266,n727,n17);
and (n1267,n731,n22);
nand (n1268,n1269,n1270,n1271);
nand (n1269,n1148,n1162);
nand (n1270,n1166,n1162);
nand (n1271,n1148,n1166);
nand (n1272,n1273,n1274,n1275);
nand (n1273,n1086,n1117);
nand (n1274,n1146,n1117);
nand (n1275,n1086,n1146);
nor (n1276,n1277,n1281);
nand (n1277,n1278,n1279,n1280);
nand (n1278,n1178,n1212);
nand (n1279,n1272,n1212);
nand (n1280,n1178,n1272);
xor (n1281,n1282,n1291);
xor (n1282,n1283,n1287);
nand (n1283,n1284,n1285,n1286);
nand (n1284,n1180,n1184);
nand (n1285,n1208,n1184);
nand (n1286,n1180,n1208);
nand (n1287,n1288,n1289,n1290);
nand (n1288,n1214,n1236);
nand (n1289,n1268,n1236);
nand (n1290,n1214,n1268);
xor (n1291,n1292,n1353);
xor (n1292,n1293,n1317);
xor (n1293,n1294,n1313);
xor (n1294,n1295,n1299);
nand (n1295,n1296,n1297,n1298);
nand (n1296,n1244,n1248);
nand (n1297,n1252,n1248);
nand (n1298,n1244,n1252);
xor (n1299,n1300,n1309);
xor (n1300,n1301,n1305);
xor (n1301,n1302,n34);
or (n1302,n1303,n1304);
and (n1303,n16,n57);
and (n1304,n21,n61);
xor (n1305,n1306,n39);
or (n1306,n1307,n1308);
and (n1307,n135,n32);
and (n1308,n107,n37);
xor (n1309,n1310,n88);
or (n1310,n1311,n1312);
and (n1311,n111,n82);
and (n1312,n185,n86);
nand (n1313,n1314,n1315,n1316);
nand (n1314,n1258,n1263);
nand (n1315,n1264,n1263);
nand (n1316,n1258,n1264);
xor (n1317,n1318,n1339);
xor (n1318,n1319,n1335);
xor (n1319,n1320,n1334);
xor (n1320,n1321,n1325);
xor (n1321,n1322,n19);
or (n1322,n1323,n1324);
and (n1323,n189,n99);
and (n1324,n193,n102);
xor (n1325,n1326,n1330);
xnor (n1326,n1327,n347);
nor (n1327,n1328,n1329);
and (n1328,n43,n742);
and (n1329,n147,n744);
xor (n1330,n1331,n222);
or (n1331,n1332,n1333);
and (n1332,n48,n345);
and (n1333,n56,n349);
and (n1334,n25,n1259);
nand (n1335,n1336,n1337,n1338);
nand (n1336,n1186,n1190);
nand (n1337,n1194,n1190);
nand (n1338,n1186,n1194);
xor (n1339,n1340,n1349);
xor (n1340,n1341,n1345);
xor (n1341,n1342,n24);
or (n1342,n1343,n1344);
and (n1343,n329,n17);
and (n1344,n727,n22);
xor (n1345,n1346,n25);
or (n1346,n1347,n1348);
and (n1347,n756,n190);
and (n1348,n770,n194);
xor (n1349,n1350,n114);
or (n1350,n1351,n1352);
and (n1351,n731,n108);
and (n1352,n733,n112);
xor (n1353,n1354,n1383);
xor (n1354,n1355,n1379);
xor (n1355,n1356,n1375);
xor (n1356,n1357,n1361);
nand (n1357,n1358,n1359,n1360);
nand (n1358,n1196,n1200);
nand (n1359,n1204,n1200);
nand (n1360,n1196,n1204);
xor (n1361,n1362,n1371);
xor (n1362,n1363,n1367);
xor (n1363,n1364,n46);
or (n1364,n1365,n1366);
and (n1365,n36,n121);
and (n1366,n72,n125);
xor (n1367,n1368,n123);
or (n1368,n1369,n1370);
and (n1369,n60,n220);
and (n1370,n31,n224);
xor (n1371,n1372,n51);
or (n1372,n1373,n1374);
and (n1373,n81,n44);
and (n1374,n85,n49);
nand (n1375,n1376,n1377,n1378);
nand (n1376,n1226,n1230);
nand (n1377,n1232,n1230);
nand (n1378,n1226,n1232);
nand (n1379,n1380,n1381,n1382);
nand (n1380,n1216,n1220);
nand (n1381,n1224,n1220);
nand (n1382,n1216,n1224);
nand (n1383,n1384,n1385,n1386);
nand (n1384,n1238,n1242);
nand (n1385,n1256,n1242);
nand (n1386,n1238,n1256);
nor (n1387,n1388,n1660);
nor (n1388,n1389,n1636);
nor (n1389,n1390,n1634);
nor (n1390,n1391,n1609);
nand (n1391,n1392,n1571);
nand (n1392,n1393,n1518,n1570);
nand (n1393,n1394,n1445);
xor (n1394,n1395,n1432);
xor (n1395,n1396,n1417);
nand (n1396,n1397,n1411,n1416);
nand (n1397,n1398,n1407);
and (n1398,n1399,n1403);
xnor (n1399,n1400,n347);
nor (n1400,n1401,n1402);
and (n1401,n21,n742);
and (n1402,n16,n744);
xor (n1403,n1404,n222);
or (n1404,n1405,n1406);
and (n1405,n135,n345);
and (n1406,n107,n349);
xor (n1407,n1408,n34);
or (n1408,n1409,n1410);
and (n1409,n727,n57);
and (n1410,n731,n61);
nand (n1411,n1412,n1407);
xor (n1412,n1413,n39);
or (n1413,n1414,n1415);
and (n1414,n733,n32);
and (n1415,n756,n37);
nand (n1416,n1398,n1412);
xor (n1417,n1418,n1427);
xor (n1418,n1419,n1423);
xor (n1419,n1420,n46);
or (n1420,n1421,n1422);
and (n1421,n111,n121);
and (n1422,n185,n125);
xor (n1423,n1424,n123);
or (n1424,n1425,n1426);
and (n1425,n135,n220);
and (n1426,n107,n224);
and (n1427,n1428,n88);
xnor (n1428,n1429,n347);
nor (n1429,n1430,n1431);
and (n1430,n16,n742);
and (n1431,n85,n744);
nand (n1432,n1433,n1439,n1444);
nand (n1433,n1434,n1438);
xor (n1434,n1435,n123);
or (n1435,n1436,n1437);
and (n1436,n107,n220);
and (n1437,n111,n224);
xor (n1438,n1428,n88);
nand (n1439,n1440,n1438);
xor (n1440,n1441,n51);
or (n1441,n1442,n1443);
and (n1442,n193,n44);
and (n1443,n329,n49);
nand (n1444,n1434,n1440);
xor (n1445,n1446,n1482);
xor (n1446,n1447,n1458);
xor (n1447,n1448,n1454);
xor (n1448,n1449,n1453);
xor (n1449,n1450,n51);
or (n1450,n1451,n1452);
and (n1451,n189,n44);
and (n1452,n193,n49);
xor (n1453,n857,n861);
xor (n1454,n1455,n34);
or (n1455,n1456,n1457);
and (n1456,n329,n57);
and (n1457,n727,n61);
xor (n1458,n1459,n1468);
xor (n1459,n1460,n1464);
xor (n1460,n1461,n39);
or (n1461,n1462,n1463);
and (n1462,n731,n32);
and (n1463,n733,n37);
xor (n1464,n1465,n88);
or (n1465,n1466,n1467);
and (n1466,n756,n82);
and (n1467,n770,n86);
nand (n1468,n1469,n1476,n1481);
nand (n1469,n1470,n1474);
xor (n1470,n1471,n222);
or (n1471,n1472,n1473);
and (n1472,n21,n345);
and (n1473,n135,n349);
xnor (n1474,n1475,n88);
nand (n1475,n770,n82);
nand (n1476,n1477,n1474);
xor (n1477,n1478,n46);
or (n1478,n1479,n1480);
and (n1479,n185,n121);
and (n1480,n189,n125);
nand (n1481,n1470,n1477);
nand (n1482,n1483,n1503,n1517);
nand (n1483,n1484,n1486);
xor (n1484,n1485,n1477);
xor (n1485,n1470,n1474);
nand (n1486,n1487,n1496,n1502);
nand (n1487,n1488,n1492);
xor (n1488,n1489,n46);
or (n1489,n1490,n1491);
and (n1490,n189,n121);
and (n1491,n193,n125);
xor (n1492,n1493,n123);
or (n1493,n1494,n1495);
and (n1494,n111,n220);
and (n1495,n185,n224);
nand (n1496,n1497,n1492);
and (n1497,n1498,n39);
xnor (n1498,n1499,n347);
nor (n1499,n1500,n1501);
and (n1500,n135,n742);
and (n1501,n21,n744);
nand (n1502,n1488,n1497);
nand (n1503,n1504,n1486);
nand (n1504,n1505,n1511,n1516);
nand (n1505,n1506,n1510);
xor (n1506,n1507,n51);
or (n1507,n1508,n1509);
and (n1508,n329,n44);
and (n1509,n727,n49);
xor (n1510,n1399,n1403);
nand (n1511,n1512,n1510);
xor (n1512,n1513,n34);
or (n1513,n1514,n1515);
and (n1514,n731,n57);
and (n1515,n733,n61);
nand (n1516,n1506,n1512);
nand (n1517,n1484,n1504);
nand (n1518,n1519,n1445);
nand (n1519,n1520,n1525,n1569);
nand (n1520,n1521,n1523);
xor (n1521,n1522,n1412);
xor (n1522,n1398,n1407);
xor (n1523,n1524,n1440);
xor (n1524,n1434,n1438);
nand (n1525,n1526,n1523);
nand (n1526,n1527,n1546,n1568);
nand (n1527,n1528,n1532);
xor (n1528,n1529,n39);
or (n1529,n1530,n1531);
and (n1530,n756,n32);
and (n1531,n770,n37);
nand (n1532,n1533,n1540,n1545);
nand (n1533,n1534,n1538);
xor (n1534,n1535,n222);
or (n1535,n1536,n1537);
and (n1536,n107,n345);
and (n1537,n111,n349);
xnor (n1538,n1539,n39);
nand (n1539,n770,n32);
nand (n1540,n1541,n1538);
xor (n1541,n1542,n46);
or (n1542,n1543,n1544);
and (n1543,n193,n121);
and (n1544,n329,n125);
nand (n1545,n1534,n1541);
nand (n1546,n1547,n1532);
nand (n1547,n1548,n1562,n1567);
nand (n1548,n1549,n1553);
xor (n1549,n1550,n123);
or (n1550,n1551,n1552);
and (n1551,n185,n220);
and (n1552,n189,n224);
and (n1553,n1554,n1558);
xnor (n1554,n1555,n347);
nor (n1555,n1556,n1557);
and (n1556,n107,n742);
and (n1557,n135,n744);
xor (n1558,n1559,n222);
or (n1559,n1560,n1561);
and (n1560,n111,n345);
and (n1561,n185,n349);
nand (n1562,n1563,n1553);
xor (n1563,n1564,n51);
or (n1564,n1565,n1566);
and (n1565,n727,n44);
and (n1566,n731,n49);
nand (n1567,n1549,n1563);
nand (n1568,n1528,n1547);
nand (n1569,n1521,n1526);
nand (n1570,n1394,n1519);
xor (n1571,n1572,n1587);
xor (n1572,n1573,n1583);
xor (n1573,n1574,n1581);
xor (n1574,n1575,n1579);
nand (n1575,n1576,n1577,n1578);
nand (n1576,n1419,n1423);
nand (n1577,n1427,n1423);
nand (n1578,n1419,n1427);
xor (n1579,n1580,n870);
xor (n1580,n856,n865);
xor (n1581,n1582,n971);
xor (n1582,n965,n969);
nand (n1583,n1584,n1585,n1586);
nand (n1584,n1447,n1458);
nand (n1585,n1482,n1458);
nand (n1586,n1447,n1482);
xor (n1587,n1588,n1597);
xor (n1588,n1589,n1593);
nand (n1589,n1590,n1591,n1592);
nand (n1590,n1460,n1464);
nand (n1591,n1468,n1464);
nand (n1592,n1460,n1468);
nand (n1593,n1594,n1595,n1596);
nand (n1594,n1396,n1417);
nand (n1595,n1432,n1417);
nand (n1596,n1396,n1432);
xor (n1597,n1598,n1607);
xor (n1598,n1599,n1603);
xor (n1599,n1600,n88);
or (n1600,n1601,n1602);
and (n1601,n733,n82);
and (n1602,n756,n86);
nand (n1603,n1604,n1605,n1606);
nand (n1604,n1449,n1453);
nand (n1605,n1454,n1453);
nand (n1606,n1449,n1454);
xor (n1607,n1608,n957);
xor (n1608,n948,n952);
nor (n1609,n1610,n1614);
nand (n1610,n1611,n1612,n1613);
nand (n1611,n1573,n1583);
nand (n1612,n1587,n1583);
nand (n1613,n1573,n1587);
xor (n1614,n1615,n1622);
xor (n1615,n1616,n1618);
xor (n1616,n1617,n878);
xor (n1617,n854,n875);
nand (n1618,n1619,n1620,n1621);
nand (n1619,n1589,n1593);
nand (n1620,n1597,n1593);
nand (n1621,n1589,n1597);
xor (n1622,n1623,n1632);
xor (n1623,n1624,n1628);
nand (n1624,n1625,n1626,n1627);
nand (n1625,n1599,n1603);
nand (n1626,n1607,n1603);
nand (n1627,n1599,n1607);
nand (n1628,n1629,n1630,n1631);
nand (n1629,n1575,n1579);
nand (n1630,n1581,n1579);
nand (n1631,n1575,n1581);
xor (n1632,n1633,n963);
xor (n1633,n946,n960);
not (n1634,n1635);
nand (n1635,n1610,n1614);
not (n1636,n1637);
nor (n1637,n1638,n1653);
nor (n1638,n1639,n1643);
nand (n1639,n1640,n1641,n1642);
nand (n1640,n1616,n1618);
nand (n1641,n1622,n1618);
nand (n1642,n1616,n1622);
xor (n1643,n1644,n1651);
xor (n1644,n1645,n1647);
xor (n1645,n1646,n944);
xor (n1646,n937,n941);
nand (n1647,n1648,n1649,n1650);
nand (n1648,n1624,n1628);
nand (n1649,n1632,n1628);
nand (n1650,n1624,n1632);
xor (n1651,n1652,n852);
xor (n1652,n798,n800);
nor (n1653,n1654,n1658);
nand (n1654,n1655,n1656,n1657);
nand (n1655,n1645,n1647);
nand (n1656,n1651,n1647);
nand (n1657,n1645,n1651);
xor (n1658,n1659,n895);
xor (n1659,n719,n796);
not (n1660,n1661);
nor (n1661,n1662,n1664);
nor (n1662,n1663,n1653);
nand (n1663,n1639,n1643);
not (n1664,n1665);
nand (n1665,n1654,n1658);
not (n1666,n1667);
nor (n1667,n1668,n1675);
nor (n1668,n1669,n1674);
nor (n1669,n1670,n1672);
nor (n1670,n1671,n1069);
nand (n1671,n717,n979);
not (n1672,n1673);
nand (n1673,n1070,n1074);
not (n1674,n1170);
not (n1675,n1676);
nor (n1676,n1677,n1679);
nor (n1677,n1678,n1276);
nand (n1678,n1172,n1176);
not (n1679,n1680);
nand (n1680,n1277,n1281);
not (n1681,n1682);
nor (n1682,n1683,n2098);
nand (n1683,n1684,n1911);
nor (n1684,n1685,n1797);
nor (n1685,n1686,n1690);
nand (n1686,n1687,n1688,n1689);
nand (n1687,n1283,n1287);
nand (n1688,n1291,n1287);
nand (n1689,n1283,n1291);
xor (n1690,n1691,n1793);
xor (n1691,n1692,n1725);
xor (n1692,n1693,n1721);
xor (n1693,n1694,n1717);
xor (n1694,n1695,n1713);
xor (n1695,n1696,n1709);
xor (n1696,n1697,n1706);
xor (n1697,n1698,n1702);
xor (n1698,n1699,n222);
or (n1699,n1700,n1701);
and (n1700,n43,n345);
and (n1701,n48,n349);
xor (n1702,n1703,n123);
or (n1703,n1704,n1705);
and (n1704,n56,n220);
and (n1705,n60,n224);
xnor (n1706,n1707,n347);
nor (n1707,n1708,n1329);
and (n1708,n147,n742);
nand (n1709,n1710,n1711,n1712);
nand (n1710,n1301,n1305);
nand (n1711,n1309,n1305);
nand (n1712,n1301,n1309);
nand (n1713,n1714,n1715,n1716);
nand (n1714,n1321,n1325);
nand (n1715,n1334,n1325);
nand (n1716,n1321,n1334);
nand (n1717,n1718,n1719,n1720);
nand (n1718,n1295,n1299);
nand (n1719,n1313,n1299);
nand (n1720,n1295,n1313);
nand (n1721,n1722,n1723,n1724);
nand (n1722,n1319,n1335);
nand (n1723,n1339,n1335);
nand (n1724,n1319,n1339);
xor (n1725,n1726,n1789);
xor (n1726,n1727,n1765);
xor (n1727,n1728,n1750);
xor (n1728,n1729,n1743);
xor (n1729,n1730,n1739);
xor (n1730,n1731,n1735);
xor (n1731,n1732,n51);
or (n1732,n1733,n1734);
and (n1733,n72,n44);
and (n1734,n81,n49);
xor (n1735,n1736,n34);
or (n1736,n1737,n1738);
and (n1737,n85,n57);
and (n1738,n16,n61);
xor (n1739,n1740,n39);
or (n1740,n1741,n1742);
and (n1741,n21,n32);
and (n1742,n135,n37);
xor (n1743,n1744,n1746);
xor (n1744,n25,n1745);
and (n1745,n1326,n1330);
xor (n1746,n1747,n24);
or (n1747,n1748,n1749);
and (n1748,n193,n17);
and (n1749,n329,n22);
xor (n1750,n1751,n1760);
xor (n1751,n1752,n1756);
xor (n1752,n1753,n88);
or (n1753,n1754,n1755);
and (n1754,n107,n82);
and (n1755,n111,n86);
xor (n1756,n1757,n19);
or (n1757,n1758,n1759);
and (n1758,n185,n99);
and (n1759,n189,n102);
xor (n1760,n25,n1761);
xor (n1761,n1762,n46);
or (n1762,n1763,n1764);
and (n1763,n31,n121);
and (n1764,n36,n125);
xor (n1765,n1766,n1775);
xor (n1766,n1767,n1771);
nand (n1767,n1768,n1769,n1770);
nand (n1768,n1341,n1345);
nand (n1769,n1349,n1345);
nand (n1770,n1341,n1349);
nand (n1771,n1772,n1773,n1774);
nand (n1772,n1357,n1361);
nand (n1773,n1375,n1361);
nand (n1774,n1357,n1375);
xor (n1775,n1776,n1785);
xor (n1776,n1777,n1781);
xor (n1777,n1778,n114);
or (n1778,n1779,n1780);
and (n1779,n727,n108);
and (n1780,n731,n112);
xor (n1781,n1782,n25);
or (n1782,n1783,n1784);
and (n1783,n733,n190);
and (n1784,n756,n194);
nand (n1785,n1786,n1787,n1788);
nand (n1786,n1363,n1367);
nand (n1787,n1371,n1367);
nand (n1788,n1363,n1371);
nand (n1789,n1790,n1791,n1792);
nand (n1790,n1355,n1379);
nand (n1791,n1383,n1379);
nand (n1792,n1355,n1383);
nand (n1793,n1794,n1795,n1796);
nand (n1794,n1293,n1317);
nand (n1795,n1353,n1317);
nand (n1796,n1293,n1353);
nor (n1797,n1798,n1802);
nand (n1798,n1799,n1800,n1801);
nand (n1799,n1692,n1725);
nand (n1800,n1793,n1725);
nand (n1801,n1692,n1793);
xor (n1802,n1803,n1812);
xor (n1803,n1804,n1808);
nand (n1804,n1805,n1806,n1807);
nand (n1805,n1694,n1717);
nand (n1806,n1721,n1717);
nand (n1807,n1694,n1721);
nand (n1808,n1809,n1810,n1811);
nand (n1809,n1727,n1765);
nand (n1810,n1789,n1765);
nand (n1811,n1727,n1789);
xor (n1812,n1813,n1870);
xor (n1813,n1814,n1845);
xor (n1814,n1815,n1831);
xor (n1815,n1816,n1820);
nand (n1816,n1817,n1818,n1819);
nand (n1817,n25,n1745);
nand (n1818,n1746,n1745);
nand (n1819,n25,n1746);
xor (n1820,n1821,n1827);
xor (n1821,n1822,n1826);
xor (n1822,n1823,n19);
or (n1823,n1824,n1825);
and (n1824,n111,n99);
and (n1825,n185,n102);
and (n1826,n25,n1761);
xor (n1827,n1828,n24);
or (n1828,n1829,n1830);
and (n1829,n189,n17);
and (n1830,n193,n22);
xor (n1831,n1832,n1841);
xor (n1832,n1833,n1837);
xor (n1833,n1834,n114);
or (n1834,n1835,n1836);
and (n1835,n329,n108);
and (n1836,n727,n112);
xor (n1837,n1838,n25);
or (n1838,n1839,n1840);
and (n1839,n731,n190);
and (n1840,n733,n194);
nand (n1841,n1842,n1843,n1844);
nand (n1842,n1698,n1702);
nand (n1843,n1706,n1702);
nand (n1844,n1698,n1706);
xor (n1845,n1846,n1855);
xor (n1846,n1847,n1851);
nand (n1847,n1848,n1849,n1850);
nand (n1848,n1777,n1781);
nand (n1849,n1785,n1781);
nand (n1850,n1777,n1785);
nand (n1851,n1852,n1853,n1854);
nand (n1852,n1696,n1709);
nand (n1853,n1713,n1709);
nand (n1854,n1696,n1713);
xor (n1855,n1856,n25);
xor (n1856,n1857,n1861);
nand (n1857,n1858,n1859,n1860);
nand (n1858,n1731,n1735);
nand (n1859,n1739,n1735);
nand (n1860,n1731,n1739);
xor (n1861,n1862,n1867);
not (n1862,n1863);
xor (n1863,n1864,n46);
or (n1864,n1865,n1866);
and (n1865,n60,n121);
and (n1866,n31,n125);
xor (n1867,n1868,n222);
or (n1868,n344,n1869);
and (n1869,n43,n349);
xor (n1870,n1871,n1907);
xor (n1871,n1872,n1876);
nand (n1872,n1873,n1874,n1875);
nand (n1873,n1729,n1743);
nand (n1874,n1750,n1743);
nand (n1875,n1729,n1750);
xor (n1876,n1877,n1896);
xor (n1877,n1878,n1882);
nand (n1878,n1879,n1880,n1881);
nand (n1879,n1752,n1756);
nand (n1880,n1760,n1756);
nand (n1881,n1752,n1760);
xor (n1882,n1883,n1892);
xor (n1883,n1884,n1888);
xor (n1884,n1885,n34);
or (n1885,n1886,n1887);
and (n1886,n81,n57);
and (n1887,n85,n61);
xor (n1888,n1889,n39);
or (n1889,n1890,n1891);
and (n1890,n16,n32);
and (n1891,n21,n37);
xor (n1892,n1893,n88);
or (n1893,n1894,n1895);
and (n1894,n135,n82);
and (n1895,n107,n86);
xor (n1896,n1897,n1903);
xor (n1897,n1898,n1902);
xor (n1898,n1899,n123);
or (n1899,n1900,n1901);
and (n1900,n48,n220);
and (n1901,n56,n224);
not (n1902,n1706);
xor (n1903,n1904,n51);
or (n1904,n1905,n1906);
and (n1905,n36,n44);
and (n1906,n72,n49);
nand (n1907,n1908,n1909,n1910);
nand (n1908,n1767,n1771);
nand (n1909,n1775,n1771);
nand (n1910,n1767,n1775);
nor (n1911,n1912,n2019);
nor (n1912,n1913,n1917);
nand (n1913,n1914,n1915,n1916);
nand (n1914,n1804,n1808);
nand (n1915,n1812,n1808);
nand (n1916,n1804,n1812);
xor (n1917,n1918,n2015);
xor (n1918,n1919,n1959);
xor (n1919,n1920,n1955);
xor (n1920,n1921,n1951);
xor (n1921,n1922,n1947);
xor (n1922,n1923,n1937);
xor (n1923,n1924,n1933);
xor (n1924,n1925,n1929);
xor (n1925,n1926,n34);
or (n1926,n1927,n1928);
and (n1927,n72,n57);
and (n1928,n81,n61);
xor (n1929,n1930,n39);
or (n1930,n1931,n1932);
and (n1931,n85,n32);
and (n1932,n16,n37);
xor (n1933,n1934,n19);
or (n1934,n1935,n1936);
and (n1935,n107,n99);
and (n1936,n111,n102);
xor (n1937,n1938,n1943);
xor (n1938,n1939,n342);
xor (n1939,n1940,n46);
or (n1940,n1941,n1942);
and (n1941,n56,n121);
and (n1942,n60,n125);
xor (n1943,n1944,n51);
or (n1944,n1945,n1946);
and (n1945,n31,n44);
and (n1946,n36,n49);
nand (n1947,n1948,n1949,n1950);
nand (n1948,n1822,n1826);
nand (n1949,n1827,n1826);
nand (n1950,n1822,n1827);
nand (n1951,n1952,n1953,n1954);
nand (n1952,n1816,n1820);
nand (n1953,n1831,n1820);
nand (n1954,n1816,n1831);
nand (n1955,n1956,n1957,n1958);
nand (n1956,n1847,n1851);
nand (n1957,n1855,n1851);
nand (n1958,n1847,n1855);
xor (n1959,n1960,n2011);
xor (n1960,n1961,n1982);
xor (n1961,n1962,n1978);
xor (n1962,n1963,n1974);
xor (n1963,n1964,n1970);
xor (n1964,n1965,n1966);
not (n1965,n383);
xor (n1966,n1967,n88);
or (n1967,n1968,n1969);
and (n1968,n21,n82);
and (n1969,n135,n86);
xor (n1970,n1971,n24);
or (n1971,n1972,n1973);
and (n1972,n185,n17);
and (n1973,n189,n22);
nand (n1974,n1975,n1976,n1977);
nand (n1975,n1833,n1837);
nand (n1976,n1841,n1837);
nand (n1977,n1833,n1841);
nand (n1978,n1979,n1980,n1981);
nand (n1979,n1857,n1861);
nand (n1980,n25,n1861);
nand (n1981,n1857,n25);
xor (n1982,n1983,n2007);
xor (n1983,n1984,n1997);
xor (n1984,n1985,n1994);
xor (n1985,n1986,n1990);
xor (n1986,n1987,n114);
or (n1987,n1988,n1989);
and (n1988,n193,n108);
and (n1989,n329,n112);
xor (n1990,n1991,n25);
or (n1991,n1992,n1993);
and (n1992,n727,n190);
and (n1993,n731,n194);
nand (n1994,n1862,n1995,n1996);
nand (n1995,n1867,n1863);
not (n1996,n1867);
xor (n1997,n1998,n2003);
xor (n1998,n25,n1999);
nand (n1999,n2000,n2001,n2002);
nand (n2000,n1898,n1902);
nand (n2001,n1903,n1902);
nand (n2002,n1898,n1903);
nand (n2003,n2004,n2005,n2006);
nand (n2004,n1884,n1888);
nand (n2005,n1892,n1888);
nand (n2006,n1884,n1892);
nand (n2007,n2008,n2009,n2010);
nand (n2008,n1878,n1882);
nand (n2009,n1896,n1882);
nand (n2010,n1878,n1896);
nand (n2011,n2012,n2013,n2014);
nand (n2012,n1872,n1876);
nand (n2013,n1907,n1876);
nand (n2014,n1872,n1907);
nand (n2015,n2016,n2017,n2018);
nand (n2016,n1814,n1845);
nand (n2017,n1870,n1845);
nand (n2018,n1814,n1870);
nor (n2019,n2020,n2024);
nand (n2020,n2021,n2022,n2023);
nand (n2021,n1919,n1959);
nand (n2022,n2015,n1959);
nand (n2023,n1919,n2015);
xor (n2024,n2025,n2034);
xor (n2025,n2026,n2030);
nand (n2026,n2027,n2028,n2029);
nand (n2027,n1921,n1951);
nand (n2028,n1955,n1951);
nand (n2029,n1921,n1955);
nand (n2030,n2031,n2032,n2033);
nand (n2031,n1961,n1982);
nand (n2032,n2011,n1982);
nand (n2033,n1961,n2011);
xor (n2034,n2035,n2066);
xor (n2035,n2036,n2040);
nand (n2036,n2037,n2038,n2039);
nand (n2037,n1984,n1997);
nand (n2038,n2007,n1997);
nand (n2039,n1984,n2007);
xor (n2040,n2041,n2054);
xor (n2041,n2042,n2046);
nand (n2042,n2043,n2044,n2045);
nand (n2043,n25,n1999);
nand (n2044,n2003,n1999);
nand (n2045,n25,n2003);
xor (n2046,n2047,n2050);
xor (n2047,n2048,n25);
xor (n2048,n2049,n341);
xor (n2049,n333,n336);
nand (n2050,n2051,n2052,n2053);
nand (n2051,n1939,n342);
nand (n2052,n1943,n342);
nand (n2053,n1939,n1943);
xor (n2054,n2055,n2062);
xor (n2055,n2056,n2058);
xor (n2056,n2057,n369);
xor (n2057,n360,n364);
nand (n2058,n2059,n2060,n2061);
nand (n2059,n1925,n1929);
nand (n2060,n1933,n1929);
nand (n2061,n1925,n1933);
nand (n2062,n2063,n2064,n2065);
nand (n2063,n1986,n1990);
nand (n2064,n1994,n1990);
nand (n2065,n1986,n1994);
xor (n2066,n2067,n2076);
xor (n2067,n2068,n2072);
nand (n2068,n2069,n2070,n2071);
nand (n2069,n1923,n1937);
nand (n2070,n1947,n1937);
nand (n2071,n1923,n1947);
nand (n2072,n2073,n2074,n2075);
nand (n2073,n1963,n1974);
nand (n2074,n1978,n1974);
nand (n2075,n1963,n1978);
xor (n2076,n2077,n2084);
xor (n2077,n2078,n2082);
nand (n2078,n2079,n2080,n2081);
nand (n2079,n1965,n1966);
nand (n2080,n1970,n1966);
nand (n2081,n1965,n1970);
xor (n2082,n2083,n388);
xor (n2083,n379,n383);
xor (n2084,n2085,n2094);
xor (n2085,n2086,n2090);
xor (n2086,n2087,n24);
or (n2087,n2088,n2089);
and (n2088,n111,n17);
and (n2089,n185,n22);
xor (n2090,n2091,n114);
or (n2091,n2092,n2093);
and (n2092,n189,n108);
and (n2093,n193,n112);
xor (n2094,n2095,n25);
or (n2095,n2096,n2097);
and (n2096,n329,n190);
and (n2097,n727,n194);
nand (n2098,n2099,n2183);
nor (n2099,n2100,n2150);
nor (n2100,n2101,n2105);
nand (n2101,n2102,n2103,n2104);
nand (n2102,n2026,n2030);
nand (n2103,n2034,n2030);
nand (n2104,n2026,n2034);
xor (n2105,n2106,n2146);
xor (n2106,n2107,n2127);
xor (n2107,n2108,n2115);
xor (n2108,n2109,n2111);
xor (n2109,n2110,n377);
xor (n2110,n358,n374);
nand (n2111,n2112,n2113,n2114);
nand (n2112,n2078,n2082);
nand (n2113,n2084,n2082);
nand (n2114,n2078,n2084);
xor (n2115,n2116,n2123);
xor (n2116,n2117,n2121);
nand (n2117,n2118,n2119,n2120);
nand (n2118,n2086,n2090);
nand (n2119,n2094,n2090);
nand (n2120,n2086,n2094);
xor (n2121,n2122,n287);
xor (n2122,n281,n285);
nand (n2123,n2124,n2125,n2126);
nand (n2124,n2048,n25);
nand (n2125,n2050,n25);
nand (n2126,n2048,n2050);
xor (n2127,n2128,n2142);
xor (n2128,n2129,n2133);
nand (n2129,n2130,n2131,n2132);
nand (n2130,n2042,n2046);
nand (n2131,n2054,n2046);
nand (n2132,n2042,n2054);
xor (n2133,n2134,n2138);
xor (n2134,n2135,n2137);
xor (n2135,n2136,n303);
xor (n2136,n294,n298);
xor (n2137,n326,n331);
nand (n2138,n2139,n2140,n2141);
nand (n2139,n2056,n2058);
nand (n2140,n2062,n2058);
nand (n2141,n2056,n2062);
nand (n2142,n2143,n2144,n2145);
nand (n2143,n2068,n2072);
nand (n2144,n2076,n2072);
nand (n2145,n2068,n2076);
nand (n2146,n2147,n2148,n2149);
nand (n2147,n2036,n2040);
nand (n2148,n2066,n2040);
nand (n2149,n2036,n2066);
nor (n2150,n2151,n2155);
nand (n2151,n2152,n2153,n2154);
nand (n2152,n2107,n2127);
nand (n2153,n2146,n2127);
nand (n2154,n2107,n2146);
xor (n2155,n2156,n2179);
xor (n2156,n2157,n2167);
xor (n2157,n2158,n2165);
xor (n2158,n2159,n2161);
xor (n2159,n2160,n274);
xor (n2160,n259,n271);
nand (n2161,n2162,n2163,n2164);
nand (n2162,n2117,n2121);
nand (n2163,n2123,n2121);
nand (n2164,n2117,n2123);
xor (n2165,n2166,n309);
xor (n2166,n279,n292);
xor (n2167,n2168,n2175);
xor (n2168,n2169,n2171);
xor (n2169,n2170,n356);
xor (n2170,n323,n353);
nand (n2171,n2172,n2173,n2174);
nand (n2172,n2135,n2137);
nand (n2173,n2138,n2137);
nand (n2174,n2135,n2138);
nand (n2175,n2176,n2177,n2178);
nand (n2176,n2109,n2111);
nand (n2177,n2115,n2111);
nand (n2178,n2109,n2115);
nand (n2179,n2180,n2181,n2182);
nand (n2180,n2129,n2133);
nand (n2181,n2142,n2133);
nand (n2182,n2129,n2142);
nor (n2183,n2184,n2201);
nor (n2184,n2185,n2189);
nand (n2185,n2186,n2187,n2188);
nand (n2186,n2157,n2167);
nand (n2187,n2179,n2167);
nand (n2188,n2157,n2179);
xor (n2189,n2190,n2197);
xor (n2190,n2191,n2195);
nand (n2191,n2192,n2193,n2194);
nand (n2192,n2159,n2161);
nand (n2193,n2165,n2161);
nand (n2194,n2159,n2165);
xor (n2195,n2196,n396);
xor (n2196,n319,n321);
nand (n2197,n2198,n2199,n2200);
nand (n2198,n2169,n2171);
nand (n2199,n2175,n2171);
nand (n2200,n2169,n2175);
nor (n2201,n2202,n2206);
nand (n2202,n2203,n2204,n2205);
nand (n2203,n2191,n2195);
nand (n2204,n2197,n2195);
nand (n2205,n2191,n2197);
xor (n2206,n2207,n317);
xor (n2207,n9,n175);
not (n2208,n2209);
nor (n2209,n2210,n2225);
nor (n2210,n2098,n2211);
nor (n2211,n2212,n2219);
nor (n2212,n2213,n2218);
nor (n2213,n2214,n2216);
nor (n2214,n2215,n1797);
nand (n2215,n1686,n1690);
not (n2216,n2217);
nand (n2217,n1798,n1802);
not (n2218,n1911);
not (n2219,n2220);
nor (n2220,n2221,n2223);
nor (n2221,n2222,n2019);
nand (n2222,n1913,n1917);
not (n2223,n2224);
nand (n2224,n2020,n2024);
not (n2225,n2226);
nor (n2226,n2227,n2234);
nor (n2227,n2228,n2233);
nor (n2228,n2229,n2231);
nor (n2229,n2230,n2150);
nand (n2230,n2101,n2105);
not (n2231,n2232);
nand (n2232,n2151,n2155);
not (n2233,n2183);
not (n2234,n2235);
nor (n2235,n2236,n2238);
nor (n2236,n2237,n2201);
nand (n2237,n2185,n2189);
not (n2238,n2239);
nand (n2239,n2202,n2206);
nand (n2240,n2241,n2660);
nand (n2241,n2242,n2553);
nor (n2242,n2243,n2538);
nor (n2243,n2244,n2409);
nand (n2244,n2245,n2386);
nor (n2245,n2246,n2363);
nor (n2246,n2247,n2336);
nand (n2247,n2248,n2293,n2335);
nand (n2248,n2249,n2261);
xor (n2249,n2250,n2256);
xor (n2250,n2251,n2252);
xor (n2251,n1554,n1558);
xor (n2252,n2253,n34);
or (n2253,n2254,n2255);
and (n2254,n756,n57);
and (n2255,n770,n61);
and (n2256,n34,n2257);
xor (n2257,n2258,n222);
or (n2258,n2259,n2260);
and (n2259,n185,n345);
and (n2260,n189,n349);
nand (n2261,n2262,n2279,n2292);
nand (n2262,n2263,n2264);
xor (n2263,n34,n2257);
nand (n2264,n2265,n2274,n2278);
nand (n2265,n2266,n2270);
xor (n2266,n2267,n46);
or (n2267,n2268,n2269);
and (n2268,n731,n121);
and (n2269,n733,n125);
xor (n2270,n2271,n123);
or (n2271,n2272,n2273);
and (n2272,n329,n220);
and (n2273,n727,n224);
nand (n2274,n2275,n2270);
and (n2275,n51,n2276);
xnor (n2276,n2277,n51);
nand (n2277,n770,n44);
nand (n2278,n2266,n2275);
nand (n2279,n2280,n2264);
xor (n2280,n2281,n2288);
xor (n2281,n2282,n2286);
xnor (n2282,n2283,n347);
nor (n2283,n2284,n2285);
and (n2284,n111,n742);
and (n2285,n107,n744);
xnor (n2286,n2287,n34);
nand (n2287,n770,n57);
xor (n2288,n2289,n46);
or (n2289,n2290,n2291);
and (n2290,n727,n121);
and (n2291,n731,n125);
nand (n2292,n2263,n2280);
nand (n2293,n2294,n2261);
xor (n2294,n2295,n2314);
xor (n2295,n2296,n2300);
nand (n2296,n2297,n2298,n2299);
nand (n2297,n2282,n2286);
nand (n2298,n2288,n2286);
nand (n2299,n2282,n2288);
xor (n2300,n2301,n2310);
xor (n2301,n2302,n2306);
xor (n2302,n2303,n46);
or (n2303,n2304,n2305);
and (n2304,n329,n121);
and (n2305,n727,n125);
xor (n2306,n2307,n123);
or (n2307,n2308,n2309);
and (n2308,n189,n220);
and (n2309,n193,n224);
xor (n2310,n2311,n51);
or (n2311,n2312,n2313);
and (n2312,n731,n44);
and (n2313,n733,n49);
nand (n2314,n2315,n2329,n2334);
nand (n2315,n2316,n2320);
xor (n2316,n2317,n123);
or (n2317,n2318,n2319);
and (n2318,n193,n220);
and (n2319,n329,n224);
and (n2320,n2321,n2325);
xnor (n2321,n2322,n347);
nor (n2322,n2323,n2324);
and (n2323,n185,n742);
and (n2324,n111,n744);
xor (n2325,n2326,n222);
or (n2326,n2327,n2328);
and (n2327,n189,n345);
and (n2328,n193,n349);
nand (n2329,n2330,n2320);
xor (n2330,n2331,n51);
or (n2331,n2332,n2333);
and (n2332,n733,n44);
and (n2333,n756,n49);
nand (n2334,n2316,n2330);
nand (n2335,n2249,n2294);
xor (n2336,n2337,n2351);
xor (n2337,n2338,n2347);
xor (n2338,n2339,n2345);
xor (n2339,n2340,n2344);
xor (n2340,n2341,n34);
or (n2341,n2342,n2343);
and (n2342,n733,n57);
and (n2343,n756,n61);
xor (n2344,n1498,n39);
xor (n2345,n2346,n1541);
xor (n2346,n1534,n1538);
nand (n2347,n2348,n2349,n2350);
nand (n2348,n2296,n2300);
nand (n2349,n2314,n2300);
nand (n2350,n2296,n2314);
xor (n2351,n2352,n2361);
xor (n2352,n2353,n2357);
nand (n2353,n2354,n2355,n2356);
nand (n2354,n2251,n2252);
nand (n2355,n2256,n2252);
nand (n2356,n2251,n2256);
nand (n2357,n2358,n2359,n2360);
nand (n2358,n2302,n2306);
nand (n2359,n2310,n2306);
nand (n2360,n2302,n2310);
xor (n2361,n2362,n1563);
xor (n2362,n1549,n1553);
nor (n2363,n2364,n2368);
nand (n2364,n2365,n2366,n2367);
nand (n2365,n2338,n2347);
nand (n2366,n2351,n2347);
nand (n2367,n2338,n2351);
xor (n2368,n2369,n2376);
xor (n2369,n2370,n2372);
xor (n2370,n2371,n1547);
xor (n2371,n1528,n1532);
nand (n2372,n2373,n2374,n2375);
nand (n2373,n2353,n2357);
nand (n2374,n2361,n2357);
nand (n2375,n2353,n2361);
xor (n2376,n2377,n2382);
xor (n2377,n2378,n2380);
xor (n2378,n2379,n1497);
xor (n2379,n1488,n1492);
xor (n2380,n2381,n1512);
xor (n2381,n1506,n1510);
nand (n2382,n2383,n2384,n2385);
nand (n2383,n2340,n2344);
nand (n2384,n2345,n2344);
nand (n2385,n2340,n2345);
nor (n2386,n2387,n2402);
nor (n2387,n2388,n2392);
nand (n2388,n2389,n2390,n2391);
nand (n2389,n2370,n2372);
nand (n2390,n2376,n2372);
nand (n2391,n2370,n2376);
xor (n2392,n2393,n2400);
xor (n2393,n2394,n2396);
xor (n2394,n2395,n1504);
xor (n2395,n1484,n1486);
nand (n2396,n2397,n2398,n2399);
nand (n2397,n2378,n2380);
nand (n2398,n2382,n2380);
nand (n2399,n2378,n2382);
xor (n2400,n2401,n1526);
xor (n2401,n1521,n1523);
nor (n2402,n2403,n2407);
nand (n2403,n2404,n2405,n2406);
nand (n2404,n2394,n2396);
nand (n2405,n2400,n2396);
nand (n2406,n2394,n2400);
xor (n2407,n2408,n1519);
xor (n2408,n1394,n1445);
nor (n2409,n2410,n2532);
nor (n2410,n2411,n2508);
nor (n2411,n2412,n2505);
nor (n2412,n2413,n2481);
nand (n2413,n2414,n2453);
or (n2414,n2415,n2439,n2452);
and (n2415,n2416,n2425);
xor (n2416,n2417,n2421);
xnor (n2417,n2418,n347);
nor (n2418,n2419,n2420);
and (n2419,n193,n742);
and (n2420,n189,n744);
xnor (n2421,n2422,n222);
nor (n2422,n2423,n2424);
and (n2423,n727,n349);
and (n2424,n329,n345);
or (n2425,n2426,n2433,n2438);
and (n2426,n2427,n2429);
not (n2427,n2428);
nand (n2428,n770,n121);
xnor (n2429,n2430,n347);
nor (n2430,n2431,n2432);
and (n2431,n329,n742);
and (n2432,n193,n744);
and (n2433,n2429,n2434);
xnor (n2434,n2435,n222);
nor (n2435,n2436,n2437);
and (n2436,n731,n349);
and (n2437,n727,n345);
and (n2438,n2427,n2434);
and (n2439,n2425,n2440);
xor (n2440,n2441,n2448);
xor (n2441,n2442,n2444);
and (n2442,n46,n2443);
xnor (n2443,n2428,n46);
xnor (n2444,n2445,n123);
nor (n2445,n2446,n2447);
and (n2446,n733,n224);
and (n2447,n731,n220);
xnor (n2448,n2449,n46);
nor (n2449,n2450,n2451);
and (n2450,n770,n125);
and (n2451,n756,n121);
and (n2452,n2416,n2440);
xor (n2453,n2454,n2470);
xor (n2454,n2455,n2459);
or (n2455,n2456,n2457,n2458);
and (n2456,n2442,n2444);
and (n2457,n2444,n2448);
and (n2458,n2442,n2448);
xor (n2459,n2460,n2466);
xor (n2460,n2461,n2462);
and (n2461,n2417,n2421);
xnor (n2462,n2463,n123);
nor (n2463,n2464,n2465);
and (n2464,n731,n224);
and (n2465,n727,n220);
xnor (n2466,n2467,n46);
nor (n2467,n2468,n2469);
and (n2468,n756,n125);
and (n2469,n733,n121);
xor (n2470,n2471,n2477);
xor (n2471,n2472,n2473);
not (n2472,n2277);
xnor (n2473,n2474,n347);
nor (n2474,n2475,n2476);
and (n2475,n189,n742);
and (n2476,n185,n744);
xnor (n2477,n2478,n222);
nor (n2478,n2479,n2480);
and (n2479,n329,n349);
and (n2480,n193,n345);
nor (n2481,n2482,n2486);
or (n2482,n2483,n2484,n2485);
and (n2483,n2455,n2459);
and (n2484,n2459,n2470);
and (n2485,n2455,n2470);
xor (n2486,n2487,n2494);
xor (n2487,n2488,n2492);
or (n2488,n2489,n2490,n2491);
and (n2489,n2461,n2462);
and (n2490,n2462,n2466);
and (n2491,n2461,n2466);
xor (n2492,n2493,n2275);
xor (n2493,n2266,n2270);
xor (n2494,n2495,n2501);
xor (n2495,n2496,n2500);
xor (n2496,n2497,n51);
or (n2497,n2498,n2499);
and (n2498,n756,n44);
and (n2499,n770,n49);
xor (n2500,n2321,n2325);
or (n2501,n2502,n2503,n2504);
and (n2502,n2472,n2473);
and (n2503,n2473,n2477);
and (n2504,n2472,n2477);
not (n2505,n2506);
not (n2506,n2507);
and (n2507,n2482,n2486);
not (n2508,n2509);
nor (n2509,n2510,n2525);
nor (n2510,n2511,n2515);
nand (n2511,n2512,n2513,n2514);
nand (n2512,n2488,n2492);
nand (n2513,n2494,n2492);
nand (n2514,n2488,n2494);
xor (n2515,n2516,n2523);
xor (n2516,n2517,n2519);
xor (n2517,n2518,n2330);
xor (n2518,n2316,n2320);
nand (n2519,n2520,n2521,n2522);
nand (n2520,n2496,n2500);
nand (n2521,n2501,n2500);
nand (n2522,n2496,n2501);
xor (n2523,n2524,n2280);
xor (n2524,n2263,n2264);
nor (n2525,n2526,n2530);
nand (n2526,n2527,n2528,n2529);
nand (n2527,n2517,n2519);
nand (n2528,n2523,n2519);
nand (n2529,n2517,n2523);
xor (n2530,n2531,n2294);
xor (n2531,n2249,n2261);
not (n2532,n2533);
nor (n2533,n2534,n2536);
nor (n2534,n2535,n2525);
nand (n2535,n2511,n2515);
not (n2536,n2537);
nand (n2537,n2526,n2530);
not (n2538,n2539);
nor (n2539,n2540,n2547);
nor (n2540,n2541,n2546);
nor (n2541,n2542,n2544);
nor (n2542,n2543,n2363);
nand (n2543,n2247,n2336);
not (n2544,n2545);
nand (n2545,n2364,n2368);
not (n2546,n2386);
not (n2547,n2548);
nor (n2548,n2549,n2551);
nor (n2549,n2550,n2402);
nand (n2550,n2388,n2392);
not (n2551,n2552);
nand (n2552,n2403,n2407);
nand (n2553,n2554,n2558);
nor (n2554,n2555,n2244);
nand (n2555,n2556,n2509);
nor (n2556,n2557,n2481);
nor (n2557,n2414,n2453);
or (n2558,n2559,n2581);
and (n2559,n2560,n2562);
xor (n2560,n2561,n2440);
xor (n2561,n2416,n2425);
or (n2562,n2563,n2577,n2580);
and (n2563,n2564,n2573);
and (n2564,n2565,n2569);
xnor (n2565,n2566,n347);
nor (n2566,n2567,n2568);
and (n2567,n727,n742);
and (n2568,n329,n744);
xnor (n2569,n2570,n222);
nor (n2570,n2571,n2572);
and (n2571,n733,n349);
and (n2572,n731,n345);
xnor (n2573,n2574,n123);
nor (n2574,n2575,n2576);
and (n2575,n756,n224);
and (n2576,n733,n220);
and (n2577,n2573,n2578);
xor (n2578,n2579,n2434);
xor (n2579,n2427,n2429);
and (n2580,n2564,n2578);
and (n2581,n2582,n2583);
xor (n2582,n2560,n2562);
or (n2583,n2584,n2599);
and (n2584,n2585,n2597);
or (n2585,n2586,n2591,n2596);
and (n2586,n2587,n2588);
xor (n2587,n2565,n2569);
and (n2588,n123,n2589);
xnor (n2589,n2590,n123);
nand (n2590,n770,n220);
and (n2591,n2588,n2592);
xnor (n2592,n2593,n123);
nor (n2593,n2594,n2595);
and (n2594,n770,n224);
and (n2595,n756,n220);
and (n2596,n2587,n2592);
xor (n2597,n2598,n2578);
xor (n2598,n2564,n2573);
and (n2599,n2600,n2601);
xor (n2600,n2585,n2597);
or (n2601,n2602,n2618);
and (n2602,n2603,n2605);
xor (n2603,n2604,n2592);
xor (n2604,n2587,n2588);
or (n2605,n2606,n2612,n2617);
and (n2606,n2607,n2608);
not (n2607,n2590);
xnor (n2608,n2609,n347);
nor (n2609,n2610,n2611);
and (n2610,n731,n742);
and (n2611,n727,n744);
and (n2612,n2608,n2613);
xnor (n2613,n2614,n222);
nor (n2614,n2615,n2616);
and (n2615,n756,n349);
and (n2616,n733,n345);
and (n2617,n2607,n2613);
and (n2618,n2619,n2620);
xor (n2619,n2603,n2605);
or (n2620,n2621,n2632);
and (n2621,n2622,n2624);
xor (n2622,n2623,n2613);
xor (n2623,n2607,n2608);
and (n2624,n2625,n2628);
and (n2625,n222,n2626);
xnor (n2626,n2627,n222);
nand (n2627,n770,n345);
xnor (n2628,n2629,n347);
nor (n2629,n2630,n2631);
and (n2630,n733,n742);
and (n2631,n731,n744);
and (n2632,n2633,n2634);
xor (n2633,n2622,n2624);
or (n2634,n2635,n2641);
and (n2635,n2636,n2640);
xnor (n2636,n2637,n222);
nor (n2637,n2638,n2639);
and (n2638,n770,n349);
and (n2639,n756,n345);
xor (n2640,n2625,n2628);
and (n2641,n2642,n2643);
xor (n2642,n2636,n2640);
or (n2643,n2644,n2650);
and (n2644,n2645,n2649);
xnor (n2645,n2646,n347);
nor (n2646,n2647,n2648);
and (n2647,n756,n742);
and (n2648,n733,n744);
not (n2649,n2627);
and (n2650,n2651,n2652);
xor (n2651,n2645,n2649);
and (n2652,n2653,n2657);
xnor (n2653,n2654,n347);
nor (n2654,n2655,n2656);
and (n2655,n770,n742);
and (n2656,n756,n744);
and (n2657,n2658,n347);
xnor (n2658,n2659,n347);
nand (n2659,n770,n744);
not (n2660,n2661);
nand (n2661,n2662,n1682);
nor (n2662,n2663,n714);
nand (n2663,n2664,n1637);
nor (n2664,n2665,n1609);
nor (n2665,n1392,n1571);
not (n2666,n2667);
nand (n2667,n2668,n560);
nor (n2668,n2669,n480);
nor (n2669,n7,n400);
nand (n2670,n2671,n2737);
not (n2671,n2672);
nor (n2672,n2673,n2733);
xor (n2673,n2674,n2729);
xor (n2674,n2675,n2709);
xor (n2675,n2676,n2705);
xor (n2676,n2677,n2691);
xor (n2677,n2678,n2687);
xor (n2678,n2679,n2683);
xor (n2679,n2680,n88);
or (n2680,n2681,n2682);
and (n2681,n43,n82);
and (n2682,n48,n86);
xor (n2683,n2684,n19);
or (n2684,n2685,n2686);
and (n2685,n56,n99);
and (n2686,n60,n102);
xor (n2687,n2688,n24);
or (n2688,n2689,n2690);
and (n2689,n31,n17);
and (n2690,n36,n22);
xor (n2691,n2692,n2701);
xor (n2692,n2693,n2697);
xor (n2693,n2694,n114);
or (n2694,n2695,n2696);
and (n2695,n72,n108);
and (n2696,n81,n112);
xor (n2697,n2698,n25);
or (n2698,n2699,n2700);
and (n2699,n85,n190);
and (n2700,n16,n194);
not (n2701,n2702);
xor (n2702,n2703,n39);
or (n2703,n657,n2704);
and (n2704,n147,n37);
nand (n2705,n2706,n2707,n2708);
nand (n2706,n675,n679);
nand (n2707,n25,n679);
nand (n2708,n675,n25);
xor (n2709,n2710,n2725);
xor (n2710,n2711,n2721);
xor (n2711,n2712,n2717);
xor (n2712,n25,n2713);
nand (n2713,n2714,n2715,n2716);
nand (n2714,n572,n655);
nand (n2715,n659,n655);
nand (n2716,n572,n659);
nand (n2717,n2718,n2719,n2720);
nand (n2718,n685,n573);
nand (n2719,n689,n573);
nand (n2720,n685,n689);
nand (n2721,n2722,n2723,n2724);
nand (n2722,n653,n663);
nand (n2723,n667,n663);
nand (n2724,n653,n667);
nand (n2725,n2726,n2727,n2728);
nand (n2726,n673,n683);
nand (n2727,n693,n683);
nand (n2728,n673,n693);
nand (n2729,n2730,n2731,n2732);
nand (n2730,n647,n651);
nand (n2731,n671,n651);
nand (n2732,n647,n671);
nand (n2733,n2734,n2735,n2736);
nand (n2734,n641,n645);
nand (n2735,n698,n645);
nand (n2736,n641,n698);
nand (n2737,n2673,n2733);
xor (n2738,n2739,n2866);
xnor (n2739,n2740,n2798);
xor (n2740,n2741,n2784);
xor (n2741,n2742,n2750);
xor (n2742,n2743,n2749);
xor (n2743,n2744,n2745);
not (n2744,n2706);
or (n2745,n2746,n2747,n2748);
not (n2746,n2714);
and (n2747,n655,n685);
and (n2748,n572,n685);
not (n2749,n2676);
or (n2750,n2751,n2772,n2783);
and (n2751,n2752,n2759);
xor (n2752,n2753,n2758);
xor (n2753,n663,n2754);
or (n2754,n2755,n2756,n2757);
and (n2755,n573,n576);
not (n2756,n669);
and (n2757,n573,n580);
xor (n2758,n654,n685);
or (n2759,n2760,n2766,n2771);
and (n2760,n599,n2761);
and (n2761,n2762,n521);
or (n2762,n2763,n2764,n2765);
and (n2763,n443,n434);
not (n2764,n518);
and (n2765,n443,n438);
and (n2766,n2761,n2767);
or (n2767,n2768,n2769,n2770);
not (n2768,n620);
and (n2769,n541,n509);
and (n2770,n537,n509);
and (n2771,n599,n2767);
and (n2772,n2759,n2773);
xor (n2773,n2774,n2781);
xor (n2774,n2775,n2776);
not (n2775,n648);
or (n2776,n2777,n2779,n2780);
and (n2777,n695,n2778);
not (n2778,n570);
and (n2779,n2778,n588);
not (n2780,n697);
xor (n2781,n2782,n674);
xor (n2782,n659,n689);
and (n2783,n2752,n2773);
xor (n2784,n2785,n2794);
xor (n2785,n2786,n2790);
or (n2786,n2787,n2788,n2789);
and (n2787,n659,n689);
and (n2788,n689,n674);
and (n2789,n659,n674);
or (n2790,n2791,n2792,n2793);
and (n2791,n663,n2754);
and (n2792,n2754,n2758);
and (n2793,n663,n2758);
or (n2794,n2795,n2796,n2797);
and (n2795,n2775,n2776);
and (n2796,n2776,n2781);
and (n2797,n2775,n2781);
or (n2798,n2799,n2830,n2865);
and (n2799,n2800,n2828);
or (n2800,n2801,n2810,n2827);
and (n2801,n2802,n2804);
xor (n2802,n2803,n588);
xor (n2803,n695,n2778);
or (n2804,n2805,n2807,n2809);
and (n2805,n2806,n499);
not (n2806,n490);
and (n2807,n499,n2808);
xor (n2808,n2762,n521);
and (n2809,n2806,n2808);
and (n2810,n2804,n2811);
or (n2811,n2812,n2823,n2826);
and (n2812,n2813,n2818);
or (n2813,n2814,n2816,n2817);
and (n2814,n454,n2815);
not (n2815,n432);
and (n2816,n2815,n419);
and (n2817,n454,n419);
or (n2818,n2819,n2821,n2822);
and (n2819,n468,n2820);
not (n2820,n415);
and (n2821,n2820,n428);
and (n2822,n468,n428);
and (n2823,n2818,n2824);
xor (n2824,n2825,n509);
xor (n2825,n537,n541);
and (n2826,n2813,n2824);
and (n2827,n2802,n2811);
xor (n2828,n2829,n2773);
xor (n2829,n2752,n2759);
and (n2830,n2828,n2831);
or (n2831,n2832,n2861,n2864);
and (n2832,n2833,n2835);
xor (n2833,n2834,n2767);
xor (n2834,n599,n2761);
or (n2835,n2836,n2857,n2860);
and (n2836,n2837,n2855);
or (n2837,n2838,n2851,n2854);
and (n2838,n2839,n2843);
or (n2839,n2840,n2841,n2842);
and (n2840,n13,n157);
and (n2841,n157,n242);
and (n2842,n13,n242);
or (n2843,n2844,n2845,n2850);
and (n2844,n26,n171);
and (n2845,n171,n2846);
or (n2846,n2847,n2848,n2849);
and (n2847,n144,n204);
not (n2848,n240);
and (n2849,n144,n200);
and (n2850,n26,n2846);
and (n2851,n2843,n2852);
xor (n2852,n2853,n419);
xor (n2853,n454,n2815);
and (n2854,n2839,n2852);
xor (n2855,n2856,n2808);
xor (n2856,n2806,n499);
and (n2857,n2855,n2858);
xor (n2858,n2859,n2824);
xor (n2859,n2813,n2818);
and (n2860,n2837,n2858);
and (n2861,n2835,n2862);
xor (n2862,n2863,n2811);
xor (n2863,n2802,n2804);
and (n2864,n2833,n2862);
and (n2865,n2800,n2831);
or (n2866,n2867,n2947);
and (n2867,n2868,n2870);
xor (n2868,n2869,n2831);
xor (n2869,n2800,n2828);
or (n2870,n2871,n2873);
xor (n2871,n2872,n2862);
xor (n2872,n2833,n2835);
or (n2873,n2874,n2897,n2946);
and (n2874,n2875,n2895);
or (n2875,n2876,n2891,n2894);
and (n2876,n2877,n2879);
xor (n2877,n2878,n428);
xor (n2878,n468,n2820);
or (n2879,n2880,n2887,n2890);
and (n2880,n141,n2881);
or (n2881,n2882,n2884,n2886);
and (n2882,n232,n2883);
not (n2883,n198);
and (n2884,n2883,n2885);
not (n2885,n180);
and (n2886,n232,n2885);
and (n2887,n2881,n2888);
xor (n2888,n2889,n242);
xor (n2889,n13,n157);
and (n2890,n141,n2888);
and (n2891,n2879,n2892);
xor (n2892,n2893,n2852);
xor (n2893,n2839,n2843);
and (n2894,n2877,n2892);
xor (n2895,n2896,n2858);
xor (n2896,n2837,n2855);
and (n2897,n2895,n2898);
or (n2898,n2899,n2910,n2945);
and (n2899,n2900,n2908);
or (n2900,n2901,n2904,n2907);
and (n2901,n2902,n64);
xor (n2902,n2903,n2846);
xor (n2903,n26,n171);
and (n2904,n64,n2905);
xor (n2905,n2906,n2888);
xor (n2906,n141,n2881);
and (n2907,n2902,n2905);
xor (n2908,n2909,n2892);
xor (n2909,n2877,n2879);
and (n2910,n2908,n2911);
or (n2911,n2912,n2941,n2944);
and (n2912,n2913,n2926);
or (n2913,n2914,n2924,n2925);
and (n2914,n2915,n277);
or (n2915,n2916,n2921,n2923);
and (n2916,n2917,n271);
or (n2917,n2918,n2919,n2920);
and (n2918,n216,n261);
not (n2919,n265);
and (n2920,n216,n266);
and (n2921,n271,n2922);
not (n2922,n274);
and (n2923,n2917,n2922);
not (n2924,n312);
and (n2925,n2915,n313);
or (n2926,n2927,n2934,n2940);
and (n2927,n2928,n2932);
or (n2928,n2929,n2930,n2931);
and (n2929,n217,n213);
not (n2930,n231);
and (n2931,n217,n227);
xor (n2932,n2933,n2885);
xor (n2933,n232,n2883);
and (n2934,n2932,n2935);
or (n2935,n2936,n2937,n2939);
and (n2936,n216,n354);
and (n2937,n354,n2938);
not (n2938,n2162);
and (n2939,n216,n2938);
and (n2940,n2928,n2935);
and (n2941,n2926,n2942);
xor (n2942,n2943,n2905);
xor (n2943,n2902,n64);
and (n2944,n2913,n2942);
and (n2945,n2900,n2911);
and (n2946,n2875,n2898);
and (n2947,n2948,n2949);
xor (n2948,n2868,n2870);
and (n2949,n2950,n2951);
xnor (n2950,n2871,n2873);
or (n2951,n2952,n3037);
and (n2952,n2953,n2955);
xor (n2953,n2954,n2898);
xor (n2954,n2875,n2895);
or (n2955,n2956,n2958);
xor (n2956,n2957,n2911);
xor (n2957,n2900,n2908);
or (n2958,n2959,n2981,n3036);
and (n2959,n2960,n2979);
or (n2960,n2961,n2975,n2978);
and (n2961,n2962,n2964);
xor (n2962,n2963,n313);
xor (n2963,n2915,n277);
or (n2964,n2965,n2968,n2974);
and (n2965,n2966,n2165);
xor (n2966,n2967,n2922);
xor (n2967,n2917,n271);
and (n2968,n2165,n2969);
or (n2969,n2970,n2971,n2973);
not (n2970,n393);
and (n2971,n377,n2972);
not (n2972,n374);
and (n2973,n358,n2972);
and (n2974,n2966,n2969);
and (n2975,n2964,n2976);
xor (n2976,n2977,n2935);
xor (n2977,n2928,n2932);
and (n2978,n2962,n2976);
xor (n2979,n2980,n2942);
xor (n2980,n2913,n2926);
and (n2981,n2979,n2982);
or (n2982,n2983,n2998,n3035);
and (n2983,n2984,n2996);
or (n2984,n2985,n2992,n2995);
and (n2985,n2986,n2990);
or (n2986,n2987,n2988,n2989);
and (n2987,n325,n2135);
and (n2988,n2135,n2116);
and (n2989,n325,n2116);
xor (n2990,n2991,n2938);
xor (n2991,n216,n354);
and (n2992,n2990,n2993);
and (n2993,n2111,n2994);
not (n2994,n2109);
and (n2995,n2986,n2993);
xor (n2996,n2997,n2976);
xor (n2997,n2962,n2964);
and (n2998,n2996,n2999);
or (n2999,n3000,n3020,n3034);
and (n3000,n3001,n3018);
or (n3001,n3002,n3007,n3017);
and (n3002,n3003,n2138);
or (n3003,n3004,n3005,n3006);
and (n3004,n342,n333);
not (n3005,n332);
and (n3006,n342,n336);
and (n3007,n2138,n3008);
or (n3008,n3009,n3014,n3016);
and (n3009,n341,n3010);
or (n3010,n3011,n3012,n3013);
and (n3011,n341,n1939);
not (n3012,n2053);
and (n3013,n341,n1943);
and (n3014,n3010,n3015);
not (n3015,n2048);
and (n3016,n341,n3015);
and (n3017,n3003,n3008);
xor (n3018,n3019,n2969);
xor (n3019,n2966,n2165);
and (n3020,n3018,n3021);
or (n3021,n3022,n3026,n3033);
and (n3022,n3023,n3025);
xor (n3023,n3024,n2116);
xor (n3024,n325,n2135);
not (n3025,n2108);
and (n3026,n3025,n3027);
or (n3027,n3028,n3031,n3032);
and (n3028,n3029,n2054);
and (n3029,n1923,n3030);
not (n3030,n1937);
and (n3031,n2054,n2076);
and (n3032,n3029,n2076);
and (n3033,n3023,n3027);
and (n3034,n3001,n3021);
and (n3035,n2984,n2999);
and (n3036,n2960,n2982);
and (n3037,n3038,n3039);
xor (n3038,n2953,n2955);
and (n3039,n3040,n3041);
xnor (n3040,n2956,n2958);
or (n3041,n3042,n3246);
and (n3042,n3043,n3045);
xor (n3043,n3044,n2982);
xor (n3044,n2960,n2979);
or (n3045,n3046,n3121,n3245);
and (n3046,n3047,n3119);
or (n3047,n3048,n3115,n3118);
and (n3048,n3049,n3051);
xor (n3049,n3050,n2993);
xor (n3050,n2986,n2990);
or (n3051,n3052,n3086,n3114);
and (n3052,n3053,n3084);
or (n3053,n3054,n3072,n3083);
and (n3054,n3055,n3064);
and (n3055,n3056,n1963);
or (n3056,n3057,n3062,n3063);
and (n3057,n3058,n1833);
or (n3058,n3059,n3060,n3061);
and (n3059,n1902,n1698);
not (n3060,n1842);
and (n3061,n1902,n1702);
not (n3062,n1975);
and (n3063,n3058,n1837);
or (n3064,n3065,n3070,n3071);
and (n3065,n2003,n3066);
or (n3066,n3067,n3068,n3069);
and (n3067,n1902,n1822);
not (n3068,n1950);
and (n3069,n1902,n1827);
and (n3070,n3066,n1984);
and (n3071,n2003,n1984);
and (n3072,n3064,n3073);
or (n3073,n3074,n3080,n3082);
and (n3074,n3075,n3076);
not (n3075,n1922);
or (n3076,n3077,n3078,n3079);
and (n3077,n1706,n1898);
not (n3078,n2002);
and (n3079,n1706,n1903);
and (n3080,n3076,n3081);
not (n3081,n1979);
and (n3082,n3075,n3081);
and (n3083,n3055,n3073);
xor (n3084,n3085,n3008);
xor (n3085,n3003,n2138);
and (n3086,n3084,n3087);
or (n3087,n3088,n3110,n3113);
and (n3088,n3089,n3091);
xor (n3089,n3090,n3015);
xor (n3090,n341,n3010);
or (n3091,n3092,n3101,n3109);
and (n3092,n3093,n3100);
or (n3093,n3094,n3096,n3099);
and (n3094,n1882,n3095);
not (n3095,n1879);
and (n3096,n3095,n3097);
xor (n3097,n3098,n1827);
xor (n3098,n1902,n1822);
and (n3099,n1882,n3097);
xor (n3100,n3056,n1963);
and (n3101,n3100,n3102);
or (n3102,n3103,n3107,n3108);
and (n3103,n3104,n3105);
not (n3104,n1896);
xor (n3105,n3106,n1837);
xor (n3106,n3058,n1833);
and (n3107,n3105,n1856);
and (n3108,n3104,n1856);
and (n3109,n3093,n3102);
and (n3110,n3091,n3111);
xor (n3111,n3112,n2076);
xor (n3112,n3029,n2054);
and (n3113,n3089,n3111);
and (n3114,n3053,n3087);
and (n3115,n3051,n3116);
xor (n3116,n3117,n3021);
xor (n3117,n3001,n3018);
and (n3118,n3049,n3116);
xor (n3119,n3120,n2999);
xor (n3120,n2984,n2996);
and (n3121,n3119,n3122);
or (n3122,n3123,n3156,n3244);
and (n3123,n3124,n3154);
or (n3124,n3125,n3150,n3153);
and (n3125,n3126,n3128);
xor (n3126,n3127,n3027);
xor (n3127,n3023,n3025);
or (n3128,n3129,n3146,n3149);
and (n3129,n3130,n3132);
xor (n3130,n3131,n3073);
xor (n3131,n3055,n3064);
or (n3132,n3133,n3138,n3145);
and (n3133,n3134,n3136);
xor (n3134,n3135,n1984);
xor (n3135,n2003,n3066);
xor (n3136,n3137,n3081);
xor (n3137,n3075,n3076);
and (n3138,n3136,n3139);
and (n3139,n1847,n3140);
or (n3140,n3141,n3142,n3144);
not (n3141,n1853);
and (n3142,n1713,n3143);
not (n3143,n1696);
and (n3144,n1709,n3143);
and (n3145,n3134,n3139);
and (n3146,n3132,n3147);
xor (n3147,n3148,n3111);
xor (n3148,n3089,n3091);
and (n3149,n3130,n3147);
and (n3150,n3128,n3151);
xor (n3151,n3152,n3087);
xor (n3152,n3053,n3084);
and (n3153,n3126,n3151);
xor (n3154,n3155,n3116);
xor (n3155,n3049,n3051);
and (n3156,n3154,n3157);
or (n3157,n3158,n3215,n3243);
and (n3158,n3159,n3161);
xor (n3159,n3160,n3151);
xor (n3160,n3126,n3128);
or (n3161,n3162,n3194,n3214);
and (n3162,n3163,n3192);
or (n3163,n3164,n3177,n3191);
and (n3164,n3165,n3175);
or (n3165,n3166,n3173,n3174);
and (n3166,n3167,n3171);
or (n3167,n3168,n3169,n3170);
and (n3168,n1761,n1746);
and (n3169,n1746,n1729);
and (n3170,n1761,n1729);
xor (n3171,n3172,n3097);
xor (n3172,n1882,n3095);
and (n3173,n3171,n1907);
and (n3174,n3167,n1907);
xor (n3175,n3176,n3102);
xor (n3176,n3093,n3100);
and (n3177,n3175,n3178);
or (n3178,n3179,n3188,n3190);
and (n3179,n3180,n3186);
or (n3180,n3181,n3182,n3185);
and (n3181,n1751,n1745);
and (n3182,n1745,n3183);
xor (n3183,n3184,n1729);
xor (n3184,n1761,n1746);
and (n3185,n1751,n3183);
xor (n3186,n3187,n1856);
xor (n3187,n3104,n3105);
and (n3188,n3186,n3189);
xor (n3189,n1847,n3140);
and (n3190,n3180,n3189);
and (n3191,n3165,n3178);
xor (n3192,n3193,n3147);
xor (n3193,n3130,n3132);
and (n3194,n3192,n3195);
or (n3195,n3196,n3210,n3213);
and (n3196,n3197,n3199);
xor (n3197,n3198,n3139);
xor (n3198,n3134,n3136);
or (n3199,n3200,n3208,n3209);
and (n3200,n3201,n3203);
xor (n3201,n3202,n1907);
xor (n3202,n3167,n3171);
or (n3203,n3204,n3205,n3207);
not (n3204,n1806);
and (n3205,n1721,n3206);
not (n3206,n1694);
and (n3207,n1717,n3206);
and (n3208,n3203,n1808);
and (n3209,n3201,n1808);
and (n3210,n3199,n3211);
xor (n3211,n3212,n3178);
xor (n3212,n3165,n3175);
and (n3213,n3197,n3211);
and (n3214,n3163,n3195);
and (n3215,n3161,n3216);
or (n3216,n3217,n3219);
xor (n3217,n3218,n3195);
xor (n3218,n3163,n3192);
or (n3219,n3220,n3236,n3242);
and (n3220,n3221,n3234);
or (n3221,n3222,n3230,n3233);
and (n3222,n3223,n3225);
xor (n3223,n3224,n3189);
xor (n3224,n3180,n3186);
or (n3225,n3226,n3228,n3229);
and (n3226,n3227,n1793);
not (n3227,n1692);
not (n3228,n1800);
and (n3229,n3227,n1725);
and (n3230,n3225,n3231);
xor (n3231,n3232,n1808);
xor (n3232,n3201,n3203);
and (n3233,n3223,n3231);
xor (n3234,n3235,n3211);
xor (n3235,n3197,n3199);
and (n3236,n3234,n3237);
or (n3237,n3238,n3240);
or (n3238,n1686,n3239);
not (n3239,n1690);
xor (n3240,n3241,n3231);
xor (n3241,n3223,n3225);
and (n3242,n3221,n3237);
and (n3243,n3159,n3216);
and (n3244,n3124,n3157);
and (n3245,n3047,n3122);
and (n3246,n3247,n3248);
xor (n3247,n3043,n3045);
and (n3248,n3249,n3251);
xor (n3249,n3250,n3122);
xor (n3250,n3047,n3119);
or (n3251,n3252,n3254);
xor (n3252,n3253,n3157);
xor (n3253,n3124,n3154);
and (n3254,n3255,n3256);
not (n3255,n3252);
and (n3256,n3257,n3259);
xor (n3257,n3258,n3216);
xor (n3258,n3159,n3161);
and (n3259,n3260,n3261);
xnor (n3260,n3217,n3219);
and (n3261,n3262,n3264);
xor (n3262,n3263,n3237);
xor (n3263,n3221,n3234);
and (n3264,n3265,n3266);
xnor (n3265,n3238,n3240);
and (n3266,n3267,n3270);
not (n3267,n3268);
nand (n3268,n3269,n2215);
not (n3269,n1685);
nand (n3270,n712,n3271);
nand (n3271,n2662,n2241);
endmodule
