module top (out,n20,n22,n27,n33,n39,n48,n50,n57,n66
        ,n74,n75,n83,n89,n96,n102,n111,n118,n133,n138
        ,n144,n161,n187,n196,n251,n380,n454,n518,n564,n591);
output out;
input n20;
input n22;
input n27;
input n33;
input n39;
input n48;
input n50;
input n57;
input n66;
input n74;
input n75;
input n83;
input n89;
input n96;
input n102;
input n111;
input n118;
input n133;
input n138;
input n144;
input n161;
input n187;
input n196;
input n251;
input n380;
input n454;
input n518;
input n564;
input n591;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n21;
wire n23;
wire n24;
wire n25;
wire n26;
wire n28;
wire n29;
wire n30;
wire n31;
wire n32;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n49;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n134;
wire n135;
wire n136;
wire n137;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
xor (out,n0,n1171);
nand (n0,n1,n1170);
or (n1,n2,n352);
not (n2,n3);
nand (n3,n4,n350);
nand (n4,n5,n301);
not (n5,n6);
or (n6,n7,n300);
and (n7,n8,n237);
xor (n8,n9,n156);
xor (n9,n10,n120);
xor (n10,n11,n93);
or (n11,n12,n92);
and (n12,n13,n68);
xor (n13,n14,n42);
nand (n14,n15,n35);
or (n15,n16,n24);
not (n16,n17);
nor (n17,n18,n23);
and (n18,n19,n21);
not (n19,n20);
not (n21,n22);
and (n23,n22,n20);
nand (n24,n25,n29);
nand (n25,n26,n28);
or (n26,n27,n21);
nand (n28,n21,n27);
not (n29,n30);
nand (n30,n31,n34);
or (n31,n32,n27);
not (n32,n33);
nand (n34,n32,n27);
nand (n35,n36,n30);
not (n36,n37);
nor (n37,n38,n40);
and (n38,n21,n39);
and (n40,n22,n41);
not (n41,n39);
nand (n42,n43,n62);
or (n43,n44,n52);
not (n44,n45);
nor (n45,n46,n51);
and (n46,n47,n49);
not (n47,n48);
not (n49,n50);
and (n51,n50,n48);
not (n52,n53);
and (n53,n54,n59);
not (n54,n55);
nand (n55,n56,n58);
or (n56,n57,n21);
nand (n58,n57,n21);
nand (n59,n60,n61);
or (n60,n57,n49);
nand (n61,n49,n57);
nand (n62,n55,n63);
nand (n63,n64,n67);
or (n64,n50,n65);
not (n65,n66);
or (n67,n49,n66);
nand (n68,n69,n86);
or (n69,n70,n81);
nand (n70,n71,n78);
nor (n71,n72,n76);
and (n72,n73,n75);
not (n73,n74);
and (n76,n74,n77);
not (n77,n75);
nand (n78,n79,n80);
or (n79,n75,n32);
nand (n80,n32,n75);
nor (n81,n82,n84);
and (n82,n32,n83);
and (n84,n33,n85);
not (n85,n83);
or (n86,n71,n87);
nor (n87,n88,n90);
and (n88,n32,n89);
and (n90,n33,n91);
not (n91,n89);
and (n92,n14,n42);
nand (n93,n94,n97);
not (n94,n95);
not (n95,n96);
nor (n97,n98,n113);
and (n98,n99,n108);
nor (n99,n100,n104);
nand (n100,n101,n103);
or (n101,n95,n102);
nand (n103,n95,n102);
nor (n104,n105,n106);
and (n105,n73,n102);
and (n106,n74,n107);
not (n107,n102);
nor (n108,n109,n112);
and (n109,n110,n73);
not (n110,n111);
and (n112,n74,n111);
nor (n113,n114,n115);
not (n114,n100);
nor (n115,n116,n119);
and (n116,n117,n74);
not (n117,n118);
and (n119,n118,n73);
xor (n120,n121,n152);
xor (n121,n122,n129);
nand (n122,n123,n125);
or (n123,n124,n52);
not (n124,n63);
nand (n125,n55,n126);
nor (n126,n127,n128);
and (n127,n19,n49);
and (n128,n50,n20);
nand (n129,n130,n139);
or (n130,n131,n136);
nor (n131,n132,n134);
and (n132,n49,n133);
and (n134,n50,n135);
not (n135,n133);
not (n136,n137);
xor (n137,n48,n138);
nand (n139,n140,n147);
not (n140,n141);
nor (n141,n142,n145);
and (n142,n143,n144);
not (n143,n138);
and (n145,n138,n146);
not (n146,n144);
not (n147,n148);
nand (n148,n131,n149);
nand (n149,n150,n151);
or (n150,n135,n138);
nand (n151,n135,n138);
nand (n152,n153,n155);
or (n153,n154,n115);
not (n154,n99);
or (n155,n114,n73);
xor (n156,n157,n206);
xor (n157,n158,n178);
xor (n158,n159,n169);
xor (n159,n160,n162);
and (n160,n138,n161);
nand (n162,n163,n164);
or (n163,n24,n37);
or (n164,n29,n165);
not (n165,n166);
nor (n166,n167,n168);
and (n167,n22,n83);
and (n168,n85,n21);
not (n169,n170);
nand (n170,n171,n172);
or (n171,n87,n70);
nand (n172,n173,n177);
not (n173,n174);
nor (n174,n175,n176);
and (n175,n110,n33);
and (n176,n111,n32);
not (n177,n71);
or (n178,n179,n205);
and (n179,n180,n188);
xor (n180,n181,n186);
nand (n181,n182,n185);
or (n182,n148,n183);
not (n183,n184);
xor (n184,n161,n138);
or (n185,n131,n141);
and (n186,n138,n187);
and (n188,n189,n198);
nand (n189,n190,n197);
or (n190,n191,n194);
nor (n191,n192,n193);
and (n192,n95,n118);
and (n193,n96,n117);
nand (n194,n96,n195);
not (n195,n196);
or (n197,n95,n195);
nand (n198,n199,n204);
or (n199,n200,n154);
not (n200,n201);
nor (n201,n202,n203);
and (n202,n74,n89);
and (n203,n91,n73);
nand (n204,n100,n108);
and (n205,n181,n186);
or (n206,n207,n236);
and (n207,n208,n235);
xor (n208,n209,n233);
or (n209,n210,n232);
and (n210,n211,n226);
xor (n211,n212,n219);
nand (n212,n213,n218);
or (n213,n214,n24);
not (n214,n215);
nor (n215,n216,n217);
and (n216,n65,n21);
and (n217,n22,n66);
nand (n218,n30,n17);
nand (n219,n220,n225);
or (n220,n221,n52);
not (n221,n222);
nand (n222,n223,n224);
or (n223,n50,n146);
or (n224,n49,n144);
nand (n225,n55,n45);
nand (n226,n227,n231);
or (n227,n70,n228);
nor (n228,n229,n230);
and (n229,n32,n39);
and (n230,n33,n41);
or (n231,n81,n71);
and (n232,n212,n219);
nand (n233,n234,n93);
or (n234,n94,n97);
xor (n235,n13,n68);
and (n236,n209,n233);
or (n237,n238,n299);
and (n238,n239,n254);
xor (n239,n240,n241);
xor (n240,n180,n188);
or (n241,n242,n253);
and (n242,n243,n252);
xor (n243,n244,n250);
nand (n244,n245,n248);
or (n245,n246,n148);
not (n246,n247);
xor (n247,n187,n138);
nand (n248,n249,n184);
not (n249,n131);
and (n250,n138,n251);
xor (n252,n189,n198);
and (n253,n244,n250);
or (n254,n255,n298);
and (n255,n256,n297);
xor (n256,n257,n272);
and (n257,n258,n265);
nand (n258,n259,n264);
or (n259,n194,n260);
not (n260,n261);
nor (n261,n262,n263);
and (n262,n111,n96);
and (n263,n110,n95);
or (n264,n191,n195);
nand (n265,n266,n271);
or (n266,n267,n154);
not (n267,n268);
nand (n268,n269,n270);
or (n269,n74,n85);
or (n270,n73,n83);
nand (n271,n100,n201);
or (n272,n273,n296);
and (n273,n274,n290);
xor (n274,n275,n282);
nand (n275,n276,n281);
or (n276,n277,n24);
not (n277,n278);
nor (n278,n279,n280);
and (n279,n47,n21);
and (n280,n48,n22);
nand (n281,n30,n215);
nand (n282,n283,n289);
or (n283,n284,n52);
not (n284,n285);
nor (n285,n286,n288);
and (n286,n287,n49);
not (n287,n161);
and (n288,n161,n50);
nand (n289,n55,n222);
nand (n290,n291,n295);
or (n291,n70,n292);
nor (n292,n293,n294);
and (n293,n32,n20);
and (n294,n33,n19);
or (n295,n71,n228);
and (n296,n275,n282);
xor (n297,n211,n226);
and (n298,n257,n272);
and (n299,n240,n241);
and (n300,n9,n156);
not (n301,n302);
xor (n302,n303,n347);
xor (n303,n304,n307);
or (n304,n305,n306);
and (n305,n10,n120);
and (n306,n11,n93);
xor (n307,n308,n329);
xor (n308,n309,n326);
xor (n309,n310,n319);
xor (n310,n311,n313);
nand (n311,n312,n74);
or (n312,n99,n100);
nand (n313,n314,n315);
or (n314,n70,n174);
or (n315,n71,n316);
nor (n316,n317,n318);
and (n317,n32,n118);
and (n318,n33,n117);
nand (n319,n320,n322);
or (n320,n52,n321);
not (n321,n126);
or (n322,n54,n323);
nor (n323,n324,n325);
and (n324,n49,n39);
and (n325,n41,n50);
or (n326,n327,n328);
and (n327,n159,n169);
and (n328,n160,n162);
xor (n329,n330,n334);
xor (n330,n170,n331);
or (n331,n332,n333);
and (n332,n121,n152);
and (n333,n122,n129);
xor (n334,n335,n346);
xor (n335,n336,n340);
nand (n336,n337,n338);
or (n337,n136,n148);
nand (n338,n249,n339);
xor (n339,n66,n138);
nand (n340,n341,n342);
or (n341,n165,n24);
nand (n342,n30,n343);
nor (n343,n344,n345);
and (n344,n91,n21);
and (n345,n22,n89);
and (n346,n138,n144);
or (n347,n348,n349);
and (n348,n157,n206);
and (n349,n158,n178);
not (n350,n351);
nor (n351,n5,n301);
not (n352,n353);
nand (n353,n354,n1156);
or (n354,n355,n639);
not (n355,n356);
and (n356,n357,n431,n500);
not (n357,n358);
nor (n358,n359,n360);
xor (n359,n8,n237);
or (n360,n361,n430);
and (n361,n362,n365);
xor (n362,n363,n364);
xor (n363,n208,n235);
xor (n364,n239,n254);
or (n365,n366,n429);
and (n366,n367,n383);
xor (n367,n368,n369);
xor (n368,n243,n252);
or (n369,n370,n382);
and (n370,n371,n381);
xor (n371,n372,n379);
nand (n372,n373,n378);
or (n373,n374,n148);
nor (n374,n375,n376);
and (n375,n251,n143);
and (n376,n138,n377);
not (n377,n251);
nand (n378,n249,n247);
and (n379,n138,n380);
xor (n381,n258,n265);
and (n382,n372,n379);
or (n383,n384,n428);
and (n384,n385,n427);
xor (n385,n386,n402);
and (n386,n387,n395);
nand (n387,n388,n389);
or (n388,n195,n260);
nand (n389,n390,n394);
not (n390,n391);
nor (n391,n392,n393);
and (n392,n95,n89);
and (n393,n96,n91);
not (n394,n194);
nand (n395,n396,n397);
or (n396,n114,n267);
nand (n397,n398,n99);
not (n398,n399);
nor (n399,n400,n401);
and (n400,n73,n39);
and (n401,n74,n41);
or (n402,n403,n426);
and (n403,n404,n420);
xor (n404,n405,n412);
nand (n405,n406,n411);
or (n406,n407,n24);
not (n407,n408);
nor (n408,n409,n410);
and (n409,n146,n21);
and (n410,n22,n144);
nand (n411,n278,n30);
nand (n412,n413,n419);
or (n413,n414,n52);
not (n414,n415);
nand (n415,n416,n418);
or (n416,n50,n417);
not (n417,n187);
or (n418,n49,n187);
nand (n419,n55,n285);
nand (n420,n421,n425);
or (n421,n70,n422);
nor (n422,n423,n424);
and (n423,n66,n32);
and (n424,n33,n65);
or (n425,n292,n71);
and (n426,n405,n412);
xor (n427,n274,n290);
and (n428,n386,n402);
and (n429,n368,n369);
and (n430,n363,n364);
not (n431,n432);
nor (n432,n433,n434);
xor (n433,n362,n365);
or (n434,n435,n499);
and (n435,n436,n439);
xor (n436,n437,n438);
xor (n437,n256,n297);
xor (n438,n367,n383);
or (n439,n440,n498);
and (n440,n441,n457);
xor (n441,n442,n443);
xor (n442,n371,n381);
or (n443,n444,n456);
and (n444,n445,n455);
xor (n445,n446,n453);
nand (n446,n447,n452);
or (n447,n148,n448);
nor (n448,n449,n450);
and (n449,n380,n143);
and (n450,n138,n451);
not (n451,n380);
or (n452,n374,n131);
and (n453,n138,n454);
xor (n455,n387,n395);
and (n456,n446,n453);
or (n457,n458,n497);
and (n458,n459,n496);
xor (n459,n460,n473);
and (n460,n461,n467);
nand (n461,n462,n466);
or (n462,n194,n463);
nor (n463,n464,n465);
and (n464,n95,n83);
and (n465,n96,n85);
or (n466,n391,n195);
nand (n467,n468,n472);
or (n468,n154,n469);
nor (n469,n470,n471);
and (n470,n73,n20);
and (n471,n74,n19);
or (n472,n114,n399);
or (n473,n474,n495);
and (n474,n475,n489);
xor (n475,n476,n483);
nand (n476,n477,n482);
or (n477,n478,n24);
not (n478,n479);
nor (n479,n480,n481);
and (n480,n287,n21);
and (n481,n22,n161);
nand (n482,n30,n408);
nand (n483,n484,n488);
or (n484,n52,n485);
nor (n485,n486,n487);
and (n486,n49,n251);
and (n487,n50,n377);
nand (n488,n55,n415);
nand (n489,n490,n494);
or (n490,n70,n491);
nor (n491,n492,n493);
and (n492,n48,n32);
and (n493,n33,n47);
or (n494,n71,n422);
and (n495,n476,n483);
xor (n496,n404,n420);
and (n497,n460,n473);
and (n498,n442,n443);
and (n499,n437,n438);
nor (n500,n501,n634);
nor (n501,n502,n568);
xor (n502,n503,n567);
xor (n503,n504,n505);
xor (n504,n385,n427);
or (n505,n506,n566);
and (n506,n507,n521);
xor (n507,n508,n509);
xor (n508,n445,n455);
or (n509,n510,n520);
and (n510,n511,n519);
xor (n511,n512,n517);
nand (n512,n513,n516);
or (n513,n514,n148);
not (n514,n515);
xor (n515,n454,n138);
or (n516,n131,n448);
and (n517,n138,n518);
xor (n519,n461,n467);
and (n520,n512,n517);
and (n521,n522,n546);
or (n522,n523,n545);
and (n523,n524,n539);
xor (n524,n525,n533);
nand (n525,n526,n531);
or (n526,n527,n154);
not (n527,n528);
nand (n528,n529,n530);
or (n529,n74,n65);
or (n530,n73,n66);
nand (n531,n532,n100);
not (n532,n469);
nand (n533,n534,n538);
or (n534,n24,n535);
nor (n535,n536,n537);
and (n536,n21,n187);
and (n537,n22,n417);
or (n538,n29,n478);
nand (n539,n540,n544);
or (n540,n52,n541);
nor (n541,n542,n543);
and (n542,n49,n380);
and (n543,n50,n451);
or (n544,n54,n485);
and (n545,n525,n533);
or (n546,n547,n565);
and (n547,n548,n563);
xor (n548,n549,n555);
nand (n549,n550,n554);
or (n550,n70,n551);
nor (n551,n552,n553);
and (n552,n32,n144);
and (n553,n33,n146);
or (n554,n491,n71);
nand (n555,n556,n557);
or (n556,n514,n131);
nand (n557,n558,n147);
not (n558,n559);
nor (n559,n560,n561);
and (n560,n518,n143);
and (n561,n562,n138);
not (n562,n518);
and (n563,n138,n564);
and (n565,n549,n555);
and (n566,n508,n509);
xor (n567,n441,n457);
or (n568,n569,n633);
and (n569,n570,n573);
xor (n570,n571,n572);
xor (n571,n459,n496);
xor (n572,n507,n521);
or (n573,n574,n632);
and (n574,n575,n578);
xor (n575,n576,n577);
xor (n576,n475,n489);
xor (n577,n511,n519);
or (n578,n579,n631);
and (n579,n580,n605);
xor (n580,n581,n587);
nand (n581,n582,n586);
or (n582,n194,n583);
nor (n583,n584,n585);
and (n584,n95,n39);
and (n585,n96,n41);
or (n586,n463,n195);
or (n587,n588,n604);
and (n588,n589,n598);
xor (n589,n590,n592);
and (n590,n138,n591);
nand (n592,n593,n594);
or (n593,n114,n527);
nand (n594,n99,n595);
nand (n595,n596,n597);
or (n596,n74,n47);
or (n597,n73,n48);
nand (n598,n599,n603);
or (n599,n24,n600);
nor (n600,n601,n602);
and (n601,n21,n251);
and (n602,n22,n377);
or (n603,n535,n29);
and (n604,n590,n592);
or (n605,n606,n630);
and (n606,n607,n623);
xor (n607,n608,n617);
nand (n608,n609,n615);
or (n609,n610,n52);
not (n610,n611);
nor (n611,n612,n614);
and (n612,n613,n49);
not (n613,n454);
and (n614,n50,n454);
nand (n615,n616,n55);
not (n616,n541);
nand (n617,n618,n622);
or (n618,n619,n194);
nor (n619,n620,n621);
and (n620,n95,n20);
and (n621,n96,n19);
or (n622,n583,n195);
nand (n623,n624,n629);
or (n624,n148,n625);
nor (n625,n626,n627);
and (n626,n143,n564);
and (n627,n138,n628);
not (n628,n564);
or (n629,n131,n559);
and (n630,n608,n617);
and (n631,n581,n587);
and (n632,n576,n577);
and (n633,n571,n572);
nor (n634,n635,n636);
xor (n635,n436,n439);
or (n636,n637,n638);
and (n637,n503,n567);
and (n638,n504,n505);
not (n639,n640);
nand (n640,n641,n863);
not (n641,n642);
nand (n642,n643,n856);
or (n643,n644,n834);
not (n644,n645);
nand (n645,n646,n833);
or (n646,n647,n782);
nor (n647,n648,n728);
xor (n648,n649,n694);
xor (n649,n650,n651);
xor (n650,n580,n605);
or (n651,n652,n693);
and (n652,n653,n656);
xor (n653,n654,n655);
xor (n654,n607,n623);
xor (n655,n589,n598);
or (n656,n657,n692);
and (n657,n658,n675);
xor (n658,n659,n666);
nand (n659,n660,n665);
or (n660,n148,n661);
nor (n661,n662,n663);
and (n662,n591,n143);
and (n663,n664,n138);
not (n664,n591);
or (n665,n131,n625);
nand (n666,n667,n671);
or (n667,n70,n668);
nor (n668,n669,n670);
and (n669,n32,n187);
and (n670,n33,n417);
or (n671,n71,n672);
nor (n672,n673,n674);
and (n673,n32,n161);
and (n674,n33,n287);
nand (n675,n676,n691);
or (n676,n677,n683);
not (n677,n678);
nand (n678,n679,n138);
nand (n679,n680,n681);
or (n680,n50,n133);
nand (n681,n682,n664);
or (n682,n135,n49);
not (n683,n684);
nand (n684,n685,n690);
or (n685,n686,n154);
not (n686,n687);
nand (n687,n688,n689);
or (n688,n74,n146);
or (n689,n73,n144);
nand (n690,n100,n595);
or (n691,n684,n678);
and (n692,n659,n666);
and (n693,n654,n655);
xor (n694,n695,n698);
xor (n695,n696,n697);
xor (n696,n548,n563);
xor (n697,n524,n539);
or (n698,n699,n727);
and (n699,n700,n705);
xor (n700,n701,n704);
nand (n701,n702,n703);
or (n702,n70,n672);
or (n703,n71,n551);
nor (n704,n683,n678);
or (n705,n706,n726);
and (n706,n707,n720);
xor (n707,n708,n714);
nand (n708,n709,n713);
or (n709,n24,n710);
nor (n710,n711,n712);
and (n711,n21,n380);
and (n712,n22,n451);
or (n713,n29,n600);
nand (n714,n715,n719);
or (n715,n52,n716);
nor (n716,n717,n718);
and (n717,n49,n518);
and (n718,n50,n562);
or (n719,n54,n610);
nand (n720,n721,n725);
or (n721,n722,n194);
nor (n722,n723,n724);
and (n723,n95,n66);
and (n724,n96,n65);
or (n725,n619,n195);
and (n726,n708,n714);
and (n727,n701,n704);
or (n728,n729,n781);
and (n729,n730,n780);
xor (n730,n731,n732);
xor (n731,n700,n705);
or (n732,n733,n779);
and (n733,n734,n778);
xor (n734,n735,n754);
or (n735,n736,n753);
and (n736,n737,n745);
xor (n737,n738,n739);
nor (n738,n131,n664);
nand (n739,n740,n744);
or (n740,n741,n154);
nor (n741,n742,n743);
and (n742,n287,n74);
and (n743,n161,n73);
nand (n744,n687,n100);
nand (n745,n746,n751);
or (n746,n747,n24);
not (n747,n748);
nand (n748,n749,n750);
or (n749,n22,n613);
or (n750,n21,n454);
nand (n751,n752,n30);
not (n752,n710);
and (n753,n738,n739);
or (n754,n755,n777);
and (n755,n756,n771);
xor (n756,n757,n765);
nand (n757,n758,n763);
or (n758,n759,n52);
not (n759,n760);
nand (n760,n761,n762);
or (n761,n50,n628);
or (n762,n49,n564);
nand (n763,n764,n55);
not (n764,n716);
nand (n765,n766,n770);
or (n766,n767,n194);
nor (n767,n768,n769);
and (n768,n95,n48);
and (n769,n96,n47);
or (n770,n722,n195);
nand (n771,n772,n776);
or (n772,n70,n773);
nor (n773,n774,n775);
and (n774,n32,n251);
and (n775,n33,n377);
or (n776,n71,n668);
and (n777,n757,n765);
xor (n778,n707,n720);
and (n779,n735,n754);
xor (n780,n653,n656);
and (n781,n731,n732);
nand (n782,n783,n784);
xor (n783,n730,n780);
or (n784,n785,n832);
and (n785,n786,n789);
xor (n786,n787,n788);
xor (n787,n658,n675);
xor (n788,n734,n778);
or (n789,n790,n831);
and (n790,n791,n830);
xor (n791,n792,n806);
and (n792,n793,n799);
and (n793,n794,n50);
nand (n794,n795,n796);
or (n795,n22,n57);
nand (n796,n797,n664);
or (n797,n798,n21);
not (n798,n57);
nand (n799,n800,n805);
or (n800,n801,n154);
not (n801,n802);
nand (n802,n803,n804);
or (n803,n74,n417);
or (n804,n73,n187);
or (n805,n114,n741);
or (n806,n807,n829);
and (n807,n808,n822);
xor (n808,n809,n815);
nand (n809,n810,n811);
or (n810,n29,n747);
or (n811,n812,n24);
nor (n812,n813,n814);
and (n813,n562,n22);
and (n814,n518,n21);
nand (n815,n816,n821);
or (n816,n817,n52);
not (n817,n818);
nand (n818,n819,n820);
or (n819,n50,n664);
or (n820,n49,n591);
nand (n821,n760,n55);
nand (n822,n823,n828);
or (n823,n824,n194);
not (n824,n825);
nor (n825,n826,n827);
and (n826,n146,n95);
and (n827,n96,n144);
or (n828,n767,n195);
and (n829,n809,n815);
xor (n830,n737,n745);
and (n831,n792,n806);
and (n832,n787,n788);
nand (n833,n648,n728);
not (n834,n835);
nor (n835,n836,n851);
nor (n836,n837,n848);
xor (n837,n838,n845);
xor (n838,n839,n844);
nand (n839,n840,n842);
or (n840,n546,n841);
not (n841,n522);
or (n842,n522,n843);
not (n843,n546);
xor (n844,n575,n578);
or (n845,n846,n847);
and (n846,n695,n698);
and (n847,n696,n697);
or (n848,n849,n850);
and (n849,n649,n694);
and (n850,n650,n651);
nor (n851,n852,n853);
xor (n852,n570,n573);
or (n853,n854,n855);
and (n854,n838,n845);
and (n855,n839,n844);
nor (n856,n857,n862);
and (n857,n858,n859);
not (n858,n851);
nor (n859,n860,n861);
not (n860,n837);
not (n861,n848);
and (n862,n852,n853);
nand (n863,n835,n864,n1153);
nand (n864,n865,n1141,n1152);
nand (n865,n866,n904,n1003);
nand (n866,n867,n869);
not (n867,n868);
xor (n868,n786,n789);
not (n869,n870);
or (n870,n871,n903);
and (n871,n872,n902);
xor (n872,n873,n874);
xor (n873,n756,n771);
or (n874,n875,n901);
and (n875,n876,n884);
xor (n876,n877,n883);
nand (n877,n878,n882);
or (n878,n70,n879);
nor (n879,n880,n881);
and (n880,n32,n380);
and (n881,n33,n451);
or (n882,n773,n71);
xor (n883,n793,n799);
or (n884,n885,n900);
and (n885,n886,n894);
xor (n886,n887,n888);
and (n887,n55,n591);
nand (n888,n889,n890);
or (n889,n195,n824);
or (n890,n891,n194);
nor (n891,n892,n893);
and (n892,n95,n161);
and (n893,n96,n287);
nand (n894,n895,n899);
or (n895,n24,n896);
nor (n896,n897,n898);
and (n897,n21,n564);
and (n898,n22,n628);
or (n899,n29,n812);
and (n900,n887,n888);
and (n901,n877,n883);
xor (n902,n791,n830);
and (n903,n873,n874);
nor (n904,n905,n998);
not (n905,n906);
nor (n906,n907,n971);
nor (n907,n908,n943);
xor (n908,n909,n942);
xor (n909,n910,n911);
xor (n910,n808,n822);
or (n911,n912,n941);
and (n912,n913,n927);
xor (n913,n914,n921);
nand (n914,n915,n920);
or (n915,n916,n154);
not (n916,n917);
nand (n917,n918,n919);
or (n918,n74,n377);
or (n919,n73,n251);
nand (n920,n100,n802);
nand (n921,n922,n926);
or (n922,n70,n923);
nor (n923,n924,n925);
and (n924,n454,n32);
and (n925,n33,n613);
or (n926,n71,n879);
and (n927,n928,n934);
nor (n928,n929,n21);
nor (n929,n930,n932);
and (n930,n931,n664);
nand (n931,n33,n27);
and (n932,n32,n933);
not (n933,n27);
nand (n934,n935,n940);
or (n935,n194,n936);
not (n936,n937);
nor (n937,n938,n939);
and (n938,n96,n187);
and (n939,n417,n95);
or (n940,n891,n195);
and (n941,n914,n921);
xor (n942,n876,n884);
or (n943,n944,n970);
and (n944,n945,n969);
xor (n945,n946,n968);
or (n946,n947,n967);
and (n947,n948,n961);
xor (n948,n949,n955);
nand (n949,n950,n954);
or (n950,n24,n951);
nor (n951,n952,n953);
and (n952,n21,n591);
and (n953,n22,n664);
or (n954,n896,n29);
nand (n955,n956,n957);
or (n956,n916,n114);
nand (n957,n99,n958);
nand (n958,n959,n960);
or (n959,n74,n451);
or (n960,n73,n380);
nand (n961,n962,n966);
or (n962,n70,n963);
nor (n963,n964,n965);
and (n964,n32,n518);
and (n965,n33,n562);
or (n966,n71,n923);
and (n967,n949,n955);
xor (n968,n886,n894);
xor (n969,n913,n927);
and (n970,n946,n968);
nor (n971,n972,n973);
xor (n972,n945,n969);
or (n973,n974,n997);
and (n974,n975,n996);
xor (n975,n976,n977);
xor (n976,n928,n934);
or (n977,n978,n995);
and (n978,n979,n988);
xor (n979,n980,n981);
and (n980,n30,n591);
nand (n981,n982,n983);
or (n982,n195,n936);
or (n983,n984,n194);
not (n984,n985);
nand (n985,n986,n987);
or (n986,n251,n95);
nand (n987,n95,n251);
nand (n988,n989,n994);
or (n989,n990,n154);
not (n990,n991);
nor (n991,n992,n993);
and (n992,n74,n454);
and (n993,n613,n73);
nand (n994,n100,n958);
and (n995,n980,n981);
xor (n996,n948,n961);
and (n997,n976,n977);
nor (n998,n999,n1000);
xor (n999,n872,n902);
or (n1000,n1001,n1002);
and (n1001,n909,n942);
and (n1002,n910,n911);
or (n1003,n1004,n1140);
and (n1004,n1005,n1032);
xor (n1005,n1006,n1031);
or (n1006,n1007,n1030);
and (n1007,n1008,n1029);
xor (n1008,n1009,n1015);
nand (n1009,n1010,n1014);
or (n1010,n70,n1011);
nor (n1011,n1012,n1013);
and (n1012,n32,n564);
and (n1013,n33,n628);
or (n1014,n71,n963);
and (n1015,n1016,n1023);
nand (n1016,n1017,n1022);
or (n1017,n194,n1018);
not (n1018,n1019);
nor (n1019,n1020,n1021);
and (n1020,n96,n380);
and (n1021,n451,n95);
nand (n1022,n985,n196);
not (n1023,n1024);
nand (n1024,n1025,n33);
nand (n1025,n1026,n1027);
or (n1026,n74,n75);
nand (n1027,n1028,n664);
or (n1028,n77,n73);
xor (n1029,n979,n988);
and (n1030,n1009,n1015);
xor (n1031,n975,n996);
or (n1032,n1033,n1139);
and (n1033,n1034,n1058);
xor (n1034,n1035,n1057);
or (n1035,n1036,n1056);
and (n1036,n1037,n1052);
xor (n1037,n1038,n1045);
nand (n1038,n1039,n1044);
or (n1039,n1040,n154);
not (n1040,n1041);
nand (n1041,n1042,n1043);
or (n1042,n74,n562);
or (n1043,n73,n518);
nand (n1044,n100,n991);
nand (n1045,n1046,n1051);
or (n1046,n1047,n70);
not (n1047,n1048);
nand (n1048,n1049,n1050);
or (n1049,n664,n33);
or (n1050,n32,n591);
or (n1051,n71,n1011);
nand (n1052,n1053,n1055);
or (n1053,n1023,n1054);
not (n1054,n1016);
or (n1055,n1016,n1024);
and (n1056,n1038,n1045);
xor (n1057,n1008,n1029);
or (n1058,n1059,n1138);
and (n1059,n1060,n1081);
xor (n1060,n1061,n1080);
or (n1061,n1062,n1079);
and (n1062,n1063,n1072);
xor (n1063,n1064,n1065);
nor (n1064,n71,n664);
nand (n1065,n1066,n1071);
or (n1066,n1067,n154);
not (n1067,n1068);
nor (n1068,n1069,n1070);
and (n1069,n628,n73);
and (n1070,n74,n564);
nand (n1071,n100,n1041);
nand (n1072,n1073,n1078);
or (n1073,n194,n1074);
not (n1074,n1075);
nor (n1075,n1076,n1077);
and (n1076,n613,n95);
and (n1077,n96,n454);
or (n1078,n1018,n195);
and (n1079,n1064,n1065);
xor (n1080,n1037,n1052);
or (n1081,n1082,n1137);
and (n1082,n1083,n1136);
xor (n1083,n1084,n1097);
nor (n1084,n1085,n1092);
not (n1085,n1086);
nand (n1086,n1087,n1088);
or (n1087,n195,n1074);
nand (n1088,n1089,n394);
nor (n1089,n1090,n1091);
and (n1090,n562,n95);
and (n1091,n96,n518);
nand (n1092,n1093,n74);
nand (n1093,n1094,n1095);
or (n1094,n102,n96);
or (n1095,n1096,n591);
and (n1096,n96,n102);
nand (n1097,n1098,n1135);
or (n1098,n1099,n1123);
not (n1099,n1100);
nand (n1100,n1101,n1122);
or (n1101,n1102,n1111);
nor (n1102,n1103,n1104);
and (n1103,n100,n591);
nand (n1104,n1105,n1107);
or (n1105,n195,n1106);
not (n1106,n1089);
nand (n1107,n1108,n394);
nand (n1108,n1109,n1110);
or (n1109,n628,n96);
or (n1110,n95,n564);
nand (n1111,n1112,n1115);
not (n1112,n1113);
nand (n1113,n1114,n96);
nand (n1114,n591,n196);
nand (n1115,n1116,n1118);
or (n1116,n195,n1117);
not (n1117,n1108);
nand (n1118,n1119,n394);
nor (n1119,n1120,n1121);
and (n1120,n664,n95);
and (n1121,n96,n591);
nand (n1122,n1103,n1104);
not (n1123,n1124);
nand (n1124,n1125,n1129);
nor (n1125,n1126,n1127);
and (n1126,n1092,n1086);
and (n1127,n1128,n1085);
not (n1128,n1092);
nor (n1129,n1130,n1134);
and (n1130,n99,n1131);
nand (n1131,n1132,n1133);
or (n1132,n74,n664);
or (n1133,n73,n591);
and (n1134,n100,n1068);
or (n1135,n1125,n1129);
xor (n1136,n1063,n1072);
and (n1137,n1084,n1097);
and (n1138,n1061,n1080);
and (n1139,n1035,n1057);
and (n1140,n1006,n1031);
nand (n1141,n1142,n866);
nand (n1142,n1143,n1151);
or (n1143,n998,n1144);
nand (n1144,n1145,n1150);
or (n1145,n1146,n1148);
not (n1146,n1147);
nand (n1147,n972,n973);
not (n1148,n1149);
nand (n1149,n908,n943);
not (n1150,n907);
nand (n1151,n999,n1000);
nand (n1152,n868,n870);
nor (n1153,n1154,n647);
not (n1154,n1155);
or (n1155,n784,n783);
not (n1156,n1157);
nand (n1157,n1158,n1166);
or (n1158,n1159,n1164);
not (n1159,n1160);
nand (n1160,n1161,n1163);
or (n1161,n634,n1162);
nand (n1162,n502,n568);
nand (n1163,n635,n636);
not (n1164,n1165);
nor (n1165,n358,n432);
nor (n1166,n1167,n1169);
and (n1167,n357,n1168);
and (n1168,n433,n434);
and (n1169,n359,n360);
or (n1170,n353,n3);
xor (n1171,n1172,n2021);
xor (n1172,n1173,n2020);
xor (n1173,n1174,n1995);
xor (n1174,n1175,n1994);
xor (n1175,n1176,n1962);
xor (n1176,n1177,n1961);
xor (n1177,n1178,n1922);
xor (n1178,n1179,n167);
xor (n1179,n1180,n1877);
xor (n1180,n1181,n1876);
xor (n1181,n1182,n1826);
xor (n1182,n1183,n128);
xor (n1183,n1184,n1770);
xor (n1184,n1185,n1769);
xor (n1185,n1186,n1708);
xor (n1186,n1187,n1707);
or (n1187,n1188,n1644);
and (n1188,n1189,n346);
or (n1189,n1190,n1581);
and (n1190,n1191,n160);
or (n1191,n1192,n1517);
and (n1192,n1193,n186);
or (n1193,n1194,n1452);
and (n1194,n1195,n250);
or (n1195,n1196,n1388);
and (n1196,n1197,n379);
or (n1197,n1198,n1326);
and (n1198,n1199,n453);
or (n1199,n1200,n1262);
and (n1200,n1201,n517);
and (n1201,n563,n1202);
or (n1202,n1203,n1205);
and (n1203,n590,n1204);
and (n1204,n133,n564);
and (n1205,n1206,n1207);
xor (n1206,n590,n1204);
or (n1207,n1208,n1211);
and (n1208,n1209,n1210);
and (n1209,n133,n591);
and (n1210,n50,n564);
and (n1211,n1212,n1213);
xor (n1212,n1209,n1210);
or (n1213,n1214,n1217);
and (n1214,n1215,n1216);
and (n1215,n50,n591);
and (n1216,n57,n564);
and (n1217,n1218,n1219);
xor (n1218,n1215,n1216);
or (n1219,n1220,n1223);
and (n1220,n1221,n1222);
and (n1221,n57,n591);
and (n1222,n22,n564);
and (n1223,n1224,n1225);
xor (n1224,n1221,n1222);
or (n1225,n1226,n1229);
and (n1226,n1227,n1228);
and (n1227,n22,n591);
and (n1228,n27,n564);
and (n1229,n1230,n1231);
xor (n1230,n1227,n1228);
or (n1231,n1232,n1235);
and (n1232,n1233,n1234);
and (n1233,n27,n591);
and (n1234,n33,n564);
and (n1235,n1236,n1237);
xor (n1236,n1233,n1234);
or (n1237,n1238,n1241);
and (n1238,n1239,n1240);
and (n1239,n33,n591);
and (n1240,n75,n564);
and (n1241,n1242,n1243);
xor (n1242,n1239,n1240);
or (n1243,n1244,n1246);
and (n1244,n1245,n1070);
and (n1245,n75,n591);
and (n1246,n1247,n1248);
xor (n1247,n1245,n1070);
or (n1248,n1249,n1252);
and (n1249,n1250,n1251);
and (n1250,n74,n591);
and (n1251,n102,n564);
and (n1252,n1253,n1254);
xor (n1253,n1250,n1251);
or (n1254,n1255,n1258);
and (n1255,n1256,n1257);
and (n1256,n102,n591);
and (n1257,n96,n564);
and (n1258,n1259,n1260);
xor (n1259,n1256,n1257);
and (n1260,n1121,n1261);
and (n1261,n196,n564);
and (n1262,n1263,n1264);
xor (n1263,n1201,n517);
or (n1264,n1265,n1268);
and (n1265,n1266,n1267);
xor (n1266,n563,n1202);
and (n1267,n133,n518);
and (n1268,n1269,n1270);
xor (n1269,n1266,n1267);
or (n1270,n1271,n1274);
and (n1271,n1272,n1273);
xor (n1272,n1206,n1207);
and (n1273,n50,n518);
and (n1274,n1275,n1276);
xor (n1275,n1272,n1273);
or (n1276,n1277,n1280);
and (n1277,n1278,n1279);
xor (n1278,n1212,n1213);
and (n1279,n57,n518);
and (n1280,n1281,n1282);
xor (n1281,n1278,n1279);
or (n1282,n1283,n1286);
and (n1283,n1284,n1285);
xor (n1284,n1218,n1219);
and (n1285,n22,n518);
and (n1286,n1287,n1288);
xor (n1287,n1284,n1285);
or (n1288,n1289,n1292);
and (n1289,n1290,n1291);
xor (n1290,n1224,n1225);
and (n1291,n27,n518);
and (n1292,n1293,n1294);
xor (n1293,n1290,n1291);
or (n1294,n1295,n1298);
and (n1295,n1296,n1297);
xor (n1296,n1230,n1231);
and (n1297,n33,n518);
and (n1298,n1299,n1300);
xor (n1299,n1296,n1297);
or (n1300,n1301,n1304);
and (n1301,n1302,n1303);
xor (n1302,n1236,n1237);
and (n1303,n75,n518);
and (n1304,n1305,n1306);
xor (n1305,n1302,n1303);
or (n1306,n1307,n1310);
and (n1307,n1308,n1309);
xor (n1308,n1242,n1243);
and (n1309,n74,n518);
and (n1310,n1311,n1312);
xor (n1311,n1308,n1309);
or (n1312,n1313,n1316);
and (n1313,n1314,n1315);
xor (n1314,n1247,n1248);
and (n1315,n102,n518);
and (n1316,n1317,n1318);
xor (n1317,n1314,n1315);
or (n1318,n1319,n1321);
and (n1319,n1320,n1091);
xor (n1320,n1253,n1254);
and (n1321,n1322,n1323);
xor (n1322,n1320,n1091);
and (n1323,n1324,n1325);
xor (n1324,n1259,n1260);
and (n1325,n196,n518);
and (n1326,n1327,n1328);
xor (n1327,n1199,n453);
or (n1328,n1329,n1332);
and (n1329,n1330,n1331);
xor (n1330,n1263,n1264);
and (n1331,n133,n454);
and (n1332,n1333,n1334);
xor (n1333,n1330,n1331);
or (n1334,n1335,n1337);
and (n1335,n1336,n614);
xor (n1336,n1269,n1270);
and (n1337,n1338,n1339);
xor (n1338,n1336,n614);
or (n1339,n1340,n1343);
and (n1340,n1341,n1342);
xor (n1341,n1275,n1276);
and (n1342,n57,n454);
and (n1343,n1344,n1345);
xor (n1344,n1341,n1342);
or (n1345,n1346,n1349);
and (n1346,n1347,n1348);
xor (n1347,n1281,n1282);
and (n1348,n22,n454);
and (n1349,n1350,n1351);
xor (n1350,n1347,n1348);
or (n1351,n1352,n1355);
and (n1352,n1353,n1354);
xor (n1353,n1287,n1288);
and (n1354,n27,n454);
and (n1355,n1356,n1357);
xor (n1356,n1353,n1354);
or (n1357,n1358,n1361);
and (n1358,n1359,n1360);
xor (n1359,n1293,n1294);
and (n1360,n33,n454);
and (n1361,n1362,n1363);
xor (n1362,n1359,n1360);
or (n1363,n1364,n1367);
and (n1364,n1365,n1366);
xor (n1365,n1299,n1300);
and (n1366,n75,n454);
and (n1367,n1368,n1369);
xor (n1368,n1365,n1366);
or (n1369,n1370,n1372);
and (n1370,n1371,n992);
xor (n1371,n1305,n1306);
and (n1372,n1373,n1374);
xor (n1373,n1371,n992);
or (n1374,n1375,n1378);
and (n1375,n1376,n1377);
xor (n1376,n1311,n1312);
and (n1377,n102,n454);
and (n1378,n1379,n1380);
xor (n1379,n1376,n1377);
or (n1380,n1381,n1383);
and (n1381,n1382,n1077);
xor (n1382,n1317,n1318);
and (n1383,n1384,n1385);
xor (n1384,n1382,n1077);
and (n1385,n1386,n1387);
xor (n1386,n1322,n1323);
and (n1387,n196,n454);
and (n1388,n1389,n1390);
xor (n1389,n1197,n379);
or (n1390,n1391,n1394);
and (n1391,n1392,n1393);
xor (n1392,n1327,n1328);
and (n1393,n133,n380);
and (n1394,n1395,n1396);
xor (n1395,n1392,n1393);
or (n1396,n1397,n1400);
and (n1397,n1398,n1399);
xor (n1398,n1333,n1334);
and (n1399,n50,n380);
and (n1400,n1401,n1402);
xor (n1401,n1398,n1399);
or (n1402,n1403,n1406);
and (n1403,n1404,n1405);
xor (n1404,n1338,n1339);
and (n1405,n57,n380);
and (n1406,n1407,n1408);
xor (n1407,n1404,n1405);
or (n1408,n1409,n1412);
and (n1409,n1410,n1411);
xor (n1410,n1344,n1345);
and (n1411,n22,n380);
and (n1412,n1413,n1414);
xor (n1413,n1410,n1411);
or (n1414,n1415,n1418);
and (n1415,n1416,n1417);
xor (n1416,n1350,n1351);
and (n1417,n27,n380);
and (n1418,n1419,n1420);
xor (n1419,n1416,n1417);
or (n1420,n1421,n1424);
and (n1421,n1422,n1423);
xor (n1422,n1356,n1357);
and (n1423,n33,n380);
and (n1424,n1425,n1426);
xor (n1425,n1422,n1423);
or (n1426,n1427,n1430);
and (n1427,n1428,n1429);
xor (n1428,n1362,n1363);
and (n1429,n75,n380);
and (n1430,n1431,n1432);
xor (n1431,n1428,n1429);
or (n1432,n1433,n1436);
and (n1433,n1434,n1435);
xor (n1434,n1368,n1369);
and (n1435,n74,n380);
and (n1436,n1437,n1438);
xor (n1437,n1434,n1435);
or (n1438,n1439,n1442);
and (n1439,n1440,n1441);
xor (n1440,n1373,n1374);
and (n1441,n102,n380);
and (n1442,n1443,n1444);
xor (n1443,n1440,n1441);
or (n1444,n1445,n1447);
and (n1445,n1446,n1020);
xor (n1446,n1379,n1380);
and (n1447,n1448,n1449);
xor (n1448,n1446,n1020);
and (n1449,n1450,n1451);
xor (n1450,n1384,n1385);
and (n1451,n196,n380);
and (n1452,n1453,n1454);
xor (n1453,n1195,n250);
or (n1454,n1455,n1458);
and (n1455,n1456,n1457);
xor (n1456,n1389,n1390);
and (n1457,n133,n251);
and (n1458,n1459,n1460);
xor (n1459,n1456,n1457);
or (n1460,n1461,n1464);
and (n1461,n1462,n1463);
xor (n1462,n1395,n1396);
and (n1463,n50,n251);
and (n1464,n1465,n1466);
xor (n1465,n1462,n1463);
or (n1466,n1467,n1470);
and (n1467,n1468,n1469);
xor (n1468,n1401,n1402);
and (n1469,n57,n251);
and (n1470,n1471,n1472);
xor (n1471,n1468,n1469);
or (n1472,n1473,n1476);
and (n1473,n1474,n1475);
xor (n1474,n1407,n1408);
and (n1475,n22,n251);
and (n1476,n1477,n1478);
xor (n1477,n1474,n1475);
or (n1478,n1479,n1482);
and (n1479,n1480,n1481);
xor (n1480,n1413,n1414);
and (n1481,n27,n251);
and (n1482,n1483,n1484);
xor (n1483,n1480,n1481);
or (n1484,n1485,n1488);
and (n1485,n1486,n1487);
xor (n1486,n1419,n1420);
and (n1487,n33,n251);
and (n1488,n1489,n1490);
xor (n1489,n1486,n1487);
or (n1490,n1491,n1494);
and (n1491,n1492,n1493);
xor (n1492,n1425,n1426);
and (n1493,n75,n251);
and (n1494,n1495,n1496);
xor (n1495,n1492,n1493);
or (n1496,n1497,n1500);
and (n1497,n1498,n1499);
xor (n1498,n1431,n1432);
and (n1499,n74,n251);
and (n1500,n1501,n1502);
xor (n1501,n1498,n1499);
or (n1502,n1503,n1506);
and (n1503,n1504,n1505);
xor (n1504,n1437,n1438);
and (n1505,n102,n251);
and (n1506,n1507,n1508);
xor (n1507,n1504,n1505);
or (n1508,n1509,n1512);
and (n1509,n1510,n1511);
xor (n1510,n1443,n1444);
and (n1511,n96,n251);
and (n1512,n1513,n1514);
xor (n1513,n1510,n1511);
and (n1514,n1515,n1516);
xor (n1515,n1448,n1449);
and (n1516,n196,n251);
and (n1517,n1518,n1519);
xor (n1518,n1193,n186);
or (n1519,n1520,n1523);
and (n1520,n1521,n1522);
xor (n1521,n1453,n1454);
and (n1522,n133,n187);
and (n1523,n1524,n1525);
xor (n1524,n1521,n1522);
or (n1525,n1526,n1529);
and (n1526,n1527,n1528);
xor (n1527,n1459,n1460);
and (n1528,n50,n187);
and (n1529,n1530,n1531);
xor (n1530,n1527,n1528);
or (n1531,n1532,n1535);
and (n1532,n1533,n1534);
xor (n1533,n1465,n1466);
and (n1534,n57,n187);
and (n1535,n1536,n1537);
xor (n1536,n1533,n1534);
or (n1537,n1538,n1541);
and (n1538,n1539,n1540);
xor (n1539,n1471,n1472);
and (n1540,n22,n187);
and (n1541,n1542,n1543);
xor (n1542,n1539,n1540);
or (n1543,n1544,n1547);
and (n1544,n1545,n1546);
xor (n1545,n1477,n1478);
and (n1546,n27,n187);
and (n1547,n1548,n1549);
xor (n1548,n1545,n1546);
or (n1549,n1550,n1553);
and (n1550,n1551,n1552);
xor (n1551,n1483,n1484);
and (n1552,n33,n187);
and (n1553,n1554,n1555);
xor (n1554,n1551,n1552);
or (n1555,n1556,n1559);
and (n1556,n1557,n1558);
xor (n1557,n1489,n1490);
and (n1558,n75,n187);
and (n1559,n1560,n1561);
xor (n1560,n1557,n1558);
or (n1561,n1562,n1565);
and (n1562,n1563,n1564);
xor (n1563,n1495,n1496);
and (n1564,n74,n187);
and (n1565,n1566,n1567);
xor (n1566,n1563,n1564);
or (n1567,n1568,n1571);
and (n1568,n1569,n1570);
xor (n1569,n1501,n1502);
and (n1570,n102,n187);
and (n1571,n1572,n1573);
xor (n1572,n1569,n1570);
or (n1573,n1574,n1576);
and (n1574,n1575,n938);
xor (n1575,n1507,n1508);
and (n1576,n1577,n1578);
xor (n1577,n1575,n938);
and (n1578,n1579,n1580);
xor (n1579,n1513,n1514);
and (n1580,n196,n187);
and (n1581,n1582,n1583);
xor (n1582,n1191,n160);
or (n1583,n1584,n1587);
and (n1584,n1585,n1586);
xor (n1585,n1518,n1519);
and (n1586,n133,n161);
and (n1587,n1588,n1589);
xor (n1588,n1585,n1586);
or (n1589,n1590,n1592);
and (n1590,n1591,n288);
xor (n1591,n1524,n1525);
and (n1592,n1593,n1594);
xor (n1593,n1591,n288);
or (n1594,n1595,n1598);
and (n1595,n1596,n1597);
xor (n1596,n1530,n1531);
and (n1597,n57,n161);
and (n1598,n1599,n1600);
xor (n1599,n1596,n1597);
or (n1600,n1601,n1603);
and (n1601,n1602,n481);
xor (n1602,n1536,n1537);
and (n1603,n1604,n1605);
xor (n1604,n1602,n481);
or (n1605,n1606,n1609);
and (n1606,n1607,n1608);
xor (n1607,n1542,n1543);
and (n1608,n27,n161);
and (n1609,n1610,n1611);
xor (n1610,n1607,n1608);
or (n1611,n1612,n1615);
and (n1612,n1613,n1614);
xor (n1613,n1548,n1549);
and (n1614,n33,n161);
and (n1615,n1616,n1617);
xor (n1616,n1613,n1614);
or (n1617,n1618,n1621);
and (n1618,n1619,n1620);
xor (n1619,n1554,n1555);
and (n1620,n75,n161);
and (n1621,n1622,n1623);
xor (n1622,n1619,n1620);
or (n1623,n1624,n1627);
and (n1624,n1625,n1626);
xor (n1625,n1560,n1561);
and (n1626,n74,n161);
and (n1627,n1628,n1629);
xor (n1628,n1625,n1626);
or (n1629,n1630,n1633);
and (n1630,n1631,n1632);
xor (n1631,n1566,n1567);
and (n1632,n102,n161);
and (n1633,n1634,n1635);
xor (n1634,n1631,n1632);
or (n1635,n1636,n1639);
and (n1636,n1637,n1638);
xor (n1637,n1572,n1573);
and (n1638,n96,n161);
and (n1639,n1640,n1641);
xor (n1640,n1637,n1638);
and (n1641,n1642,n1643);
xor (n1642,n1577,n1578);
and (n1643,n196,n161);
and (n1644,n1645,n1646);
xor (n1645,n1189,n346);
or (n1646,n1647,n1650);
and (n1647,n1648,n1649);
xor (n1648,n1582,n1583);
and (n1649,n133,n144);
and (n1650,n1651,n1652);
xor (n1651,n1648,n1649);
or (n1652,n1653,n1656);
and (n1653,n1654,n1655);
xor (n1654,n1588,n1589);
and (n1655,n50,n144);
and (n1656,n1657,n1658);
xor (n1657,n1654,n1655);
or (n1658,n1659,n1662);
and (n1659,n1660,n1661);
xor (n1660,n1593,n1594);
and (n1661,n57,n144);
and (n1662,n1663,n1664);
xor (n1663,n1660,n1661);
or (n1664,n1665,n1667);
and (n1665,n1666,n410);
xor (n1666,n1599,n1600);
and (n1667,n1668,n1669);
xor (n1668,n1666,n410);
or (n1669,n1670,n1673);
and (n1670,n1671,n1672);
xor (n1671,n1604,n1605);
and (n1672,n27,n144);
and (n1673,n1674,n1675);
xor (n1674,n1671,n1672);
or (n1675,n1676,n1679);
and (n1676,n1677,n1678);
xor (n1677,n1610,n1611);
and (n1678,n33,n144);
and (n1679,n1680,n1681);
xor (n1680,n1677,n1678);
or (n1681,n1682,n1685);
and (n1682,n1683,n1684);
xor (n1683,n1616,n1617);
and (n1684,n75,n144);
and (n1685,n1686,n1687);
xor (n1686,n1683,n1684);
or (n1687,n1688,n1691);
and (n1688,n1689,n1690);
xor (n1689,n1622,n1623);
and (n1690,n74,n144);
and (n1691,n1692,n1693);
xor (n1692,n1689,n1690);
or (n1693,n1694,n1697);
and (n1694,n1695,n1696);
xor (n1695,n1628,n1629);
and (n1696,n102,n144);
and (n1697,n1698,n1699);
xor (n1698,n1695,n1696);
or (n1699,n1700,n1702);
and (n1700,n1701,n827);
xor (n1701,n1634,n1635);
and (n1702,n1703,n1704);
xor (n1703,n1701,n827);
and (n1704,n1705,n1706);
xor (n1705,n1640,n1641);
and (n1706,n196,n144);
and (n1707,n138,n48);
or (n1708,n1709,n1712);
and (n1709,n1710,n1711);
xor (n1710,n1645,n1646);
and (n1711,n133,n48);
and (n1712,n1713,n1714);
xor (n1713,n1710,n1711);
or (n1714,n1715,n1717);
and (n1715,n1716,n51);
xor (n1716,n1651,n1652);
and (n1717,n1718,n1719);
xor (n1718,n1716,n51);
or (n1719,n1720,n1723);
and (n1720,n1721,n1722);
xor (n1721,n1657,n1658);
and (n1722,n57,n48);
and (n1723,n1724,n1725);
xor (n1724,n1721,n1722);
or (n1725,n1726,n1728);
and (n1726,n1727,n280);
xor (n1727,n1663,n1664);
and (n1728,n1729,n1730);
xor (n1729,n1727,n280);
or (n1730,n1731,n1734);
and (n1731,n1732,n1733);
xor (n1732,n1668,n1669);
and (n1733,n27,n48);
and (n1734,n1735,n1736);
xor (n1735,n1732,n1733);
or (n1736,n1737,n1740);
and (n1737,n1738,n1739);
xor (n1738,n1674,n1675);
and (n1739,n33,n48);
and (n1740,n1741,n1742);
xor (n1741,n1738,n1739);
or (n1742,n1743,n1746);
and (n1743,n1744,n1745);
xor (n1744,n1680,n1681);
and (n1745,n75,n48);
and (n1746,n1747,n1748);
xor (n1747,n1744,n1745);
or (n1748,n1749,n1752);
and (n1749,n1750,n1751);
xor (n1750,n1686,n1687);
and (n1751,n74,n48);
and (n1752,n1753,n1754);
xor (n1753,n1750,n1751);
or (n1754,n1755,n1758);
and (n1755,n1756,n1757);
xor (n1756,n1692,n1693);
and (n1757,n102,n48);
and (n1758,n1759,n1760);
xor (n1759,n1756,n1757);
or (n1760,n1761,n1764);
and (n1761,n1762,n1763);
xor (n1762,n1698,n1699);
and (n1763,n96,n48);
and (n1764,n1765,n1766);
xor (n1765,n1762,n1763);
and (n1766,n1767,n1768);
xor (n1767,n1703,n1704);
and (n1768,n196,n48);
and (n1769,n133,n66);
or (n1770,n1771,n1774);
and (n1771,n1772,n1773);
xor (n1772,n1713,n1714);
and (n1773,n50,n66);
and (n1774,n1775,n1776);
xor (n1775,n1772,n1773);
or (n1776,n1777,n1780);
and (n1777,n1778,n1779);
xor (n1778,n1718,n1719);
and (n1779,n57,n66);
and (n1780,n1781,n1782);
xor (n1781,n1778,n1779);
or (n1782,n1783,n1785);
and (n1783,n1784,n217);
xor (n1784,n1724,n1725);
and (n1785,n1786,n1787);
xor (n1786,n1784,n217);
or (n1787,n1788,n1791);
and (n1788,n1789,n1790);
xor (n1789,n1729,n1730);
and (n1790,n27,n66);
and (n1791,n1792,n1793);
xor (n1792,n1789,n1790);
or (n1793,n1794,n1797);
and (n1794,n1795,n1796);
xor (n1795,n1735,n1736);
and (n1796,n33,n66);
and (n1797,n1798,n1799);
xor (n1798,n1795,n1796);
or (n1799,n1800,n1803);
and (n1800,n1801,n1802);
xor (n1801,n1741,n1742);
and (n1802,n75,n66);
and (n1803,n1804,n1805);
xor (n1804,n1801,n1802);
or (n1805,n1806,n1809);
and (n1806,n1807,n1808);
xor (n1807,n1747,n1748);
and (n1808,n74,n66);
and (n1809,n1810,n1811);
xor (n1810,n1807,n1808);
or (n1811,n1812,n1815);
and (n1812,n1813,n1814);
xor (n1813,n1753,n1754);
and (n1814,n102,n66);
and (n1815,n1816,n1817);
xor (n1816,n1813,n1814);
or (n1817,n1818,n1821);
and (n1818,n1819,n1820);
xor (n1819,n1759,n1760);
and (n1820,n96,n66);
and (n1821,n1822,n1823);
xor (n1822,n1819,n1820);
and (n1823,n1824,n1825);
xor (n1824,n1765,n1766);
and (n1825,n196,n66);
or (n1826,n1827,n1830);
and (n1827,n1828,n1829);
xor (n1828,n1775,n1776);
and (n1829,n57,n20);
and (n1830,n1831,n1832);
xor (n1831,n1828,n1829);
or (n1832,n1833,n1835);
and (n1833,n1834,n23);
xor (n1834,n1781,n1782);
and (n1835,n1836,n1837);
xor (n1836,n1834,n23);
or (n1837,n1838,n1841);
and (n1838,n1839,n1840);
xor (n1839,n1786,n1787);
and (n1840,n27,n20);
and (n1841,n1842,n1843);
xor (n1842,n1839,n1840);
or (n1843,n1844,n1847);
and (n1844,n1845,n1846);
xor (n1845,n1792,n1793);
and (n1846,n33,n20);
and (n1847,n1848,n1849);
xor (n1848,n1845,n1846);
or (n1849,n1850,n1853);
and (n1850,n1851,n1852);
xor (n1851,n1798,n1799);
and (n1852,n75,n20);
and (n1853,n1854,n1855);
xor (n1854,n1851,n1852);
or (n1855,n1856,n1859);
and (n1856,n1857,n1858);
xor (n1857,n1804,n1805);
and (n1858,n74,n20);
and (n1859,n1860,n1861);
xor (n1860,n1857,n1858);
or (n1861,n1862,n1865);
and (n1862,n1863,n1864);
xor (n1863,n1810,n1811);
and (n1864,n102,n20);
and (n1865,n1866,n1867);
xor (n1866,n1863,n1864);
or (n1867,n1868,n1871);
and (n1868,n1869,n1870);
xor (n1869,n1816,n1817);
and (n1870,n96,n20);
and (n1871,n1872,n1873);
xor (n1872,n1869,n1870);
and (n1873,n1874,n1875);
xor (n1874,n1822,n1823);
and (n1875,n196,n20);
and (n1876,n57,n39);
or (n1877,n1878,n1881);
and (n1878,n1879,n1880);
xor (n1879,n1831,n1832);
and (n1880,n22,n39);
and (n1881,n1882,n1883);
xor (n1882,n1879,n1880);
or (n1883,n1884,n1887);
and (n1884,n1885,n1886);
xor (n1885,n1836,n1837);
and (n1886,n27,n39);
and (n1887,n1888,n1889);
xor (n1888,n1885,n1886);
or (n1889,n1890,n1893);
and (n1890,n1891,n1892);
xor (n1891,n1842,n1843);
and (n1892,n33,n39);
and (n1893,n1894,n1895);
xor (n1894,n1891,n1892);
or (n1895,n1896,n1899);
and (n1896,n1897,n1898);
xor (n1897,n1848,n1849);
and (n1898,n75,n39);
and (n1899,n1900,n1901);
xor (n1900,n1897,n1898);
or (n1901,n1902,n1905);
and (n1902,n1903,n1904);
xor (n1903,n1854,n1855);
and (n1904,n74,n39);
and (n1905,n1906,n1907);
xor (n1906,n1903,n1904);
or (n1907,n1908,n1911);
and (n1908,n1909,n1910);
xor (n1909,n1860,n1861);
and (n1910,n102,n39);
and (n1911,n1912,n1913);
xor (n1912,n1909,n1910);
or (n1913,n1914,n1917);
and (n1914,n1915,n1916);
xor (n1915,n1866,n1867);
and (n1916,n96,n39);
and (n1917,n1918,n1919);
xor (n1918,n1915,n1916);
and (n1919,n1920,n1921);
xor (n1920,n1872,n1873);
and (n1921,n196,n39);
or (n1922,n1923,n1926);
and (n1923,n1924,n1925);
xor (n1924,n1882,n1883);
and (n1925,n27,n83);
and (n1926,n1927,n1928);
xor (n1927,n1924,n1925);
or (n1928,n1929,n1932);
and (n1929,n1930,n1931);
xor (n1930,n1888,n1889);
and (n1931,n33,n83);
and (n1932,n1933,n1934);
xor (n1933,n1930,n1931);
or (n1934,n1935,n1938);
and (n1935,n1936,n1937);
xor (n1936,n1894,n1895);
and (n1937,n75,n83);
and (n1938,n1939,n1940);
xor (n1939,n1936,n1937);
or (n1940,n1941,n1944);
and (n1941,n1942,n1943);
xor (n1942,n1900,n1901);
and (n1943,n74,n83);
and (n1944,n1945,n1946);
xor (n1945,n1942,n1943);
or (n1946,n1947,n1950);
and (n1947,n1948,n1949);
xor (n1948,n1906,n1907);
and (n1949,n102,n83);
and (n1950,n1951,n1952);
xor (n1951,n1948,n1949);
or (n1952,n1953,n1956);
and (n1953,n1954,n1955);
xor (n1954,n1912,n1913);
and (n1955,n96,n83);
and (n1956,n1957,n1958);
xor (n1957,n1954,n1955);
and (n1958,n1959,n1960);
xor (n1959,n1918,n1919);
and (n1960,n196,n83);
and (n1961,n27,n89);
or (n1962,n1963,n1966);
and (n1963,n1964,n1965);
xor (n1964,n1927,n1928);
and (n1965,n33,n89);
and (n1966,n1967,n1968);
xor (n1967,n1964,n1965);
or (n1968,n1969,n1972);
and (n1969,n1970,n1971);
xor (n1970,n1933,n1934);
and (n1971,n75,n89);
and (n1972,n1973,n1974);
xor (n1973,n1970,n1971);
or (n1974,n1975,n1977);
and (n1975,n1976,n202);
xor (n1976,n1939,n1940);
and (n1977,n1978,n1979);
xor (n1978,n1976,n202);
or (n1979,n1980,n1983);
and (n1980,n1981,n1982);
xor (n1981,n1945,n1946);
and (n1982,n102,n89);
and (n1983,n1984,n1985);
xor (n1984,n1981,n1982);
or (n1985,n1986,n1989);
and (n1986,n1987,n1988);
xor (n1987,n1951,n1952);
and (n1988,n96,n89);
and (n1989,n1990,n1991);
xor (n1990,n1987,n1988);
and (n1991,n1992,n1993);
xor (n1992,n1957,n1958);
and (n1993,n196,n89);
and (n1994,n33,n111);
or (n1995,n1996,n1999);
and (n1996,n1997,n1998);
xor (n1997,n1967,n1968);
and (n1998,n75,n111);
and (n1999,n2000,n2001);
xor (n2000,n1997,n1998);
or (n2001,n2002,n2004);
and (n2002,n2003,n112);
xor (n2003,n1973,n1974);
and (n2004,n2005,n2006);
xor (n2005,n2003,n112);
or (n2006,n2007,n2010);
and (n2007,n2008,n2009);
xor (n2008,n1978,n1979);
and (n2009,n102,n111);
and (n2010,n2011,n2012);
xor (n2011,n2008,n2009);
or (n2012,n2013,n2015);
and (n2013,n2014,n262);
xor (n2014,n1984,n1985);
and (n2015,n2016,n2017);
xor (n2016,n2014,n262);
and (n2017,n2018,n2019);
xor (n2018,n1990,n1991);
and (n2019,n196,n111);
and (n2020,n75,n118);
or (n2021,n2022,n2025);
and (n2022,n2023,n2024);
xor (n2023,n2000,n2001);
and (n2024,n74,n118);
and (n2025,n2026,n2027);
xor (n2026,n2023,n2024);
or (n2027,n2028,n2031);
and (n2028,n2029,n2030);
xor (n2029,n2005,n2006);
and (n2030,n102,n118);
and (n2031,n2032,n2033);
xor (n2032,n2029,n2030);
or (n2033,n2034,n2037);
and (n2034,n2035,n2036);
xor (n2035,n2011,n2012);
and (n2036,n96,n118);
and (n2037,n2038,n2039);
xor (n2038,n2035,n2036);
and (n2039,n2040,n2041);
xor (n2040,n2016,n2017);
and (n2041,n196,n118);
endmodule
