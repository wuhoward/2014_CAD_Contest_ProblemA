module top (out,n19,n24,n25,n26,n28,n29,n40,n43,n46
        ,n49,n52,n55,n58,n61,n64,n67,n70,n73,n76
        ,n79,n82,n85,n88,n91,n94,n97,n100,n103,n106
        ,n108,n111,n119,n145,n150,n153,n156,n159,n162,n165
        ,n168,n171,n174,n177,n180,n183,n186,n189,n192,n195
        ,n198,n201,n204,n207,n210,n218,n578,n617,n622,n634
        ,n1052,n1077);
output out;
input n19;
input n24;
input n25;
input n26;
input n28;
input n29;
input n40;
input n43;
input n46;
input n49;
input n52;
input n55;
input n58;
input n61;
input n64;
input n67;
input n70;
input n73;
input n76;
input n79;
input n82;
input n85;
input n88;
input n91;
input n94;
input n97;
input n100;
input n103;
input n106;
input n108;
input n111;
input n119;
input n145;
input n150;
input n153;
input n156;
input n159;
input n162;
input n165;
input n168;
input n171;
input n174;
input n177;
input n180;
input n183;
input n186;
input n189;
input n192;
input n195;
input n198;
input n201;
input n204;
input n207;
input n210;
input n218;
input n578;
input n617;
input n622;
input n634;
input n1052;
input n1077;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n20;
wire n21;
wire n22;
wire n23;
wire n27;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n41;
wire n42;
wire n44;
wire n45;
wire n47;
wire n48;
wire n50;
wire n51;
wire n53;
wire n54;
wire n56;
wire n57;
wire n59;
wire n60;
wire n62;
wire n63;
wire n65;
wire n66;
wire n68;
wire n69;
wire n71;
wire n72;
wire n74;
wire n75;
wire n77;
wire n78;
wire n80;
wire n81;
wire n83;
wire n84;
wire n86;
wire n87;
wire n89;
wire n90;
wire n92;
wire n93;
wire n95;
wire n96;
wire n98;
wire n99;
wire n101;
wire n102;
wire n104;
wire n105;
wire n107;
wire n109;
wire n110;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n146;
wire n147;
wire n148;
wire n149;
wire n151;
wire n152;
wire n154;
wire n155;
wire n157;
wire n158;
wire n160;
wire n161;
wire n163;
wire n164;
wire n166;
wire n167;
wire n169;
wire n170;
wire n172;
wire n173;
wire n175;
wire n176;
wire n178;
wire n179;
wire n181;
wire n182;
wire n184;
wire n185;
wire n187;
wire n188;
wire n190;
wire n191;
wire n193;
wire n194;
wire n196;
wire n197;
wire n199;
wire n200;
wire n202;
wire n203;
wire n205;
wire n206;
wire n208;
wire n209;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n618;
wire n619;
wire n620;
wire n621;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2988;
wire n2989;
wire n2990;
wire n2991;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2996;
wire n2997;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3003;
wire n3004;
wire n3005;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3010;
wire n3011;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3038;
wire n3039;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
wire n3056;
wire n3057;
wire n3058;
wire n3059;
wire n3060;
wire n3061;
wire n3062;
wire n3063;
wire n3064;
wire n3065;
wire n3066;
wire n3067;
wire n3068;
wire n3069;
wire n3070;
wire n3071;
wire n3072;
wire n3073;
wire n3074;
wire n3075;
wire n3076;
wire n3077;
wire n3078;
wire n3079;
wire n3080;
wire n3081;
wire n3082;
wire n3083;
wire n3084;
wire n3085;
wire n3086;
wire n3087;
wire n3088;
wire n3089;
wire n3090;
wire n3091;
wire n3092;
wire n3093;
wire n3094;
wire n3095;
wire n3096;
wire n3097;
wire n3098;
wire n3099;
wire n3100;
wire n3101;
wire n3102;
wire n3103;
wire n3104;
wire n3105;
wire n3106;
wire n3107;
wire n3108;
wire n3109;
wire n3110;
wire n3111;
wire n3112;
wire n3113;
wire n3114;
wire n3115;
wire n3116;
wire n3117;
wire n3118;
wire n3119;
wire n3120;
wire n3121;
wire n3122;
wire n3123;
wire n3124;
wire n3125;
wire n3126;
wire n3127;
wire n3128;
wire n3129;
wire n3130;
wire n3131;
wire n3132;
wire n3133;
wire n3134;
wire n3135;
wire n3136;
wire n3137;
wire n3138;
wire n3139;
wire n3140;
wire n3141;
wire n3142;
wire n3143;
wire n3144;
wire n3145;
wire n3146;
wire n3147;
wire n3148;
wire n3149;
wire n3150;
wire n3151;
wire n3152;
wire n3153;
wire n3154;
wire n3155;
wire n3156;
wire n3157;
wire n3158;
wire n3159;
wire n3160;
wire n3161;
wire n3162;
wire n3163;
wire n3164;
wire n3165;
wire n3166;
wire n3167;
wire n3168;
wire n3169;
wire n3170;
wire n3171;
wire n3172;
wire n3173;
wire n3174;
wire n3175;
wire n3176;
wire n3177;
wire n3178;
wire n3179;
wire n3180;
wire n3181;
wire n3182;
wire n3183;
wire n3184;
wire n3185;
wire n3186;
wire n3187;
wire n3188;
wire n3189;
wire n3190;
wire n3191;
wire n3192;
wire n3193;
wire n3194;
wire n3195;
wire n3196;
wire n3197;
wire n3198;
wire n3199;
wire n3200;
wire n3201;
wire n3202;
wire n3203;
wire n3204;
wire n3205;
wire n3206;
wire n3207;
wire n3208;
wire n3209;
wire n3210;
wire n3211;
wire n3212;
wire n3213;
wire n3214;
wire n3215;
wire n3216;
wire n3217;
wire n3218;
wire n3219;
wire n3220;
wire n3221;
wire n3222;
wire n3223;
wire n3224;
wire n3225;
wire n3226;
wire n3227;
wire n3228;
wire n3229;
wire n3230;
wire n3231;
wire n3232;
wire n3233;
wire n3234;
wire n3235;
wire n3236;
wire n3237;
wire n3238;
wire n3239;
wire n3240;
wire n3241;
wire n3242;
wire n3243;
wire n3244;
wire n3245;
wire n3246;
wire n3247;
wire n3248;
wire n3249;
wire n3250;
wire n3251;
wire n3252;
wire n3253;
wire n3254;
wire n3255;
wire n3256;
wire n3257;
wire n3258;
wire n3259;
wire n3260;
wire n3261;
wire n3262;
wire n3263;
wire n3264;
wire n3265;
wire n3266;
wire n3267;
wire n3268;
wire n3269;
wire n3270;
wire n3271;
wire n3272;
wire n3273;
wire n3274;
wire n3275;
wire n3276;
wire n3277;
wire n3278;
wire n3279;
wire n3280;
wire n3281;
wire n3282;
wire n3283;
wire n3284;
wire n3285;
wire n3286;
wire n3287;
wire n3288;
wire n3289;
wire n3290;
wire n3291;
wire n3292;
wire n3293;
wire n3294;
wire n3295;
wire n3296;
wire n3297;
wire n3298;
wire n3299;
wire n3300;
wire n3301;
wire n3302;
wire n3303;
wire n3304;
wire n3305;
wire n3306;
wire n3307;
wire n3308;
wire n3309;
wire n3310;
wire n3311;
wire n3312;
wire n3313;
wire n3314;
wire n3315;
wire n3316;
wire n3317;
wire n3318;
wire n3319;
wire n3320;
wire n3321;
wire n3322;
wire n3323;
wire n3324;
wire n3325;
wire n3326;
wire n3327;
wire n3328;
wire n3329;
wire n3330;
wire n3331;
wire n3332;
wire n3333;
wire n3334;
wire n3335;
wire n3336;
wire n3337;
wire n3338;
wire n3339;
wire n3340;
wire n3341;
wire n3342;
wire n3343;
wire n3344;
wire n3345;
wire n3346;
wire n3347;
wire n3348;
wire n3349;
wire n3350;
wire n3351;
wire n3352;
wire n3353;
wire n3354;
wire n3355;
wire n3356;
wire n3357;
wire n3358;
wire n3359;
wire n3360;
wire n3361;
wire n3362;
wire n3363;
wire n3364;
wire n3365;
wire n3366;
wire n3367;
wire n3368;
wire n3369;
wire n3370;
wire n3371;
wire n3372;
wire n3373;
wire n3374;
wire n3375;
wire n3376;
wire n3377;
wire n3378;
wire n3379;
wire n3380;
wire n3381;
wire n3382;
wire n3383;
wire n3384;
wire n3385;
wire n3386;
wire n3387;
wire n3388;
wire n3389;
wire n3390;
wire n3391;
wire n3392;
wire n3393;
wire n3394;
wire n3395;
wire n3396;
wire n3397;
wire n3398;
wire n3399;
wire n3400;
wire n3401;
wire n3402;
wire n3403;
wire n3404;
wire n3405;
wire n3406;
wire n3407;
wire n3408;
wire n3409;
wire n3410;
wire n3411;
wire n3412;
wire n3413;
wire n3414;
wire n3415;
wire n3416;
wire n3417;
wire n3418;
wire n3419;
wire n3420;
wire n3421;
wire n3422;
wire n3423;
wire n3424;
wire n3425;
wire n3426;
wire n3427;
wire n3428;
wire n3429;
wire n3430;
wire n3431;
wire n3432;
wire n3433;
wire n3434;
wire n3435;
wire n3436;
wire n3437;
wire n3438;
wire n3439;
wire n3440;
wire n3441;
wire n3442;
wire n3443;
wire n3444;
wire n3445;
wire n3446;
wire n3447;
wire n3448;
wire n3449;
wire n3450;
wire n3451;
wire n3452;
wire n3453;
wire n3454;
wire n3455;
wire n3456;
wire n3457;
wire n3458;
wire n3459;
wire n3460;
wire n3461;
wire n3462;
wire n3463;
wire n3464;
wire n3465;
wire n3466;
wire n3467;
wire n3468;
wire n3469;
wire n3470;
wire n3471;
wire n3472;
wire n3473;
wire n3474;
wire n3475;
wire n3476;
wire n3477;
wire n3478;
wire n3479;
wire n3480;
wire n3481;
wire n3482;
wire n3483;
wire n3484;
wire n3485;
wire n3486;
wire n3487;
wire n3488;
wire n3489;
wire n3490;
wire n3491;
wire n3492;
wire n3493;
wire n3494;
wire n3495;
wire n3496;
wire n3497;
wire n3498;
wire n3499;
wire n3500;
wire n3501;
wire n3502;
wire n3503;
wire n3504;
wire n3505;
wire n3506;
wire n3507;
wire n3508;
wire n3509;
wire n3510;
wire n3511;
wire n3512;
wire n3513;
wire n3514;
wire n3515;
wire n3516;
wire n3517;
wire n3518;
wire n3519;
wire n3520;
wire n3521;
wire n3522;
wire n3523;
wire n3524;
wire n3525;
wire n3526;
wire n3527;
wire n3528;
wire n3529;
wire n3530;
wire n3531;
wire n3532;
wire n3533;
wire n3534;
wire n3535;
wire n3536;
wire n3537;
wire n3538;
wire n3539;
wire n3540;
wire n3541;
wire n3542;
wire n3543;
wire n3544;
wire n3545;
wire n3546;
wire n3547;
wire n3548;
wire n3549;
wire n3550;
wire n3551;
wire n3552;
wire n3553;
wire n3554;
wire n3555;
wire n3556;
wire n3557;
wire n3558;
wire n3559;
wire n3560;
wire n3561;
wire n3562;
wire n3563;
wire n3564;
wire n3565;
wire n3566;
wire n3567;
wire n3568;
wire n3569;
wire n3570;
wire n3571;
wire n3572;
wire n3573;
wire n3574;
wire n3575;
wire n3576;
wire n3577;
wire n3578;
wire n3579;
wire n3580;
wire n3581;
wire n3582;
wire n3583;
wire n3584;
wire n3585;
wire n3586;
wire n3587;
wire n3588;
wire n3589;
wire n3590;
wire n3591;
wire n3592;
wire n3593;
wire n3594;
wire n3595;
wire n3596;
wire n3597;
wire n3598;
wire n3599;
wire n3600;
wire n3601;
wire n3602;
wire n3603;
wire n3604;
wire n3605;
wire n3606;
wire n3607;
wire n3608;
wire n3609;
wire n3610;
wire n3611;
wire n3612;
wire n3613;
wire n3614;
wire n3615;
wire n3616;
wire n3617;
wire n3618;
wire n3619;
wire n3620;
wire n3621;
wire n3622;
wire n3623;
wire n3624;
wire n3625;
wire n3626;
wire n3627;
wire n3628;
wire n3629;
wire n3630;
wire n3631;
wire n3632;
wire n3633;
wire n3634;
wire n3635;
wire n3636;
wire n3637;
wire n3638;
wire n3639;
wire n3640;
wire n3641;
wire n3642;
wire n3643;
wire n3644;
wire n3645;
wire n3646;
wire n3647;
wire n3648;
wire n3649;
wire n3650;
wire n3651;
wire n3652;
wire n3653;
wire n3654;
wire n3655;
wire n3656;
wire n3657;
wire n3658;
wire n3659;
wire n3660;
wire n3661;
wire n3662;
wire n3663;
wire n3664;
wire n3665;
wire n3666;
wire n3667;
wire n3668;
wire n3669;
wire n3670;
wire n3671;
wire n3672;
wire n3673;
wire n3674;
wire n3675;
wire n3676;
wire n3677;
wire n3678;
wire n3679;
wire n3680;
wire n3681;
wire n3682;
wire n3683;
wire n3684;
wire n3685;
wire n3686;
wire n3687;
wire n3688;
wire n3689;
wire n3690;
wire n3691;
wire n3692;
wire n3693;
wire n3694;
wire n3695;
wire n3696;
wire n3697;
wire n3698;
wire n3699;
wire n3700;
wire n3701;
wire n3702;
wire n3703;
wire n3704;
wire n3705;
wire n3706;
wire n3707;
wire n3708;
wire n3709;
wire n3710;
wire n3711;
wire n3712;
wire n3713;
wire n3714;
wire n3715;
wire n3716;
wire n3717;
wire n3718;
wire n3719;
wire n3720;
wire n3721;
wire n3722;
wire n3723;
wire n3724;
wire n3725;
wire n3726;
wire n3727;
wire n3728;
wire n3729;
wire n3730;
wire n3731;
wire n3732;
wire n3733;
wire n3734;
wire n3735;
wire n3736;
wire n3737;
wire n3738;
wire n3739;
wire n3740;
wire n3741;
wire n3742;
wire n3743;
wire n3744;
wire n3745;
wire n3746;
wire n3747;
wire n3748;
wire n3749;
wire n3750;
wire n3751;
wire n3752;
wire n3753;
wire n3754;
wire n3755;
wire n3756;
wire n3757;
wire n3758;
wire n3759;
wire n3760;
wire n3761;
wire n3762;
wire n3763;
wire n3764;
wire n3765;
wire n3766;
wire n3767;
wire n3768;
wire n3769;
wire n3770;
wire n3771;
wire n3772;
wire n3773;
wire n3774;
wire n3775;
wire n3776;
wire n3777;
wire n3778;
wire n3779;
wire n3780;
wire n3781;
wire n3782;
wire n3783;
wire n3784;
wire n3785;
wire n3786;
wire n3787;
wire n3788;
wire n3789;
wire n3790;
wire n3791;
wire n3792;
wire n3793;
wire n3794;
wire n3795;
wire n3796;
wire n3797;
wire n3798;
wire n3799;
wire n3800;
wire n3801;
wire n3802;
wire n3803;
wire n3804;
wire n3805;
wire n3806;
wire n3807;
wire n3808;
wire n3809;
wire n3810;
wire n3811;
wire n3812;
wire n3813;
wire n3814;
wire n3815;
wire n3816;
wire n3817;
wire n3818;
wire n3819;
wire n3820;
wire n3821;
wire n3822;
wire n3823;
wire n3824;
wire n3825;
wire n3826;
wire n3827;
wire n3828;
wire n3829;
wire n3830;
wire n3831;
wire n3832;
wire n3833;
wire n3834;
wire n3835;
wire n3836;
wire n3837;
wire n3838;
wire n3839;
wire n3840;
wire n3841;
wire n3842;
wire n3843;
wire n3844;
wire n3845;
wire n3846;
wire n3847;
wire n3848;
wire n3849;
wire n3850;
wire n3851;
wire n3852;
wire n3853;
wire n3854;
wire n3855;
wire n3856;
wire n3857;
wire n3858;
wire n3859;
wire n3860;
wire n3861;
wire n3862;
wire n3863;
wire n3864;
wire n3865;
wire n3866;
wire n3867;
wire n3868;
wire n3869;
wire n3870;
wire n3871;
wire n3872;
wire n3873;
wire n3874;
wire n3875;
wire n3876;
wire n3877;
wire n3878;
wire n3879;
wire n3880;
wire n3881;
wire n3882;
wire n3883;
wire n3884;
wire n3885;
wire n3886;
wire n3887;
wire n3888;
wire n3889;
wire n3890;
wire n3891;
wire n3892;
wire n3893;
wire n3894;
wire n3895;
wire n3896;
wire n3897;
wire n3898;
wire n3899;
wire n3900;
wire n3901;
wire n3902;
wire n3903;
wire n3904;
wire n3905;
wire n3906;
wire n3907;
wire n3908;
wire n3909;
wire n3910;
wire n3911;
wire n3912;
wire n3913;
wire n3914;
wire n3915;
wire n3916;
wire n3917;
wire n3918;
wire n3919;
wire n3920;
wire n3921;
wire n3922;
wire n3923;
wire n3924;
wire n3925;
wire n3926;
wire n3927;
wire n3928;
wire n3929;
wire n3930;
wire n3931;
wire n3932;
wire n3933;
wire n3934;
wire n3935;
wire n3936;
wire n3937;
wire n3938;
wire n3939;
wire n3940;
wire n3941;
wire n3942;
wire n3943;
wire n3944;
wire n3945;
wire n3946;
wire n3947;
wire n3948;
wire n3949;
wire n3950;
wire n3951;
wire n3952;
wire n3953;
wire n3954;
wire n3955;
wire n3956;
wire n3957;
wire n3958;
wire n3959;
wire n3960;
wire n3961;
wire n3962;
wire n3963;
wire n3964;
wire n3965;
wire n3966;
wire n3967;
wire n3968;
wire n3969;
wire n3970;
wire n3971;
wire n3972;
wire n3973;
wire n3974;
wire n3975;
wire n3976;
wire n3977;
wire n3978;
wire n3979;
wire n3980;
wire n3981;
wire n3982;
wire n3983;
wire n3984;
wire n3985;
wire n3986;
wire n3987;
wire n3988;
wire n3989;
wire n3990;
wire n3991;
wire n3992;
wire n3993;
wire n3994;
wire n3995;
wire n3996;
wire n3997;
wire n3998;
wire n3999;
wire n4000;
wire n4001;
wire n4002;
wire n4003;
wire n4004;
wire n4005;
wire n4006;
wire n4007;
wire n4008;
wire n4009;
wire n4010;
wire n4011;
wire n4012;
wire n4013;
wire n4014;
wire n4015;
wire n4016;
wire n4017;
wire n4018;
wire n4019;
wire n4020;
wire n4021;
wire n4022;
wire n4023;
wire n4024;
wire n4025;
wire n4026;
wire n4027;
wire n4028;
wire n4029;
wire n4030;
wire n4031;
wire n4032;
wire n4033;
wire n4034;
wire n4035;
wire n4036;
wire n4037;
wire n4038;
wire n4039;
wire n4040;
wire n4041;
wire n4042;
wire n4043;
wire n4044;
wire n4045;
wire n4046;
wire n4047;
wire n4048;
wire n4049;
wire n4050;
wire n4051;
wire n4052;
wire n4053;
wire n4054;
wire n4055;
wire n4056;
wire n4057;
wire n4058;
wire n4059;
wire n4060;
wire n4061;
wire n4062;
wire n4063;
wire n4064;
wire n4065;
wire n4066;
wire n4067;
wire n4068;
wire n4069;
wire n4070;
wire n4071;
wire n4072;
wire n4073;
wire n4074;
wire n4075;
wire n4076;
wire n4077;
wire n4078;
wire n4079;
wire n4080;
wire n4081;
wire n4082;
wire n4083;
wire n4084;
wire n4085;
wire n4086;
wire n4087;
wire n4088;
wire n4089;
wire n4090;
wire n4091;
wire n4092;
wire n4093;
wire n4094;
wire n4095;
wire n4096;
wire n4097;
wire n4098;
wire n4099;
wire n4100;
wire n4101;
wire n4102;
wire n4103;
wire n4104;
wire n4105;
wire n4106;
wire n4107;
wire n4108;
wire n4109;
wire n4110;
wire n4111;
wire n4112;
wire n4113;
wire n4114;
wire n4115;
wire n4116;
wire n4117;
wire n4118;
wire n4119;
wire n4120;
wire n4121;
wire n4122;
wire n4123;
wire n4124;
wire n4125;
wire n4126;
wire n4127;
wire n4128;
wire n4129;
wire n4130;
wire n4131;
wire n4132;
wire n4133;
wire n4134;
wire n4135;
wire n4136;
wire n4137;
wire n4138;
wire n4139;
wire n4140;
wire n4141;
wire n4142;
wire n4143;
wire n4144;
wire n4145;
wire n4146;
wire n4147;
wire n4148;
wire n4149;
wire n4150;
wire n4151;
wire n4152;
wire n4153;
wire n4154;
wire n4155;
wire n4156;
wire n4157;
wire n4158;
wire n4159;
wire n4160;
wire n4161;
wire n4162;
wire n4163;
wire n4164;
wire n4165;
wire n4166;
wire n4167;
wire n4168;
wire n4169;
wire n4170;
wire n4171;
wire n4172;
wire n4173;
wire n4174;
wire n4175;
wire n4176;
wire n4177;
wire n4178;
wire n4179;
wire n4180;
wire n4181;
wire n4182;
wire n4183;
wire n4184;
wire n4185;
wire n4186;
wire n4187;
wire n4188;
wire n4189;
wire n4190;
wire n4191;
wire n4192;
wire n4193;
wire n4194;
wire n4195;
wire n4196;
wire n4197;
wire n4198;
wire n4199;
wire n4200;
wire n4201;
wire n4202;
wire n4203;
wire n4204;
wire n4205;
wire n4206;
wire n4207;
wire n4208;
wire n4209;
wire n4210;
wire n4211;
wire n4212;
wire n4213;
wire n4214;
wire n4215;
wire n4216;
wire n4217;
wire n4218;
wire n4219;
wire n4220;
wire n4221;
wire n4222;
wire n4223;
wire n4224;
wire n4225;
wire n4226;
wire n4227;
wire n4228;
wire n4229;
wire n4230;
wire n4231;
wire n4232;
wire n4233;
wire n4234;
wire n4235;
wire n4236;
wire n4237;
wire n4238;
wire n4239;
wire n4240;
wire n4241;
wire n4242;
wire n4243;
wire n4244;
wire n4245;
wire n4246;
wire n4247;
wire n4248;
wire n4249;
wire n4250;
wire n4251;
wire n4252;
wire n4253;
wire n4254;
wire n4255;
wire n4256;
wire n4257;
wire n4258;
wire n4259;
wire n4260;
wire n4261;
wire n4262;
wire n4263;
wire n4264;
wire n4265;
wire n4266;
wire n4267;
wire n4268;
wire n4269;
wire n4270;
wire n4271;
wire n4272;
wire n4273;
wire n4274;
wire n4275;
wire n4276;
wire n4277;
wire n4278;
wire n4279;
wire n4280;
wire n4281;
wire n4282;
wire n4283;
wire n4284;
wire n4285;
wire n4286;
wire n4287;
wire n4288;
wire n4289;
wire n4290;
wire n4291;
wire n4292;
wire n4293;
wire n4294;
wire n4295;
wire n4296;
wire n4297;
wire n4298;
wire n4299;
wire n4300;
wire n4301;
wire n4302;
wire n4303;
wire n4304;
wire n4305;
wire n4306;
wire n4307;
wire n4308;
wire n4309;
wire n4310;
wire n4311;
wire n4312;
wire n4313;
wire n4314;
wire n4315;
wire n4316;
wire n4317;
wire n4318;
wire n4319;
wire n4320;
wire n4321;
wire n4322;
wire n4323;
wire n4324;
wire n4325;
wire n4326;
wire n4327;
wire n4328;
wire n4329;
wire n4330;
wire n4331;
wire n4332;
wire n4333;
wire n4334;
wire n4335;
wire n4336;
wire n4337;
wire n4338;
wire n4339;
wire n4340;
wire n4341;
wire n4342;
wire n4343;
wire n4344;
wire n4345;
wire n4346;
wire n4347;
wire n4348;
wire n4349;
wire n4350;
wire n4351;
wire n4352;
wire n4353;
wire n4354;
wire n4355;
wire n4356;
wire n4357;
wire n4358;
wire n4359;
wire n4360;
wire n4361;
wire n4362;
wire n4363;
wire n4364;
wire n4365;
wire n4366;
wire n4367;
wire n4368;
wire n4369;
wire n4370;
wire n4371;
wire n4372;
wire n4373;
wire n4374;
wire n4375;
wire n4376;
wire n4377;
wire n4378;
wire n4379;
wire n4380;
wire n4381;
wire n4382;
wire n4383;
wire n4384;
wire n4385;
wire n4386;
wire n4387;
wire n4388;
wire n4389;
wire n4390;
wire n4391;
wire n4392;
wire n4393;
wire n4394;
wire n4395;
wire n4396;
wire n4397;
wire n4398;
wire n4399;
wire n4400;
wire n4401;
wire n4402;
wire n4403;
wire n4404;
wire n4405;
wire n4406;
wire n4407;
wire n4408;
wire n4409;
wire n4410;
wire n4411;
wire n4412;
wire n4413;
wire n4414;
wire n4415;
wire n4416;
wire n4417;
wire n4418;
wire n4419;
wire n4420;
wire n4421;
wire n4422;
wire n4423;
wire n4424;
wire n4425;
wire n4426;
wire n4427;
wire n4428;
wire n4429;
wire n4430;
wire n4431;
wire n4432;
wire n4433;
wire n4434;
wire n4435;
wire n4436;
wire n4437;
wire n4438;
wire n4439;
wire n4440;
wire n4441;
wire n4442;
wire n4443;
wire n4444;
wire n4445;
wire n4446;
wire n4447;
wire n4448;
wire n4449;
wire n4450;
wire n4451;
wire n4452;
wire n4453;
wire n4454;
wire n4455;
wire n4456;
wire n4457;
wire n4458;
wire n4459;
wire n4460;
wire n4461;
wire n4462;
wire n4463;
wire n4464;
wire n4465;
wire n4466;
wire n4467;
wire n4468;
wire n4469;
wire n4470;
wire n4471;
wire n4472;
wire n4473;
wire n4474;
wire n4475;
wire n4476;
wire n4477;
wire n4478;
wire n4479;
wire n4480;
xor (out,n0,n2542);
xor (n0,n1,n1185);
xor (n1,n2,n1034);
or (n2,n3,n1033);
and (n3,n4,n972);
xor (n4,n5,n664);
xor (n5,n6,n595);
xor (n6,n7,n467);
or (n7,n8,n466);
and (n8,n9,n366);
xor (n9,n10,n260);
xor (n10,n11,n224);
xor (n11,n12,n120);
nor (n12,n13,n117);
and (n13,n14,n115);
nand (n14,n15,n112);
not (n15,n16);
wire s0n16,s1n16,notn16;
or (n16,s0n16,s1n16);
not(notn16,n109);
and (s0n16,notn16,n17);
and (s1n16,n109,n36);
wire s0n17,s1n17,notn17;
or (n17,s0n17,s1n17);
not(notn17,n20);
and (s0n17,notn17,1'b0);
and (s1n17,n20,n19);
or (n20,n21,n32);
or (n21,n22,n30);
nor (n22,n23,n25,n26,n27,n29);
not (n23,n24);
not (n27,n28);
nor (n30,n24,n31,n26,n27,n29);
not (n31,n25);
or (n32,n33,n35);
and (n33,n23,n25,n26,n27,n34);
not (n34,n29);
nor (n35,n23,n31,n26,n27,n29);
xor (n36,n37,n38);
not (n37,n19);
and (n38,n39,n41);
not (n39,n40);
and (n41,n42,n44);
not (n42,n43);
and (n44,n45,n47);
not (n45,n46);
and (n47,n48,n50);
not (n48,n49);
and (n50,n51,n53);
not (n51,n52);
and (n53,n54,n56);
not (n54,n55);
and (n56,n57,n59);
not (n57,n58);
and (n59,n60,n62);
not (n60,n61);
and (n62,n63,n65);
not (n63,n64);
and (n65,n66,n68);
not (n66,n67);
and (n68,n69,n71);
not (n69,n70);
and (n71,n72,n74);
not (n72,n73);
and (n74,n75,n77);
not (n75,n76);
and (n77,n78,n80);
not (n78,n79);
and (n80,n81,n83);
not (n81,n82);
and (n83,n84,n86);
not (n84,n85);
and (n86,n87,n89);
not (n87,n88);
and (n89,n90,n92);
not (n90,n91);
and (n92,n93,n95);
not (n93,n94);
and (n95,n96,n98);
not (n96,n97);
and (n98,n99,n101);
not (n99,n100);
and (n101,n102,n104);
not (n102,n103);
and (n104,n105,n107);
not (n105,n106);
not (n107,n108);
and (n109,n110,n111);
or (n110,n22,n33);
wire s0n112,s1n112,notn112;
or (n112,s0n112,s1n112);
not(notn112,n109);
and (s0n112,notn112,n113);
and (s1n112,n109,n114);
wire s0n113,s1n113,notn113;
or (n113,s0n113,s1n113);
not(notn113,n20);
and (s0n113,notn113,1'b0);
and (s1n113,n20,n40);
xor (n114,n39,n41);
nand (n115,n16,n116);
not (n116,n112);
not (n117,n118);
wire s0n118,s1n118,notn118;
or (n118,s0n118,s1n118);
not(notn118,n20);
and (s0n118,notn118,1'b0);
and (s1n118,n20,n119);
nand (n120,n121,n213);
or (n121,n122,n141);
nand (n122,n123,n134);
nor (n123,n124,n132);
and (n124,n125,n129);
not (n125,n126);
wire s0n126,s1n126,notn126;
or (n126,s0n126,s1n126);
not(notn126,n109);
and (s0n126,notn126,n127);
and (s1n126,n109,n128);
wire s0n127,s1n127,notn127;
or (n127,s0n127,s1n127);
not(notn127,n20);
and (s0n127,notn127,1'b0);
and (s1n127,n20,n106);
xor (n128,n105,n107);
wire s0n129,s1n129,notn129;
or (n129,s0n129,s1n129);
not(notn129,n109);
and (s0n129,notn129,n130);
and (s1n129,n109,n131);
wire s0n130,s1n130,notn130;
or (n130,s0n130,s1n130);
not(notn130,n20);
and (s0n130,notn130,1'b0);
and (s1n130,n20,n103);
xor (n131,n102,n104);
and (n132,n126,n133);
not (n133,n129);
nand (n134,n135,n140);
or (n135,n136,n129);
not (n136,n137);
wire s0n137,s1n137,notn137;
or (n137,s0n137,s1n137);
not(notn137,n109);
and (s0n137,notn137,n138);
and (s1n137,n109,n139);
wire s0n138,s1n138,notn138;
or (n138,s0n138,s1n138);
not(notn138,n20);
and (s0n138,notn138,1'b0);
and (s1n138,n20,n100);
xor (n139,n99,n101);
nand (n140,n136,n129);
nor (n141,n142,n211);
and (n142,n143,n136);
wire s0n143,s1n143,notn143;
or (n143,s0n143,s1n143);
not(notn143,n209);
and (s0n143,notn143,n144);
and (s1n143,n209,n146);
wire s0n144,s1n144,notn144;
or (n144,s0n144,s1n144);
not(notn144,n20);
and (s0n144,notn144,1'b0);
and (s1n144,n20,n145);
xor (n146,n147,n148);
not (n147,n145);
and (n148,n149,n151);
not (n149,n150);
and (n151,n152,n154);
not (n152,n153);
and (n154,n155,n157);
not (n155,n156);
and (n157,n158,n160);
not (n158,n159);
and (n160,n161,n163);
not (n161,n162);
and (n163,n164,n166);
not (n164,n165);
and (n166,n167,n169);
not (n167,n168);
and (n169,n170,n172);
not (n170,n171);
and (n172,n173,n175);
not (n173,n174);
and (n175,n176,n178);
not (n176,n177);
and (n178,n179,n181);
not (n179,n180);
and (n181,n182,n184);
not (n182,n183);
and (n184,n185,n187);
not (n185,n186);
and (n187,n188,n190);
not (n188,n189);
and (n190,n191,n193);
not (n191,n192);
and (n193,n194,n196);
not (n194,n195);
and (n196,n197,n199);
not (n197,n198);
and (n199,n200,n202);
not (n200,n201);
and (n202,n203,n205);
not (n203,n204);
and (n205,n206,n208);
not (n206,n207);
not (n208,n119);
and (n209,n110,n210);
and (n211,n212,n137);
not (n212,n143);
or (n213,n123,n214);
nor (n214,n215,n222);
and (n215,n216,n136);
wire s0n216,s1n216,notn216;
or (n216,s0n216,s1n216);
not(notn216,n209);
and (s0n216,notn216,n217);
and (s1n216,n209,n219);
wire s0n217,s1n217,notn217;
or (n217,s0n217,s1n217);
not(notn217,n20);
and (s0n217,notn217,1'b0);
and (s1n217,n20,n218);
xor (n219,n220,n221);
not (n220,n218);
and (n221,n147,n148);
and (n222,n223,n137);
not (n223,n216);
nand (n224,n225,n252);
or (n225,n226,n245);
nand (n226,n227,n238);
or (n227,n228,n235);
and (n228,n229,n232);
wire s0n229,s1n229,notn229;
or (n229,s0n229,s1n229);
not(notn229,n109);
and (s0n229,notn229,n230);
and (s1n229,n109,n231);
wire s0n230,s1n230,notn230;
or (n230,s0n230,s1n230);
not(notn230,n20);
and (s0n230,notn230,1'b0);
and (s1n230,n20,n94);
xor (n231,n93,n95);
wire s0n232,s1n232,notn232;
or (n232,s0n232,s1n232);
not(notn232,n109);
and (s0n232,notn232,n233);
and (s1n232,n109,n234);
wire s0n233,s1n233,notn233;
or (n233,s0n233,s1n233);
not(notn233,n20);
and (s0n233,notn233,1'b0);
and (s1n233,n20,n91);
xor (n234,n90,n92);
and (n235,n236,n237);
not (n236,n229);
not (n237,n232);
nor (n238,n239,n243);
and (n239,n240,n232);
wire s0n240,s1n240,notn240;
or (n240,s0n240,s1n240);
not(notn240,n109);
and (s0n240,notn240,n241);
and (s1n240,n109,n242);
wire s0n241,s1n241,notn241;
or (n241,s0n241,s1n241);
not(notn241,n20);
and (s0n241,notn241,1'b0);
and (s1n241,n20,n88);
xor (n242,n87,n89);
and (n243,n244,n237);
not (n244,n240);
nor (n245,n246,n250);
and (n246,n247,n244);
wire s0n247,s1n247,notn247;
or (n247,s0n247,s1n247);
not(notn247,n209);
and (s0n247,notn247,n248);
and (s1n247,n209,n249);
wire s0n248,s1n248,notn248;
or (n248,s0n248,s1n248);
not(notn248,n20);
and (s0n248,notn248,1'b0);
and (s1n248,n20,n159);
xor (n249,n158,n160);
and (n250,n251,n240);
not (n251,n247);
or (n252,n253,n227);
nor (n253,n254,n258);
and (n254,n255,n244);
wire s0n255,s1n255,notn255;
or (n255,s0n255,s1n255);
not(notn255,n209);
and (s0n255,notn255,n256);
and (s1n255,n209,n257);
wire s0n256,s1n256,notn256;
or (n256,s0n256,s1n256);
not(notn256,n20);
and (s0n256,notn256,1'b0);
and (s1n256,n20,n156);
xor (n257,n155,n157);
and (n258,n259,n240);
not (n259,n255);
xor (n260,n261,n333);
xor (n261,n262,n300);
nand (n262,n263,n291);
or (n263,n264,n284);
not (n264,n265);
nor (n265,n266,n276);
nand (n266,n267,n275);
or (n267,n268,n272);
not (n268,n269);
wire s0n269,s1n269,notn269;
or (n269,s0n269,s1n269);
not(notn269,n109);
and (s0n269,notn269,n270);
and (s1n269,n109,n271);
wire s0n270,s1n270,notn270;
or (n270,s0n270,s1n270);
not(notn270,n20);
and (s0n270,notn270,1'b0);
and (s1n270,n20,n70);
xor (n271,n69,n71);
wire s0n272,s1n272,notn272;
or (n272,s0n272,s1n272);
not(notn272,n109);
and (s0n272,notn272,n273);
and (s1n272,n109,n274);
wire s0n273,s1n273,notn273;
or (n273,s0n273,s1n273);
not(notn273,n20);
and (s0n273,notn273,1'b0);
and (s1n273,n20,n67);
xor (n274,n66,n68);
nand (n275,n268,n272);
nor (n276,n277,n282);
and (n277,n278,n272);
not (n278,n279);
wire s0n279,s1n279,notn279;
or (n279,s0n279,s1n279);
not(notn279,n109);
and (s0n279,notn279,n280);
and (s1n279,n109,n281);
wire s0n280,s1n280,notn280;
or (n280,s0n280,s1n280);
not(notn280,n20);
and (s0n280,notn280,1'b0);
and (s1n280,n20,n64);
xor (n281,n63,n65);
and (n282,n283,n279);
not (n283,n272);
nor (n284,n285,n289);
and (n285,n278,n286);
wire s0n286,s1n286,notn286;
or (n286,s0n286,s1n286);
not(notn286,n209);
and (s0n286,notn286,n287);
and (s1n286,n209,n288);
wire s0n287,s1n287,notn287;
or (n287,s0n287,s1n287);
not(notn287,n20);
and (s0n287,notn287,1'b0);
and (s1n287,n20,n183);
xor (n288,n182,n184);
and (n289,n279,n290);
not (n290,n286);
or (n291,n292,n293);
not (n292,n266);
nor (n293,n294,n298);
and (n294,n278,n295);
wire s0n295,s1n295,notn295;
or (n295,s0n295,s1n295);
not(notn295,n209);
and (s0n295,notn295,n296);
and (s1n295,n209,n297);
wire s0n296,s1n296,notn296;
or (n296,s0n296,s1n296);
not(notn296,n20);
and (s0n296,notn296,1'b0);
and (s1n296,n20,n180);
xor (n297,n179,n181);
and (n298,n279,n299);
not (n299,n295);
nand (n300,n301,n325);
or (n301,n302,n318);
not (n302,n303);
and (n303,n304,n311);
nor (n304,n305,n310);
and (n305,n279,n306);
not (n306,n307);
wire s0n307,s1n307,notn307;
or (n307,s0n307,s1n307);
not(notn307,n109);
and (s0n307,notn307,n308);
and (s1n307,n109,n309);
wire s0n308,s1n308,notn308;
or (n308,s0n308,s1n308);
not(notn308,n20);
and (s0n308,notn308,1'b0);
and (s1n308,n20,n61);
xor (n309,n60,n62);
and (n310,n278,n307);
nand (n311,n312,n316);
or (n312,n306,n313);
wire s0n313,s1n313,notn313;
or (n313,s0n313,s1n313);
not(notn313,n109);
and (s0n313,notn313,n314);
and (s1n313,n109,n315);
wire s0n314,s1n314,notn314;
or (n314,s0n314,s1n314);
not(notn314,n20);
and (s0n314,notn314,1'b0);
and (s1n314,n20,n58);
xor (n315,n57,n59);
or (n316,n317,n307);
not (n317,n313);
nor (n318,n319,n323);
and (n319,n317,n320);
wire s0n320,s1n320,notn320;
or (n320,s0n320,s1n320);
not(notn320,n209);
and (s0n320,notn320,n321);
and (s1n320,n209,n322);
wire s0n321,s1n321,notn321;
or (n321,s0n321,s1n321);
not(notn321,n20);
and (s0n321,notn321,1'b0);
and (s1n321,n20,n189);
xor (n322,n188,n190);
and (n323,n313,n324);
not (n324,n320);
or (n325,n326,n304);
nor (n326,n327,n331);
and (n327,n317,n328);
wire s0n328,s1n328,notn328;
or (n328,s0n328,s1n328);
not(notn328,n209);
and (s0n328,notn328,n329);
and (s1n328,n209,n330);
wire s0n329,s1n329,notn329;
or (n329,s0n329,s1n329);
not(notn329,n20);
and (s0n329,notn329,1'b0);
and (s1n329,n20,n186);
xor (n330,n185,n187);
and (n331,n313,n332);
not (n332,n328);
nand (n333,n334,n358);
or (n334,n335,n351);
nand (n335,n336,n347);
nor (n336,n337,n344);
and (n337,n338,n341);
wire s0n338,s1n338,notn338;
or (n338,s0n338,s1n338);
not(notn338,n109);
and (s0n338,notn338,n339);
and (s1n338,n109,n340);
wire s0n339,s1n339,notn339;
or (n339,s0n339,s1n339);
not(notn339,n20);
and (s0n339,notn339,1'b0);
and (s1n339,n20,n85);
xor (n340,n84,n86);
wire s0n341,s1n341,notn341;
or (n341,s0n341,s1n341);
not(notn341,n109);
and (s0n341,notn341,n342);
and (s1n341,n109,n343);
wire s0n342,s1n342,notn342;
or (n342,s0n342,s1n342);
not(notn342,n20);
and (s0n342,notn342,1'b0);
and (s1n342,n20,n82);
xor (n343,n81,n83);
and (n344,n345,n346);
not (n345,n338);
not (n346,n341);
not (n347,n348);
nor (n348,n349,n350);
and (n349,n240,n338);
and (n350,n244,n345);
nor (n351,n352,n356);
and (n352,n346,n353);
wire s0n353,s1n353,notn353;
or (n353,s0n353,s1n353);
not(notn353,n209);
and (s0n353,notn353,n354);
and (s1n353,n209,n355);
wire s0n354,s1n354,notn354;
or (n354,s0n354,s1n354);
not(notn354,n20);
and (s0n354,notn354,1'b0);
and (s1n354,n20,n165);
xor (n355,n164,n166);
and (n356,n341,n357);
not (n357,n353);
or (n358,n359,n347);
nor (n359,n360,n364);
and (n360,n346,n361);
wire s0n361,s1n361,notn361;
or (n361,s0n361,s1n361);
not(notn361,n209);
and (s0n361,notn361,n362);
and (s1n361,n209,n363);
wire s0n362,s1n362,notn362;
or (n362,s0n362,s1n362);
not(notn362,n20);
and (s0n362,notn362,1'b0);
and (s1n362,n20,n162);
xor (n363,n161,n163);
and (n364,n341,n365);
not (n365,n361);
xor (n366,n367,n434);
xor (n367,n368,n401);
nand (n368,n369,n392);
or (n369,n370,n385);
or (n370,n371,n378);
nor (n371,n372,n376);
and (n372,n268,n373);
wire s0n373,s1n373,notn373;
or (n373,s0n373,s1n373);
not(notn373,n109);
and (s0n373,notn373,n374);
and (s1n373,n109,n375);
wire s0n374,s1n374,notn374;
or (n374,s0n374,s1n374);
not(notn374,n20);
and (s0n374,notn374,1'b0);
and (s1n374,n20,n73);
xor (n375,n72,n74);
and (n376,n377,n269);
not (n377,n373);
nor (n378,n379,n383);
and (n379,n373,n380);
wire s0n380,s1n380,notn380;
or (n380,s0n380,s1n380);
not(notn380,n109);
and (s0n380,notn380,n381);
and (s1n380,n109,n382);
wire s0n381,s1n381,notn381;
or (n381,s0n381,s1n381);
not(notn381,n20);
and (s0n381,notn381,1'b0);
and (s1n381,n20,n76);
xor (n382,n75,n77);
and (n383,n377,n384);
not (n384,n380);
nor (n385,n386,n390);
and (n386,n268,n387);
wire s0n387,s1n387,notn387;
or (n387,s0n387,s1n387);
not(notn387,n209);
and (s0n387,notn387,n388);
and (s1n387,n209,n389);
wire s0n388,s1n388,notn388;
or (n388,s0n388,s1n388);
not(notn388,n20);
and (s0n388,notn388,1'b0);
and (s1n388,n20,n177);
xor (n389,n176,n178);
and (n390,n269,n391);
not (n391,n387);
or (n392,n393,n394);
not (n393,n378);
nor (n394,n395,n399);
and (n395,n268,n396);
wire s0n396,s1n396,notn396;
or (n396,s0n396,s1n396);
not(notn396,n209);
and (s0n396,notn396,n397);
and (s1n396,n209,n398);
wire s0n397,s1n397,notn397;
or (n397,s0n397,s1n397);
not(notn397,n20);
and (s0n397,notn397,1'b0);
and (s1n397,n20,n174);
xor (n398,n173,n175);
and (n399,n269,n400);
not (n400,n396);
nand (n401,n402,n425);
or (n402,n403,n418);
or (n403,n404,n411);
nor (n404,n405,n409);
and (n405,n406,n313);
wire s0n406,s1n406,notn406;
or (n406,s0n406,s1n406);
not(notn406,n109);
and (s0n406,notn406,n407);
and (s1n406,n109,n408);
wire s0n407,s1n407,notn407;
or (n407,s0n407,s1n407);
not(notn407,n20);
and (s0n407,notn407,1'b0);
and (s1n407,n20,n55);
xor (n408,n54,n56);
and (n409,n410,n317);
not (n410,n406);
nor (n411,n412,n417);
and (n412,n406,n413);
not (n413,n414);
wire s0n414,s1n414,notn414;
or (n414,s0n414,s1n414);
not(notn414,n109);
and (s0n414,notn414,n415);
and (s1n414,n109,n416);
wire s0n415,s1n415,notn415;
or (n415,s0n415,s1n415);
not(notn415,n20);
and (s0n415,notn415,1'b0);
and (s1n415,n20,n52);
xor (n416,n51,n53);
and (n417,n410,n414);
nor (n418,n419,n423);
and (n419,n420,n413);
wire s0n420,s1n420,notn420;
or (n420,s0n420,s1n420);
not(notn420,n209);
and (s0n420,notn420,n421);
and (s1n420,n209,n422);
wire s0n421,s1n421,notn421;
or (n421,s0n421,s1n421);
not(notn421,n20);
and (s0n421,notn421,1'b0);
and (s1n421,n20,n195);
xor (n422,n194,n196);
and (n423,n424,n414);
not (n424,n420);
or (n425,n426,n427);
not (n426,n404);
nor (n427,n428,n432);
and (n428,n413,n429);
wire s0n429,s1n429,notn429;
or (n429,s0n429,s1n429);
not(notn429,n209);
and (s0n429,notn429,n430);
and (s1n429,n209,n431);
wire s0n430,s1n430,notn430;
or (n430,s0n430,s1n430);
not(notn430,n20);
and (s0n430,notn430,1'b0);
and (s1n430,n20,n192);
xor (n431,n191,n193);
and (n432,n414,n433);
not (n433,n429);
nand (n434,n435,n458);
or (n435,n436,n451);
nand (n436,n437,n444);
nor (n437,n438,n442);
and (n438,n413,n439);
wire s0n439,s1n439,notn439;
or (n439,s0n439,s1n439);
not(notn439,n109);
and (s0n439,notn439,n440);
and (s1n439,n109,n441);
wire s0n440,s1n440,notn440;
or (n440,s0n440,s1n440);
not(notn440,n20);
and (s0n440,notn440,1'b0);
and (s1n440,n20,n49);
xor (n441,n48,n50);
and (n442,n414,n443);
not (n443,n439);
nand (n444,n445,n449);
or (n445,n443,n446);
wire s0n446,s1n446,notn446;
or (n446,s0n446,s1n446);
not(notn446,n109);
and (s0n446,notn446,n447);
and (s1n446,n109,n448);
wire s0n447,s1n447,notn447;
or (n447,s0n447,s1n447);
not(notn447,n20);
and (s0n447,notn447,1'b0);
and (s1n447,n20,n46);
xor (n448,n45,n47);
or (n449,n439,n450);
not (n450,n446);
nor (n451,n452,n456);
and (n452,n453,n450);
wire s0n453,s1n453,notn453;
or (n453,s0n453,s1n453);
not(notn453,n209);
and (s0n453,notn453,n454);
and (s1n453,n209,n455);
wire s0n454,s1n454,notn454;
or (n454,s0n454,s1n454);
not(notn454,n20);
and (s0n454,notn454,1'b0);
and (s1n454,n20,n201);
xor (n455,n200,n202);
and (n456,n457,n446);
not (n457,n453);
or (n458,n437,n459);
nor (n459,n460,n464);
and (n460,n450,n461);
wire s0n461,s1n461,notn461;
or (n461,s0n461,s1n461);
not(notn461,n209);
and (s0n461,notn461,n462);
and (s1n461,n209,n463);
wire s0n462,s1n462,notn462;
or (n462,s0n462,s1n462);
not(notn462,n20);
and (s0n462,notn462,1'b0);
and (s1n462,n20,n198);
xor (n463,n197,n199);
and (n464,n446,n465);
not (n465,n461);
and (n466,n10,n260);
xor (n467,n468,n536);
xor (n468,n469,n493);
xor (n469,n470,n487);
xor (n470,n471,n481);
nand (n471,n472,n473);
or (n472,n226,n253);
or (n473,n474,n227);
nor (n474,n475,n479);
and (n475,n476,n244);
wire s0n476,s1n476,notn476;
or (n476,s0n476,s1n476);
not(notn476,n209);
and (s0n476,notn476,n477);
and (s1n476,n209,n478);
wire s0n477,s1n477,notn477;
or (n477,s0n477,s1n477);
not(notn477,n20);
and (s0n477,notn477,1'b0);
and (s1n477,n20,n153);
xor (n478,n152,n154);
and (n479,n480,n240);
not (n480,n476);
nand (n481,n482,n483);
or (n482,n264,n293);
or (n483,n292,n484);
nor (n484,n485,n486);
and (n485,n278,n387);
and (n486,n279,n391);
nand (n487,n488,n489);
or (n488,n302,n326);
or (n489,n490,n304);
nor (n490,n491,n492);
and (n491,n317,n286);
and (n492,n313,n290);
xor (n493,n494,n530);
xor (n494,n495,n520);
nand (n495,n496,n516);
or (n496,n497,n509);
nand (n497,n498,n505);
not (n498,n499);
nand (n499,n500,n504);
or (n500,n136,n501);
wire s0n501,s1n501,notn501;
or (n501,s0n501,s1n501);
not(notn501,n109);
and (s0n501,notn501,n502);
and (s1n501,n109,n503);
wire s0n502,s1n502,notn502;
or (n502,s0n502,s1n502);
not(notn502,n20);
and (s0n502,notn502,1'b0);
and (s1n502,n20,n97);
xor (n503,n96,n98);
nand (n504,n501,n136);
nor (n505,n506,n508);
and (n506,n236,n507);
not (n507,n501);
and (n508,n229,n501);
nor (n509,n510,n514);
and (n510,n511,n236);
wire s0n511,s1n511,notn511;
or (n511,s0n511,s1n511);
not(notn511,n209);
and (s0n511,notn511,n512);
and (s1n511,n209,n513);
wire s0n512,s1n512,notn512;
or (n512,s0n512,s1n512);
not(notn512,n20);
and (s0n512,notn512,1'b0);
and (s1n512,n20,n150);
xor (n513,n149,n151);
and (n514,n515,n229);
not (n515,n511);
or (n516,n517,n498);
nor (n517,n518,n519);
and (n518,n143,n236);
and (n519,n212,n229);
nand (n520,n521,n522);
or (n521,n370,n394);
or (n522,n393,n523);
nor (n523,n524,n528);
and (n524,n268,n525);
wire s0n525,s1n525,notn525;
or (n525,s0n525,s1n525);
not(notn525,n209);
and (s0n525,notn525,n526);
and (s1n525,n209,n527);
wire s0n526,s1n526,notn526;
or (n526,s0n526,s1n526);
not(notn526,n20);
and (s0n526,notn526,1'b0);
and (s1n526,n20,n171);
xor (n527,n170,n172);
and (n528,n269,n529);
not (n529,n525);
nand (n530,n531,n532);
or (n531,n403,n427);
or (n532,n426,n533);
nor (n533,n534,n535);
and (n534,n413,n320);
and (n535,n414,n324);
xor (n536,n537,n569);
xor (n537,n538,n544);
nand (n538,n539,n540);
or (n539,n436,n459);
or (n540,n437,n541);
nor (n541,n542,n543);
and (n542,n450,n420);
and (n543,n424,n446);
nand (n544,n545,n565);
or (n545,n546,n558);
or (n546,n547,n555);
not (n547,n548);
and (n548,n549,n554);
nand (n549,n550,n446);
not (n550,n551);
wire s0n551,s1n551,notn551;
or (n551,s0n551,s1n551);
not(notn551,n109);
and (s0n551,notn551,n552);
and (s1n551,n109,n553);
wire s0n552,s1n552,notn552;
or (n552,s0n552,s1n552);
not(notn552,n20);
and (s0n552,notn552,1'b0);
and (s1n552,n20,n43);
xor (n553,n42,n44);
nand (n554,n551,n450);
nor (n555,n556,n557);
and (n556,n551,n116);
and (n557,n550,n112);
nor (n558,n559,n563);
and (n559,n560,n116);
wire s0n560,s1n560,notn560;
or (n560,s0n560,s1n560);
not(notn560,n209);
and (s0n560,notn560,n561);
and (s1n560,n209,n562);
wire s0n561,s1n561,notn561;
or (n561,s0n561,s1n561);
not(notn561,n20);
and (s0n561,notn561,1'b0);
and (s1n561,n20,n204);
xor (n562,n203,n205);
and (n563,n564,n112);
not (n564,n560);
or (n565,n548,n566);
nor (n566,n567,n568);
and (n567,n453,n116);
and (n568,n457,n112);
nand (n569,n570,n587);
or (n570,n571,n584);
nand (n571,n572,n13);
or (n572,n573,n582);
not (n573,n574);
nand (n574,n16,n575);
not (n575,n576);
wire s0n576,s1n576,notn576;
or (n576,s0n576,s1n576);
not(notn576,n109);
and (s0n576,notn576,n577);
and (s1n576,n109,n579);
wire s0n577,s1n577,notn577;
or (n577,s0n577,s1n577);
not(notn577,n20);
and (s0n577,notn577,1'b0);
and (s1n577,n20,n578);
xor (n579,n580,n581);
not (n580,n578);
and (n581,n37,n38);
not (n582,n583);
nand (n583,n15,n576);
nor (n584,n585,n586);
and (n585,n576,n117);
and (n586,n575,n118);
or (n587,n13,n588);
nor (n588,n589,n593);
and (n589,n590,n575);
wire s0n590,s1n590,notn590;
or (n590,s0n590,s1n590);
not(notn590,n209);
and (s0n590,notn590,n591);
and (s1n590,n209,n592);
wire s0n591,s1n591,notn591;
or (n591,s0n591,s1n591);
not(notn591,n20);
and (s0n591,notn591,1'b0);
and (s1n591,n20,n207);
xor (n592,n206,n208);
and (n593,n594,n576);
not (n594,n590);
xor (n595,n596,n603);
xor (n596,n597,n600);
or (n597,n598,n599);
and (n598,n11,n224);
and (n599,n12,n120);
or (n600,n601,n602);
and (n601,n367,n434);
and (n602,n368,n401);
xor (n603,n604,n640);
xor (n604,n605,n611);
nand (n605,n606,n607);
or (n606,n335,n359);
or (n607,n608,n347);
nor (n608,n609,n610);
and (n609,n247,n346);
and (n610,n251,n341);
nand (n611,n612,n629);
or (n612,n613,n626);
nor (n613,n614,n624);
and (n614,n615,n125);
wire s0n615,s1n615,notn615;
or (n615,s0n615,s1n615);
not(notn615,n209);
and (s0n615,notn615,n616);
and (s1n615,n209,n618);
wire s0n616,s1n616,notn616;
or (n616,s0n616,s1n616);
not(notn616,n20);
and (s0n616,notn616,1'b0);
and (s1n616,n20,n617);
xor (n618,n619,n620);
not (n619,n617);
and (n620,n621,n623);
not (n621,n622);
and (n623,n220,n221);
and (n624,n625,n126);
not (n625,n615);
nand (n626,n126,n627);
not (n627,n628);
wire s0n628,s1n628,notn628;
or (n628,s0n628,s1n628);
not(notn628,n20);
and (s0n628,notn628,1'b0);
and (s1n628,n20,n108);
or (n629,n630,n627);
nor (n630,n631,n638);
and (n631,n632,n125);
wire s0n632,s1n632,notn632;
or (n632,s0n632,s1n632);
not(notn632,n209);
and (s0n632,notn632,n633);
and (s1n632,n209,n635);
wire s0n633,s1n633,notn633;
or (n633,s0n633,s1n633);
not(notn633,n20);
and (s0n633,notn633,1'b0);
and (s1n633,n20,n634);
xor (n635,n636,n637);
not (n636,n634);
and (n637,n619,n620);
and (n638,n639,n126);
not (n639,n632);
nand (n640,n641,n660);
or (n641,n642,n653);
nand (n642,n643,n650);
or (n643,n644,n648);
and (n644,n645,n341);
wire s0n645,s1n645,notn645;
or (n645,s0n645,s1n645);
not(notn645,n109);
and (s0n645,notn645,n646);
and (s1n645,n109,n647);
wire s0n646,s1n646,notn646;
or (n646,s0n646,s1n646);
not(notn646,n20);
and (s0n646,notn646,1'b0);
and (s1n646,n20,n79);
xor (n647,n78,n80);
and (n648,n649,n346);
not (n649,n645);
nand (n650,n651,n652);
or (n651,n649,n380);
or (n652,n384,n645);
nor (n653,n654,n658);
and (n654,n384,n655);
wire s0n655,s1n655,notn655;
or (n655,s0n655,s1n655);
not(notn655,n209);
and (s0n655,notn655,n656);
and (s1n655,n209,n657);
wire s0n656,s1n656,notn656;
or (n656,s0n656,s1n656);
not(notn656,n20);
and (s0n656,notn656,1'b0);
and (s1n656,n20,n168);
xor (n657,n167,n169);
and (n658,n380,n659);
not (n659,n655);
or (n660,n643,n661);
nor (n661,n662,n663);
and (n662,n384,n353);
and (n663,n380,n357);
or (n664,n665,n971);
and (n665,n666,n893);
xor (n666,n667,n803);
or (n667,n668,n802);
and (n668,n669,n720);
xor (n669,n670,n690);
xor (n670,n671,n684);
xor (n671,n672,n678);
nand (n672,n673,n677);
or (n673,n226,n674);
nor (n674,n675,n676);
and (n675,n361,n244);
and (n676,n365,n240);
or (n677,n245,n227);
nand (n678,n679,n683);
or (n679,n264,n680);
nor (n680,n681,n682);
and (n681,n278,n328);
and (n682,n279,n332);
or (n683,n292,n284);
nand (n684,n685,n689);
or (n685,n302,n686);
nor (n686,n687,n688);
and (n687,n317,n429);
and (n688,n313,n433);
or (n689,n318,n304);
xor (n690,n691,n707);
xor (n691,n692,n698);
nand (n692,n693,n697);
or (n693,n436,n694);
nor (n694,n695,n696);
and (n695,n560,n450);
and (n696,n564,n446);
or (n697,n437,n451);
nand (n698,n699,n703);
or (n699,n546,n700);
nor (n700,n701,n702);
and (n701,n112,n117);
and (n702,n116,n118);
or (n703,n548,n704);
nor (n704,n705,n706);
and (n705,n590,n116);
and (n706,n594,n112);
xor (n707,n708,n714);
nor (n708,n709,n116);
nor (n709,n710,n713);
and (n710,n711,n450);
not (n711,n712);
and (n712,n118,n551);
and (n713,n550,n117);
nand (n714,n715,n719);
or (n715,n122,n716);
nor (n716,n717,n718);
and (n717,n511,n136);
and (n718,n515,n137);
or (n719,n141,n123);
or (n720,n721,n801);
and (n721,n722,n770);
xor (n722,n723,n739);
and (n723,n724,n730);
nor (n724,n725,n450);
nor (n725,n726,n729);
and (n726,n727,n413);
not (n727,n728);
and (n728,n118,n439);
and (n729,n443,n117);
nand (n730,n731,n735);
or (n731,n122,n732);
nor (n732,n733,n734);
and (n733,n255,n136);
and (n734,n259,n137);
or (n735,n123,n736);
nor (n736,n737,n738);
and (n737,n476,n136);
and (n738,n480,n137);
or (n739,n740,n769);
and (n740,n741,n760);
xor (n741,n742,n751);
nand (n742,n743,n747);
or (n743,n335,n744);
nor (n744,n745,n746);
and (n745,n346,n396);
and (n746,n341,n400);
or (n747,n748,n347);
nor (n748,n749,n750);
and (n749,n346,n525);
and (n750,n341,n529);
nand (n751,n752,n756);
or (n752,n753,n626);
nor (n753,n754,n755);
and (n754,n511,n125);
and (n755,n515,n126);
or (n756,n757,n627);
nor (n757,n758,n759);
and (n758,n143,n125);
and (n759,n212,n126);
nand (n760,n761,n765);
or (n761,n497,n762);
nor (n762,n763,n764);
and (n763,n361,n236);
and (n764,n365,n229);
or (n765,n766,n498);
nor (n766,n767,n768);
and (n767,n247,n236);
and (n768,n251,n229);
and (n769,n742,n751);
or (n770,n771,n800);
and (n771,n772,n791);
xor (n772,n773,n782);
nand (n773,n774,n778);
or (n774,n226,n775);
nor (n775,n776,n777);
and (n776,n655,n244);
and (n777,n659,n240);
or (n778,n227,n779);
nor (n779,n780,n781);
and (n780,n353,n244);
and (n781,n357,n240);
nand (n782,n783,n787);
or (n783,n264,n784);
nor (n784,n785,n786);
and (n785,n278,n429);
and (n786,n279,n433);
or (n787,n788,n292);
nor (n788,n789,n790);
and (n789,n278,n320);
and (n790,n279,n324);
nand (n791,n792,n796);
or (n792,n302,n793);
nor (n793,n794,n795);
and (n794,n317,n461);
and (n795,n313,n465);
or (n796,n797,n304);
nor (n797,n798,n799);
and (n798,n317,n420);
and (n799,n313,n424);
and (n800,n773,n782);
and (n801,n723,n739);
and (n802,n670,n690);
xor (n803,n804,n846);
xor (n804,n805,n808);
or (n805,n806,n807);
and (n806,n691,n707);
and (n807,n692,n698);
xor (n808,n809,n814);
xor (n809,n810,n813);
nand (n810,n811,n812);
or (n811,n546,n704);
or (n812,n548,n558);
and (n813,n708,n714);
or (n814,n815,n845);
and (n815,n816,n836);
xor (n816,n817,n823);
nand (n817,n818,n822);
or (n818,n335,n819);
nor (n819,n820,n821);
and (n820,n346,n655);
and (n821,n341,n659);
or (n822,n351,n347);
nand (n823,n824,n828);
or (n824,n825,n626);
nor (n825,n826,n827);
and (n826,n216,n125);
and (n827,n223,n126);
or (n828,n829,n627);
nor (n829,n830,n834);
and (n830,n831,n125);
wire s0n831,s1n831,notn831;
or (n831,s0n831,s1n831);
not(notn831,n209);
and (s0n831,notn831,n832);
and (s1n831,n209,n833);
wire s0n832,s1n832,notn832;
or (n832,s0n832,s1n832);
not(notn832,n20);
and (s0n832,notn832,1'b0);
and (s1n832,n20,n622);
xor (n833,n621,n623);
and (n834,n835,n126);
not (n835,n831);
nand (n836,n837,n841);
or (n837,n497,n838);
nor (n838,n839,n840);
and (n839,n255,n236);
and (n840,n259,n229);
or (n841,n842,n498);
nor (n842,n843,n844);
and (n843,n476,n236);
and (n844,n480,n229);
and (n845,n817,n823);
or (n846,n847,n892);
and (n847,n848,n879);
xor (n848,n849,n868);
or (n849,n850,n867);
and (n850,n851,n858);
xor (n851,n852,n855);
nand (n852,n853,n854);
or (n853,n757,n626);
or (n854,n825,n627);
nand (n855,n856,n857);
or (n856,n497,n766);
or (n857,n838,n498);
nand (n858,n859,n863);
or (n859,n642,n860);
nor (n860,n861,n862);
and (n861,n384,n387);
and (n862,n380,n391);
or (n863,n643,n864);
nor (n864,n865,n866);
and (n865,n384,n396);
and (n866,n380,n400);
and (n867,n852,n855);
or (n868,n869,n878);
and (n869,n870,n875);
xor (n870,n871,n872);
nor (n871,n548,n117);
nand (n872,n873,n874);
or (n873,n122,n736);
or (n874,n123,n716);
nand (n875,n876,n877);
or (n876,n226,n779);
or (n877,n227,n674);
and (n878,n871,n872);
or (n879,n880,n891);
and (n880,n881,n888);
xor (n881,n882,n885);
nand (n882,n883,n884);
or (n883,n264,n788);
or (n884,n292,n680);
nand (n885,n886,n887);
or (n886,n302,n797);
or (n887,n686,n304);
nand (n888,n889,n890);
or (n889,n335,n748);
or (n890,n819,n347);
and (n891,n882,n885);
and (n892,n849,n868);
or (n893,n894,n970);
and (n894,n895,n931);
xor (n895,n896,n930);
or (n896,n897,n929);
and (n897,n898,n928);
xor (n898,n899,n927);
or (n899,n900,n926);
and (n900,n901,n917);
xor (n901,n902,n908);
nand (n902,n903,n907);
or (n903,n642,n904);
nor (n904,n905,n906);
and (n905,n384,n295);
and (n906,n380,n299);
or (n907,n643,n860);
nand (n908,n909,n913);
or (n909,n370,n910);
nor (n910,n911,n912);
and (n911,n268,n328);
and (n912,n269,n332);
or (n913,n393,n914);
nor (n914,n915,n916);
and (n915,n268,n286);
and (n916,n269,n290);
nand (n917,n918,n922);
or (n918,n403,n919);
nor (n919,n920,n921);
and (n920,n560,n413);
and (n921,n564,n414);
or (n922,n426,n923);
nor (n923,n924,n925);
and (n924,n453,n413);
and (n925,n457,n414);
and (n926,n902,n908);
xor (n927,n851,n858);
xor (n928,n881,n888);
and (n929,n899,n927);
xor (n930,n848,n879);
xor (n931,n932,n954);
xor (n932,n933,n953);
xor (n933,n934,n947);
xor (n934,n935,n941);
nand (n935,n936,n937);
or (n936,n642,n864);
or (n937,n643,n938);
nor (n938,n939,n940);
and (n939,n384,n525);
and (n940,n380,n529);
nand (n941,n942,n946);
or (n942,n370,n943);
nor (n943,n944,n945);
and (n944,n268,n295);
and (n945,n269,n299);
or (n946,n393,n385);
nand (n947,n948,n952);
or (n948,n403,n949);
nor (n949,n950,n951);
and (n950,n413,n461);
and (n951,n414,n465);
or (n952,n426,n418);
xor (n953,n816,n836);
or (n954,n955,n969);
and (n955,n956,n963);
xor (n956,n957,n960);
nand (n957,n958,n959);
or (n958,n370,n914);
or (n959,n393,n943);
nand (n960,n961,n962);
or (n961,n403,n923);
or (n962,n426,n949);
nand (n963,n964,n968);
or (n964,n436,n965);
nor (n965,n966,n967);
and (n966,n590,n450);
and (n967,n594,n446);
or (n968,n437,n694);
and (n969,n957,n960);
and (n970,n896,n930);
and (n971,n667,n803);
xor (n972,n973,n1024);
xor (n973,n974,n977);
or (n974,n975,n976);
and (n975,n804,n846);
and (n976,n805,n808);
xor (n977,n978,n1003);
xor (n978,n979,n982);
or (n979,n980,n981);
and (n980,n809,n814);
and (n981,n810,n813);
or (n982,n983,n1002);
and (n983,n984,n991);
xor (n984,n985,n988);
or (n985,n986,n987);
and (n986,n671,n684);
and (n987,n672,n678);
or (n988,n989,n990);
and (n989,n934,n947);
and (n990,n935,n941);
xor (n991,n992,n999);
xor (n992,n993,n996);
nand (n993,n994,n995);
or (n994,n829,n626);
or (n995,n613,n627);
nand (n996,n997,n998);
or (n997,n497,n842);
or (n998,n498,n509);
nand (n999,n1000,n1001);
or (n1000,n642,n938);
or (n1001,n643,n653);
and (n1002,n985,n988);
xor (n1003,n1004,n1021);
xor (n1004,n1005,n1018);
xor (n1005,n1006,n1012);
nor (n1006,n1007,n575);
nor (n1007,n1008,n1011);
and (n1008,n1009,n116);
not (n1009,n1010);
and (n1010,n118,n16);
and (n1011,n15,n117);
nand (n1012,n1013,n1014);
or (n1013,n122,n214);
or (n1014,n123,n1015);
nor (n1015,n1016,n1017);
and (n1016,n831,n136);
and (n1017,n835,n137);
or (n1018,n1019,n1020);
and (n1019,n261,n333);
and (n1020,n262,n300);
or (n1021,n1022,n1023);
and (n1022,n992,n999);
and (n1023,n993,n996);
or (n1024,n1025,n1032);
and (n1025,n1026,n1031);
xor (n1026,n1027,n1030);
or (n1027,n1028,n1029);
and (n1028,n932,n954);
and (n1029,n933,n953);
xor (n1030,n9,n366);
xor (n1031,n984,n991);
and (n1032,n1027,n1030);
and (n1033,n5,n664);
xor (n1034,n1035,n1158);
xor (n1035,n1036,n1155);
xor (n1036,n1037,n1098);
xor (n1037,n1038,n1095);
xor (n1038,n1039,n1070);
xor (n1039,n1040,n1043);
or (n1040,n1041,n1042);
and (n1041,n494,n530);
and (n1042,n495,n520);
xor (n1043,n1044,n1064);
xor (n1044,n1045,n1058);
nand (n1045,n1046,n1047);
or (n1046,n630,n626);
or (n1047,n1048,n627);
nor (n1048,n1049,n1056);
and (n1049,n1050,n125);
wire s0n1050,s1n1050,notn1050;
or (n1050,s0n1050,s1n1050);
not(notn1050,n209);
and (s0n1050,notn1050,n1051);
and (s1n1050,n209,n1053);
wire s0n1051,s1n1051,notn1051;
or (n1051,s0n1051,s1n1051);
not(notn1051,n20);
and (s0n1051,notn1051,1'b0);
and (s1n1051,n20,n1052);
xor (n1053,n1054,n1055);
not (n1054,n1052);
and (n1055,n636,n637);
and (n1056,n1057,n126);
not (n1057,n1050);
nand (n1058,n1059,n1060);
or (n1059,n642,n661);
or (n1060,n643,n1061);
nor (n1061,n1062,n1063);
and (n1062,n384,n361);
and (n1063,n380,n365);
nand (n1064,n1065,n1066);
or (n1065,n497,n517);
or (n1066,n1067,n498);
nor (n1067,n1068,n1069);
and (n1068,n216,n236);
and (n1069,n223,n229);
xor (n1070,n1071,n1089);
xor (n1071,n1072,n1083);
nor (n1072,n1073,n117);
nor (n1073,n1074,n1081);
and (n1074,n575,n1075);
wire s0n1075,s1n1075,notn1075;
or (n1075,s0n1075,s1n1075);
not(notn1075,n109);
and (s0n1075,notn1075,n1076);
and (s1n1075,n109,n1078);
wire s0n1076,s1n1076,notn1076;
or (n1076,s0n1076,s1n1076);
not(notn1076,n20);
and (s0n1076,notn1076,1'b0);
and (s1n1076,n20,n1077);
xor (n1078,n1079,n1080);
not (n1079,n1077);
and (n1080,n580,n581);
and (n1081,n576,n1082);
not (n1082,n1075);
nand (n1083,n1084,n1085);
or (n1084,n122,n1015);
or (n1085,n1086,n123);
nor (n1086,n1087,n1088);
and (n1087,n615,n136);
and (n1088,n625,n137);
nand (n1089,n1090,n1091);
or (n1090,n226,n474);
or (n1091,n1092,n227);
nor (n1092,n1093,n1094);
and (n1093,n511,n244);
and (n1094,n515,n240);
or (n1095,n1096,n1097);
and (n1096,n468,n536);
and (n1097,n469,n493);
xor (n1098,n1099,n1135);
xor (n1099,n1100,n1120);
xor (n1100,n1101,n1114);
xor (n1101,n1102,n1108);
nand (n1102,n1103,n1104);
or (n1103,n264,n484);
or (n1104,n292,n1105);
nor (n1105,n1106,n1107);
and (n1106,n278,n396);
and (n1107,n279,n400);
nand (n1108,n1109,n1110);
or (n1109,n302,n490);
or (n1110,n304,n1111);
nor (n1111,n1112,n1113);
and (n1112,n317,n295);
and (n1113,n313,n299);
nand (n1114,n1115,n1116);
or (n1115,n335,n608);
or (n1116,n1117,n347);
nor (n1117,n1118,n1119);
and (n1118,n255,n346);
and (n1119,n259,n341);
xor (n1120,n1121,n1134);
xor (n1121,n1122,n1128);
nand (n1122,n1123,n1124);
or (n1123,n546,n566);
or (n1124,n548,n1125);
nor (n1125,n1126,n1127);
and (n1126,n116,n461);
and (n1127,n465,n112);
nand (n1128,n1129,n1130);
or (n1129,n571,n588);
or (n1130,n1131,n13);
nor (n1131,n1132,n1133);
and (n1132,n560,n575);
and (n1133,n564,n576);
and (n1134,n1006,n1012);
xor (n1135,n1136,n1149);
xor (n1136,n1137,n1143);
nand (n1137,n1138,n1139);
or (n1138,n370,n523);
or (n1139,n393,n1140);
nor (n1140,n1141,n1142);
and (n1141,n268,n655);
and (n1142,n269,n659);
nand (n1143,n1144,n1145);
or (n1144,n403,n533);
or (n1145,n426,n1146);
nor (n1146,n1147,n1148);
and (n1147,n413,n328);
and (n1148,n414,n332);
nand (n1149,n1150,n1151);
or (n1150,n436,n541);
or (n1151,n437,n1152);
nor (n1152,n1153,n1154);
and (n1153,n450,n429);
and (n1154,n433,n446);
or (n1155,n1156,n1157);
and (n1156,n973,n1024);
and (n1157,n974,n977);
xor (n1158,n1159,n1166);
xor (n1159,n1160,n1163);
or (n1160,n1161,n1162);
and (n1161,n978,n1003);
and (n1162,n979,n982);
or (n1163,n1164,n1165);
and (n1164,n6,n595);
and (n1165,n7,n467);
xor (n1166,n1167,n1182);
xor (n1167,n1168,n1171);
or (n1168,n1169,n1170);
and (n1169,n1004,n1021);
and (n1170,n1005,n1018);
xor (n1171,n1172,n1179);
xor (n1172,n1173,n1176);
or (n1173,n1174,n1175);
and (n1174,n470,n487);
and (n1175,n471,n481);
or (n1176,n1177,n1178);
and (n1177,n604,n640);
and (n1178,n605,n611);
or (n1179,n1180,n1181);
and (n1180,n537,n569);
and (n1181,n538,n544);
or (n1182,n1183,n1184);
and (n1183,n596,n603);
and (n1184,n597,n600);
nand (n1185,n1186,n2536);
or (n1186,n1187,n2518,n2531);
nor (n1187,n1188,n2517);
and (n1188,n1189,n2496);
or (n1189,n1190,n2495);
and (n1190,n1191,n1545);
xor (n1191,n1192,n1518);
or (n1192,n1193,n1517);
and (n1193,n1194,n1432);
xor (n1194,n1195,n1319);
xor (n1195,n1196,n1289);
xor (n1196,n1197,n1228);
xor (n1197,n1198,n1206);
xor (n1198,n1199,n1205);
nand (n1199,n1200,n1204);
or (n1200,n436,n1201);
nor (n1201,n1202,n1203);
and (n1202,n446,n117);
and (n1203,n450,n118);
or (n1204,n437,n965);
xor (n1205,n724,n730);
or (n1206,n1207,n1227);
and (n1207,n1208,n1221);
xor (n1208,n1209,n1215);
nand (n1209,n1210,n1214);
or (n1210,n335,n1211);
nor (n1211,n1212,n1213);
and (n1212,n346,n387);
and (n1213,n341,n391);
or (n1214,n744,n347);
nand (n1215,n1216,n1220);
or (n1216,n497,n1217);
nor (n1217,n1218,n1219);
and (n1218,n353,n236);
and (n1219,n357,n229);
or (n1220,n498,n762);
nand (n1221,n1222,n1226);
or (n1222,n642,n1223);
nor (n1223,n1224,n1225);
and (n1224,n384,n286);
and (n1225,n380,n290);
or (n1226,n643,n904);
and (n1227,n1209,n1215);
or (n1228,n1229,n1288);
and (n1229,n1230,n1287);
xor (n1230,n1231,n1262);
or (n1231,n1232,n1261);
and (n1232,n1233,n1252);
xor (n1233,n1234,n1243);
nand (n1234,n1235,n1239);
or (n1235,n226,n1236);
nor (n1236,n1237,n1238);
and (n1237,n396,n244);
and (n1238,n400,n240);
or (n1239,n227,n1240);
nor (n1240,n1241,n1242);
and (n1241,n525,n244);
and (n1242,n529,n240);
nand (n1243,n1244,n1248);
or (n1244,n264,n1245);
nor (n1245,n1246,n1247);
and (n1246,n278,n461);
and (n1247,n465,n279);
or (n1248,n292,n1249);
nor (n1249,n1250,n1251);
and (n1250,n420,n278);
and (n1251,n424,n279);
nand (n1252,n1253,n1257);
or (n1253,n302,n1254);
nor (n1254,n1255,n1256);
and (n1255,n560,n317);
and (n1256,n564,n313);
or (n1257,n1258,n304);
nor (n1258,n1259,n1260);
and (n1259,n453,n317);
and (n1260,n457,n313);
and (n1261,n1234,n1243);
or (n1262,n1263,n1286);
and (n1263,n1264,n1280);
xor (n1264,n1265,n1274);
nand (n1265,n1266,n1270);
or (n1266,n122,n1267);
nor (n1267,n1268,n1269);
and (n1268,n136,n361);
and (n1269,n365,n137);
or (n1270,n1271,n123);
nor (n1271,n1272,n1273);
and (n1272,n247,n136);
and (n1273,n251,n137);
nand (n1274,n1275,n1279);
or (n1275,n335,n1276);
nor (n1276,n1277,n1278);
and (n1277,n346,n295);
and (n1278,n341,n299);
or (n1279,n1211,n347);
nand (n1280,n1281,n1285);
or (n1281,n497,n1282);
nor (n1282,n1283,n1284);
and (n1283,n655,n236);
and (n1284,n659,n229);
or (n1285,n498,n1217);
and (n1286,n1265,n1274);
xor (n1287,n1208,n1221);
and (n1288,n1231,n1262);
xor (n1289,n1290,n1318);
xor (n1290,n1291,n1305);
or (n1291,n1292,n1304);
and (n1292,n1293,n1301);
xor (n1293,n1294,n1295);
nor (n1294,n437,n117);
nand (n1295,n1296,n1300);
or (n1296,n1297,n626);
nor (n1297,n1298,n1299);
and (n1298,n476,n125);
and (n1299,n480,n126);
or (n1300,n753,n627);
nand (n1301,n1302,n1303);
or (n1302,n226,n1240);
or (n1303,n227,n775);
and (n1304,n1294,n1295);
or (n1305,n1306,n1317);
and (n1306,n1307,n1314);
xor (n1307,n1308,n1311);
nand (n1308,n1309,n1310);
or (n1309,n264,n1249);
or (n1310,n784,n292);
nand (n1311,n1312,n1313);
or (n1312,n302,n1258);
or (n1313,n793,n304);
nand (n1314,n1315,n1316);
or (n1315,n122,n1271);
or (n1316,n123,n732);
and (n1317,n1308,n1311);
xor (n1318,n741,n760);
xor (n1319,n1320,n1382);
xor (n1320,n1321,n1355);
or (n1321,n1322,n1354);
and (n1322,n1323,n1326);
xor (n1323,n1324,n1325);
xor (n1324,n1293,n1301);
xor (n1325,n1307,n1314);
or (n1326,n1327,n1353);
and (n1327,n1328,n1344);
xor (n1328,n1329,n1335);
nand (n1329,n1330,n1334);
or (n1330,n642,n1331);
nor (n1331,n1332,n1333);
and (n1332,n384,n328);
and (n1333,n380,n332);
or (n1334,n643,n1223);
nand (n1335,n1336,n1340);
or (n1336,n370,n1337);
nor (n1337,n1338,n1339);
and (n1338,n268,n429);
and (n1339,n269,n433);
or (n1340,n1341,n393);
nor (n1341,n1342,n1343);
and (n1342,n268,n320);
and (n1343,n269,n324);
nand (n1344,n1345,n1349);
or (n1345,n403,n1346);
nor (n1346,n1347,n1348);
and (n1347,n414,n117);
and (n1348,n413,n118);
or (n1349,n426,n1350);
nor (n1350,n1351,n1352);
and (n1351,n590,n413);
and (n1352,n594,n414);
and (n1353,n1329,n1335);
and (n1354,n1324,n1325);
xor (n1355,n1356,n1359);
xor (n1356,n1357,n1358);
xor (n1357,n772,n791);
xor (n1358,n901,n917);
or (n1359,n1360,n1381);
and (n1360,n1361,n1368);
xor (n1361,n1362,n1365);
nand (n1362,n1363,n1364);
or (n1363,n370,n1341);
or (n1364,n393,n910);
nand (n1365,n1366,n1367);
or (n1366,n403,n1350);
or (n1367,n426,n919);
and (n1368,n1369,n1375);
nor (n1369,n1370,n413);
nor (n1370,n1371,n1374);
and (n1371,n1372,n317);
not (n1372,n1373);
and (n1373,n118,n406);
and (n1374,n410,n117);
nand (n1375,n1376,n1380);
or (n1376,n1377,n626);
nor (n1377,n1378,n1379);
and (n1378,n255,n125);
and (n1379,n259,n126);
or (n1380,n1297,n627);
and (n1381,n1362,n1365);
or (n1382,n1383,n1431);
and (n1383,n1384,n1430);
xor (n1384,n1385,n1386);
xor (n1385,n1361,n1368);
or (n1386,n1387,n1429);
and (n1387,n1388,n1407);
xor (n1388,n1389,n1390);
xor (n1389,n1369,n1375);
or (n1390,n1391,n1406);
and (n1391,n1392,n1400);
xor (n1392,n1393,n1394);
nor (n1393,n426,n117);
nand (n1394,n1395,n1399);
or (n1395,n1396,n626);
nor (n1396,n1397,n1398);
and (n1397,n247,n125);
and (n1398,n251,n126);
or (n1399,n1377,n627);
nand (n1400,n1401,n1402);
or (n1401,n1236,n227);
or (n1402,n226,n1403);
nor (n1403,n1404,n1405);
and (n1404,n387,n244);
and (n1405,n391,n240);
and (n1406,n1393,n1394);
or (n1407,n1408,n1428);
and (n1408,n1409,n1422);
xor (n1409,n1410,n1416);
nand (n1410,n1411,n1415);
or (n1411,n264,n1412);
nor (n1412,n1413,n1414);
and (n1413,n453,n278);
and (n1414,n457,n279);
or (n1415,n1245,n292);
nand (n1416,n1417,n1421);
or (n1417,n302,n1418);
nor (n1418,n1419,n1420);
and (n1419,n590,n317);
and (n1420,n594,n313);
or (n1421,n1254,n304);
nand (n1422,n1423,n1427);
or (n1423,n122,n1424);
nor (n1424,n1425,n1426);
and (n1425,n136,n353);
and (n1426,n357,n137);
or (n1427,n123,n1267);
and (n1428,n1410,n1416);
and (n1429,n1389,n1390);
xor (n1430,n1230,n1287);
and (n1431,n1385,n1386);
or (n1432,n1433,n1516);
and (n1433,n1434,n1464);
xor (n1434,n1435,n1463);
or (n1435,n1436,n1462);
and (n1436,n1437,n1461);
xor (n1437,n1438,n1460);
or (n1438,n1439,n1459);
and (n1439,n1440,n1453);
xor (n1440,n1441,n1447);
nand (n1441,n1442,n1446);
or (n1442,n335,n1443);
nor (n1443,n1444,n1445);
and (n1444,n346,n286);
and (n1445,n341,n290);
or (n1446,n1276,n347);
nand (n1447,n1448,n1452);
or (n1448,n497,n1449);
nor (n1449,n1450,n1451);
and (n1450,n525,n236);
and (n1451,n529,n229);
or (n1452,n498,n1282);
nand (n1453,n1454,n1458);
or (n1454,n642,n1455);
nor (n1455,n1456,n1457);
and (n1456,n384,n320);
and (n1457,n380,n324);
or (n1458,n643,n1331);
and (n1459,n1441,n1447);
xor (n1460,n1264,n1280);
xor (n1461,n1233,n1252);
and (n1462,n1438,n1460);
xor (n1463,n1323,n1326);
or (n1464,n1465,n1515);
and (n1465,n1466,n1514);
xor (n1466,n1467,n1468);
xor (n1467,n1328,n1344);
or (n1468,n1469,n1513);
and (n1469,n1470,n1490);
xor (n1470,n1471,n1477);
nand (n1471,n1472,n1476);
or (n1472,n370,n1473);
nor (n1473,n1474,n1475);
and (n1474,n268,n420);
and (n1475,n269,n424);
or (n1476,n1337,n393);
and (n1477,n1478,n1484);
nor (n1478,n1479,n317);
nor (n1479,n1480,n1483);
and (n1480,n278,n1481);
not (n1481,n1482);
and (n1482,n118,n307);
and (n1483,n306,n117);
nand (n1484,n1485,n1489);
or (n1485,n1486,n626);
nor (n1486,n1487,n1488);
and (n1487,n361,n125);
and (n1488,n365,n126);
or (n1489,n1396,n627);
or (n1490,n1491,n1512);
and (n1491,n1492,n1505);
xor (n1492,n1493,n1499);
nand (n1493,n1494,n1498);
or (n1494,n226,n1495);
nor (n1495,n1496,n1497);
and (n1496,n295,n244);
and (n1497,n299,n240);
or (n1498,n1403,n227);
nand (n1499,n1500,n1504);
or (n1500,n264,n1501);
nor (n1501,n1502,n1503);
and (n1502,n560,n278);
and (n1503,n564,n279);
or (n1504,n292,n1412);
nand (n1505,n1506,n1511);
or (n1506,n1507,n302);
not (n1507,n1508);
nand (n1508,n1509,n1510);
or (n1509,n317,n118);
or (n1510,n313,n117);
or (n1511,n1418,n304);
and (n1512,n1493,n1499);
and (n1513,n1471,n1477);
xor (n1514,n1388,n1407);
and (n1515,n1467,n1468);
and (n1516,n1435,n1463);
and (n1517,n1195,n1319);
xor (n1518,n1519,n1542);
xor (n1519,n1520,n1529);
xor (n1520,n1521,n1526);
xor (n1521,n1522,n1523);
xor (n1522,n722,n770);
or (n1523,n1524,n1525);
and (n1524,n1290,n1318);
and (n1525,n1291,n1305);
or (n1526,n1527,n1528);
and (n1527,n1356,n1359);
and (n1528,n1357,n1358);
xor (n1529,n1530,n1539);
xor (n1530,n1531,n1532);
xor (n1531,n898,n928);
xor (n1532,n1533,n1536);
xor (n1533,n1534,n1535);
xor (n1534,n870,n875);
xor (n1535,n956,n963);
or (n1536,n1537,n1538);
and (n1537,n1198,n1206);
and (n1538,n1199,n1205);
or (n1539,n1540,n1541);
and (n1540,n1196,n1289);
and (n1541,n1197,n1228);
or (n1542,n1543,n1544);
and (n1543,n1320,n1382);
and (n1544,n1321,n1355);
nand (n1545,n1546,n2489);
or (n1546,n1547,n2482);
nand (n1547,n1548,n2471);
not (n1548,n1549);
nor (n1549,n1550,n2460);
nor (n1550,n1551,n2409);
nand (n1551,n1552,n2283);
or (n1552,n1553,n2282);
and (n1553,n1554,n1872);
xor (n1554,n1555,n1786);
or (n1555,n1556,n1785);
and (n1556,n1557,n1734);
xor (n1557,n1558,n1641);
xor (n1558,n1559,n1610);
xor (n1559,n1560,n1581);
xor (n1560,n1561,n1572);
xor (n1561,n1562,n1563);
nor (n1562,n292,n117);
nand (n1563,n1564,n1568);
or (n1564,n1565,n626);
nor (n1565,n1566,n1567);
and (n1566,n125,n525);
and (n1567,n529,n126);
or (n1568,n1569,n627);
nor (n1569,n1570,n1571);
and (n1570,n655,n125);
and (n1571,n659,n126);
nand (n1572,n1573,n1577);
or (n1573,n122,n1574);
nor (n1574,n1575,n1576);
and (n1575,n136,n387);
and (n1576,n391,n137);
or (n1577,n123,n1578);
nor (n1578,n1579,n1580);
and (n1579,n396,n136);
and (n1580,n400,n137);
or (n1581,n1582,n1609);
and (n1582,n1583,n1599);
xor (n1583,n1584,n1590);
nand (n1584,n1585,n1589);
or (n1585,n122,n1586);
nor (n1586,n1587,n1588);
and (n1587,n136,n295);
and (n1588,n299,n137);
or (n1589,n123,n1574);
nand (n1590,n1591,n1595);
or (n1591,n226,n1592);
nor (n1592,n1593,n1594);
and (n1593,n429,n244);
and (n1594,n433,n240);
or (n1595,n227,n1596);
nor (n1596,n1597,n1598);
and (n1597,n320,n244);
and (n1598,n324,n240);
nand (n1599,n1600,n1605);
or (n1600,n1601,n335);
not (n1601,n1602);
nand (n1602,n1603,n1604);
or (n1603,n341,n465);
or (n1604,n346,n461);
or (n1605,n1606,n347);
nor (n1606,n1607,n1608);
and (n1607,n346,n420);
and (n1608,n341,n424);
and (n1609,n1584,n1590);
or (n1610,n1611,n1640);
and (n1611,n1612,n1631);
xor (n1612,n1613,n1622);
nand (n1613,n1614,n1618);
or (n1614,n497,n1615);
nor (n1615,n1616,n1617);
and (n1616,n328,n236);
and (n1617,n332,n229);
or (n1618,n1619,n498);
nor (n1619,n1620,n1621);
and (n1620,n286,n236);
and (n1621,n290,n229);
nand (n1622,n1623,n1627);
or (n1623,n642,n1624);
nor (n1624,n1625,n1626);
and (n1625,n560,n384);
and (n1626,n564,n380);
or (n1627,n1628,n643);
nor (n1628,n1629,n1630);
and (n1629,n453,n384);
and (n1630,n457,n380);
nand (n1631,n1632,n1636);
or (n1632,n393,n1633);
nor (n1633,n1634,n1635);
and (n1634,n590,n268);
and (n1635,n594,n269);
or (n1636,n370,n1637);
nor (n1637,n1638,n1639);
and (n1638,n269,n117);
and (n1639,n268,n118);
and (n1640,n1613,n1622);
xor (n1641,n1642,n1690);
xor (n1642,n1643,n1670);
xor (n1643,n1644,n1657);
xor (n1644,n1645,n1651);
nand (n1645,n1646,n1647);
or (n1646,n642,n1628);
or (n1647,n1648,n643);
nor (n1648,n1649,n1650);
and (n1649,n384,n461);
and (n1650,n380,n465);
nand (n1651,n1652,n1653);
or (n1652,n370,n1633);
or (n1653,n1654,n393);
nor (n1654,n1655,n1656);
and (n1655,n560,n268);
and (n1656,n564,n269);
and (n1657,n1658,n1664);
nand (n1658,n1659,n1663);
or (n1659,n1660,n626);
nor (n1660,n1661,n1662);
and (n1661,n125,n396);
and (n1662,n400,n126);
or (n1663,n1565,n627);
nor (n1664,n1665,n268);
nor (n1665,n1666,n1669);
and (n1666,n384,n1667);
not (n1667,n1668);
and (n1668,n118,n373);
and (n1669,n377,n117);
xor (n1670,n1671,n1684);
xor (n1671,n1672,n1678);
nand (n1672,n1673,n1674);
or (n1673,n226,n1596);
or (n1674,n1675,n227);
nor (n1675,n1676,n1677);
and (n1676,n328,n244);
and (n1677,n332,n240);
nand (n1678,n1679,n1680);
or (n1679,n335,n1606);
or (n1680,n1681,n347);
nor (n1681,n1682,n1683);
and (n1682,n346,n429);
and (n1683,n341,n433);
nand (n1684,n1685,n1689);
or (n1685,n498,n1686);
nor (n1686,n1687,n1688);
and (n1687,n295,n236);
and (n1688,n299,n229);
or (n1689,n497,n1619);
or (n1690,n1691,n1733);
and (n1691,n1692,n1711);
xor (n1692,n1693,n1694);
xor (n1693,n1658,n1664);
or (n1694,n1695,n1710);
and (n1695,n1696,n1704);
xor (n1696,n1697,n1698);
nor (n1697,n393,n117);
nand (n1698,n1699,n1703);
or (n1699,n1700,n626);
nor (n1700,n1701,n1702);
and (n1701,n125,n387);
and (n1702,n391,n126);
or (n1703,n1660,n627);
nand (n1704,n1705,n1706);
or (n1705,n123,n1586);
or (n1706,n122,n1707);
nor (n1707,n1708,n1709);
and (n1708,n286,n136);
and (n1709,n290,n137);
and (n1710,n1697,n1698);
or (n1711,n1712,n1732);
and (n1712,n1713,n1726);
xor (n1713,n1714,n1720);
nand (n1714,n1715,n1719);
or (n1715,n226,n1716);
nor (n1716,n1717,n1718);
and (n1717,n420,n244);
and (n1718,n424,n240);
or (n1719,n1592,n227);
nand (n1720,n1721,n1722);
or (n1721,n347,n1601);
or (n1722,n335,n1723);
nor (n1723,n1724,n1725);
and (n1724,n346,n453);
and (n1725,n341,n457);
nand (n1726,n1727,n1728);
or (n1727,n643,n1624);
or (n1728,n642,n1729);
nor (n1729,n1730,n1731);
and (n1730,n590,n384);
and (n1731,n594,n380);
and (n1732,n1714,n1720);
and (n1733,n1693,n1694);
or (n1734,n1735,n1784);
and (n1735,n1736,n1739);
xor (n1736,n1737,n1738);
xor (n1737,n1612,n1631);
xor (n1738,n1583,n1599);
or (n1739,n1740,n1783);
and (n1740,n1741,n1761);
xor (n1741,n1742,n1748);
nand (n1742,n1743,n1747);
or (n1743,n497,n1744);
nor (n1744,n1745,n1746);
and (n1745,n320,n236);
and (n1746,n324,n229);
or (n1747,n498,n1615);
and (n1748,n1749,n1755);
nand (n1749,n1750,n1754);
or (n1750,n1751,n626);
nor (n1751,n1752,n1753);
and (n1752,n295,n125);
and (n1753,n299,n126);
or (n1754,n1700,n627);
nor (n1755,n1756,n384);
nor (n1756,n1757,n1760);
and (n1757,n346,n1758);
not (n1758,n1759);
and (n1759,n118,n645);
and (n1760,n649,n117);
or (n1761,n1762,n1782);
and (n1762,n1763,n1776);
xor (n1763,n1764,n1770);
nand (n1764,n1765,n1769);
or (n1765,n122,n1766);
nor (n1766,n1767,n1768);
and (n1767,n328,n136);
and (n1768,n332,n137);
or (n1769,n123,n1707);
nand (n1770,n1771,n1775);
or (n1771,n226,n1772);
nor (n1772,n1773,n1774);
and (n1773,n461,n244);
and (n1774,n465,n240);
or (n1775,n1716,n227);
nand (n1776,n1777,n1781);
or (n1777,n335,n1778);
nor (n1778,n1779,n1780);
and (n1779,n560,n346);
and (n1780,n564,n341);
or (n1781,n1723,n347);
and (n1782,n1764,n1770);
and (n1783,n1742,n1748);
and (n1784,n1737,n1738);
and (n1785,n1558,n1641);
xor (n1786,n1787,n1820);
xor (n1787,n1788,n1817);
xor (n1788,n1789,n1796);
xor (n1789,n1790,n1793);
or (n1790,n1791,n1792);
and (n1791,n1671,n1684);
and (n1792,n1672,n1678);
or (n1793,n1794,n1795);
and (n1794,n1644,n1657);
and (n1795,n1645,n1651);
xor (n1796,n1797,n1810);
xor (n1797,n1798,n1804);
nand (n1798,n1799,n1800);
or (n1799,n335,n1681);
or (n1800,n1801,n347);
nor (n1801,n1802,n1803);
and (n1802,n346,n320);
and (n1803,n341,n324);
nand (n1804,n1805,n1806);
or (n1805,n497,n1686);
or (n1806,n498,n1807);
nor (n1807,n1808,n1809);
and (n1808,n387,n236);
and (n1809,n391,n229);
nand (n1810,n1811,n1816);
or (n1811,n643,n1812);
not (n1812,n1813);
nand (n1813,n1814,n1815);
or (n1814,n424,n380);
or (n1815,n384,n420);
or (n1816,n642,n1648);
or (n1817,n1818,n1819);
and (n1818,n1642,n1690);
and (n1819,n1643,n1670);
xor (n1820,n1821,n1848);
xor (n1821,n1822,n1845);
xor (n1822,n1823,n1839);
xor (n1823,n1824,n1830);
nand (n1824,n1825,n1826);
or (n1825,n122,n1578);
or (n1826,n123,n1827);
nor (n1827,n1828,n1829);
and (n1828,n136,n525);
and (n1829,n529,n137);
nand (n1830,n1831,n1835);
or (n1831,n264,n1832);
nor (n1832,n1833,n1834);
and (n1833,n279,n117);
and (n1834,n278,n118);
or (n1835,n1836,n292);
nor (n1836,n1837,n1838);
and (n1837,n590,n278);
and (n1838,n594,n279);
nand (n1839,n1840,n1844);
or (n1840,n1841,n227);
nor (n1841,n1842,n1843);
and (n1842,n286,n244);
and (n1843,n290,n240);
or (n1844,n226,n1675);
or (n1845,n1846,n1847);
and (n1846,n1559,n1610);
and (n1847,n1560,n1581);
xor (n1848,n1849,n1869);
xor (n1849,n1850,n1856);
nand (n1850,n1851,n1852);
or (n1851,n370,n1654);
or (n1852,n1853,n393);
nor (n1853,n1854,n1855);
and (n1854,n453,n268);
and (n1855,n457,n269);
xor (n1856,n1857,n1863);
nand (n1857,n1858,n1859);
or (n1858,n1569,n626);
or (n1859,n1860,n627);
nor (n1860,n1861,n1862);
and (n1861,n353,n125);
and (n1862,n357,n126);
nor (n1863,n1864,n278);
nor (n1864,n1865,n1868);
and (n1865,n268,n1866);
not (n1866,n1867);
and (n1867,n118,n272);
and (n1868,n283,n117);
or (n1869,n1870,n1871);
and (n1870,n1561,n1572);
and (n1871,n1562,n1563);
or (n1872,n1873,n2281);
and (n1873,n1874,n1905);
xor (n1874,n1875,n1904);
or (n1875,n1876,n1903);
and (n1876,n1877,n1902);
xor (n1877,n1878,n1901);
or (n1878,n1879,n1900);
and (n1879,n1880,n1883);
xor (n1880,n1881,n1882);
xor (n1881,n1696,n1704);
xor (n1882,n1713,n1726);
or (n1883,n1884,n1899);
and (n1884,n1885,n1898);
xor (n1885,n1886,n1892);
nand (n1886,n1887,n1891);
or (n1887,n642,n1888);
nor (n1888,n1889,n1890);
and (n1889,n380,n117);
and (n1890,n384,n118);
or (n1891,n1729,n643);
nand (n1892,n1893,n1897);
or (n1893,n497,n1894);
nor (n1894,n1895,n1896);
and (n1895,n429,n236);
and (n1896,n433,n229);
or (n1897,n1744,n498);
xor (n1898,n1749,n1755);
and (n1899,n1886,n1892);
and (n1900,n1881,n1882);
xor (n1901,n1692,n1711);
xor (n1902,n1736,n1739);
and (n1903,n1878,n1901);
xor (n1904,n1557,n1734);
nand (n1905,n1906,n2278,n2280);
or (n1906,n1907,n2273);
nand (n1907,n1908,n2262);
or (n1908,n1909,n2261);
and (n1909,n1910,n2031);
xor (n1910,n1911,n2016);
or (n1911,n1912,n2015);
and (n1912,n1913,n1981);
xor (n1913,n1914,n1936);
xor (n1914,n1915,n1930);
xor (n1915,n1916,n1923);
nand (n1916,n1917,n1922);
or (n1917,n226,n1918);
not (n1918,n1919);
nor (n1919,n1920,n1921);
and (n1920,n244,n457);
and (n1921,n453,n240);
or (n1922,n1772,n227);
nand (n1923,n1924,n1929);
or (n1924,n1925,n335);
not (n1925,n1926);
nand (n1926,n1927,n1928);
or (n1927,n594,n341);
or (n1928,n590,n346);
or (n1929,n1778,n347);
nand (n1930,n1931,n1935);
or (n1931,n497,n1932);
nor (n1932,n1933,n1934);
and (n1933,n420,n236);
and (n1934,n424,n229);
or (n1935,n498,n1894);
or (n1936,n1937,n1980);
and (n1937,n1938,n1960);
xor (n1938,n1939,n1945);
nand (n1939,n1940,n1944);
or (n1940,n497,n1941);
nor (n1941,n1942,n1943);
and (n1942,n461,n236);
and (n1943,n465,n229);
or (n1944,n1932,n498);
xor (n1945,n1946,n1952);
nor (n1946,n1947,n346);
nor (n1947,n1948,n1951);
and (n1948,n1949,n244);
not (n1949,n1950);
and (n1950,n118,n338);
and (n1951,n345,n117);
nand (n1952,n1953,n1956);
or (n1953,n626,n1954);
not (n1954,n1955);
xnor (n1955,n328,n125);
or (n1956,n1957,n627);
nor (n1957,n1958,n1959);
and (n1958,n125,n286);
and (n1959,n290,n126);
or (n1960,n1961,n1979);
and (n1961,n1962,n1970);
xor (n1962,n1963,n1964);
nor (n1963,n347,n117);
nand (n1964,n1965,n1966);
or (n1965,n627,n1954);
or (n1966,n1967,n626);
nor (n1967,n1968,n1969);
and (n1968,n125,n320);
and (n1969,n324,n126);
nand (n1970,n1971,n1975);
or (n1971,n226,n1972);
nor (n1972,n1973,n1974);
and (n1973,n590,n244);
and (n1974,n594,n240);
or (n1975,n1976,n227);
nor (n1976,n1977,n1978);
and (n1977,n560,n244);
and (n1978,n564,n240);
and (n1979,n1963,n1964);
and (n1980,n1939,n1945);
xor (n1981,n1982,n1996);
xor (n1982,n1983,n1984);
and (n1983,n1946,n1952);
xor (n1984,n1985,n1990);
xor (n1985,n1986,n1987);
nor (n1986,n643,n117);
nand (n1987,n1988,n1989);
or (n1988,n1957,n626);
or (n1989,n1751,n627);
nand (n1990,n1991,n1995);
or (n1991,n122,n1992);
nor (n1992,n1993,n1994);
and (n1993,n320,n136);
and (n1994,n324,n137);
or (n1995,n123,n1766);
or (n1996,n1997,n2014);
and (n1997,n1998,n2008);
xor (n1998,n1999,n2005);
nand (n1999,n2000,n2004);
or (n2000,n122,n2001);
nor (n2001,n2002,n2003);
and (n2002,n136,n429);
and (n2003,n433,n137);
or (n2004,n1992,n123);
nand (n2005,n2006,n2007);
or (n2006,n227,n1918);
or (n2007,n1976,n226);
nand (n2008,n2009,n2010);
or (n2009,n347,n1925);
or (n2010,n335,n2011);
nor (n2011,n2012,n2013);
and (n2012,n341,n117);
and (n2013,n346,n118);
and (n2014,n1999,n2005);
and (n2015,n1914,n1936);
xor (n2016,n2017,n2022);
xor (n2017,n2018,n2019);
xor (n2018,n1763,n1776);
or (n2019,n2020,n2021);
and (n2020,n1982,n1996);
and (n2021,n1983,n1984);
xor (n2022,n2023,n2030);
xor (n2023,n2024,n2027);
or (n2024,n2025,n2026);
and (n2025,n1985,n1990);
and (n2026,n1986,n1987);
or (n2027,n2028,n2029);
and (n2028,n1915,n1930);
and (n2029,n1916,n1923);
xor (n2030,n1885,n1898);
or (n2031,n2032,n2260);
and (n2032,n2033,n2070);
xor (n2033,n2034,n2069);
or (n2034,n2035,n2068);
and (n2035,n2036,n2067);
xor (n2036,n2037,n2066);
or (n2037,n2038,n2065);
and (n2038,n2039,n2052);
xor (n2039,n2040,n2046);
nand (n2040,n2041,n2045);
or (n2041,n122,n2042);
nor (n2042,n2043,n2044);
and (n2043,n420,n136);
and (n2044,n137,n424);
or (n2045,n2001,n123);
nand (n2046,n2047,n2051);
or (n2047,n497,n2048);
nor (n2048,n2049,n2050);
and (n2049,n453,n236);
and (n2050,n457,n229);
or (n2051,n1941,n498);
and (n2052,n2053,n2059);
nor (n2053,n2054,n244);
nor (n2054,n2055,n2058);
and (n2055,n2056,n236);
not (n2056,n2057);
and (n2057,n118,n232);
and (n2058,n237,n117);
nand (n2059,n2060,n2064);
or (n2060,n2061,n626);
nor (n2061,n2062,n2063);
and (n2062,n125,n429);
and (n2063,n433,n126);
or (n2064,n1967,n627);
and (n2065,n2040,n2046);
xor (n2066,n1998,n2008);
xor (n2067,n1938,n1960);
and (n2068,n2037,n2066);
xor (n2069,n1913,n1981);
nand (n2070,n2071,n2257,n2259);
or (n2071,n2072,n2130);
nand (n2072,n2073,n2125);
not (n2073,n2074);
nor (n2074,n2075,n2101);
xor (n2075,n2076,n2100);
xor (n2076,n2077,n2099);
or (n2077,n2078,n2098);
and (n2078,n2079,n2092);
xor (n2079,n2080,n2086);
nand (n2080,n2081,n2085);
or (n2081,n226,n2082);
nor (n2082,n2083,n2084);
and (n2083,n240,n117);
and (n2084,n244,n118);
or (n2085,n1972,n227);
nand (n2086,n2087,n2091);
or (n2087,n2088,n122);
nor (n2088,n2089,n2090);
and (n2089,n137,n465);
and (n2090,n136,n461);
or (n2091,n2042,n123);
nand (n2092,n2093,n2097);
or (n2093,n497,n2094);
nor (n2094,n2095,n2096);
and (n2095,n560,n236);
and (n2096,n564,n229);
or (n2097,n2048,n498);
and (n2098,n2080,n2086);
xor (n2099,n1962,n1970);
xor (n2100,n2039,n2052);
or (n2101,n2102,n2124);
and (n2102,n2103,n2123);
xor (n2103,n2104,n2105);
xor (n2104,n2053,n2059);
or (n2105,n2106,n2122);
and (n2106,n2107,n2116);
xor (n2107,n2108,n2109);
nor (n2108,n227,n117);
nand (n2109,n2110,n2115);
or (n2110,n2111,n626);
not (n2111,n2112);
nand (n2112,n2113,n2114);
or (n2113,n126,n424);
nand (n2114,n424,n126);
or (n2115,n2061,n627);
nand (n2116,n2117,n2121);
or (n2117,n122,n2118);
nor (n2118,n2119,n2120);
and (n2119,n136,n453);
and (n2120,n137,n457);
or (n2121,n2088,n123);
and (n2122,n2108,n2109);
xor (n2123,n2079,n2092);
and (n2124,n2104,n2105);
or (n2125,n2126,n2127);
xor (n2126,n2036,n2067);
or (n2127,n2128,n2129);
and (n2128,n2076,n2100);
and (n2129,n2077,n2099);
nor (n2130,n2131,n2256);
and (n2131,n2132,n2251);
or (n2132,n2133,n2250);
and (n2133,n2134,n2175);
xor (n2134,n2135,n2168);
or (n2135,n2136,n2167);
and (n2136,n2137,n2153);
xor (n2137,n2138,n2144);
nand (n2138,n2139,n2143);
or (n2139,n122,n2140);
nor (n2140,n2141,n2142);
and (n2141,n137,n564);
and (n2142,n136,n560);
or (n2143,n2118,n123);
or (n2144,n2145,n2149);
nor (n2145,n2146,n498);
nor (n2146,n2147,n2148);
and (n2147,n236,n590);
and (n2148,n229,n594);
nor (n2149,n497,n2150);
nor (n2150,n2151,n2152);
and (n2151,n229,n117);
and (n2152,n236,n118);
xor (n2153,n2154,n2160);
nor (n2154,n2155,n236);
nor (n2155,n2156,n2159);
and (n2156,n2157,n136);
not (n2157,n2158);
and (n2158,n118,n501);
and (n2159,n507,n117);
nand (n2160,n2161,n2166);
or (n2161,n626,n2162);
not (n2162,n2163);
nand (n2163,n2164,n2165);
or (n2164,n125,n461);
nand (n2165,n461,n125);
nand (n2166,n2112,n628);
and (n2167,n2138,n2144);
xor (n2168,n2169,n2174);
xor (n2169,n2170,n2173);
nand (n2170,n2171,n2172);
or (n2171,n497,n2146);
or (n2172,n2094,n498);
and (n2173,n2154,n2160);
xor (n2174,n2107,n2116);
or (n2175,n2176,n2249);
and (n2176,n2177,n2197);
xor (n2177,n2178,n2196);
or (n2178,n2179,n2195);
and (n2179,n2180,n2189);
xor (n2180,n2181,n2182);
and (n2181,n499,n118);
nand (n2182,n2183,n2188);
or (n2183,n626,n2184);
not (n2184,n2185);
nand (n2185,n2186,n2187);
or (n2186,n126,n457);
nand (n2187,n457,n126);
nand (n2188,n2163,n628);
nand (n2189,n2190,n2194);
or (n2190,n122,n2191);
nor (n2191,n2192,n2193);
and (n2192,n136,n590);
and (n2193,n137,n594);
or (n2194,n2140,n123);
and (n2195,n2181,n2182);
xor (n2196,n2137,n2153);
or (n2197,n2198,n2248);
and (n2198,n2199,n2216);
xor (n2199,n2200,n2215);
and (n2200,n2201,n2207);
and (n2201,n2202,n137);
nand (n2202,n2203,n2206);
nand (n2203,n2204,n125);
not (n2204,n2205);
and (n2205,n118,n129);
nand (n2206,n133,n117);
nand (n2207,n2208,n2209);
or (n2208,n627,n2184);
nand (n2209,n2210,n2214);
not (n2210,n2211);
nor (n2211,n2212,n2213);
and (n2212,n564,n126);
and (n2213,n560,n125);
not (n2214,n626);
xor (n2215,n2180,n2189);
or (n2216,n2217,n2247);
and (n2217,n2218,n2226);
xor (n2218,n2219,n2225);
nand (n2219,n2220,n2224);
or (n2220,n122,n2221);
nor (n2221,n2222,n2223);
and (n2222,n137,n117);
and (n2223,n136,n118);
or (n2224,n2191,n123);
xor (n2225,n2201,n2207);
or (n2226,n2227,n2246);
and (n2227,n2228,n2236);
xor (n2228,n2229,n2230);
nor (n2229,n123,n117);
nand (n2230,n2231,n2235);
or (n2231,n2232,n626);
or (n2232,n2233,n2234);
and (n2233,n125,n594);
and (n2234,n590,n126);
or (n2235,n2211,n627);
nor (n2236,n2237,n2244);
nor (n2237,n2238,n2240);
and (n2238,n2239,n628);
not (n2239,n2232);
and (n2240,n2241,n2214);
nand (n2241,n2242,n2243);
or (n2242,n125,n118);
or (n2243,n126,n117);
or (n2244,n125,n2245);
and (n2245,n118,n628);
and (n2246,n2229,n2230);
and (n2247,n2219,n2225);
and (n2248,n2200,n2215);
and (n2249,n2178,n2196);
and (n2250,n2135,n2168);
or (n2251,n2252,n2253);
xor (n2252,n2103,n2123);
or (n2253,n2254,n2255);
and (n2254,n2169,n2174);
and (n2255,n2170,n2173);
and (n2256,n2252,n2253);
nand (n2257,n2125,n2258);
and (n2258,n2075,n2101);
nand (n2259,n2126,n2127);
and (n2260,n2034,n2069);
and (n2261,n1911,n2016);
or (n2262,n2263,n2270);
xor (n2263,n2264,n2269);
xor (n2264,n2265,n2266);
xor (n2265,n1741,n1761);
or (n2266,n2267,n2268);
and (n2267,n2023,n2030);
and (n2268,n2024,n2027);
xor (n2269,n1880,n1883);
or (n2270,n2271,n2272);
and (n2271,n2017,n2022);
and (n2272,n2018,n2019);
nor (n2273,n2274,n2275);
xor (n2274,n1877,n1902);
or (n2275,n2276,n2277);
and (n2276,n2264,n2269);
and (n2277,n2265,n2266);
or (n2278,n2273,n2279);
nand (n2279,n2263,n2270);
nand (n2280,n2274,n2275);
and (n2281,n1875,n1904);
and (n2282,n1555,n1786);
nor (n2283,n2284,n2404);
nor (n2284,n2285,n2395);
xor (n2285,n2286,n2350);
xor (n2286,n2287,n2325);
xor (n2287,n2288,n2310);
xor (n2288,n2289,n2290);
xor (n2289,n1492,n1505);
xor (n2290,n2291,n2304);
xor (n2291,n2292,n2298);
nand (n2292,n2293,n2297);
or (n2293,n122,n2294);
nor (n2294,n2295,n2296);
and (n2295,n136,n655);
and (n2296,n659,n137);
or (n2297,n123,n1424);
nand (n2298,n2299,n2303);
or (n2299,n335,n2300);
nor (n2300,n2301,n2302);
and (n2301,n346,n328);
and (n2302,n341,n332);
or (n2303,n1443,n347);
nand (n2304,n2305,n2309);
or (n2305,n2306,n497);
nor (n2306,n2307,n2308);
and (n2307,n396,n236);
and (n2308,n400,n229);
or (n2309,n498,n1449);
xor (n2310,n2311,n2324);
xor (n2311,n2312,n2318);
nand (n2312,n2313,n2317);
or (n2313,n642,n2314);
nor (n2314,n2315,n2316);
and (n2315,n384,n429);
and (n2316,n380,n433);
or (n2317,n1455,n643);
nand (n2318,n2319,n2323);
or (n2319,n370,n2320);
nor (n2320,n2321,n2322);
and (n2321,n268,n461);
and (n2322,n465,n269);
or (n2323,n393,n1473);
xor (n2324,n1478,n1484);
or (n2325,n2326,n2349);
and (n2326,n2327,n2334);
xor (n2327,n2328,n2331);
or (n2328,n2329,n2330);
and (n2329,n1849,n1869);
and (n2330,n1850,n1856);
or (n2331,n2332,n2333);
and (n2332,n1789,n1796);
and (n2333,n1790,n1793);
xor (n2334,n2335,n2346);
xor (n2335,n2336,n2337);
and (n2336,n1857,n1863);
xor (n2337,n2338,n2343);
xor (n2338,n2339,n2340);
nor (n2339,n304,n117);
nand (n2340,n2341,n2342);
or (n2341,n1860,n626);
or (n2342,n1486,n627);
nand (n2343,n2344,n2345);
or (n2344,n122,n1827);
or (n2345,n123,n2294);
or (n2346,n2347,n2348);
and (n2347,n1823,n1839);
and (n2348,n1824,n1830);
and (n2349,n2328,n2331);
xor (n2350,n2351,n2386);
xor (n2351,n2352,n2355);
or (n2352,n2353,n2354);
and (n2353,n2335,n2346);
and (n2354,n2336,n2337);
xor (n2355,n2356,n2373);
xor (n2356,n2357,n2360);
or (n2357,n2358,n2359);
and (n2358,n2338,n2343);
and (n2359,n2339,n2340);
or (n2360,n2361,n2372);
and (n2361,n2362,n2369);
xor (n2362,n2363,n2366);
nand (n2363,n2364,n2365);
or (n2364,n497,n1807);
or (n2365,n498,n2306);
nand (n2366,n2367,n2368);
or (n2367,n1812,n642);
or (n2368,n2314,n643);
nand (n2369,n2370,n2371);
or (n2370,n370,n1853);
or (n2371,n2320,n393);
and (n2372,n2363,n2366);
or (n2373,n2374,n2385);
and (n2374,n2375,n2382);
xor (n2375,n2376,n2379);
nand (n2376,n2377,n2378);
or (n2377,n264,n1836);
or (n2378,n1501,n292);
nand (n2379,n2380,n2381);
or (n2380,n226,n1841);
or (n2381,n1495,n227);
nand (n2382,n2383,n2384);
or (n2383,n335,n1801);
or (n2384,n2300,n347);
and (n2385,n2376,n2379);
or (n2386,n2387,n2394);
and (n2387,n2388,n2393);
xor (n2388,n2389,n2392);
or (n2389,n2390,n2391);
and (n2390,n1797,n1810);
and (n2391,n1798,n1804);
xor (n2392,n2362,n2369);
xor (n2393,n2375,n2382);
and (n2394,n2389,n2392);
or (n2395,n2396,n2403);
and (n2396,n2397,n2402);
xor (n2397,n2398,n2399);
xor (n2398,n2388,n2393);
or (n2399,n2400,n2401);
and (n2400,n1821,n1848);
and (n2401,n1822,n1845);
xor (n2402,n2327,n2334);
and (n2403,n2398,n2399);
nor (n2404,n2405,n2406);
xor (n2405,n2397,n2402);
or (n2406,n2407,n2408);
and (n2407,n1787,n1820);
and (n2408,n1788,n1817);
or (n2409,n2410,n2455);
nor (n2410,n2411,n2446);
xor (n2411,n2412,n2431);
xor (n2412,n2413,n2414);
xor (n2413,n1466,n1514);
or (n2414,n2415,n2430);
and (n2415,n2416,n2423);
xor (n2416,n2417,n2420);
or (n2417,n2418,n2419);
and (n2418,n2356,n2373);
and (n2419,n2357,n2360);
or (n2420,n2421,n2422);
and (n2421,n2288,n2310);
and (n2422,n2289,n2290);
xor (n2423,n2424,n2429);
xor (n2424,n2425,n2428);
or (n2425,n2426,n2427);
and (n2426,n2291,n2304);
and (n2427,n2292,n2298);
xor (n2428,n1440,n1453);
xor (n2429,n1392,n1400);
and (n2430,n2417,n2420);
xor (n2431,n2432,n2437);
xor (n2432,n2433,n2436);
or (n2433,n2434,n2435);
and (n2434,n2424,n2429);
and (n2435,n2425,n2428);
xor (n2436,n1437,n1461);
or (n2437,n2438,n2445);
and (n2438,n2439,n2444);
xor (n2439,n2440,n2441);
xor (n2440,n1409,n1422);
or (n2441,n2442,n2443);
and (n2442,n2311,n2324);
and (n2443,n2312,n2318);
xor (n2444,n1470,n1490);
and (n2445,n2440,n2441);
or (n2446,n2447,n2454);
and (n2447,n2448,n2453);
xor (n2448,n2449,n2450);
xor (n2449,n2439,n2444);
or (n2450,n2451,n2452);
and (n2451,n2351,n2386);
and (n2452,n2352,n2355);
xor (n2453,n2416,n2423);
and (n2454,n2449,n2450);
nor (n2455,n2456,n2459);
or (n2456,n2457,n2458);
and (n2457,n2286,n2350);
and (n2458,n2287,n2325);
xor (n2459,n2448,n2453);
nand (n2460,n2461,n2470);
or (n2461,n2462,n2410);
nor (n2462,n2463,n2469);
and (n2463,n2464,n2468);
nand (n2464,n2465,n2467);
or (n2465,n2284,n2466);
nand (n2466,n2405,n2406);
nand (n2467,n2285,n2395);
not (n2468,n2455);
and (n2469,n2456,n2459);
nand (n2470,n2411,n2446);
or (n2471,n2472,n2479);
xor (n2472,n2473,n2478);
xor (n2473,n2474,n2475);
xor (n2474,n1384,n1430);
or (n2475,n2476,n2477);
and (n2476,n2432,n2437);
and (n2477,n2433,n2436);
xor (n2478,n1434,n1464);
or (n2479,n2480,n2481);
and (n2480,n2412,n2431);
and (n2481,n2413,n2414);
and (n2482,n2483,n2485);
not (n2483,n2484);
xor (n2484,n1194,n1432);
not (n2485,n2486);
or (n2486,n2487,n2488);
and (n2487,n2473,n2478);
and (n2488,n2474,n2475);
nor (n2489,n2490,n2494);
and (n2490,n2491,n2492);
not (n2491,n2482);
not (n2492,n2493);
nand (n2493,n2472,n2479);
nor (n2494,n2483,n2485);
and (n2495,n1192,n1518);
nand (n2496,n2497,n2501);
not (n2497,n2498);
or (n2498,n2499,n2500);
and (n2499,n1519,n1542);
and (n2500,n1520,n1529);
not (n2501,n2502);
xor (n2502,n2503,n2508);
xor (n2503,n2504,n2505);
xor (n2504,n895,n931);
or (n2505,n2506,n2507);
and (n2506,n1530,n1539);
and (n2507,n1531,n1532);
xor (n2508,n2509,n2514);
xor (n2509,n2510,n2511);
xor (n2510,n669,n720);
or (n2511,n2512,n2513);
and (n2512,n1533,n1536);
and (n2513,n1534,n1535);
or (n2514,n2515,n2516);
and (n2515,n1521,n1526);
and (n2516,n1522,n1523);
nor (n2517,n2501,n2497);
and (n2518,n2519,n2529);
not (n2519,n2520);
or (n2520,n2521,n2528);
and (n2521,n2522,n2525);
xor (n2522,n2523,n2524);
xor (n2523,n1026,n1031);
xor (n2524,n666,n893);
or (n2525,n2526,n2527);
and (n2526,n2509,n2514);
and (n2527,n2510,n2511);
and (n2528,n2523,n2524);
not (n2529,n2530);
xor (n2530,n4,n972);
nor (n2531,n2532,n2533);
xor (n2532,n2522,n2525);
or (n2533,n2534,n2535);
and (n2534,n2503,n2508);
and (n2535,n2504,n2505);
nor (n2536,n2537,n2541);
and (n2537,n2538,n2539);
not (n2538,n2518);
not (n2539,n2540);
nand (n2540,n2532,n2533);
nor (n2541,n2519,n2529);
xor (n2542,n2543,n4480);
xor (n2543,n2544,n4477);
xor (n2544,n2545,n4476);
xor (n2545,n2546,n4468);
xor (n2546,n2547,n4467);
xor (n2547,n2548,n4452);
xor (n2548,n2549,n4451);
xor (n2549,n2550,n4431);
xor (n2550,n2551,n4430);
xor (n2551,n2552,n4403);
xor (n2552,n2553,n4402);
xor (n2553,n2554,n4370);
xor (n2554,n2555,n4369);
xor (n2555,n2556,n4330);
xor (n2556,n2557,n4329);
xor (n2557,n2558,n4285);
xor (n2558,n2559,n4284);
xor (n2559,n2560,n4233);
xor (n2560,n2561,n4232);
xor (n2561,n2562,n4176);
xor (n2562,n2563,n4175);
xor (n2563,n2564,n4112);
xor (n2564,n2565,n4111);
xor (n2565,n2566,n4043);
xor (n2566,n2567,n4042);
xor (n2567,n2568,n3967);
xor (n2568,n2569,n3966);
xor (n2569,n2570,n3886);
xor (n2570,n2571,n3885);
xor (n2571,n2572,n3798);
xor (n2572,n2573,n3797);
xor (n2573,n2574,n3705);
xor (n2574,n2575,n3704);
xor (n2575,n2576,n3605);
xor (n2576,n2577,n3604);
xor (n2577,n2578,n3500);
xor (n2578,n2579,n3499);
xor (n2579,n2580,n3389);
xor (n2580,n2581,n3388);
xor (n2581,n2582,n3272);
xor (n2582,n2583,n3271);
xor (n2583,n2584,n3148);
xor (n2584,n2585,n3147);
xor (n2585,n2586,n3019);
xor (n2586,n2587,n3018);
xor (n2587,n2588,n2883);
xor (n2588,n2589,n2882);
xor (n2589,n2590,n2742);
xor (n2590,n2591,n2741);
xor (n2591,n2592,n2595);
xor (n2592,n2593,n2594);
and (n2593,n1050,n628);
and (n2594,n632,n126);
or (n2595,n2596,n2599);
and (n2596,n2597,n2598);
and (n2597,n632,n628);
and (n2598,n615,n126);
and (n2599,n2600,n2601);
xor (n2600,n2597,n2598);
or (n2601,n2602,n2605);
and (n2602,n2603,n2604);
and (n2603,n615,n628);
and (n2604,n831,n126);
and (n2605,n2606,n2607);
xor (n2606,n2603,n2604);
or (n2607,n2608,n2611);
and (n2608,n2609,n2610);
and (n2609,n831,n628);
and (n2610,n216,n126);
and (n2611,n2612,n2613);
xor (n2612,n2609,n2610);
or (n2613,n2614,n2617);
and (n2614,n2615,n2616);
and (n2615,n216,n628);
and (n2616,n143,n126);
and (n2617,n2618,n2619);
xor (n2618,n2615,n2616);
or (n2619,n2620,n2623);
and (n2620,n2621,n2622);
and (n2621,n143,n628);
and (n2622,n511,n126);
and (n2623,n2624,n2625);
xor (n2624,n2621,n2622);
or (n2625,n2626,n2629);
and (n2626,n2627,n2628);
and (n2627,n511,n628);
and (n2628,n476,n126);
and (n2629,n2630,n2631);
xor (n2630,n2627,n2628);
or (n2631,n2632,n2635);
and (n2632,n2633,n2634);
and (n2633,n476,n628);
and (n2634,n255,n126);
and (n2635,n2636,n2637);
xor (n2636,n2633,n2634);
or (n2637,n2638,n2641);
and (n2638,n2639,n2640);
and (n2639,n255,n628);
and (n2640,n247,n126);
and (n2641,n2642,n2643);
xor (n2642,n2639,n2640);
or (n2643,n2644,n2647);
and (n2644,n2645,n2646);
and (n2645,n247,n628);
and (n2646,n361,n126);
and (n2647,n2648,n2649);
xor (n2648,n2645,n2646);
or (n2649,n2650,n2653);
and (n2650,n2651,n2652);
and (n2651,n361,n628);
and (n2652,n353,n126);
and (n2653,n2654,n2655);
xor (n2654,n2651,n2652);
or (n2655,n2656,n2659);
and (n2656,n2657,n2658);
and (n2657,n353,n628);
and (n2658,n655,n126);
and (n2659,n2660,n2661);
xor (n2660,n2657,n2658);
or (n2661,n2662,n2665);
and (n2662,n2663,n2664);
and (n2663,n655,n628);
and (n2664,n525,n126);
and (n2665,n2666,n2667);
xor (n2666,n2663,n2664);
or (n2667,n2668,n2671);
and (n2668,n2669,n2670);
and (n2669,n525,n628);
and (n2670,n396,n126);
and (n2671,n2672,n2673);
xor (n2672,n2669,n2670);
or (n2673,n2674,n2677);
and (n2674,n2675,n2676);
and (n2675,n396,n628);
and (n2676,n387,n126);
and (n2677,n2678,n2679);
xor (n2678,n2675,n2676);
or (n2679,n2680,n2683);
and (n2680,n2681,n2682);
and (n2681,n387,n628);
and (n2682,n295,n126);
and (n2683,n2684,n2685);
xor (n2684,n2681,n2682);
or (n2685,n2686,n2689);
and (n2686,n2687,n2688);
and (n2687,n295,n628);
and (n2688,n286,n126);
and (n2689,n2690,n2691);
xor (n2690,n2687,n2688);
or (n2691,n2692,n2695);
and (n2692,n2693,n2694);
and (n2693,n286,n628);
and (n2694,n328,n126);
and (n2695,n2696,n2697);
xor (n2696,n2693,n2694);
or (n2697,n2698,n2701);
and (n2698,n2699,n2700);
and (n2699,n328,n628);
and (n2700,n320,n126);
and (n2701,n2702,n2703);
xor (n2702,n2699,n2700);
or (n2703,n2704,n2707);
and (n2704,n2705,n2706);
and (n2705,n320,n628);
and (n2706,n429,n126);
and (n2707,n2708,n2709);
xor (n2708,n2705,n2706);
or (n2709,n2710,n2713);
and (n2710,n2711,n2712);
and (n2711,n429,n628);
and (n2712,n420,n126);
and (n2713,n2714,n2715);
xor (n2714,n2711,n2712);
or (n2715,n2716,n2719);
and (n2716,n2717,n2718);
and (n2717,n420,n628);
and (n2718,n461,n126);
and (n2719,n2720,n2721);
xor (n2720,n2717,n2718);
or (n2721,n2722,n2725);
and (n2722,n2723,n2724);
and (n2723,n461,n628);
and (n2724,n453,n126);
and (n2725,n2726,n2727);
xor (n2726,n2723,n2724);
or (n2727,n2728,n2731);
and (n2728,n2729,n2730);
and (n2729,n453,n628);
and (n2730,n560,n126);
and (n2731,n2732,n2733);
xor (n2732,n2729,n2730);
or (n2733,n2734,n2736);
and (n2734,n2735,n2234);
and (n2735,n560,n628);
and (n2736,n2737,n2738);
xor (n2737,n2735,n2234);
and (n2738,n2739,n2740);
and (n2739,n590,n628);
and (n2740,n118,n126);
and (n2741,n615,n129);
or (n2742,n2743,n2746);
and (n2743,n2744,n2745);
xor (n2744,n2600,n2601);
and (n2745,n831,n129);
and (n2746,n2747,n2748);
xor (n2747,n2744,n2745);
or (n2748,n2749,n2752);
and (n2749,n2750,n2751);
xor (n2750,n2606,n2607);
and (n2751,n216,n129);
and (n2752,n2753,n2754);
xor (n2753,n2750,n2751);
or (n2754,n2755,n2758);
and (n2755,n2756,n2757);
xor (n2756,n2612,n2613);
and (n2757,n143,n129);
and (n2758,n2759,n2760);
xor (n2759,n2756,n2757);
or (n2760,n2761,n2764);
and (n2761,n2762,n2763);
xor (n2762,n2618,n2619);
and (n2763,n511,n129);
and (n2764,n2765,n2766);
xor (n2765,n2762,n2763);
or (n2766,n2767,n2770);
and (n2767,n2768,n2769);
xor (n2768,n2624,n2625);
and (n2769,n476,n129);
and (n2770,n2771,n2772);
xor (n2771,n2768,n2769);
or (n2772,n2773,n2776);
and (n2773,n2774,n2775);
xor (n2774,n2630,n2631);
and (n2775,n255,n129);
and (n2776,n2777,n2778);
xor (n2777,n2774,n2775);
or (n2778,n2779,n2782);
and (n2779,n2780,n2781);
xor (n2780,n2636,n2637);
and (n2781,n247,n129);
and (n2782,n2783,n2784);
xor (n2783,n2780,n2781);
or (n2784,n2785,n2788);
and (n2785,n2786,n2787);
xor (n2786,n2642,n2643);
and (n2787,n361,n129);
and (n2788,n2789,n2790);
xor (n2789,n2786,n2787);
or (n2790,n2791,n2794);
and (n2791,n2792,n2793);
xor (n2792,n2648,n2649);
and (n2793,n353,n129);
and (n2794,n2795,n2796);
xor (n2795,n2792,n2793);
or (n2796,n2797,n2800);
and (n2797,n2798,n2799);
xor (n2798,n2654,n2655);
and (n2799,n655,n129);
and (n2800,n2801,n2802);
xor (n2801,n2798,n2799);
or (n2802,n2803,n2806);
and (n2803,n2804,n2805);
xor (n2804,n2660,n2661);
and (n2805,n525,n129);
and (n2806,n2807,n2808);
xor (n2807,n2804,n2805);
or (n2808,n2809,n2812);
and (n2809,n2810,n2811);
xor (n2810,n2666,n2667);
and (n2811,n396,n129);
and (n2812,n2813,n2814);
xor (n2813,n2810,n2811);
or (n2814,n2815,n2818);
and (n2815,n2816,n2817);
xor (n2816,n2672,n2673);
and (n2817,n387,n129);
and (n2818,n2819,n2820);
xor (n2819,n2816,n2817);
or (n2820,n2821,n2824);
and (n2821,n2822,n2823);
xor (n2822,n2678,n2679);
and (n2823,n295,n129);
and (n2824,n2825,n2826);
xor (n2825,n2822,n2823);
or (n2826,n2827,n2830);
and (n2827,n2828,n2829);
xor (n2828,n2684,n2685);
and (n2829,n286,n129);
and (n2830,n2831,n2832);
xor (n2831,n2828,n2829);
or (n2832,n2833,n2836);
and (n2833,n2834,n2835);
xor (n2834,n2690,n2691);
and (n2835,n328,n129);
and (n2836,n2837,n2838);
xor (n2837,n2834,n2835);
or (n2838,n2839,n2842);
and (n2839,n2840,n2841);
xor (n2840,n2696,n2697);
and (n2841,n320,n129);
and (n2842,n2843,n2844);
xor (n2843,n2840,n2841);
or (n2844,n2845,n2848);
and (n2845,n2846,n2847);
xor (n2846,n2702,n2703);
and (n2847,n429,n129);
and (n2848,n2849,n2850);
xor (n2849,n2846,n2847);
or (n2850,n2851,n2854);
and (n2851,n2852,n2853);
xor (n2852,n2708,n2709);
and (n2853,n420,n129);
and (n2854,n2855,n2856);
xor (n2855,n2852,n2853);
or (n2856,n2857,n2860);
and (n2857,n2858,n2859);
xor (n2858,n2714,n2715);
and (n2859,n461,n129);
and (n2860,n2861,n2862);
xor (n2861,n2858,n2859);
or (n2862,n2863,n2866);
and (n2863,n2864,n2865);
xor (n2864,n2720,n2721);
and (n2865,n453,n129);
and (n2866,n2867,n2868);
xor (n2867,n2864,n2865);
or (n2868,n2869,n2872);
and (n2869,n2870,n2871);
xor (n2870,n2726,n2727);
and (n2871,n560,n129);
and (n2872,n2873,n2874);
xor (n2873,n2870,n2871);
or (n2874,n2875,n2878);
and (n2875,n2876,n2877);
xor (n2876,n2732,n2733);
and (n2877,n590,n129);
and (n2878,n2879,n2880);
xor (n2879,n2876,n2877);
and (n2880,n2881,n2205);
xor (n2881,n2737,n2738);
and (n2882,n831,n137);
or (n2883,n2884,n2887);
and (n2884,n2885,n2886);
xor (n2885,n2747,n2748);
and (n2886,n216,n137);
and (n2887,n2888,n2889);
xor (n2888,n2885,n2886);
or (n2889,n2890,n2893);
and (n2890,n2891,n2892);
xor (n2891,n2753,n2754);
and (n2892,n143,n137);
and (n2893,n2894,n2895);
xor (n2894,n2891,n2892);
or (n2895,n2896,n2899);
and (n2896,n2897,n2898);
xor (n2897,n2759,n2760);
and (n2898,n511,n137);
and (n2899,n2900,n2901);
xor (n2900,n2897,n2898);
or (n2901,n2902,n2905);
and (n2902,n2903,n2904);
xor (n2903,n2765,n2766);
and (n2904,n476,n137);
and (n2905,n2906,n2907);
xor (n2906,n2903,n2904);
or (n2907,n2908,n2911);
and (n2908,n2909,n2910);
xor (n2909,n2771,n2772);
and (n2910,n255,n137);
and (n2911,n2912,n2913);
xor (n2912,n2909,n2910);
or (n2913,n2914,n2917);
and (n2914,n2915,n2916);
xor (n2915,n2777,n2778);
and (n2916,n247,n137);
and (n2917,n2918,n2919);
xor (n2918,n2915,n2916);
or (n2919,n2920,n2923);
and (n2920,n2921,n2922);
xor (n2921,n2783,n2784);
and (n2922,n361,n137);
and (n2923,n2924,n2925);
xor (n2924,n2921,n2922);
or (n2925,n2926,n2929);
and (n2926,n2927,n2928);
xor (n2927,n2789,n2790);
and (n2928,n353,n137);
and (n2929,n2930,n2931);
xor (n2930,n2927,n2928);
or (n2931,n2932,n2935);
and (n2932,n2933,n2934);
xor (n2933,n2795,n2796);
and (n2934,n655,n137);
and (n2935,n2936,n2937);
xor (n2936,n2933,n2934);
or (n2937,n2938,n2941);
and (n2938,n2939,n2940);
xor (n2939,n2801,n2802);
and (n2940,n525,n137);
and (n2941,n2942,n2943);
xor (n2942,n2939,n2940);
or (n2943,n2944,n2947);
and (n2944,n2945,n2946);
xor (n2945,n2807,n2808);
and (n2946,n396,n137);
and (n2947,n2948,n2949);
xor (n2948,n2945,n2946);
or (n2949,n2950,n2953);
and (n2950,n2951,n2952);
xor (n2951,n2813,n2814);
and (n2952,n387,n137);
and (n2953,n2954,n2955);
xor (n2954,n2951,n2952);
or (n2955,n2956,n2959);
and (n2956,n2957,n2958);
xor (n2957,n2819,n2820);
and (n2958,n295,n137);
and (n2959,n2960,n2961);
xor (n2960,n2957,n2958);
or (n2961,n2962,n2965);
and (n2962,n2963,n2964);
xor (n2963,n2825,n2826);
and (n2964,n286,n137);
and (n2965,n2966,n2967);
xor (n2966,n2963,n2964);
or (n2967,n2968,n2971);
and (n2968,n2969,n2970);
xor (n2969,n2831,n2832);
and (n2970,n328,n137);
and (n2971,n2972,n2973);
xor (n2972,n2969,n2970);
or (n2973,n2974,n2977);
and (n2974,n2975,n2976);
xor (n2975,n2837,n2838);
and (n2976,n320,n137);
and (n2977,n2978,n2979);
xor (n2978,n2975,n2976);
or (n2979,n2980,n2983);
and (n2980,n2981,n2982);
xor (n2981,n2843,n2844);
and (n2982,n429,n137);
and (n2983,n2984,n2985);
xor (n2984,n2981,n2982);
or (n2985,n2986,n2989);
and (n2986,n2987,n2988);
xor (n2987,n2849,n2850);
and (n2988,n420,n137);
and (n2989,n2990,n2991);
xor (n2990,n2987,n2988);
or (n2991,n2992,n2995);
and (n2992,n2993,n2994);
xor (n2993,n2855,n2856);
and (n2994,n461,n137);
and (n2995,n2996,n2997);
xor (n2996,n2993,n2994);
or (n2997,n2998,n3001);
and (n2998,n2999,n3000);
xor (n2999,n2861,n2862);
and (n3000,n453,n137);
and (n3001,n3002,n3003);
xor (n3002,n2999,n3000);
or (n3003,n3004,n3007);
and (n3004,n3005,n3006);
xor (n3005,n2867,n2868);
and (n3006,n560,n137);
and (n3007,n3008,n3009);
xor (n3008,n3005,n3006);
or (n3009,n3010,n3013);
and (n3010,n3011,n3012);
xor (n3011,n2873,n2874);
and (n3012,n590,n137);
and (n3013,n3014,n3015);
xor (n3014,n3011,n3012);
and (n3015,n3016,n3017);
xor (n3016,n2879,n2880);
and (n3017,n118,n137);
and (n3018,n216,n501);
or (n3019,n3020,n3023);
and (n3020,n3021,n3022);
xor (n3021,n2888,n2889);
and (n3022,n143,n501);
and (n3023,n3024,n3025);
xor (n3024,n3021,n3022);
or (n3025,n3026,n3029);
and (n3026,n3027,n3028);
xor (n3027,n2894,n2895);
and (n3028,n511,n501);
and (n3029,n3030,n3031);
xor (n3030,n3027,n3028);
or (n3031,n3032,n3035);
and (n3032,n3033,n3034);
xor (n3033,n2900,n2901);
and (n3034,n476,n501);
and (n3035,n3036,n3037);
xor (n3036,n3033,n3034);
or (n3037,n3038,n3041);
and (n3038,n3039,n3040);
xor (n3039,n2906,n2907);
and (n3040,n255,n501);
and (n3041,n3042,n3043);
xor (n3042,n3039,n3040);
or (n3043,n3044,n3047);
and (n3044,n3045,n3046);
xor (n3045,n2912,n2913);
and (n3046,n247,n501);
and (n3047,n3048,n3049);
xor (n3048,n3045,n3046);
or (n3049,n3050,n3053);
and (n3050,n3051,n3052);
xor (n3051,n2918,n2919);
and (n3052,n361,n501);
and (n3053,n3054,n3055);
xor (n3054,n3051,n3052);
or (n3055,n3056,n3059);
and (n3056,n3057,n3058);
xor (n3057,n2924,n2925);
and (n3058,n353,n501);
and (n3059,n3060,n3061);
xor (n3060,n3057,n3058);
or (n3061,n3062,n3065);
and (n3062,n3063,n3064);
xor (n3063,n2930,n2931);
and (n3064,n655,n501);
and (n3065,n3066,n3067);
xor (n3066,n3063,n3064);
or (n3067,n3068,n3071);
and (n3068,n3069,n3070);
xor (n3069,n2936,n2937);
and (n3070,n525,n501);
and (n3071,n3072,n3073);
xor (n3072,n3069,n3070);
or (n3073,n3074,n3077);
and (n3074,n3075,n3076);
xor (n3075,n2942,n2943);
and (n3076,n396,n501);
and (n3077,n3078,n3079);
xor (n3078,n3075,n3076);
or (n3079,n3080,n3083);
and (n3080,n3081,n3082);
xor (n3081,n2948,n2949);
and (n3082,n387,n501);
and (n3083,n3084,n3085);
xor (n3084,n3081,n3082);
or (n3085,n3086,n3089);
and (n3086,n3087,n3088);
xor (n3087,n2954,n2955);
and (n3088,n295,n501);
and (n3089,n3090,n3091);
xor (n3090,n3087,n3088);
or (n3091,n3092,n3095);
and (n3092,n3093,n3094);
xor (n3093,n2960,n2961);
and (n3094,n286,n501);
and (n3095,n3096,n3097);
xor (n3096,n3093,n3094);
or (n3097,n3098,n3101);
and (n3098,n3099,n3100);
xor (n3099,n2966,n2967);
and (n3100,n328,n501);
and (n3101,n3102,n3103);
xor (n3102,n3099,n3100);
or (n3103,n3104,n3107);
and (n3104,n3105,n3106);
xor (n3105,n2972,n2973);
and (n3106,n320,n501);
and (n3107,n3108,n3109);
xor (n3108,n3105,n3106);
or (n3109,n3110,n3113);
and (n3110,n3111,n3112);
xor (n3111,n2978,n2979);
and (n3112,n429,n501);
and (n3113,n3114,n3115);
xor (n3114,n3111,n3112);
or (n3115,n3116,n3119);
and (n3116,n3117,n3118);
xor (n3117,n2984,n2985);
and (n3118,n420,n501);
and (n3119,n3120,n3121);
xor (n3120,n3117,n3118);
or (n3121,n3122,n3125);
and (n3122,n3123,n3124);
xor (n3123,n2990,n2991);
and (n3124,n461,n501);
and (n3125,n3126,n3127);
xor (n3126,n3123,n3124);
or (n3127,n3128,n3131);
and (n3128,n3129,n3130);
xor (n3129,n2996,n2997);
and (n3130,n453,n501);
and (n3131,n3132,n3133);
xor (n3132,n3129,n3130);
or (n3133,n3134,n3137);
and (n3134,n3135,n3136);
xor (n3135,n3002,n3003);
and (n3136,n560,n501);
and (n3137,n3138,n3139);
xor (n3138,n3135,n3136);
or (n3139,n3140,n3143);
and (n3140,n3141,n3142);
xor (n3141,n3008,n3009);
and (n3142,n590,n501);
and (n3143,n3144,n3145);
xor (n3144,n3141,n3142);
and (n3145,n3146,n2158);
xor (n3146,n3014,n3015);
and (n3147,n143,n229);
or (n3148,n3149,n3152);
and (n3149,n3150,n3151);
xor (n3150,n3024,n3025);
and (n3151,n511,n229);
and (n3152,n3153,n3154);
xor (n3153,n3150,n3151);
or (n3154,n3155,n3158);
and (n3155,n3156,n3157);
xor (n3156,n3030,n3031);
and (n3157,n476,n229);
and (n3158,n3159,n3160);
xor (n3159,n3156,n3157);
or (n3160,n3161,n3164);
and (n3161,n3162,n3163);
xor (n3162,n3036,n3037);
and (n3163,n255,n229);
and (n3164,n3165,n3166);
xor (n3165,n3162,n3163);
or (n3166,n3167,n3170);
and (n3167,n3168,n3169);
xor (n3168,n3042,n3043);
and (n3169,n247,n229);
and (n3170,n3171,n3172);
xor (n3171,n3168,n3169);
or (n3172,n3173,n3176);
and (n3173,n3174,n3175);
xor (n3174,n3048,n3049);
and (n3175,n361,n229);
and (n3176,n3177,n3178);
xor (n3177,n3174,n3175);
or (n3178,n3179,n3182);
and (n3179,n3180,n3181);
xor (n3180,n3054,n3055);
and (n3181,n353,n229);
and (n3182,n3183,n3184);
xor (n3183,n3180,n3181);
or (n3184,n3185,n3188);
and (n3185,n3186,n3187);
xor (n3186,n3060,n3061);
and (n3187,n655,n229);
and (n3188,n3189,n3190);
xor (n3189,n3186,n3187);
or (n3190,n3191,n3194);
and (n3191,n3192,n3193);
xor (n3192,n3066,n3067);
and (n3193,n525,n229);
and (n3194,n3195,n3196);
xor (n3195,n3192,n3193);
or (n3196,n3197,n3200);
and (n3197,n3198,n3199);
xor (n3198,n3072,n3073);
and (n3199,n396,n229);
and (n3200,n3201,n3202);
xor (n3201,n3198,n3199);
or (n3202,n3203,n3206);
and (n3203,n3204,n3205);
xor (n3204,n3078,n3079);
and (n3205,n387,n229);
and (n3206,n3207,n3208);
xor (n3207,n3204,n3205);
or (n3208,n3209,n3212);
and (n3209,n3210,n3211);
xor (n3210,n3084,n3085);
and (n3211,n295,n229);
and (n3212,n3213,n3214);
xor (n3213,n3210,n3211);
or (n3214,n3215,n3218);
and (n3215,n3216,n3217);
xor (n3216,n3090,n3091);
and (n3217,n286,n229);
and (n3218,n3219,n3220);
xor (n3219,n3216,n3217);
or (n3220,n3221,n3224);
and (n3221,n3222,n3223);
xor (n3222,n3096,n3097);
and (n3223,n328,n229);
and (n3224,n3225,n3226);
xor (n3225,n3222,n3223);
or (n3226,n3227,n3230);
and (n3227,n3228,n3229);
xor (n3228,n3102,n3103);
and (n3229,n320,n229);
and (n3230,n3231,n3232);
xor (n3231,n3228,n3229);
or (n3232,n3233,n3236);
and (n3233,n3234,n3235);
xor (n3234,n3108,n3109);
and (n3235,n429,n229);
and (n3236,n3237,n3238);
xor (n3237,n3234,n3235);
or (n3238,n3239,n3242);
and (n3239,n3240,n3241);
xor (n3240,n3114,n3115);
and (n3241,n420,n229);
and (n3242,n3243,n3244);
xor (n3243,n3240,n3241);
or (n3244,n3245,n3248);
and (n3245,n3246,n3247);
xor (n3246,n3120,n3121);
and (n3247,n461,n229);
and (n3248,n3249,n3250);
xor (n3249,n3246,n3247);
or (n3250,n3251,n3254);
and (n3251,n3252,n3253);
xor (n3252,n3126,n3127);
and (n3253,n453,n229);
and (n3254,n3255,n3256);
xor (n3255,n3252,n3253);
or (n3256,n3257,n3260);
and (n3257,n3258,n3259);
xor (n3258,n3132,n3133);
and (n3259,n560,n229);
and (n3260,n3261,n3262);
xor (n3261,n3258,n3259);
or (n3262,n3263,n3266);
and (n3263,n3264,n3265);
xor (n3264,n3138,n3139);
and (n3265,n590,n229);
and (n3266,n3267,n3268);
xor (n3267,n3264,n3265);
and (n3268,n3269,n3270);
xor (n3269,n3144,n3145);
and (n3270,n118,n229);
and (n3271,n511,n232);
or (n3272,n3273,n3276);
and (n3273,n3274,n3275);
xor (n3274,n3153,n3154);
and (n3275,n476,n232);
and (n3276,n3277,n3278);
xor (n3277,n3274,n3275);
or (n3278,n3279,n3282);
and (n3279,n3280,n3281);
xor (n3280,n3159,n3160);
and (n3281,n255,n232);
and (n3282,n3283,n3284);
xor (n3283,n3280,n3281);
or (n3284,n3285,n3288);
and (n3285,n3286,n3287);
xor (n3286,n3165,n3166);
and (n3287,n247,n232);
and (n3288,n3289,n3290);
xor (n3289,n3286,n3287);
or (n3290,n3291,n3294);
and (n3291,n3292,n3293);
xor (n3292,n3171,n3172);
and (n3293,n361,n232);
and (n3294,n3295,n3296);
xor (n3295,n3292,n3293);
or (n3296,n3297,n3300);
and (n3297,n3298,n3299);
xor (n3298,n3177,n3178);
and (n3299,n353,n232);
and (n3300,n3301,n3302);
xor (n3301,n3298,n3299);
or (n3302,n3303,n3306);
and (n3303,n3304,n3305);
xor (n3304,n3183,n3184);
and (n3305,n655,n232);
and (n3306,n3307,n3308);
xor (n3307,n3304,n3305);
or (n3308,n3309,n3312);
and (n3309,n3310,n3311);
xor (n3310,n3189,n3190);
and (n3311,n525,n232);
and (n3312,n3313,n3314);
xor (n3313,n3310,n3311);
or (n3314,n3315,n3318);
and (n3315,n3316,n3317);
xor (n3316,n3195,n3196);
and (n3317,n396,n232);
and (n3318,n3319,n3320);
xor (n3319,n3316,n3317);
or (n3320,n3321,n3324);
and (n3321,n3322,n3323);
xor (n3322,n3201,n3202);
and (n3323,n387,n232);
and (n3324,n3325,n3326);
xor (n3325,n3322,n3323);
or (n3326,n3327,n3330);
and (n3327,n3328,n3329);
xor (n3328,n3207,n3208);
and (n3329,n295,n232);
and (n3330,n3331,n3332);
xor (n3331,n3328,n3329);
or (n3332,n3333,n3336);
and (n3333,n3334,n3335);
xor (n3334,n3213,n3214);
and (n3335,n286,n232);
and (n3336,n3337,n3338);
xor (n3337,n3334,n3335);
or (n3338,n3339,n3342);
and (n3339,n3340,n3341);
xor (n3340,n3219,n3220);
and (n3341,n328,n232);
and (n3342,n3343,n3344);
xor (n3343,n3340,n3341);
or (n3344,n3345,n3348);
and (n3345,n3346,n3347);
xor (n3346,n3225,n3226);
and (n3347,n320,n232);
and (n3348,n3349,n3350);
xor (n3349,n3346,n3347);
or (n3350,n3351,n3354);
and (n3351,n3352,n3353);
xor (n3352,n3231,n3232);
and (n3353,n429,n232);
and (n3354,n3355,n3356);
xor (n3355,n3352,n3353);
or (n3356,n3357,n3360);
and (n3357,n3358,n3359);
xor (n3358,n3237,n3238);
and (n3359,n420,n232);
and (n3360,n3361,n3362);
xor (n3361,n3358,n3359);
or (n3362,n3363,n3366);
and (n3363,n3364,n3365);
xor (n3364,n3243,n3244);
and (n3365,n461,n232);
and (n3366,n3367,n3368);
xor (n3367,n3364,n3365);
or (n3368,n3369,n3372);
and (n3369,n3370,n3371);
xor (n3370,n3249,n3250);
and (n3371,n453,n232);
and (n3372,n3373,n3374);
xor (n3373,n3370,n3371);
or (n3374,n3375,n3378);
and (n3375,n3376,n3377);
xor (n3376,n3255,n3256);
and (n3377,n560,n232);
and (n3378,n3379,n3380);
xor (n3379,n3376,n3377);
or (n3380,n3381,n3384);
and (n3381,n3382,n3383);
xor (n3382,n3261,n3262);
and (n3383,n590,n232);
and (n3384,n3385,n3386);
xor (n3385,n3382,n3383);
and (n3386,n3387,n2057);
xor (n3387,n3267,n3268);
and (n3388,n476,n240);
or (n3389,n3390,n3393);
and (n3390,n3391,n3392);
xor (n3391,n3277,n3278);
and (n3392,n255,n240);
and (n3393,n3394,n3395);
xor (n3394,n3391,n3392);
or (n3395,n3396,n3399);
and (n3396,n3397,n3398);
xor (n3397,n3283,n3284);
and (n3398,n247,n240);
and (n3399,n3400,n3401);
xor (n3400,n3397,n3398);
or (n3401,n3402,n3405);
and (n3402,n3403,n3404);
xor (n3403,n3289,n3290);
and (n3404,n361,n240);
and (n3405,n3406,n3407);
xor (n3406,n3403,n3404);
or (n3407,n3408,n3411);
and (n3408,n3409,n3410);
xor (n3409,n3295,n3296);
and (n3410,n353,n240);
and (n3411,n3412,n3413);
xor (n3412,n3409,n3410);
or (n3413,n3414,n3417);
and (n3414,n3415,n3416);
xor (n3415,n3301,n3302);
and (n3416,n655,n240);
and (n3417,n3418,n3419);
xor (n3418,n3415,n3416);
or (n3419,n3420,n3423);
and (n3420,n3421,n3422);
xor (n3421,n3307,n3308);
and (n3422,n525,n240);
and (n3423,n3424,n3425);
xor (n3424,n3421,n3422);
or (n3425,n3426,n3429);
and (n3426,n3427,n3428);
xor (n3427,n3313,n3314);
and (n3428,n396,n240);
and (n3429,n3430,n3431);
xor (n3430,n3427,n3428);
or (n3431,n3432,n3435);
and (n3432,n3433,n3434);
xor (n3433,n3319,n3320);
and (n3434,n387,n240);
and (n3435,n3436,n3437);
xor (n3436,n3433,n3434);
or (n3437,n3438,n3441);
and (n3438,n3439,n3440);
xor (n3439,n3325,n3326);
and (n3440,n295,n240);
and (n3441,n3442,n3443);
xor (n3442,n3439,n3440);
or (n3443,n3444,n3447);
and (n3444,n3445,n3446);
xor (n3445,n3331,n3332);
and (n3446,n286,n240);
and (n3447,n3448,n3449);
xor (n3448,n3445,n3446);
or (n3449,n3450,n3453);
and (n3450,n3451,n3452);
xor (n3451,n3337,n3338);
and (n3452,n328,n240);
and (n3453,n3454,n3455);
xor (n3454,n3451,n3452);
or (n3455,n3456,n3459);
and (n3456,n3457,n3458);
xor (n3457,n3343,n3344);
and (n3458,n320,n240);
and (n3459,n3460,n3461);
xor (n3460,n3457,n3458);
or (n3461,n3462,n3465);
and (n3462,n3463,n3464);
xor (n3463,n3349,n3350);
and (n3464,n429,n240);
and (n3465,n3466,n3467);
xor (n3466,n3463,n3464);
or (n3467,n3468,n3471);
and (n3468,n3469,n3470);
xor (n3469,n3355,n3356);
and (n3470,n420,n240);
and (n3471,n3472,n3473);
xor (n3472,n3469,n3470);
or (n3473,n3474,n3477);
and (n3474,n3475,n3476);
xor (n3475,n3361,n3362);
and (n3476,n461,n240);
and (n3477,n3478,n3479);
xor (n3478,n3475,n3476);
or (n3479,n3480,n3482);
and (n3480,n3481,n1921);
xor (n3481,n3367,n3368);
and (n3482,n3483,n3484);
xor (n3483,n3481,n1921);
or (n3484,n3485,n3488);
and (n3485,n3486,n3487);
xor (n3486,n3373,n3374);
and (n3487,n560,n240);
and (n3488,n3489,n3490);
xor (n3489,n3486,n3487);
or (n3490,n3491,n3494);
and (n3491,n3492,n3493);
xor (n3492,n3379,n3380);
and (n3493,n590,n240);
and (n3494,n3495,n3496);
xor (n3495,n3492,n3493);
and (n3496,n3497,n3498);
xor (n3497,n3385,n3386);
and (n3498,n118,n240);
and (n3499,n255,n338);
or (n3500,n3501,n3504);
and (n3501,n3502,n3503);
xor (n3502,n3394,n3395);
and (n3503,n247,n338);
and (n3504,n3505,n3506);
xor (n3505,n3502,n3503);
or (n3506,n3507,n3510);
and (n3507,n3508,n3509);
xor (n3508,n3400,n3401);
and (n3509,n361,n338);
and (n3510,n3511,n3512);
xor (n3511,n3508,n3509);
or (n3512,n3513,n3516);
and (n3513,n3514,n3515);
xor (n3514,n3406,n3407);
and (n3515,n353,n338);
and (n3516,n3517,n3518);
xor (n3517,n3514,n3515);
or (n3518,n3519,n3522);
and (n3519,n3520,n3521);
xor (n3520,n3412,n3413);
and (n3521,n655,n338);
and (n3522,n3523,n3524);
xor (n3523,n3520,n3521);
or (n3524,n3525,n3528);
and (n3525,n3526,n3527);
xor (n3526,n3418,n3419);
and (n3527,n525,n338);
and (n3528,n3529,n3530);
xor (n3529,n3526,n3527);
or (n3530,n3531,n3534);
and (n3531,n3532,n3533);
xor (n3532,n3424,n3425);
and (n3533,n396,n338);
and (n3534,n3535,n3536);
xor (n3535,n3532,n3533);
or (n3536,n3537,n3540);
and (n3537,n3538,n3539);
xor (n3538,n3430,n3431);
and (n3539,n387,n338);
and (n3540,n3541,n3542);
xor (n3541,n3538,n3539);
or (n3542,n3543,n3546);
and (n3543,n3544,n3545);
xor (n3544,n3436,n3437);
and (n3545,n295,n338);
and (n3546,n3547,n3548);
xor (n3547,n3544,n3545);
or (n3548,n3549,n3552);
and (n3549,n3550,n3551);
xor (n3550,n3442,n3443);
and (n3551,n286,n338);
and (n3552,n3553,n3554);
xor (n3553,n3550,n3551);
or (n3554,n3555,n3558);
and (n3555,n3556,n3557);
xor (n3556,n3448,n3449);
and (n3557,n328,n338);
and (n3558,n3559,n3560);
xor (n3559,n3556,n3557);
or (n3560,n3561,n3564);
and (n3561,n3562,n3563);
xor (n3562,n3454,n3455);
and (n3563,n320,n338);
and (n3564,n3565,n3566);
xor (n3565,n3562,n3563);
or (n3566,n3567,n3570);
and (n3567,n3568,n3569);
xor (n3568,n3460,n3461);
and (n3569,n429,n338);
and (n3570,n3571,n3572);
xor (n3571,n3568,n3569);
or (n3572,n3573,n3576);
and (n3573,n3574,n3575);
xor (n3574,n3466,n3467);
and (n3575,n420,n338);
and (n3576,n3577,n3578);
xor (n3577,n3574,n3575);
or (n3578,n3579,n3582);
and (n3579,n3580,n3581);
xor (n3580,n3472,n3473);
and (n3581,n461,n338);
and (n3582,n3583,n3584);
xor (n3583,n3580,n3581);
or (n3584,n3585,n3588);
and (n3585,n3586,n3587);
xor (n3586,n3478,n3479);
and (n3587,n453,n338);
and (n3588,n3589,n3590);
xor (n3589,n3586,n3587);
or (n3590,n3591,n3594);
and (n3591,n3592,n3593);
xor (n3592,n3483,n3484);
and (n3593,n560,n338);
and (n3594,n3595,n3596);
xor (n3595,n3592,n3593);
or (n3596,n3597,n3600);
and (n3597,n3598,n3599);
xor (n3598,n3489,n3490);
and (n3599,n590,n338);
and (n3600,n3601,n3602);
xor (n3601,n3598,n3599);
and (n3602,n3603,n1950);
xor (n3603,n3495,n3496);
and (n3604,n247,n341);
or (n3605,n3606,n3609);
and (n3606,n3607,n3608);
xor (n3607,n3505,n3506);
and (n3608,n361,n341);
and (n3609,n3610,n3611);
xor (n3610,n3607,n3608);
or (n3611,n3612,n3615);
and (n3612,n3613,n3614);
xor (n3613,n3511,n3512);
and (n3614,n353,n341);
and (n3615,n3616,n3617);
xor (n3616,n3613,n3614);
or (n3617,n3618,n3621);
and (n3618,n3619,n3620);
xor (n3619,n3517,n3518);
and (n3620,n655,n341);
and (n3621,n3622,n3623);
xor (n3622,n3619,n3620);
or (n3623,n3624,n3627);
and (n3624,n3625,n3626);
xor (n3625,n3523,n3524);
and (n3626,n525,n341);
and (n3627,n3628,n3629);
xor (n3628,n3625,n3626);
or (n3629,n3630,n3633);
and (n3630,n3631,n3632);
xor (n3631,n3529,n3530);
and (n3632,n396,n341);
and (n3633,n3634,n3635);
xor (n3634,n3631,n3632);
or (n3635,n3636,n3639);
and (n3636,n3637,n3638);
xor (n3637,n3535,n3536);
and (n3638,n387,n341);
and (n3639,n3640,n3641);
xor (n3640,n3637,n3638);
or (n3641,n3642,n3645);
and (n3642,n3643,n3644);
xor (n3643,n3541,n3542);
and (n3644,n295,n341);
and (n3645,n3646,n3647);
xor (n3646,n3643,n3644);
or (n3647,n3648,n3651);
and (n3648,n3649,n3650);
xor (n3649,n3547,n3548);
and (n3650,n286,n341);
and (n3651,n3652,n3653);
xor (n3652,n3649,n3650);
or (n3653,n3654,n3657);
and (n3654,n3655,n3656);
xor (n3655,n3553,n3554);
and (n3656,n328,n341);
and (n3657,n3658,n3659);
xor (n3658,n3655,n3656);
or (n3659,n3660,n3663);
and (n3660,n3661,n3662);
xor (n3661,n3559,n3560);
and (n3662,n320,n341);
and (n3663,n3664,n3665);
xor (n3664,n3661,n3662);
or (n3665,n3666,n3669);
and (n3666,n3667,n3668);
xor (n3667,n3565,n3566);
and (n3668,n429,n341);
and (n3669,n3670,n3671);
xor (n3670,n3667,n3668);
or (n3671,n3672,n3675);
and (n3672,n3673,n3674);
xor (n3673,n3571,n3572);
and (n3674,n420,n341);
and (n3675,n3676,n3677);
xor (n3676,n3673,n3674);
or (n3677,n3678,n3681);
and (n3678,n3679,n3680);
xor (n3679,n3577,n3578);
and (n3680,n461,n341);
and (n3681,n3682,n3683);
xor (n3682,n3679,n3680);
or (n3683,n3684,n3687);
and (n3684,n3685,n3686);
xor (n3685,n3583,n3584);
and (n3686,n453,n341);
and (n3687,n3688,n3689);
xor (n3688,n3685,n3686);
or (n3689,n3690,n3693);
and (n3690,n3691,n3692);
xor (n3691,n3589,n3590);
and (n3692,n560,n341);
and (n3693,n3694,n3695);
xor (n3694,n3691,n3692);
or (n3695,n3696,n3699);
and (n3696,n3697,n3698);
xor (n3697,n3595,n3596);
and (n3698,n590,n341);
and (n3699,n3700,n3701);
xor (n3700,n3697,n3698);
and (n3701,n3702,n3703);
xor (n3702,n3601,n3602);
and (n3703,n118,n341);
and (n3704,n361,n645);
or (n3705,n3706,n3709);
and (n3706,n3707,n3708);
xor (n3707,n3610,n3611);
and (n3708,n353,n645);
and (n3709,n3710,n3711);
xor (n3710,n3707,n3708);
or (n3711,n3712,n3715);
and (n3712,n3713,n3714);
xor (n3713,n3616,n3617);
and (n3714,n655,n645);
and (n3715,n3716,n3717);
xor (n3716,n3713,n3714);
or (n3717,n3718,n3721);
and (n3718,n3719,n3720);
xor (n3719,n3622,n3623);
and (n3720,n525,n645);
and (n3721,n3722,n3723);
xor (n3722,n3719,n3720);
or (n3723,n3724,n3727);
and (n3724,n3725,n3726);
xor (n3725,n3628,n3629);
and (n3726,n396,n645);
and (n3727,n3728,n3729);
xor (n3728,n3725,n3726);
or (n3729,n3730,n3733);
and (n3730,n3731,n3732);
xor (n3731,n3634,n3635);
and (n3732,n387,n645);
and (n3733,n3734,n3735);
xor (n3734,n3731,n3732);
or (n3735,n3736,n3739);
and (n3736,n3737,n3738);
xor (n3737,n3640,n3641);
and (n3738,n295,n645);
and (n3739,n3740,n3741);
xor (n3740,n3737,n3738);
or (n3741,n3742,n3745);
and (n3742,n3743,n3744);
xor (n3743,n3646,n3647);
and (n3744,n286,n645);
and (n3745,n3746,n3747);
xor (n3746,n3743,n3744);
or (n3747,n3748,n3751);
and (n3748,n3749,n3750);
xor (n3749,n3652,n3653);
and (n3750,n328,n645);
and (n3751,n3752,n3753);
xor (n3752,n3749,n3750);
or (n3753,n3754,n3757);
and (n3754,n3755,n3756);
xor (n3755,n3658,n3659);
and (n3756,n320,n645);
and (n3757,n3758,n3759);
xor (n3758,n3755,n3756);
or (n3759,n3760,n3763);
and (n3760,n3761,n3762);
xor (n3761,n3664,n3665);
and (n3762,n429,n645);
and (n3763,n3764,n3765);
xor (n3764,n3761,n3762);
or (n3765,n3766,n3769);
and (n3766,n3767,n3768);
xor (n3767,n3670,n3671);
and (n3768,n420,n645);
and (n3769,n3770,n3771);
xor (n3770,n3767,n3768);
or (n3771,n3772,n3775);
and (n3772,n3773,n3774);
xor (n3773,n3676,n3677);
and (n3774,n461,n645);
and (n3775,n3776,n3777);
xor (n3776,n3773,n3774);
or (n3777,n3778,n3781);
and (n3778,n3779,n3780);
xor (n3779,n3682,n3683);
and (n3780,n453,n645);
and (n3781,n3782,n3783);
xor (n3782,n3779,n3780);
or (n3783,n3784,n3787);
and (n3784,n3785,n3786);
xor (n3785,n3688,n3689);
and (n3786,n560,n645);
and (n3787,n3788,n3789);
xor (n3788,n3785,n3786);
or (n3789,n3790,n3793);
and (n3790,n3791,n3792);
xor (n3791,n3694,n3695);
and (n3792,n590,n645);
and (n3793,n3794,n3795);
xor (n3794,n3791,n3792);
and (n3795,n3796,n1759);
xor (n3796,n3700,n3701);
and (n3797,n353,n380);
or (n3798,n3799,n3802);
and (n3799,n3800,n3801);
xor (n3800,n3710,n3711);
and (n3801,n655,n380);
and (n3802,n3803,n3804);
xor (n3803,n3800,n3801);
or (n3804,n3805,n3808);
and (n3805,n3806,n3807);
xor (n3806,n3716,n3717);
and (n3807,n525,n380);
and (n3808,n3809,n3810);
xor (n3809,n3806,n3807);
or (n3810,n3811,n3814);
and (n3811,n3812,n3813);
xor (n3812,n3722,n3723);
and (n3813,n396,n380);
and (n3814,n3815,n3816);
xor (n3815,n3812,n3813);
or (n3816,n3817,n3820);
and (n3817,n3818,n3819);
xor (n3818,n3728,n3729);
and (n3819,n387,n380);
and (n3820,n3821,n3822);
xor (n3821,n3818,n3819);
or (n3822,n3823,n3826);
and (n3823,n3824,n3825);
xor (n3824,n3734,n3735);
and (n3825,n295,n380);
and (n3826,n3827,n3828);
xor (n3827,n3824,n3825);
or (n3828,n3829,n3832);
and (n3829,n3830,n3831);
xor (n3830,n3740,n3741);
and (n3831,n286,n380);
and (n3832,n3833,n3834);
xor (n3833,n3830,n3831);
or (n3834,n3835,n3838);
and (n3835,n3836,n3837);
xor (n3836,n3746,n3747);
and (n3837,n328,n380);
and (n3838,n3839,n3840);
xor (n3839,n3836,n3837);
or (n3840,n3841,n3844);
and (n3841,n3842,n3843);
xor (n3842,n3752,n3753);
and (n3843,n320,n380);
and (n3844,n3845,n3846);
xor (n3845,n3842,n3843);
or (n3846,n3847,n3850);
and (n3847,n3848,n3849);
xor (n3848,n3758,n3759);
and (n3849,n429,n380);
and (n3850,n3851,n3852);
xor (n3851,n3848,n3849);
or (n3852,n3853,n3856);
and (n3853,n3854,n3855);
xor (n3854,n3764,n3765);
and (n3855,n420,n380);
and (n3856,n3857,n3858);
xor (n3857,n3854,n3855);
or (n3858,n3859,n3862);
and (n3859,n3860,n3861);
xor (n3860,n3770,n3771);
and (n3861,n461,n380);
and (n3862,n3863,n3864);
xor (n3863,n3860,n3861);
or (n3864,n3865,n3868);
and (n3865,n3866,n3867);
xor (n3866,n3776,n3777);
and (n3867,n453,n380);
and (n3868,n3869,n3870);
xor (n3869,n3866,n3867);
or (n3870,n3871,n3874);
and (n3871,n3872,n3873);
xor (n3872,n3782,n3783);
and (n3873,n560,n380);
and (n3874,n3875,n3876);
xor (n3875,n3872,n3873);
or (n3876,n3877,n3880);
and (n3877,n3878,n3879);
xor (n3878,n3788,n3789);
and (n3879,n590,n380);
and (n3880,n3881,n3882);
xor (n3881,n3878,n3879);
and (n3882,n3883,n3884);
xor (n3883,n3794,n3795);
and (n3884,n118,n380);
and (n3885,n655,n373);
or (n3886,n3887,n3890);
and (n3887,n3888,n3889);
xor (n3888,n3803,n3804);
and (n3889,n525,n373);
and (n3890,n3891,n3892);
xor (n3891,n3888,n3889);
or (n3892,n3893,n3896);
and (n3893,n3894,n3895);
xor (n3894,n3809,n3810);
and (n3895,n396,n373);
and (n3896,n3897,n3898);
xor (n3897,n3894,n3895);
or (n3898,n3899,n3902);
and (n3899,n3900,n3901);
xor (n3900,n3815,n3816);
and (n3901,n387,n373);
and (n3902,n3903,n3904);
xor (n3903,n3900,n3901);
or (n3904,n3905,n3908);
and (n3905,n3906,n3907);
xor (n3906,n3821,n3822);
and (n3907,n295,n373);
and (n3908,n3909,n3910);
xor (n3909,n3906,n3907);
or (n3910,n3911,n3914);
and (n3911,n3912,n3913);
xor (n3912,n3827,n3828);
and (n3913,n286,n373);
and (n3914,n3915,n3916);
xor (n3915,n3912,n3913);
or (n3916,n3917,n3920);
and (n3917,n3918,n3919);
xor (n3918,n3833,n3834);
and (n3919,n328,n373);
and (n3920,n3921,n3922);
xor (n3921,n3918,n3919);
or (n3922,n3923,n3926);
and (n3923,n3924,n3925);
xor (n3924,n3839,n3840);
and (n3925,n320,n373);
and (n3926,n3927,n3928);
xor (n3927,n3924,n3925);
or (n3928,n3929,n3932);
and (n3929,n3930,n3931);
xor (n3930,n3845,n3846);
and (n3931,n429,n373);
and (n3932,n3933,n3934);
xor (n3933,n3930,n3931);
or (n3934,n3935,n3938);
and (n3935,n3936,n3937);
xor (n3936,n3851,n3852);
and (n3937,n420,n373);
and (n3938,n3939,n3940);
xor (n3939,n3936,n3937);
or (n3940,n3941,n3944);
and (n3941,n3942,n3943);
xor (n3942,n3857,n3858);
and (n3943,n461,n373);
and (n3944,n3945,n3946);
xor (n3945,n3942,n3943);
or (n3946,n3947,n3950);
and (n3947,n3948,n3949);
xor (n3948,n3863,n3864);
and (n3949,n453,n373);
and (n3950,n3951,n3952);
xor (n3951,n3948,n3949);
or (n3952,n3953,n3956);
and (n3953,n3954,n3955);
xor (n3954,n3869,n3870);
and (n3955,n560,n373);
and (n3956,n3957,n3958);
xor (n3957,n3954,n3955);
or (n3958,n3959,n3962);
and (n3959,n3960,n3961);
xor (n3960,n3875,n3876);
and (n3961,n590,n373);
and (n3962,n3963,n3964);
xor (n3963,n3960,n3961);
and (n3964,n3965,n1668);
xor (n3965,n3881,n3882);
and (n3966,n525,n269);
or (n3967,n3968,n3971);
and (n3968,n3969,n3970);
xor (n3969,n3891,n3892);
and (n3970,n396,n269);
and (n3971,n3972,n3973);
xor (n3972,n3969,n3970);
or (n3973,n3974,n3977);
and (n3974,n3975,n3976);
xor (n3975,n3897,n3898);
and (n3976,n387,n269);
and (n3977,n3978,n3979);
xor (n3978,n3975,n3976);
or (n3979,n3980,n3983);
and (n3980,n3981,n3982);
xor (n3981,n3903,n3904);
and (n3982,n295,n269);
and (n3983,n3984,n3985);
xor (n3984,n3981,n3982);
or (n3985,n3986,n3989);
and (n3986,n3987,n3988);
xor (n3987,n3909,n3910);
and (n3988,n286,n269);
and (n3989,n3990,n3991);
xor (n3990,n3987,n3988);
or (n3991,n3992,n3995);
and (n3992,n3993,n3994);
xor (n3993,n3915,n3916);
and (n3994,n328,n269);
and (n3995,n3996,n3997);
xor (n3996,n3993,n3994);
or (n3997,n3998,n4001);
and (n3998,n3999,n4000);
xor (n3999,n3921,n3922);
and (n4000,n320,n269);
and (n4001,n4002,n4003);
xor (n4002,n3999,n4000);
or (n4003,n4004,n4007);
and (n4004,n4005,n4006);
xor (n4005,n3927,n3928);
and (n4006,n429,n269);
and (n4007,n4008,n4009);
xor (n4008,n4005,n4006);
or (n4009,n4010,n4013);
and (n4010,n4011,n4012);
xor (n4011,n3933,n3934);
and (n4012,n420,n269);
and (n4013,n4014,n4015);
xor (n4014,n4011,n4012);
or (n4015,n4016,n4019);
and (n4016,n4017,n4018);
xor (n4017,n3939,n3940);
and (n4018,n461,n269);
and (n4019,n4020,n4021);
xor (n4020,n4017,n4018);
or (n4021,n4022,n4025);
and (n4022,n4023,n4024);
xor (n4023,n3945,n3946);
and (n4024,n453,n269);
and (n4025,n4026,n4027);
xor (n4026,n4023,n4024);
or (n4027,n4028,n4031);
and (n4028,n4029,n4030);
xor (n4029,n3951,n3952);
and (n4030,n560,n269);
and (n4031,n4032,n4033);
xor (n4032,n4029,n4030);
or (n4033,n4034,n4037);
and (n4034,n4035,n4036);
xor (n4035,n3957,n3958);
and (n4036,n590,n269);
and (n4037,n4038,n4039);
xor (n4038,n4035,n4036);
and (n4039,n4040,n4041);
xor (n4040,n3963,n3964);
and (n4041,n118,n269);
and (n4042,n396,n272);
or (n4043,n4044,n4047);
and (n4044,n4045,n4046);
xor (n4045,n3972,n3973);
and (n4046,n387,n272);
and (n4047,n4048,n4049);
xor (n4048,n4045,n4046);
or (n4049,n4050,n4053);
and (n4050,n4051,n4052);
xor (n4051,n3978,n3979);
and (n4052,n295,n272);
and (n4053,n4054,n4055);
xor (n4054,n4051,n4052);
or (n4055,n4056,n4059);
and (n4056,n4057,n4058);
xor (n4057,n3984,n3985);
and (n4058,n286,n272);
and (n4059,n4060,n4061);
xor (n4060,n4057,n4058);
or (n4061,n4062,n4065);
and (n4062,n4063,n4064);
xor (n4063,n3990,n3991);
and (n4064,n328,n272);
and (n4065,n4066,n4067);
xor (n4066,n4063,n4064);
or (n4067,n4068,n4071);
and (n4068,n4069,n4070);
xor (n4069,n3996,n3997);
and (n4070,n320,n272);
and (n4071,n4072,n4073);
xor (n4072,n4069,n4070);
or (n4073,n4074,n4077);
and (n4074,n4075,n4076);
xor (n4075,n4002,n4003);
and (n4076,n429,n272);
and (n4077,n4078,n4079);
xor (n4078,n4075,n4076);
or (n4079,n4080,n4083);
and (n4080,n4081,n4082);
xor (n4081,n4008,n4009);
and (n4082,n420,n272);
and (n4083,n4084,n4085);
xor (n4084,n4081,n4082);
or (n4085,n4086,n4089);
and (n4086,n4087,n4088);
xor (n4087,n4014,n4015);
and (n4088,n461,n272);
and (n4089,n4090,n4091);
xor (n4090,n4087,n4088);
or (n4091,n4092,n4095);
and (n4092,n4093,n4094);
xor (n4093,n4020,n4021);
and (n4094,n453,n272);
and (n4095,n4096,n4097);
xor (n4096,n4093,n4094);
or (n4097,n4098,n4101);
and (n4098,n4099,n4100);
xor (n4099,n4026,n4027);
and (n4100,n560,n272);
and (n4101,n4102,n4103);
xor (n4102,n4099,n4100);
or (n4103,n4104,n4107);
and (n4104,n4105,n4106);
xor (n4105,n4032,n4033);
and (n4106,n590,n272);
and (n4107,n4108,n4109);
xor (n4108,n4105,n4106);
and (n4109,n4110,n1867);
xor (n4110,n4038,n4039);
and (n4111,n387,n279);
or (n4112,n4113,n4116);
and (n4113,n4114,n4115);
xor (n4114,n4048,n4049);
and (n4115,n295,n279);
and (n4116,n4117,n4118);
xor (n4117,n4114,n4115);
or (n4118,n4119,n4122);
and (n4119,n4120,n4121);
xor (n4120,n4054,n4055);
and (n4121,n286,n279);
and (n4122,n4123,n4124);
xor (n4123,n4120,n4121);
or (n4124,n4125,n4128);
and (n4125,n4126,n4127);
xor (n4126,n4060,n4061);
and (n4127,n328,n279);
and (n4128,n4129,n4130);
xor (n4129,n4126,n4127);
or (n4130,n4131,n4134);
and (n4131,n4132,n4133);
xor (n4132,n4066,n4067);
and (n4133,n320,n279);
and (n4134,n4135,n4136);
xor (n4135,n4132,n4133);
or (n4136,n4137,n4140);
and (n4137,n4138,n4139);
xor (n4138,n4072,n4073);
and (n4139,n429,n279);
and (n4140,n4141,n4142);
xor (n4141,n4138,n4139);
or (n4142,n4143,n4146);
and (n4143,n4144,n4145);
xor (n4144,n4078,n4079);
and (n4145,n420,n279);
and (n4146,n4147,n4148);
xor (n4147,n4144,n4145);
or (n4148,n4149,n4152);
and (n4149,n4150,n4151);
xor (n4150,n4084,n4085);
and (n4151,n461,n279);
and (n4152,n4153,n4154);
xor (n4153,n4150,n4151);
or (n4154,n4155,n4158);
and (n4155,n4156,n4157);
xor (n4156,n4090,n4091);
and (n4157,n453,n279);
and (n4158,n4159,n4160);
xor (n4159,n4156,n4157);
or (n4160,n4161,n4164);
and (n4161,n4162,n4163);
xor (n4162,n4096,n4097);
and (n4163,n560,n279);
and (n4164,n4165,n4166);
xor (n4165,n4162,n4163);
or (n4166,n4167,n4170);
and (n4167,n4168,n4169);
xor (n4168,n4102,n4103);
and (n4169,n590,n279);
and (n4170,n4171,n4172);
xor (n4171,n4168,n4169);
and (n4172,n4173,n4174);
xor (n4173,n4108,n4109);
and (n4174,n118,n279);
and (n4175,n295,n307);
or (n4176,n4177,n4180);
and (n4177,n4178,n4179);
xor (n4178,n4117,n4118);
and (n4179,n286,n307);
and (n4180,n4181,n4182);
xor (n4181,n4178,n4179);
or (n4182,n4183,n4186);
and (n4183,n4184,n4185);
xor (n4184,n4123,n4124);
and (n4185,n328,n307);
and (n4186,n4187,n4188);
xor (n4187,n4184,n4185);
or (n4188,n4189,n4192);
and (n4189,n4190,n4191);
xor (n4190,n4129,n4130);
and (n4191,n320,n307);
and (n4192,n4193,n4194);
xor (n4193,n4190,n4191);
or (n4194,n4195,n4198);
and (n4195,n4196,n4197);
xor (n4196,n4135,n4136);
and (n4197,n429,n307);
and (n4198,n4199,n4200);
xor (n4199,n4196,n4197);
or (n4200,n4201,n4204);
and (n4201,n4202,n4203);
xor (n4202,n4141,n4142);
and (n4203,n420,n307);
and (n4204,n4205,n4206);
xor (n4205,n4202,n4203);
or (n4206,n4207,n4210);
and (n4207,n4208,n4209);
xor (n4208,n4147,n4148);
and (n4209,n461,n307);
and (n4210,n4211,n4212);
xor (n4211,n4208,n4209);
or (n4212,n4213,n4216);
and (n4213,n4214,n4215);
xor (n4214,n4153,n4154);
and (n4215,n453,n307);
and (n4216,n4217,n4218);
xor (n4217,n4214,n4215);
or (n4218,n4219,n4222);
and (n4219,n4220,n4221);
xor (n4220,n4159,n4160);
and (n4221,n560,n307);
and (n4222,n4223,n4224);
xor (n4223,n4220,n4221);
or (n4224,n4225,n4228);
and (n4225,n4226,n4227);
xor (n4226,n4165,n4166);
and (n4227,n590,n307);
and (n4228,n4229,n4230);
xor (n4229,n4226,n4227);
and (n4230,n4231,n1482);
xor (n4231,n4171,n4172);
and (n4232,n286,n313);
or (n4233,n4234,n4237);
and (n4234,n4235,n4236);
xor (n4235,n4181,n4182);
and (n4236,n328,n313);
and (n4237,n4238,n4239);
xor (n4238,n4235,n4236);
or (n4239,n4240,n4243);
and (n4240,n4241,n4242);
xor (n4241,n4187,n4188);
and (n4242,n320,n313);
and (n4243,n4244,n4245);
xor (n4244,n4241,n4242);
or (n4245,n4246,n4249);
and (n4246,n4247,n4248);
xor (n4247,n4193,n4194);
and (n4248,n429,n313);
and (n4249,n4250,n4251);
xor (n4250,n4247,n4248);
or (n4251,n4252,n4255);
and (n4252,n4253,n4254);
xor (n4253,n4199,n4200);
and (n4254,n420,n313);
and (n4255,n4256,n4257);
xor (n4256,n4253,n4254);
or (n4257,n4258,n4261);
and (n4258,n4259,n4260);
xor (n4259,n4205,n4206);
and (n4260,n461,n313);
and (n4261,n4262,n4263);
xor (n4262,n4259,n4260);
or (n4263,n4264,n4267);
and (n4264,n4265,n4266);
xor (n4265,n4211,n4212);
and (n4266,n453,n313);
and (n4267,n4268,n4269);
xor (n4268,n4265,n4266);
or (n4269,n4270,n4273);
and (n4270,n4271,n4272);
xor (n4271,n4217,n4218);
and (n4272,n560,n313);
and (n4273,n4274,n4275);
xor (n4274,n4271,n4272);
or (n4275,n4276,n4279);
and (n4276,n4277,n4278);
xor (n4277,n4223,n4224);
and (n4278,n590,n313);
and (n4279,n4280,n4281);
xor (n4280,n4277,n4278);
and (n4281,n4282,n4283);
xor (n4282,n4229,n4230);
and (n4283,n118,n313);
and (n4284,n328,n406);
or (n4285,n4286,n4289);
and (n4286,n4287,n4288);
xor (n4287,n4238,n4239);
and (n4288,n320,n406);
and (n4289,n4290,n4291);
xor (n4290,n4287,n4288);
or (n4291,n4292,n4295);
and (n4292,n4293,n4294);
xor (n4293,n4244,n4245);
and (n4294,n429,n406);
and (n4295,n4296,n4297);
xor (n4296,n4293,n4294);
or (n4297,n4298,n4301);
and (n4298,n4299,n4300);
xor (n4299,n4250,n4251);
and (n4300,n420,n406);
and (n4301,n4302,n4303);
xor (n4302,n4299,n4300);
or (n4303,n4304,n4307);
and (n4304,n4305,n4306);
xor (n4305,n4256,n4257);
and (n4306,n461,n406);
and (n4307,n4308,n4309);
xor (n4308,n4305,n4306);
or (n4309,n4310,n4313);
and (n4310,n4311,n4312);
xor (n4311,n4262,n4263);
and (n4312,n453,n406);
and (n4313,n4314,n4315);
xor (n4314,n4311,n4312);
or (n4315,n4316,n4319);
and (n4316,n4317,n4318);
xor (n4317,n4268,n4269);
and (n4318,n560,n406);
and (n4319,n4320,n4321);
xor (n4320,n4317,n4318);
or (n4321,n4322,n4325);
and (n4322,n4323,n4324);
xor (n4323,n4274,n4275);
and (n4324,n590,n406);
and (n4325,n4326,n4327);
xor (n4326,n4323,n4324);
and (n4327,n4328,n1373);
xor (n4328,n4280,n4281);
and (n4329,n320,n414);
or (n4330,n4331,n4334);
and (n4331,n4332,n4333);
xor (n4332,n4290,n4291);
and (n4333,n429,n414);
and (n4334,n4335,n4336);
xor (n4335,n4332,n4333);
or (n4336,n4337,n4340);
and (n4337,n4338,n4339);
xor (n4338,n4296,n4297);
and (n4339,n420,n414);
and (n4340,n4341,n4342);
xor (n4341,n4338,n4339);
or (n4342,n4343,n4346);
and (n4343,n4344,n4345);
xor (n4344,n4302,n4303);
and (n4345,n461,n414);
and (n4346,n4347,n4348);
xor (n4347,n4344,n4345);
or (n4348,n4349,n4352);
and (n4349,n4350,n4351);
xor (n4350,n4308,n4309);
and (n4351,n453,n414);
and (n4352,n4353,n4354);
xor (n4353,n4350,n4351);
or (n4354,n4355,n4358);
and (n4355,n4356,n4357);
xor (n4356,n4314,n4315);
and (n4357,n560,n414);
and (n4358,n4359,n4360);
xor (n4359,n4356,n4357);
or (n4360,n4361,n4364);
and (n4361,n4362,n4363);
xor (n4362,n4320,n4321);
and (n4363,n590,n414);
and (n4364,n4365,n4366);
xor (n4365,n4362,n4363);
and (n4366,n4367,n4368);
xor (n4367,n4326,n4327);
and (n4368,n118,n414);
and (n4369,n429,n439);
or (n4370,n4371,n4374);
and (n4371,n4372,n4373);
xor (n4372,n4335,n4336);
and (n4373,n420,n439);
and (n4374,n4375,n4376);
xor (n4375,n4372,n4373);
or (n4376,n4377,n4380);
and (n4377,n4378,n4379);
xor (n4378,n4341,n4342);
and (n4379,n461,n439);
and (n4380,n4381,n4382);
xor (n4381,n4378,n4379);
or (n4382,n4383,n4386);
and (n4383,n4384,n4385);
xor (n4384,n4347,n4348);
and (n4385,n453,n439);
and (n4386,n4387,n4388);
xor (n4387,n4384,n4385);
or (n4388,n4389,n4392);
and (n4389,n4390,n4391);
xor (n4390,n4353,n4354);
and (n4391,n560,n439);
and (n4392,n4393,n4394);
xor (n4393,n4390,n4391);
or (n4394,n4395,n4398);
and (n4395,n4396,n4397);
xor (n4396,n4359,n4360);
and (n4397,n590,n439);
and (n4398,n4399,n4400);
xor (n4399,n4396,n4397);
and (n4400,n4401,n728);
xor (n4401,n4365,n4366);
and (n4402,n420,n446);
or (n4403,n4404,n4407);
and (n4404,n4405,n4406);
xor (n4405,n4375,n4376);
and (n4406,n461,n446);
and (n4407,n4408,n4409);
xor (n4408,n4405,n4406);
or (n4409,n4410,n4413);
and (n4410,n4411,n4412);
xor (n4411,n4381,n4382);
and (n4412,n453,n446);
and (n4413,n4414,n4415);
xor (n4414,n4411,n4412);
or (n4415,n4416,n4419);
and (n4416,n4417,n4418);
xor (n4417,n4387,n4388);
and (n4418,n560,n446);
and (n4419,n4420,n4421);
xor (n4420,n4417,n4418);
or (n4421,n4422,n4425);
and (n4422,n4423,n4424);
xor (n4423,n4393,n4394);
and (n4424,n590,n446);
and (n4425,n4426,n4427);
xor (n4426,n4423,n4424);
and (n4427,n4428,n4429);
xor (n4428,n4399,n4400);
and (n4429,n118,n446);
and (n4430,n461,n551);
or (n4431,n4432,n4435);
and (n4432,n4433,n4434);
xor (n4433,n4408,n4409);
and (n4434,n453,n551);
and (n4435,n4436,n4437);
xor (n4436,n4433,n4434);
or (n4437,n4438,n4441);
and (n4438,n4439,n4440);
xor (n4439,n4414,n4415);
and (n4440,n560,n551);
and (n4441,n4442,n4443);
xor (n4442,n4439,n4440);
or (n4443,n4444,n4447);
and (n4444,n4445,n4446);
xor (n4445,n4420,n4421);
and (n4446,n590,n551);
and (n4447,n4448,n4449);
xor (n4448,n4445,n4446);
and (n4449,n4450,n712);
xor (n4450,n4426,n4427);
and (n4451,n453,n112);
or (n4452,n4453,n4456);
and (n4453,n4454,n4455);
xor (n4454,n4436,n4437);
and (n4455,n560,n112);
and (n4456,n4457,n4458);
xor (n4457,n4454,n4455);
or (n4458,n4459,n4462);
and (n4459,n4460,n4461);
xor (n4460,n4442,n4443);
and (n4461,n590,n112);
and (n4462,n4463,n4464);
xor (n4463,n4460,n4461);
and (n4464,n4465,n4466);
xor (n4465,n4448,n4449);
and (n4466,n118,n112);
and (n4467,n560,n16);
or (n4468,n4469,n4472);
and (n4469,n4470,n4471);
xor (n4470,n4457,n4458);
and (n4471,n590,n16);
and (n4472,n4473,n4474);
xor (n4473,n4470,n4471);
and (n4474,n4475,n1010);
xor (n4475,n4463,n4464);
and (n4476,n590,n576);
and (n4477,n4478,n4479);
xor (n4478,n4473,n4474);
and (n4479,n118,n576);
and (n4480,n118,n1075);
endmodule
