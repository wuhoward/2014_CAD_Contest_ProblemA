module top (out,n4,n5,n23,n24,n30,n34,n40,n50,n51
        ,n59,n65,n77,n78,n86,n92,n106,n112,n116,n122
        ,n137,n152,n153,n161,n167,n218,n219,n329,n335,n360
        ,n408,n416,n420,n442,n476,n1431);
output out;
input n4;
input n5;
input n23;
input n24;
input n30;
input n34;
input n40;
input n50;
input n51;
input n59;
input n65;
input n77;
input n78;
input n86;
input n92;
input n106;
input n112;
input n116;
input n122;
input n137;
input n152;
input n153;
input n161;
input n167;
input n218;
input n219;
input n329;
input n335;
input n360;
input n408;
input n416;
input n420;
input n442;
input n476;
input n1431;
wire n0;
wire n1;
wire n2;
wire n3;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n25;
wire n26;
wire n27;
wire n28;
wire n29;
wire n31;
wire n32;
wire n33;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n113;
wire n114;
wire n115;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n417;
wire n418;
wire n419;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
xor (out,n0,n1433);
or (n0,n1,n1430);
and (n1,n2,n6);
nor (n2,n3,n5);
not (n3,n4);
nand (n6,n7,n1429);
or (n7,n8,n288);
not (n8,n9);
nand (n9,n10,n287);
or (n10,n11,n247);
or (n11,n12,n246);
and (n12,n13,n205);
xor (n13,n14,n127);
or (n14,n15,n126);
and (n15,n16,n68);
xor (n16,n17,n43);
nand (n17,n18,n37);
or (n18,n19,n32);
nand (n19,n20,n27);
nor (n20,n21,n25);
and (n21,n22,n24);
not (n22,n23);
and (n25,n23,n26);
not (n26,n24);
nand (n27,n28,n31);
nand (n28,n29,n24);
not (n29,n30);
nand (n31,n30,n26);
nor (n32,n33,n35);
and (n33,n29,n34);
and (n35,n30,n36);
not (n36,n34);
or (n37,n20,n38);
nor (n38,n39,n41);
and (n39,n29,n40);
and (n41,n30,n42);
not (n42,n40);
not (n43,n44);
nand (n44,n45,n62);
or (n45,n46,n57);
nand (n46,n47,n54);
nor (n47,n48,n52);
and (n48,n49,n51);
not (n49,n50);
and (n52,n50,n53);
not (n53,n51);
nand (n54,n55,n56);
or (n55,n22,n51);
nand (n56,n22,n51);
nor (n57,n58,n60);
and (n58,n22,n59);
and (n60,n23,n61);
not (n61,n59);
or (n62,n47,n63);
nor (n63,n64,n66);
and (n64,n22,n65);
and (n66,n23,n67);
not (n67,n65);
or (n68,n69,n125);
and (n69,n70,n101);
xor (n70,n71,n95);
nand (n71,n72,n89);
or (n72,n73,n84);
nand (n73,n74,n81);
or (n74,n75,n79);
and (n75,n76,n78);
not (n76,n77);
and (n79,n77,n80);
not (n80,n78);
nor (n81,n82,n83);
and (n82,n30,n76);
and (n83,n29,n77);
nor (n84,n85,n87);
and (n85,n80,n86);
and (n87,n78,n88);
not (n88,n86);
or (n89,n90,n81);
nor (n90,n91,n93);
and (n91,n92,n80);
and (n93,n78,n94);
not (n94,n92);
nand (n95,n96,n100);
or (n96,n46,n97);
nor (n97,n98,n99);
and (n98,n22,n40);
and (n99,n23,n42);
or (n100,n47,n57);
nand (n101,n102,n119);
or (n102,n103,n114);
nand (n103,n104,n109);
nor (n104,n105,n107);
and (n105,n80,n106);
and (n107,n78,n108);
not (n108,n106);
nand (n109,n110,n113);
or (n110,n111,n106);
not (n111,n112);
nand (n113,n111,n106);
nor (n114,n115,n117);
and (n115,n116,n111);
and (n117,n112,n118);
not (n118,n116);
or (n119,n120,n104);
nor (n120,n121,n123);
and (n121,n122,n111);
and (n123,n112,n124);
not (n124,n122);
and (n125,n71,n95);
and (n126,n17,n43);
xor (n127,n128,n191);
xor (n128,n129,n171);
or (n129,n130,n170);
and (n130,n131,n146);
xor (n131,n132,n140);
nand (n132,n133,n134);
or (n133,n73,n90);
or (n134,n135,n81);
nor (n135,n136,n138);
and (n136,n80,n137);
and (n138,n78,n139);
not (n139,n137);
nand (n140,n141,n142);
or (n141,n103,n120);
or (n142,n104,n143);
nor (n143,n144,n145);
and (n144,n111,n86);
and (n145,n112,n88);
nand (n146,n147,n164);
or (n147,n148,n159);
nand (n148,n149,n156);
nor (n149,n150,n154);
and (n150,n151,n153);
not (n151,n152);
and (n154,n152,n155);
not (n155,n153);
nand (n156,n157,n158);
or (n157,n153,n49);
nand (n158,n49,n153);
nor (n159,n160,n162);
and (n160,n49,n161);
and (n162,n50,n163);
not (n163,n161);
or (n164,n149,n165);
nor (n165,n166,n168);
and (n166,n49,n167);
and (n168,n50,n169);
not (n169,n167);
and (n170,n132,n140);
xor (n171,n172,n184);
xor (n172,n173,n178);
nand (n173,n174,n177);
or (n174,n175,n176);
not (n175,n149);
not (n176,n148);
not (n177,n165);
nand (n178,n179,n180);
or (n179,n46,n63);
or (n180,n47,n181);
nor (n181,n182,n183);
and (n182,n22,n161);
and (n183,n23,n163);
nand (n184,n185,n190);
or (n185,n81,n186);
not (n186,n187);
nand (n187,n188,n189);
or (n188,n78,n36);
or (n189,n80,n34);
or (n190,n73,n135);
xor (n191,n192,n44);
xor (n192,n193,n199);
nand (n193,n194,n195);
or (n194,n103,n143);
or (n195,n196,n104);
nor (n196,n197,n198);
and (n197,n111,n92);
and (n198,n112,n94);
nand (n199,n200,n201);
or (n200,n19,n38);
or (n201,n20,n202);
nor (n202,n203,n204);
and (n203,n29,n59);
and (n204,n30,n61);
or (n205,n206,n245);
and (n206,n207,n244);
xor (n207,n208,n243);
or (n208,n209,n242);
and (n209,n210,n236);
xor (n210,n211,n230);
nand (n211,n212,n226);
or (n212,n213,n225);
not (n213,n214);
nand (n214,n215,n222);
nor (n215,n216,n220);
and (n216,n217,n219);
not (n217,n218);
and (n220,n218,n221);
not (n221,n219);
nand (n222,n223,n224);
or (n223,n218,n151);
nand (n224,n151,n218);
not (n225,n215);
not (n226,n227);
nor (n227,n228,n229);
and (n228,n151,n167);
and (n229,n152,n169);
nand (n230,n231,n235);
or (n231,n148,n232);
nor (n232,n233,n234);
and (n233,n49,n65);
and (n234,n50,n67);
or (n235,n149,n159);
nand (n236,n237,n241);
or (n237,n19,n238);
nor (n238,n239,n240);
and (n239,n29,n137);
and (n240,n30,n139);
or (n241,n20,n32);
and (n242,n211,n230);
xor (n243,n131,n146);
xor (n244,n16,n68);
and (n245,n208,n243);
and (n246,n14,n127);
xor (n247,n248,n284);
xor (n248,n249,n252);
or (n249,n250,n251);
and (n250,n192,n44);
and (n251,n193,n199);
xor (n252,n253,n264);
xor (n253,n254,n261);
not (n254,n255);
nand (n255,n256,n257);
or (n256,n46,n181);
or (n257,n47,n258);
nor (n258,n259,n260);
and (n259,n22,n167);
and (n260,n23,n169);
or (n261,n262,n263);
and (n262,n172,n184);
and (n263,n173,n178);
xor (n264,n265,n278);
xor (n265,n266,n272);
nand (n266,n267,n268);
or (n267,n103,n196);
or (n268,n104,n269);
nor (n269,n270,n271);
and (n270,n111,n137);
and (n271,n112,n139);
nand (n272,n273,n274);
or (n273,n19,n202);
or (n274,n20,n275);
nor (n275,n276,n277);
and (n276,n29,n65);
and (n277,n30,n67);
nand (n278,n279,n280);
or (n279,n186,n73);
or (n280,n281,n81);
nor (n281,n282,n283);
and (n282,n80,n40);
and (n283,n78,n42);
or (n284,n285,n286);
and (n285,n128,n191);
and (n286,n129,n171);
nand (n287,n11,n247);
not (n288,n289);
nand (n289,n290,n1428);
or (n290,n291,n1423);
nor (n291,n292,n1419);
and (n292,n293,n1381);
nand (n293,n294,n1370);
or (n294,n295,n869);
nand (n295,n296,n748,n864);
nor (n296,n297,n684);
nor (n297,n298,n592);
xor (n298,n299,n544);
xor (n299,n300,n390);
xor (n300,n301,n367);
xor (n301,n302,n339);
or (n302,n303,n338);
and (n303,n304,n325);
xor (n304,n305,n316);
nand (n305,n306,n311);
or (n306,n215,n307);
not (n307,n308);
nand (n308,n309,n310);
or (n309,n152,n61);
or (n310,n151,n59);
nand (n311,n312,n213);
not (n312,n313);
nor (n313,n314,n315);
and (n314,n40,n151);
and (n315,n42,n152);
nand (n316,n317,n321);
or (n317,n19,n318);
nor (n318,n319,n320);
and (n319,n116,n29);
and (n320,n30,n118);
or (n321,n322,n20);
nor (n322,n323,n324);
and (n323,n122,n29);
and (n324,n30,n124);
nand (n325,n326,n332);
or (n326,n73,n327);
nor (n327,n328,n330);
and (n328,n329,n80);
and (n330,n78,n331);
not (n331,n329);
or (n332,n333,n81);
nor (n333,n334,n336);
and (n334,n335,n80);
and (n336,n78,n337);
not (n337,n335);
and (n338,n305,n316);
xor (n339,n340,n356);
xor (n340,n341,n350);
nand (n341,n342,n346);
or (n342,n148,n343);
nor (n343,n344,n345);
and (n344,n49,n34);
and (n345,n50,n36);
or (n346,n149,n347);
nor (n347,n348,n349);
and (n348,n49,n40);
and (n349,n50,n42);
nand (n350,n351,n352);
or (n351,n73,n333);
or (n352,n353,n81);
nor (n353,n354,n355);
and (n354,n116,n80);
and (n355,n78,n118);
nand (n356,n357,n363);
or (n357,n103,n358);
nor (n358,n359,n361);
and (n359,n360,n111);
and (n361,n112,n362);
not (n362,n360);
or (n363,n364,n104);
nor (n364,n365,n366);
and (n365,n329,n111);
and (n366,n112,n331);
xor (n367,n368,n384);
xor (n368,n369,n375);
nand (n369,n370,n371);
or (n370,n307,n214);
or (n371,n215,n372);
nor (n372,n373,n374);
and (n373,n151,n65);
and (n374,n152,n67);
nand (n375,n376,n380);
or (n376,n46,n377);
nor (n377,n378,n379);
and (n378,n22,n92);
and (n379,n23,n94);
or (n380,n47,n381);
nor (n381,n382,n383);
and (n382,n22,n137);
and (n383,n23,n139);
nand (n384,n385,n386);
or (n385,n19,n322);
or (n386,n20,n387);
nor (n387,n388,n389);
and (n388,n86,n29);
and (n389,n30,n88);
or (n390,n391,n543);
and (n391,n392,n515);
xor (n392,n393,n456);
or (n393,n394,n455);
and (n394,n395,n425);
xor (n395,n396,n403);
nand (n396,n397,n402);
or (n397,n73,n398);
not (n398,n399);
nand (n399,n400,n401);
or (n400,n362,n78);
or (n401,n80,n360);
or (n402,n327,n81);
xor (n403,n404,n411);
nor (n404,n405,n111);
nor (n405,n406,n409);
and (n406,n407,n80);
nand (n407,n408,n106);
and (n409,n410,n108);
not (n410,n408);
nand (n411,n412,n421);
or (n412,n413,n418);
nor (n413,n414,n417);
and (n414,n161,n415);
not (n415,n416);
and (n417,n163,n416);
nand (n418,n419,n416);
not (n419,n420);
or (n421,n422,n419);
nor (n422,n423,n424);
and (n423,n415,n167);
and (n424,n416,n169);
or (n425,n426,n454);
and (n426,n427,n435);
xor (n427,n428,n429);
nor (n428,n104,n410);
nand (n429,n430,n434);
or (n430,n431,n418);
nor (n431,n432,n433);
and (n432,n416,n67);
nor (n433,n416,n67);
or (n434,n413,n419);
nand (n435,n436,n450);
or (n436,n437,n447);
nand (n437,n438,n444);
not (n438,n439);
nand (n439,n440,n443);
or (n440,n441,n416);
not (n441,n442);
nand (n443,n441,n416);
nand (n444,n445,n446);
or (n445,n441,n219);
nand (n446,n219,n441);
nor (n447,n448,n449);
and (n448,n221,n40);
and (n449,n219,n42);
or (n450,n438,n451);
nor (n451,n452,n453);
and (n452,n221,n59);
and (n453,n219,n61);
and (n454,n428,n429);
and (n455,n396,n403);
xor (n456,n457,n489);
xor (n457,n458,n459);
and (n458,n404,n411);
or (n459,n460,n488);
and (n460,n461,n479);
xor (n461,n462,n468);
nand (n462,n463,n464);
or (n463,n437,n451);
or (n464,n438,n465);
nor (n465,n466,n467);
and (n466,n221,n65);
and (n467,n219,n67);
nand (n468,n469,n473);
or (n469,n103,n470);
nor (n470,n471,n472);
and (n471,n410,n112);
and (n472,n408,n111);
or (n473,n474,n104);
nor (n474,n475,n477);
and (n475,n476,n111);
and (n477,n478,n112);
not (n478,n476);
nand (n479,n480,n484);
or (n480,n148,n481);
nor (n481,n482,n483);
and (n482,n49,n92);
and (n483,n50,n94);
or (n484,n149,n485);
nor (n485,n486,n487);
and (n486,n49,n137);
and (n487,n50,n139);
and (n488,n462,n468);
or (n489,n490,n514);
and (n490,n491,n508);
xor (n491,n492,n502);
nand (n492,n493,n498);
or (n493,n47,n494);
not (n494,n495);
nor (n495,n496,n497);
and (n496,n88,n22);
and (n497,n86,n23);
or (n498,n46,n499);
nor (n499,n500,n501);
and (n500,n22,n122);
and (n501,n23,n124);
nand (n502,n503,n507);
or (n503,n214,n504);
nor (n504,n505,n506);
and (n505,n151,n34);
and (n506,n152,n36);
or (n507,n215,n313);
nand (n508,n509,n513);
or (n509,n19,n510);
nor (n510,n511,n512);
and (n511,n29,n335);
and (n512,n30,n337);
or (n513,n20,n318);
and (n514,n492,n502);
or (n515,n516,n542);
and (n516,n517,n541);
xor (n517,n518,n540);
or (n518,n519,n539);
and (n519,n520,n533);
xor (n520,n521,n527);
nand (n521,n522,n526);
or (n522,n148,n523);
nor (n523,n524,n525);
and (n524,n86,n49);
and (n525,n50,n88);
or (n526,n481,n149);
nand (n527,n528,n532);
or (n528,n46,n529);
nor (n529,n530,n531);
and (n530,n22,n116);
and (n531,n23,n118);
or (n532,n499,n47);
nand (n533,n534,n538);
or (n534,n214,n535);
nor (n535,n536,n537);
and (n536,n151,n137);
and (n537,n152,n139);
or (n538,n215,n504);
and (n539,n521,n527);
xor (n540,n491,n508);
xor (n541,n461,n479);
and (n542,n518,n540);
and (n543,n393,n456);
xor (n544,n545,n584);
xor (n545,n546,n549);
or (n546,n547,n548);
and (n547,n457,n489);
and (n548,n458,n459);
xor (n549,n550,n571);
xor (n550,n551,n561);
not (n551,n552);
nand (n552,n553,n557);
or (n553,n437,n554);
nor (n554,n555,n556);
and (n555,n221,n161);
and (n556,n219,n163);
or (n557,n438,n558);
nor (n558,n559,n560);
and (n559,n221,n167);
and (n560,n219,n169);
nand (n561,n562,n567);
not (n562,n563);
nand (n563,n564,n566);
or (n564,n565,n420);
not (n565,n418);
not (n566,n422);
not (n567,n568);
nand (n568,n569,n570);
or (n569,n437,n465);
or (n570,n438,n554);
or (n571,n572,n583);
and (n572,n573,n580);
xor (n573,n574,n577);
nand (n574,n575,n576);
or (n575,n103,n474);
or (n576,n358,n104);
nand (n577,n578,n579);
or (n578,n148,n485);
or (n579,n149,n343);
nand (n580,n581,n582);
or (n581,n46,n494);
or (n582,n377,n47);
and (n583,n574,n577);
or (n584,n585,n591);
and (n585,n586,n590);
xor (n586,n587,n588);
xor (n587,n304,n325);
nand (n588,n589,n561);
or (n589,n562,n567);
xor (n590,n573,n580);
and (n591,n587,n588);
or (n592,n593,n683);
and (n593,n594,n682);
xor (n594,n595,n596);
xor (n595,n586,n590);
or (n596,n597,n681);
and (n597,n598,n630);
xor (n598,n599,n629);
or (n599,n600,n628);
and (n600,n601,n616);
xor (n601,n602,n608);
nand (n602,n603,n607);
or (n603,n19,n604);
nor (n604,n605,n606);
and (n605,n329,n29);
and (n606,n30,n331);
or (n607,n20,n510);
nand (n608,n609,n610);
or (n609,n81,n398);
nand (n610,n611,n615);
not (n611,n612);
nor (n612,n613,n614);
and (n613,n80,n476);
and (n614,n478,n78);
not (n615,n73);
and (n616,n617,n622);
nor (n617,n618,n80);
nor (n618,n619,n621);
and (n619,n620,n29);
nand (n620,n77,n408);
and (n621,n410,n76);
nand (n622,n623,n627);
or (n623,n624,n418);
nor (n624,n625,n626);
and (n625,n415,n59);
and (n626,n416,n61);
or (n627,n431,n419);
and (n628,n602,n608);
xor (n629,n395,n425);
or (n630,n631,n680);
and (n631,n632,n679);
xor (n632,n633,n657);
or (n633,n634,n656);
and (n634,n635,n649);
xor (n635,n636,n642);
nand (n636,n637,n641);
or (n637,n437,n638);
nor (n638,n639,n640);
and (n639,n34,n221);
and (n640,n36,n219);
or (n641,n438,n447);
nand (n642,n643,n648);
or (n643,n644,n148);
not (n644,n645);
nand (n645,n646,n647);
or (n646,n50,n124);
or (n647,n49,n122);
or (n648,n523,n149);
nand (n649,n650,n655);
or (n650,n46,n651);
not (n651,n652);
nor (n652,n653,n654);
and (n653,n337,n22);
and (n654,n335,n23);
or (n655,n529,n47);
and (n656,n636,n642);
or (n657,n658,n678);
and (n658,n659,n672);
xor (n659,n660,n666);
nand (n660,n661,n665);
or (n661,n214,n662);
nor (n662,n663,n664);
and (n663,n151,n92);
and (n664,n152,n94);
or (n665,n215,n535);
nand (n666,n667,n671);
or (n667,n19,n668);
nor (n668,n669,n670);
and (n669,n360,n29);
and (n670,n30,n362);
or (n671,n604,n20);
nand (n672,n673,n677);
or (n673,n73,n674);
nor (n674,n675,n676);
and (n675,n410,n78);
and (n676,n408,n80);
or (n677,n612,n81);
and (n678,n660,n666);
xor (n679,n427,n435);
and (n680,n633,n657);
and (n681,n599,n629);
xor (n682,n392,n515);
and (n683,n595,n596);
nor (n684,n685,n747);
or (n685,n686,n746);
and (n686,n687,n745);
xor (n687,n688,n689);
xor (n688,n517,n541);
or (n689,n690,n744);
and (n690,n691,n694);
xor (n691,n692,n693);
xor (n692,n520,n533);
xor (n693,n601,n616);
or (n694,n695,n743);
and (n695,n696,n719);
xor (n696,n697,n698);
xor (n697,n617,n622);
or (n698,n699,n718);
and (n699,n700,n711);
xor (n700,n701,n703);
and (n701,n702,n408);
not (n702,n81);
nand (n703,n704,n709);
or (n704,n705,n437);
not (n705,n706);
nand (n706,n707,n708);
or (n707,n219,n139);
or (n708,n221,n137);
nand (n709,n710,n439);
not (n710,n638);
nand (n711,n712,n717);
or (n712,n148,n713);
not (n713,n714);
nand (n714,n715,n716);
or (n715,n50,n118);
or (n716,n49,n116);
or (n717,n149,n644);
and (n718,n701,n703);
or (n719,n720,n742);
and (n720,n721,n736);
xor (n721,n722,n730);
nand (n722,n723,n728);
or (n723,n724,n46);
not (n724,n725);
nand (n725,n726,n727);
or (n726,n23,n331);
or (n727,n22,n329);
nand (n728,n652,n729);
not (n729,n47);
nand (n730,n731,n732);
or (n731,n419,n624);
or (n732,n733,n418);
nor (n733,n734,n735);
and (n734,n415,n40);
and (n735,n416,n42);
nand (n736,n737,n741);
or (n737,n738,n19);
nor (n738,n739,n740);
and (n739,n476,n29);
and (n740,n30,n478);
or (n741,n668,n20);
and (n742,n722,n730);
and (n743,n697,n698);
and (n744,n692,n693);
xor (n745,n598,n630);
and (n746,n688,n689);
xor (n747,n594,n682);
or (n748,n749,n819);
or (n749,n750,n818);
and (n750,n751,n815);
xor (n751,n752,n796);
xor (n752,n753,n777);
xor (n753,n754,n757);
or (n754,n755,n756);
and (n755,n340,n356);
and (n756,n341,n350);
xor (n757,n758,n771);
xor (n758,n759,n765);
nand (n759,n760,n761);
or (n760,n19,n387);
or (n761,n762,n20);
nor (n762,n763,n764);
and (n763,n92,n29);
and (n764,n30,n94);
nand (n765,n766,n767);
or (n766,n148,n347);
or (n767,n149,n768);
nor (n768,n769,n770);
and (n769,n49,n59);
and (n770,n50,n61);
nand (n771,n772,n773);
or (n772,n73,n353);
or (n773,n774,n81);
nor (n774,n775,n776);
and (n775,n122,n80);
and (n776,n78,n124);
xor (n777,n778,n789);
xor (n778,n779,n783);
nand (n779,n780,n782);
or (n780,n439,n781);
not (n781,n437);
not (n782,n558);
nand (n783,n784,n785);
or (n784,n214,n372);
or (n785,n215,n786);
nor (n786,n787,n788);
and (n787,n151,n161);
and (n788,n152,n163);
nand (n789,n790,n795);
or (n790,n791,n47);
not (n791,n792);
nand (n792,n793,n794);
or (n793,n23,n36);
or (n794,n22,n34);
or (n795,n46,n381);
xor (n796,n797,n812);
xor (n797,n798,n809);
xor (n798,n799,n806);
xor (n799,n800,n552);
nand (n800,n801,n802);
or (n801,n103,n364);
or (n802,n803,n104);
nor (n803,n804,n805);
and (n804,n111,n335);
and (n805,n112,n337);
or (n806,n807,n808);
and (n807,n368,n384);
and (n808,n369,n375);
or (n809,n810,n811);
and (n810,n550,n571);
and (n811,n551,n561);
or (n812,n813,n814);
and (n813,n301,n367);
and (n814,n302,n339);
or (n815,n816,n817);
and (n816,n545,n584);
and (n817,n546,n549);
and (n818,n752,n796);
xor (n819,n820,n861);
xor (n820,n821,n840);
xor (n821,n822,n829);
xor (n822,n823,n826);
or (n823,n824,n825);
and (n824,n758,n771);
and (n825,n759,n765);
or (n826,n827,n828);
and (n827,n778,n789);
and (n828,n779,n783);
xor (n829,n830,n837);
xor (n830,n831,n834);
nand (n831,n832,n833);
or (n832,n19,n762);
or (n833,n20,n238);
nand (n834,n835,n836);
or (n835,n73,n774);
or (n836,n84,n81);
nand (n837,n838,n839);
or (n838,n214,n786);
or (n839,n215,n227);
xor (n840,n841,n858);
xor (n841,n842,n855);
xor (n842,n843,n851);
xor (n843,n844,n847);
nand (n844,n845,n846);
or (n845,n103,n803);
or (n846,n114,n104);
nand (n847,n848,n849);
or (n848,n791,n46);
nand (n849,n850,n729);
not (n850,n97);
not (n851,n852);
nand (n852,n853,n854);
or (n853,n148,n768);
or (n854,n149,n232);
or (n855,n856,n857);
and (n856,n799,n806);
and (n857,n800,n552);
or (n858,n859,n860);
and (n859,n753,n777);
and (n860,n754,n757);
or (n861,n862,n863);
and (n862,n797,n812);
and (n863,n798,n809);
or (n864,n865,n866);
xor (n865,n751,n815);
or (n866,n867,n868);
and (n867,n299,n544);
and (n868,n300,n390);
not (n869,n870);
or (n870,n871,n1369);
and (n871,n872,n935);
xor (n872,n873,n934);
or (n873,n874,n933);
and (n874,n875,n878);
xor (n875,n876,n877);
xor (n876,n632,n679);
xor (n877,n691,n694);
or (n878,n879,n932);
and (n879,n880,n883);
xor (n880,n881,n882);
xor (n881,n659,n672);
xor (n882,n635,n649);
or (n883,n884,n931);
and (n884,n885,n906);
xor (n885,n886,n892);
nand (n886,n887,n891);
or (n887,n214,n888);
nor (n888,n889,n890);
and (n889,n151,n86);
and (n890,n152,n88);
or (n891,n215,n662);
nor (n892,n893,n900);
not (n893,n894);
nand (n894,n895,n899);
or (n895,n896,n437);
nor (n896,n897,n898);
and (n897,n92,n221);
and (n898,n94,n219);
nand (n899,n439,n706);
nand (n900,n901,n30);
nand (n901,n902,n903);
or (n902,n408,n24);
nand (n903,n904,n22);
not (n904,n905);
and (n905,n408,n24);
or (n906,n907,n930);
and (n907,n908,n923);
xor (n908,n909,n916);
nand (n909,n910,n911);
or (n910,n149,n713);
nand (n911,n912,n176);
not (n912,n913);
nor (n913,n914,n915);
and (n914,n337,n50);
and (n915,n335,n49);
nand (n916,n917,n922);
or (n917,n918,n46);
not (n918,n919);
nor (n919,n920,n921);
and (n920,n22,n362);
and (n921,n23,n360);
nand (n922,n729,n725);
nand (n923,n924,n929);
or (n924,n925,n418);
not (n925,n926);
or (n926,n927,n928);
and (n927,n36,n416);
and (n928,n34,n415);
or (n929,n733,n419);
and (n930,n909,n916);
and (n931,n886,n892);
and (n932,n881,n882);
and (n933,n876,n877);
xor (n934,n687,n745);
or (n935,n936,n1368);
and (n936,n937,n971);
xor (n937,n938,n970);
or (n938,n939,n969);
and (n939,n940,n968);
xor (n940,n941,n942);
xor (n941,n696,n719);
or (n942,n943,n967);
and (n943,n944,n947);
xor (n944,n945,n946);
xor (n945,n721,n736);
xor (n946,n700,n711);
or (n947,n948,n966);
and (n948,n949,n962);
xor (n949,n950,n956);
nand (n950,n951,n955);
or (n951,n19,n952);
nor (n952,n953,n954);
and (n953,n410,n30);
and (n954,n408,n29);
or (n955,n738,n20);
nand (n956,n957,n961);
or (n957,n214,n958);
nor (n958,n959,n960);
and (n959,n151,n122);
and (n960,n152,n124);
or (n961,n215,n888);
nand (n962,n963,n965);
or (n963,n964,n893);
not (n964,n900);
or (n965,n894,n900);
and (n966,n950,n956);
and (n967,n945,n946);
xor (n968,n880,n883);
and (n969,n941,n942);
xor (n970,n875,n878);
nand (n971,n972,n1364);
or (n972,n973,n1342);
nor (n973,n974,n1341);
and (n974,n975,n1322);
or (n975,n976,n1321);
and (n976,n977,n1119);
xor (n977,n978,n1088);
or (n978,n979,n1087);
and (n979,n980,n1050);
xor (n980,n981,n1011);
xor (n981,n982,n1001);
xor (n982,n983,n992);
nand (n983,n984,n988);
or (n984,n148,n985);
nor (n985,n986,n987);
and (n986,n360,n49);
and (n987,n362,n50);
or (n988,n989,n149);
nor (n989,n990,n991);
and (n990,n49,n329);
and (n991,n50,n331);
nand (n992,n993,n997);
or (n993,n46,n994);
nor (n994,n995,n996);
and (n995,n410,n23);
and (n996,n408,n22);
or (n997,n998,n47);
nor (n998,n999,n1000);
and (n999,n476,n22);
and (n1000,n478,n23);
nand (n1001,n1002,n1007);
or (n1002,n418,n1003);
not (n1003,n1004);
nor (n1004,n1005,n1006);
and (n1005,n92,n416);
and (n1006,n94,n415);
or (n1007,n1008,n419);
nor (n1008,n1009,n1010);
and (n1009,n137,n415);
and (n1010,n139,n416);
or (n1011,n1012,n1049);
and (n1012,n1013,n1032);
xor (n1013,n1014,n1023);
nand (n1014,n1015,n1019);
or (n1015,n437,n1016);
nor (n1016,n1017,n1018);
and (n1017,n221,n116);
and (n1018,n219,n118);
or (n1019,n438,n1020);
nor (n1020,n1021,n1022);
and (n1021,n124,n219);
and (n1022,n122,n221);
nand (n1023,n1024,n1028);
or (n1024,n214,n1025);
nor (n1025,n1026,n1027);
and (n1026,n329,n151);
and (n1027,n152,n331);
or (n1028,n215,n1029);
nor (n1029,n1030,n1031);
and (n1030,n151,n335);
and (n1031,n152,n337);
and (n1032,n1033,n1039);
nor (n1033,n1034,n49);
nor (n1034,n1035,n1038);
and (n1035,n1036,n151);
not (n1036,n1037);
and (n1037,n408,n153);
and (n1038,n410,n155);
nand (n1039,n1040,n1045);
or (n1040,n1041,n418);
not (n1041,n1042);
nor (n1042,n1043,n1044);
and (n1043,n124,n415);
and (n1044,n122,n416);
or (n1045,n1046,n419);
nor (n1046,n1047,n1048);
and (n1047,n86,n415);
and (n1048,n88,n416);
and (n1049,n1014,n1023);
xor (n1050,n1051,n1072);
xor (n1051,n1052,n1058);
nand (n1052,n1053,n1054);
or (n1053,n214,n1029);
or (n1054,n215,n1055);
nor (n1055,n1056,n1057);
and (n1056,n151,n116);
and (n1057,n152,n118);
xor (n1058,n1059,n1064);
nor (n1059,n1060,n22);
nor (n1060,n1061,n1063);
and (n1061,n1062,n49);
nand (n1062,n408,n51);
and (n1063,n410,n53);
nand (n1064,n1065,n1070);
or (n1065,n438,n1066);
not (n1066,n1067);
nand (n1067,n1068,n1069);
or (n1068,n219,n88);
or (n1069,n221,n86);
nand (n1070,n1071,n781);
not (n1071,n1020);
or (n1072,n1073,n1086);
and (n1073,n1074,n1079);
xor (n1074,n1075,n1076);
nor (n1075,n47,n410);
nand (n1076,n1077,n1078);
or (n1077,n419,n1003);
or (n1078,n1046,n418);
nand (n1079,n1080,n1081);
or (n1080,n149,n985);
nand (n1081,n1082,n176);
not (n1082,n1083);
or (n1083,n1084,n1085);
and (n1084,n478,n49);
and (n1085,n476,n50);
and (n1086,n1075,n1076);
and (n1087,n981,n1011);
xor (n1088,n1089,n1104);
xor (n1089,n1090,n1101);
xor (n1090,n1091,n1098);
xor (n1091,n1092,n1095);
nand (n1092,n1093,n1094);
or (n1093,n47,n918);
or (n1094,n46,n998);
nand (n1095,n1096,n1097);
or (n1096,n1008,n418);
nand (n1097,n926,n420);
nand (n1098,n1099,n1100);
or (n1099,n214,n1055);
or (n1100,n215,n958);
or (n1101,n1102,n1103);
and (n1102,n1051,n1072);
and (n1103,n1052,n1058);
xor (n1104,n1105,n1110);
xor (n1105,n1106,n1107);
and (n1106,n1059,n1064);
or (n1107,n1108,n1109);
and (n1108,n982,n1001);
and (n1109,n983,n992);
xor (n1110,n1111,n1116);
xor (n1111,n1112,n1113);
nor (n1112,n20,n410);
nand (n1113,n1114,n1115);
or (n1114,n1066,n437);
or (n1115,n438,n896);
nand (n1116,n1117,n1118);
or (n1117,n148,n989);
or (n1118,n149,n913);
nand (n1119,n1120,n1317,n1320);
nand (n1120,n1121,n1175,n1310);
not (n1121,n1122);
nor (n1122,n1123,n1150);
xor (n1123,n1124,n1149);
xor (n1124,n1125,n1148);
or (n1125,n1126,n1147);
and (n1126,n1127,n1141);
xor (n1127,n1128,n1134);
nand (n1128,n1129,n1133);
or (n1129,n148,n1130);
nor (n1130,n1131,n1132);
and (n1131,n410,n50);
and (n1132,n408,n49);
or (n1133,n1083,n149);
nand (n1134,n1135,n1140);
or (n1135,n1136,n437);
not (n1136,n1137);
nor (n1137,n1138,n1139);
and (n1138,n335,n219);
and (n1139,n337,n221);
or (n1140,n438,n1016);
nand (n1141,n1142,n1146);
or (n1142,n214,n1143);
nor (n1143,n1144,n1145);
and (n1144,n360,n151);
and (n1145,n152,n362);
or (n1146,n215,n1025);
and (n1147,n1128,n1134);
xor (n1148,n1074,n1079);
xor (n1149,n1013,n1032);
or (n1150,n1151,n1174);
and (n1151,n1152,n1173);
xor (n1152,n1153,n1154);
xor (n1153,n1033,n1039);
or (n1154,n1155,n1172);
and (n1155,n1156,n1165);
xor (n1156,n1157,n1158);
and (n1157,n175,n408);
nand (n1158,n1159,n1164);
or (n1159,n418,n1160);
not (n1160,n1161);
nor (n1161,n1162,n1163);
and (n1162,n118,n415);
and (n1163,n116,n416);
nand (n1164,n1042,n420);
nand (n1165,n1166,n1171);
or (n1166,n1167,n437);
not (n1167,n1168);
nor (n1168,n1169,n1170);
and (n1169,n331,n221);
and (n1170,n329,n219);
nand (n1171,n1137,n439);
and (n1172,n1157,n1158);
xor (n1173,n1127,n1141);
and (n1174,n1153,n1154);
or (n1175,n1176,n1309);
and (n1176,n1177,n1203);
xor (n1177,n1178,n1202);
or (n1178,n1179,n1201);
and (n1179,n1180,n1200);
xor (n1180,n1181,n1187);
nand (n1181,n1182,n1186);
or (n1182,n214,n1183);
nor (n1183,n1184,n1185);
and (n1184,n151,n476);
and (n1185,n152,n478);
or (n1186,n1143,n215);
and (n1187,n1188,n1194);
and (n1188,n1189,n152);
nand (n1189,n1190,n1191);
or (n1190,n408,n218);
nand (n1191,n1192,n221);
not (n1192,n1193);
and (n1193,n408,n218);
nand (n1194,n1195,n1196);
or (n1195,n419,n1160);
or (n1196,n1197,n418);
nor (n1197,n1198,n1199);
and (n1198,n415,n335);
and (n1199,n416,n337);
xor (n1200,n1156,n1165);
and (n1201,n1181,n1187);
xor (n1202,n1152,n1173);
nand (n1203,n1204,n1308);
or (n1204,n1205,n1303);
nor (n1205,n1206,n1302);
and (n1206,n1207,n1281);
nand (n1207,n1208,n1279);
or (n1208,n1209,n1263);
not (n1209,n1210);
or (n1210,n1211,n1262);
and (n1211,n1212,n1241);
xor (n1212,n1213,n1222);
nand (n1213,n1214,n1218);
or (n1214,n437,n1215);
nor (n1215,n1216,n1217);
and (n1216,n219,n410);
and (n1217,n408,n221);
or (n1218,n438,n1219);
nor (n1219,n1220,n1221);
and (n1220,n478,n219);
and (n1221,n476,n221);
nand (n1222,n1223,n1240);
or (n1223,n1224,n1230);
not (n1224,n1225);
nand (n1225,n1226,n219);
nand (n1226,n1227,n1229);
or (n1227,n1228,n416);
and (n1228,n408,n442);
nand (n1229,n410,n441);
not (n1230,n1231);
nand (n1231,n1232,n1236);
or (n1232,n1233,n418);
or (n1233,n1234,n1235);
and (n1234,n360,n416);
and (n1235,n362,n415);
or (n1236,n1237,n419);
nor (n1237,n1238,n1239);
and (n1238,n331,n416);
and (n1239,n329,n415);
or (n1240,n1231,n1225);
or (n1241,n1242,n1261);
and (n1242,n1243,n1251);
xor (n1243,n1244,n1245);
nor (n1244,n438,n410);
nand (n1245,n1246,n1250);
or (n1246,n1247,n418);
nor (n1247,n1248,n1249);
and (n1248,n478,n416);
and (n1249,n476,n415);
or (n1250,n1233,n419);
nor (n1251,n1252,n1259);
nor (n1252,n1253,n1255);
and (n1253,n1254,n420);
not (n1254,n1247);
and (n1255,n1256,n565);
nand (n1256,n1257,n1258);
or (n1257,n410,n416);
nand (n1258,n416,n410);
or (n1259,n1260,n415);
and (n1260,n408,n420);
and (n1261,n1244,n1245);
and (n1262,n1213,n1222);
not (n1263,n1264);
nand (n1264,n1265,n1278);
not (n1265,n1266);
xor (n1266,n1267,n1275);
xor (n1267,n1268,n1269);
and (n1268,n225,n408);
nand (n1269,n1270,n1271);
or (n1270,n1219,n437);
nand (n1271,n1272,n439);
nor (n1272,n1273,n1274);
and (n1273,n362,n221);
and (n1274,n360,n219);
nand (n1275,n1276,n1277);
or (n1276,n1237,n418);
or (n1277,n1197,n419);
nand (n1278,n1224,n1231);
nand (n1279,n1280,n1266);
not (n1280,n1278);
nand (n1281,n1282,n1298);
not (n1282,n1283);
xor (n1283,n1284,n1297);
xor (n1284,n1285,n1289);
nand (n1285,n1286,n1288);
or (n1286,n1287,n437);
not (n1287,n1272);
nand (n1288,n1168,n439);
nand (n1289,n1290,n1295);
or (n1290,n1291,n214);
not (n1291,n1292);
nand (n1292,n1293,n1294);
or (n1293,n408,n151);
or (n1294,n410,n152);
nand (n1295,n1296,n225);
not (n1296,n1183);
xor (n1297,n1188,n1194);
not (n1298,n1299);
or (n1299,n1300,n1301);
and (n1300,n1267,n1275);
and (n1301,n1268,n1269);
nor (n1302,n1282,n1298);
nor (n1303,n1304,n1305);
xor (n1304,n1180,n1200);
or (n1305,n1306,n1307);
and (n1306,n1284,n1297);
and (n1307,n1285,n1289);
nand (n1308,n1304,n1305);
and (n1309,n1178,n1202);
nand (n1310,n1311,n1315);
not (n1311,n1312);
or (n1312,n1313,n1314);
and (n1313,n1124,n1149);
and (n1314,n1125,n1148);
not (n1315,n1316);
xor (n1316,n980,n1050);
nand (n1317,n1318,n1310);
not (n1318,n1319);
nand (n1319,n1123,n1150);
nand (n1320,n1316,n1312);
and (n1321,n978,n1088);
or (n1322,n1323,n1338);
xor (n1323,n1324,n1335);
xor (n1324,n1325,n1326);
xor (n1325,n949,n962);
xor (n1326,n1327,n1334);
xor (n1327,n1328,n1331);
or (n1328,n1329,n1330);
and (n1329,n1111,n1116);
and (n1330,n1112,n1113);
or (n1331,n1332,n1333);
and (n1332,n1091,n1098);
and (n1333,n1092,n1095);
xor (n1334,n908,n923);
or (n1335,n1336,n1337);
and (n1336,n1105,n1110);
and (n1337,n1106,n1107);
or (n1338,n1339,n1340);
and (n1339,n1089,n1104);
and (n1340,n1090,n1101);
and (n1341,n1323,n1338);
nand (n1342,n1343,n1357);
not (n1343,n1344);
and (n1344,n1345,n1353);
not (n1345,n1346);
xor (n1346,n1347,n1352);
xor (n1347,n1348,n1349);
xor (n1348,n885,n906);
or (n1349,n1350,n1351);
and (n1350,n1327,n1334);
and (n1351,n1328,n1331);
xor (n1352,n944,n947);
not (n1353,n1354);
or (n1354,n1355,n1356);
and (n1355,n1324,n1335);
and (n1356,n1325,n1326);
nand (n1357,n1358,n1360);
not (n1358,n1359);
xor (n1359,n940,n968);
not (n1360,n1361);
or (n1361,n1362,n1363);
and (n1362,n1347,n1352);
and (n1363,n1348,n1349);
nor (n1364,n1365,n1367);
and (n1365,n1357,n1366);
nor (n1366,n1345,n1353);
nor (n1367,n1358,n1360);
and (n1368,n938,n970);
and (n1369,n873,n934);
nor (n1370,n1371,n1380);
and (n1371,n1372,n748);
nand (n1372,n1373,n1375);
not (n1373,n1374);
and (n1374,n865,n866);
nand (n1375,n1376,n864);
nand (n1376,n1377,n1379);
or (n1377,n297,n1378);
nand (n1378,n747,n685);
nand (n1379,n298,n592);
and (n1380,n819,n749);
nor (n1381,n1382,n1406);
nor (n1382,n1383,n1386);
or (n1383,n1384,n1385);
and (n1384,n820,n861);
and (n1385,n821,n840);
xor (n1386,n1387,n1403);
xor (n1387,n1388,n1391);
or (n1388,n1389,n1390);
and (n1389,n822,n829);
and (n1390,n823,n826);
xor (n1391,n1392,n1397);
xor (n1392,n1393,n1394);
xor (n1393,n210,n236);
or (n1394,n1395,n1396);
and (n1395,n843,n851);
and (n1396,n844,n847);
xor (n1397,n1398,n1402);
xor (n1398,n852,n1399);
or (n1399,n1400,n1401);
and (n1400,n830,n837);
and (n1401,n831,n834);
xor (n1402,n70,n101);
or (n1403,n1404,n1405);
and (n1404,n841,n858);
and (n1405,n842,n855);
nor (n1406,n1407,n1410);
or (n1407,n1408,n1409);
and (n1408,n1387,n1403);
and (n1409,n1388,n1391);
xor (n1410,n1411,n1416);
xor (n1411,n1412,n1415);
or (n1412,n1413,n1414);
and (n1413,n1398,n1402);
and (n1414,n852,n1399);
xor (n1415,n207,n244);
or (n1416,n1417,n1418);
and (n1417,n1392,n1397);
and (n1418,n1393,n1394);
nand (n1419,n1420,n1422);
or (n1420,n1421,n1406);
nand (n1421,n1383,n1386);
nand (n1422,n1407,n1410);
nor (n1423,n1424,n1425);
xor (n1424,n13,n205);
or (n1425,n1426,n1427);
and (n1426,n1411,n1416);
and (n1427,n1412,n1415);
nand (n1428,n1425,n1424);
or (n1429,n289,n9);
and (n1430,n1431,n1432);
not (n1432,n2);
or (n1433,n1434,n1430);
and (n1434,n1435,n2);
xor (n1435,n1436,n2623);
xor (n1436,n1437,n2741);
xor (n1437,n1438,n2618);
xor (n1438,n1439,n2734);
xor (n1439,n1440,n2612);
xor (n1440,n1441,n2722);
xor (n1441,n1442,n2606);
xor (n1442,n1443,n2705);
xor (n1443,n1444,n2600);
xor (n1444,n1445,n2683);
xor (n1445,n1446,n2594);
xor (n1446,n1447,n2656);
xor (n1447,n1448,n2588);
xor (n1448,n1449,n2624);
xor (n1449,n1450,n2582);
xor (n1450,n1451,n2579);
xor (n1451,n1452,n2578);
xor (n1452,n1453,n2527);
xor (n1453,n1454,n2526);
xor (n1454,n1455,n2469);
xor (n1455,n1456,n2468);
xor (n1456,n1457,n2405);
xor (n1457,n1458,n2404);
xor (n1458,n1459,n2335);
xor (n1459,n1460,n2334);
xor (n1460,n1461,n2260);
xor (n1461,n1462,n2259);
xor (n1462,n1463,n2181);
xor (n1463,n1464,n2180);
xor (n1464,n1465,n1496);
xor (n1465,n1466,n1495);
xor (n1466,n1467,n1494);
xor (n1467,n1468,n1493);
xor (n1468,n1469,n1492);
xor (n1469,n1470,n1491);
xor (n1470,n1471,n1490);
xor (n1471,n1472,n1489);
xor (n1472,n1473,n1488);
xor (n1473,n1474,n1487);
xor (n1474,n1475,n1486);
xor (n1475,n1476,n1485);
xor (n1476,n1477,n1484);
xor (n1477,n1478,n1483);
xor (n1478,n1479,n1482);
xor (n1479,n1480,n1481);
and (n1480,n167,n420);
and (n1481,n167,n416);
and (n1482,n1480,n1481);
and (n1483,n167,n442);
and (n1484,n1478,n1483);
and (n1485,n167,n219);
and (n1486,n1476,n1485);
and (n1487,n167,n218);
and (n1488,n1474,n1487);
and (n1489,n167,n152);
and (n1490,n1472,n1489);
and (n1491,n167,n153);
and (n1492,n1470,n1491);
and (n1493,n167,n50);
and (n1494,n1468,n1493);
and (n1495,n167,n51);
or (n1496,n1497,n2097);
and (n1497,n1498,n2096);
xor (n1498,n1467,n1499);
or (n1499,n1500,n2014);
and (n1500,n1501,n2013);
xor (n1501,n1469,n1502);
or (n1502,n1503,n1931);
and (n1503,n1504,n1930);
xor (n1504,n1471,n1505);
or (n1505,n1506,n1847);
and (n1506,n1507,n1846);
xor (n1507,n1473,n1508);
or (n1508,n1509,n1764);
and (n1509,n1510,n1763);
xor (n1510,n1475,n1511);
or (n1511,n1512,n1683);
and (n1512,n1513,n1682);
xor (n1513,n1477,n1514);
or (n1514,n1515,n1600);
and (n1515,n1516,n1599);
xor (n1516,n1479,n1517);
or (n1517,n1518,n1520);
and (n1518,n1480,n1519);
and (n1519,n161,n416);
and (n1520,n1521,n1522);
xor (n1521,n1480,n1519);
or (n1522,n1523,n1526);
and (n1523,n1524,n1525);
and (n1524,n161,n420);
and (n1525,n65,n416);
and (n1526,n1527,n1528);
xor (n1527,n1524,n1525);
or (n1528,n1529,n1532);
and (n1529,n1530,n1531);
and (n1530,n65,n420);
and (n1531,n59,n416);
and (n1532,n1533,n1534);
xor (n1533,n1530,n1531);
or (n1534,n1535,n1538);
and (n1535,n1536,n1537);
and (n1536,n59,n420);
and (n1537,n40,n416);
and (n1538,n1539,n1540);
xor (n1539,n1536,n1537);
or (n1540,n1541,n1544);
and (n1541,n1542,n1543);
and (n1542,n40,n420);
and (n1543,n34,n416);
and (n1544,n1545,n1546);
xor (n1545,n1542,n1543);
or (n1546,n1547,n1550);
and (n1547,n1548,n1549);
and (n1548,n34,n420);
and (n1549,n137,n416);
and (n1550,n1551,n1552);
xor (n1551,n1548,n1549);
or (n1552,n1553,n1555);
and (n1553,n1554,n1005);
and (n1554,n137,n420);
and (n1555,n1556,n1557);
xor (n1556,n1554,n1005);
or (n1557,n1558,n1561);
and (n1558,n1559,n1560);
and (n1559,n92,n420);
and (n1560,n86,n416);
and (n1561,n1562,n1563);
xor (n1562,n1559,n1560);
or (n1563,n1564,n1566);
and (n1564,n1565,n1044);
and (n1565,n86,n420);
and (n1566,n1567,n1568);
xor (n1567,n1565,n1044);
or (n1568,n1569,n1571);
and (n1569,n1570,n1163);
and (n1570,n122,n420);
and (n1571,n1572,n1573);
xor (n1572,n1570,n1163);
or (n1573,n1574,n1577);
and (n1574,n1575,n1576);
and (n1575,n116,n420);
and (n1576,n335,n416);
and (n1577,n1578,n1579);
xor (n1578,n1575,n1576);
or (n1579,n1580,n1583);
and (n1580,n1581,n1582);
and (n1581,n335,n420);
and (n1582,n329,n416);
and (n1583,n1584,n1585);
xor (n1584,n1581,n1582);
or (n1585,n1586,n1588);
and (n1586,n1587,n1234);
and (n1587,n329,n420);
and (n1588,n1589,n1590);
xor (n1589,n1587,n1234);
or (n1590,n1591,n1594);
and (n1591,n1592,n1593);
and (n1592,n360,n420);
and (n1593,n476,n416);
and (n1594,n1595,n1596);
xor (n1595,n1592,n1593);
and (n1596,n1597,n1598);
and (n1597,n476,n420);
and (n1598,n408,n416);
and (n1599,n161,n442);
and (n1600,n1601,n1602);
xor (n1601,n1516,n1599);
or (n1602,n1603,n1606);
and (n1603,n1604,n1605);
xor (n1604,n1521,n1522);
and (n1605,n65,n442);
and (n1606,n1607,n1608);
xor (n1607,n1604,n1605);
or (n1608,n1609,n1612);
and (n1609,n1610,n1611);
xor (n1610,n1527,n1528);
and (n1611,n59,n442);
and (n1612,n1613,n1614);
xor (n1613,n1610,n1611);
or (n1614,n1615,n1618);
and (n1615,n1616,n1617);
xor (n1616,n1533,n1534);
and (n1617,n40,n442);
and (n1618,n1619,n1620);
xor (n1619,n1616,n1617);
or (n1620,n1621,n1624);
and (n1621,n1622,n1623);
xor (n1622,n1539,n1540);
and (n1623,n34,n442);
and (n1624,n1625,n1626);
xor (n1625,n1622,n1623);
or (n1626,n1627,n1630);
and (n1627,n1628,n1629);
xor (n1628,n1545,n1546);
and (n1629,n137,n442);
and (n1630,n1631,n1632);
xor (n1631,n1628,n1629);
or (n1632,n1633,n1636);
and (n1633,n1634,n1635);
xor (n1634,n1551,n1552);
and (n1635,n92,n442);
and (n1636,n1637,n1638);
xor (n1637,n1634,n1635);
or (n1638,n1639,n1642);
and (n1639,n1640,n1641);
xor (n1640,n1556,n1557);
and (n1641,n86,n442);
and (n1642,n1643,n1644);
xor (n1643,n1640,n1641);
or (n1644,n1645,n1648);
and (n1645,n1646,n1647);
xor (n1646,n1562,n1563);
and (n1647,n122,n442);
and (n1648,n1649,n1650);
xor (n1649,n1646,n1647);
or (n1650,n1651,n1654);
and (n1651,n1652,n1653);
xor (n1652,n1567,n1568);
and (n1653,n116,n442);
and (n1654,n1655,n1656);
xor (n1655,n1652,n1653);
or (n1656,n1657,n1660);
and (n1657,n1658,n1659);
xor (n1658,n1572,n1573);
and (n1659,n335,n442);
and (n1660,n1661,n1662);
xor (n1661,n1658,n1659);
or (n1662,n1663,n1666);
and (n1663,n1664,n1665);
xor (n1664,n1578,n1579);
and (n1665,n329,n442);
and (n1666,n1667,n1668);
xor (n1667,n1664,n1665);
or (n1668,n1669,n1672);
and (n1669,n1670,n1671);
xor (n1670,n1584,n1585);
and (n1671,n360,n442);
and (n1672,n1673,n1674);
xor (n1673,n1670,n1671);
or (n1674,n1675,n1678);
and (n1675,n1676,n1677);
xor (n1676,n1589,n1590);
and (n1677,n476,n442);
and (n1678,n1679,n1680);
xor (n1679,n1676,n1677);
and (n1680,n1681,n1228);
xor (n1681,n1595,n1596);
and (n1682,n161,n219);
and (n1683,n1684,n1685);
xor (n1684,n1513,n1682);
or (n1685,n1686,n1689);
and (n1686,n1687,n1688);
xor (n1687,n1601,n1602);
and (n1688,n65,n219);
and (n1689,n1690,n1691);
xor (n1690,n1687,n1688);
or (n1691,n1692,n1695);
and (n1692,n1693,n1694);
xor (n1693,n1607,n1608);
and (n1694,n59,n219);
and (n1695,n1696,n1697);
xor (n1696,n1693,n1694);
or (n1697,n1698,n1701);
and (n1698,n1699,n1700);
xor (n1699,n1613,n1614);
and (n1700,n40,n219);
and (n1701,n1702,n1703);
xor (n1702,n1699,n1700);
or (n1703,n1704,n1707);
and (n1704,n1705,n1706);
xor (n1705,n1619,n1620);
and (n1706,n34,n219);
and (n1707,n1708,n1709);
xor (n1708,n1705,n1706);
or (n1709,n1710,n1713);
and (n1710,n1711,n1712);
xor (n1711,n1625,n1626);
and (n1712,n137,n219);
and (n1713,n1714,n1715);
xor (n1714,n1711,n1712);
or (n1715,n1716,n1719);
and (n1716,n1717,n1718);
xor (n1717,n1631,n1632);
and (n1718,n92,n219);
and (n1719,n1720,n1721);
xor (n1720,n1717,n1718);
or (n1721,n1722,n1725);
and (n1722,n1723,n1724);
xor (n1723,n1637,n1638);
and (n1724,n86,n219);
and (n1725,n1726,n1727);
xor (n1726,n1723,n1724);
or (n1727,n1728,n1731);
and (n1728,n1729,n1730);
xor (n1729,n1643,n1644);
and (n1730,n122,n219);
and (n1731,n1732,n1733);
xor (n1732,n1729,n1730);
or (n1733,n1734,n1737);
and (n1734,n1735,n1736);
xor (n1735,n1649,n1650);
and (n1736,n116,n219);
and (n1737,n1738,n1739);
xor (n1738,n1735,n1736);
or (n1739,n1740,n1742);
and (n1740,n1741,n1138);
xor (n1741,n1655,n1656);
and (n1742,n1743,n1744);
xor (n1743,n1741,n1138);
or (n1744,n1745,n1747);
and (n1745,n1746,n1170);
xor (n1746,n1661,n1662);
and (n1747,n1748,n1749);
xor (n1748,n1746,n1170);
or (n1749,n1750,n1752);
and (n1750,n1751,n1274);
xor (n1751,n1667,n1668);
and (n1752,n1753,n1754);
xor (n1753,n1751,n1274);
or (n1754,n1755,n1758);
and (n1755,n1756,n1757);
xor (n1756,n1673,n1674);
and (n1757,n476,n219);
and (n1758,n1759,n1760);
xor (n1759,n1756,n1757);
and (n1760,n1761,n1762);
xor (n1761,n1679,n1680);
and (n1762,n408,n219);
and (n1763,n161,n218);
and (n1764,n1765,n1766);
xor (n1765,n1510,n1763);
or (n1766,n1767,n1770);
and (n1767,n1768,n1769);
xor (n1768,n1684,n1685);
and (n1769,n65,n218);
and (n1770,n1771,n1772);
xor (n1771,n1768,n1769);
or (n1772,n1773,n1776);
and (n1773,n1774,n1775);
xor (n1774,n1690,n1691);
and (n1775,n59,n218);
and (n1776,n1777,n1778);
xor (n1777,n1774,n1775);
or (n1778,n1779,n1782);
and (n1779,n1780,n1781);
xor (n1780,n1696,n1697);
and (n1781,n40,n218);
and (n1782,n1783,n1784);
xor (n1783,n1780,n1781);
or (n1784,n1785,n1788);
and (n1785,n1786,n1787);
xor (n1786,n1702,n1703);
and (n1787,n34,n218);
and (n1788,n1789,n1790);
xor (n1789,n1786,n1787);
or (n1790,n1791,n1794);
and (n1791,n1792,n1793);
xor (n1792,n1708,n1709);
and (n1793,n137,n218);
and (n1794,n1795,n1796);
xor (n1795,n1792,n1793);
or (n1796,n1797,n1800);
and (n1797,n1798,n1799);
xor (n1798,n1714,n1715);
and (n1799,n92,n218);
and (n1800,n1801,n1802);
xor (n1801,n1798,n1799);
or (n1802,n1803,n1806);
and (n1803,n1804,n1805);
xor (n1804,n1720,n1721);
and (n1805,n86,n218);
and (n1806,n1807,n1808);
xor (n1807,n1804,n1805);
or (n1808,n1809,n1812);
and (n1809,n1810,n1811);
xor (n1810,n1726,n1727);
and (n1811,n122,n218);
and (n1812,n1813,n1814);
xor (n1813,n1810,n1811);
or (n1814,n1815,n1818);
and (n1815,n1816,n1817);
xor (n1816,n1732,n1733);
and (n1817,n116,n218);
and (n1818,n1819,n1820);
xor (n1819,n1816,n1817);
or (n1820,n1821,n1824);
and (n1821,n1822,n1823);
xor (n1822,n1738,n1739);
and (n1823,n335,n218);
and (n1824,n1825,n1826);
xor (n1825,n1822,n1823);
or (n1826,n1827,n1830);
and (n1827,n1828,n1829);
xor (n1828,n1743,n1744);
and (n1829,n329,n218);
and (n1830,n1831,n1832);
xor (n1831,n1828,n1829);
or (n1832,n1833,n1836);
and (n1833,n1834,n1835);
xor (n1834,n1748,n1749);
and (n1835,n360,n218);
and (n1836,n1837,n1838);
xor (n1837,n1834,n1835);
or (n1838,n1839,n1842);
and (n1839,n1840,n1841);
xor (n1840,n1753,n1754);
and (n1841,n476,n218);
and (n1842,n1843,n1844);
xor (n1843,n1840,n1841);
and (n1844,n1845,n1193);
xor (n1845,n1759,n1760);
and (n1846,n161,n152);
and (n1847,n1848,n1849);
xor (n1848,n1507,n1846);
or (n1849,n1850,n1853);
and (n1850,n1851,n1852);
xor (n1851,n1765,n1766);
and (n1852,n65,n152);
and (n1853,n1854,n1855);
xor (n1854,n1851,n1852);
or (n1855,n1856,n1859);
and (n1856,n1857,n1858);
xor (n1857,n1771,n1772);
and (n1858,n59,n152);
and (n1859,n1860,n1861);
xor (n1860,n1857,n1858);
or (n1861,n1862,n1865);
and (n1862,n1863,n1864);
xor (n1863,n1777,n1778);
and (n1864,n40,n152);
and (n1865,n1866,n1867);
xor (n1866,n1863,n1864);
or (n1867,n1868,n1871);
and (n1868,n1869,n1870);
xor (n1869,n1783,n1784);
and (n1870,n34,n152);
and (n1871,n1872,n1873);
xor (n1872,n1869,n1870);
or (n1873,n1874,n1877);
and (n1874,n1875,n1876);
xor (n1875,n1789,n1790);
and (n1876,n137,n152);
and (n1877,n1878,n1879);
xor (n1878,n1875,n1876);
or (n1879,n1880,n1883);
and (n1880,n1881,n1882);
xor (n1881,n1795,n1796);
and (n1882,n92,n152);
and (n1883,n1884,n1885);
xor (n1884,n1881,n1882);
or (n1885,n1886,n1889);
and (n1886,n1887,n1888);
xor (n1887,n1801,n1802);
and (n1888,n86,n152);
and (n1889,n1890,n1891);
xor (n1890,n1887,n1888);
or (n1891,n1892,n1895);
and (n1892,n1893,n1894);
xor (n1893,n1807,n1808);
and (n1894,n122,n152);
and (n1895,n1896,n1897);
xor (n1896,n1893,n1894);
or (n1897,n1898,n1901);
and (n1898,n1899,n1900);
xor (n1899,n1813,n1814);
and (n1900,n116,n152);
and (n1901,n1902,n1903);
xor (n1902,n1899,n1900);
or (n1903,n1904,n1907);
and (n1904,n1905,n1906);
xor (n1905,n1819,n1820);
and (n1906,n335,n152);
and (n1907,n1908,n1909);
xor (n1908,n1905,n1906);
or (n1909,n1910,n1913);
and (n1910,n1911,n1912);
xor (n1911,n1825,n1826);
and (n1912,n329,n152);
and (n1913,n1914,n1915);
xor (n1914,n1911,n1912);
or (n1915,n1916,n1919);
and (n1916,n1917,n1918);
xor (n1917,n1831,n1832);
and (n1918,n360,n152);
and (n1919,n1920,n1921);
xor (n1920,n1917,n1918);
or (n1921,n1922,n1925);
and (n1922,n1923,n1924);
xor (n1923,n1837,n1838);
and (n1924,n476,n152);
and (n1925,n1926,n1927);
xor (n1926,n1923,n1924);
and (n1927,n1928,n1929);
xor (n1928,n1843,n1844);
and (n1929,n408,n152);
and (n1930,n161,n153);
and (n1931,n1932,n1933);
xor (n1932,n1504,n1930);
or (n1933,n1934,n1937);
and (n1934,n1935,n1936);
xor (n1935,n1848,n1849);
and (n1936,n65,n153);
and (n1937,n1938,n1939);
xor (n1938,n1935,n1936);
or (n1939,n1940,n1943);
and (n1940,n1941,n1942);
xor (n1941,n1854,n1855);
and (n1942,n59,n153);
and (n1943,n1944,n1945);
xor (n1944,n1941,n1942);
or (n1945,n1946,n1949);
and (n1946,n1947,n1948);
xor (n1947,n1860,n1861);
and (n1948,n40,n153);
and (n1949,n1950,n1951);
xor (n1950,n1947,n1948);
or (n1951,n1952,n1955);
and (n1952,n1953,n1954);
xor (n1953,n1866,n1867);
and (n1954,n34,n153);
and (n1955,n1956,n1957);
xor (n1956,n1953,n1954);
or (n1957,n1958,n1961);
and (n1958,n1959,n1960);
xor (n1959,n1872,n1873);
and (n1960,n137,n153);
and (n1961,n1962,n1963);
xor (n1962,n1959,n1960);
or (n1963,n1964,n1967);
and (n1964,n1965,n1966);
xor (n1965,n1878,n1879);
and (n1966,n92,n153);
and (n1967,n1968,n1969);
xor (n1968,n1965,n1966);
or (n1969,n1970,n1973);
and (n1970,n1971,n1972);
xor (n1971,n1884,n1885);
and (n1972,n86,n153);
and (n1973,n1974,n1975);
xor (n1974,n1971,n1972);
or (n1975,n1976,n1979);
and (n1976,n1977,n1978);
xor (n1977,n1890,n1891);
and (n1978,n122,n153);
and (n1979,n1980,n1981);
xor (n1980,n1977,n1978);
or (n1981,n1982,n1985);
and (n1982,n1983,n1984);
xor (n1983,n1896,n1897);
and (n1984,n116,n153);
and (n1985,n1986,n1987);
xor (n1986,n1983,n1984);
or (n1987,n1988,n1991);
and (n1988,n1989,n1990);
xor (n1989,n1902,n1903);
and (n1990,n335,n153);
and (n1991,n1992,n1993);
xor (n1992,n1989,n1990);
or (n1993,n1994,n1997);
and (n1994,n1995,n1996);
xor (n1995,n1908,n1909);
and (n1996,n329,n153);
and (n1997,n1998,n1999);
xor (n1998,n1995,n1996);
or (n1999,n2000,n2003);
and (n2000,n2001,n2002);
xor (n2001,n1914,n1915);
and (n2002,n360,n153);
and (n2003,n2004,n2005);
xor (n2004,n2001,n2002);
or (n2005,n2006,n2009);
and (n2006,n2007,n2008);
xor (n2007,n1920,n1921);
and (n2008,n476,n153);
and (n2009,n2010,n2011);
xor (n2010,n2007,n2008);
and (n2011,n2012,n1037);
xor (n2012,n1926,n1927);
and (n2013,n161,n50);
and (n2014,n2015,n2016);
xor (n2015,n1501,n2013);
or (n2016,n2017,n2020);
and (n2017,n2018,n2019);
xor (n2018,n1932,n1933);
and (n2019,n65,n50);
and (n2020,n2021,n2022);
xor (n2021,n2018,n2019);
or (n2022,n2023,n2026);
and (n2023,n2024,n2025);
xor (n2024,n1938,n1939);
and (n2025,n59,n50);
and (n2026,n2027,n2028);
xor (n2027,n2024,n2025);
or (n2028,n2029,n2032);
and (n2029,n2030,n2031);
xor (n2030,n1944,n1945);
and (n2031,n40,n50);
and (n2032,n2033,n2034);
xor (n2033,n2030,n2031);
or (n2034,n2035,n2038);
and (n2035,n2036,n2037);
xor (n2036,n1950,n1951);
and (n2037,n34,n50);
and (n2038,n2039,n2040);
xor (n2039,n2036,n2037);
or (n2040,n2041,n2044);
and (n2041,n2042,n2043);
xor (n2042,n1956,n1957);
and (n2043,n137,n50);
and (n2044,n2045,n2046);
xor (n2045,n2042,n2043);
or (n2046,n2047,n2050);
and (n2047,n2048,n2049);
xor (n2048,n1962,n1963);
and (n2049,n92,n50);
and (n2050,n2051,n2052);
xor (n2051,n2048,n2049);
or (n2052,n2053,n2056);
and (n2053,n2054,n2055);
xor (n2054,n1968,n1969);
and (n2055,n86,n50);
and (n2056,n2057,n2058);
xor (n2057,n2054,n2055);
or (n2058,n2059,n2062);
and (n2059,n2060,n2061);
xor (n2060,n1974,n1975);
and (n2061,n122,n50);
and (n2062,n2063,n2064);
xor (n2063,n2060,n2061);
or (n2064,n2065,n2068);
and (n2065,n2066,n2067);
xor (n2066,n1980,n1981);
and (n2067,n116,n50);
and (n2068,n2069,n2070);
xor (n2069,n2066,n2067);
or (n2070,n2071,n2074);
and (n2071,n2072,n2073);
xor (n2072,n1986,n1987);
and (n2073,n335,n50);
and (n2074,n2075,n2076);
xor (n2075,n2072,n2073);
or (n2076,n2077,n2080);
and (n2077,n2078,n2079);
xor (n2078,n1992,n1993);
and (n2079,n329,n50);
and (n2080,n2081,n2082);
xor (n2081,n2078,n2079);
or (n2082,n2083,n2086);
and (n2083,n2084,n2085);
xor (n2084,n1998,n1999);
and (n2085,n360,n50);
and (n2086,n2087,n2088);
xor (n2087,n2084,n2085);
or (n2088,n2089,n2091);
and (n2089,n2090,n1085);
xor (n2090,n2004,n2005);
and (n2091,n2092,n2093);
xor (n2092,n2090,n1085);
and (n2093,n2094,n2095);
xor (n2094,n2010,n2011);
and (n2095,n408,n50);
and (n2096,n161,n51);
and (n2097,n2098,n2099);
xor (n2098,n1498,n2096);
or (n2099,n2100,n2103);
and (n2100,n2101,n2102);
xor (n2101,n2015,n2016);
and (n2102,n65,n51);
and (n2103,n2104,n2105);
xor (n2104,n2101,n2102);
or (n2105,n2106,n2109);
and (n2106,n2107,n2108);
xor (n2107,n2021,n2022);
and (n2108,n59,n51);
and (n2109,n2110,n2111);
xor (n2110,n2107,n2108);
or (n2111,n2112,n2115);
and (n2112,n2113,n2114);
xor (n2113,n2027,n2028);
and (n2114,n40,n51);
and (n2115,n2116,n2117);
xor (n2116,n2113,n2114);
or (n2117,n2118,n2121);
and (n2118,n2119,n2120);
xor (n2119,n2033,n2034);
and (n2120,n34,n51);
and (n2121,n2122,n2123);
xor (n2122,n2119,n2120);
or (n2123,n2124,n2127);
and (n2124,n2125,n2126);
xor (n2125,n2039,n2040);
and (n2126,n137,n51);
and (n2127,n2128,n2129);
xor (n2128,n2125,n2126);
or (n2129,n2130,n2133);
and (n2130,n2131,n2132);
xor (n2131,n2045,n2046);
and (n2132,n92,n51);
and (n2133,n2134,n2135);
xor (n2134,n2131,n2132);
or (n2135,n2136,n2139);
and (n2136,n2137,n2138);
xor (n2137,n2051,n2052);
and (n2138,n86,n51);
and (n2139,n2140,n2141);
xor (n2140,n2137,n2138);
or (n2141,n2142,n2145);
and (n2142,n2143,n2144);
xor (n2143,n2057,n2058);
and (n2144,n122,n51);
and (n2145,n2146,n2147);
xor (n2146,n2143,n2144);
or (n2147,n2148,n2151);
and (n2148,n2149,n2150);
xor (n2149,n2063,n2064);
and (n2150,n116,n51);
and (n2151,n2152,n2153);
xor (n2152,n2149,n2150);
or (n2153,n2154,n2157);
and (n2154,n2155,n2156);
xor (n2155,n2069,n2070);
and (n2156,n335,n51);
and (n2157,n2158,n2159);
xor (n2158,n2155,n2156);
or (n2159,n2160,n2163);
and (n2160,n2161,n2162);
xor (n2161,n2075,n2076);
and (n2162,n329,n51);
and (n2163,n2164,n2165);
xor (n2164,n2161,n2162);
or (n2165,n2166,n2169);
and (n2166,n2167,n2168);
xor (n2167,n2081,n2082);
and (n2168,n360,n51);
and (n2169,n2170,n2171);
xor (n2170,n2167,n2168);
or (n2171,n2172,n2175);
and (n2172,n2173,n2174);
xor (n2173,n2087,n2088);
and (n2174,n476,n51);
and (n2175,n2176,n2177);
xor (n2176,n2173,n2174);
and (n2177,n2178,n2179);
xor (n2178,n2092,n2093);
not (n2179,n1062);
and (n2180,n161,n23);
or (n2181,n2182,n2185);
and (n2182,n2183,n2184);
xor (n2183,n2098,n2099);
and (n2184,n65,n23);
and (n2185,n2186,n2187);
xor (n2186,n2183,n2184);
or (n2187,n2188,n2191);
and (n2188,n2189,n2190);
xor (n2189,n2104,n2105);
and (n2190,n59,n23);
and (n2191,n2192,n2193);
xor (n2192,n2189,n2190);
or (n2193,n2194,n2197);
and (n2194,n2195,n2196);
xor (n2195,n2110,n2111);
and (n2196,n40,n23);
and (n2197,n2198,n2199);
xor (n2198,n2195,n2196);
or (n2199,n2200,n2203);
and (n2200,n2201,n2202);
xor (n2201,n2116,n2117);
and (n2202,n34,n23);
and (n2203,n2204,n2205);
xor (n2204,n2201,n2202);
or (n2205,n2206,n2209);
and (n2206,n2207,n2208);
xor (n2207,n2122,n2123);
and (n2208,n137,n23);
and (n2209,n2210,n2211);
xor (n2210,n2207,n2208);
or (n2211,n2212,n2215);
and (n2212,n2213,n2214);
xor (n2213,n2128,n2129);
and (n2214,n92,n23);
and (n2215,n2216,n2217);
xor (n2216,n2213,n2214);
or (n2217,n2218,n2220);
and (n2218,n2219,n497);
xor (n2219,n2134,n2135);
and (n2220,n2221,n2222);
xor (n2221,n2219,n497);
or (n2222,n2223,n2226);
and (n2223,n2224,n2225);
xor (n2224,n2140,n2141);
and (n2225,n122,n23);
and (n2226,n2227,n2228);
xor (n2227,n2224,n2225);
or (n2228,n2229,n2232);
and (n2229,n2230,n2231);
xor (n2230,n2146,n2147);
and (n2231,n116,n23);
and (n2232,n2233,n2234);
xor (n2233,n2230,n2231);
or (n2234,n2235,n2237);
and (n2235,n2236,n654);
xor (n2236,n2152,n2153);
and (n2237,n2238,n2239);
xor (n2238,n2236,n654);
or (n2239,n2240,n2243);
and (n2240,n2241,n2242);
xor (n2241,n2158,n2159);
and (n2242,n329,n23);
and (n2243,n2244,n2245);
xor (n2244,n2241,n2242);
or (n2245,n2246,n2248);
and (n2246,n2247,n921);
xor (n2247,n2164,n2165);
and (n2248,n2249,n2250);
xor (n2249,n2247,n921);
or (n2250,n2251,n2254);
and (n2251,n2252,n2253);
xor (n2252,n2170,n2171);
and (n2253,n476,n23);
and (n2254,n2255,n2256);
xor (n2255,n2252,n2253);
and (n2256,n2257,n2258);
xor (n2257,n2176,n2177);
and (n2258,n408,n23);
and (n2259,n65,n24);
or (n2260,n2261,n2264);
and (n2261,n2262,n2263);
xor (n2262,n2186,n2187);
and (n2263,n59,n24);
and (n2264,n2265,n2266);
xor (n2265,n2262,n2263);
or (n2266,n2267,n2270);
and (n2267,n2268,n2269);
xor (n2268,n2192,n2193);
and (n2269,n40,n24);
and (n2270,n2271,n2272);
xor (n2271,n2268,n2269);
or (n2272,n2273,n2276);
and (n2273,n2274,n2275);
xor (n2274,n2198,n2199);
and (n2275,n34,n24);
and (n2276,n2277,n2278);
xor (n2277,n2274,n2275);
or (n2278,n2279,n2282);
and (n2279,n2280,n2281);
xor (n2280,n2204,n2205);
and (n2281,n137,n24);
and (n2282,n2283,n2284);
xor (n2283,n2280,n2281);
or (n2284,n2285,n2288);
and (n2285,n2286,n2287);
xor (n2286,n2210,n2211);
and (n2287,n92,n24);
and (n2288,n2289,n2290);
xor (n2289,n2286,n2287);
or (n2290,n2291,n2294);
and (n2291,n2292,n2293);
xor (n2292,n2216,n2217);
and (n2293,n86,n24);
and (n2294,n2295,n2296);
xor (n2295,n2292,n2293);
or (n2296,n2297,n2300);
and (n2297,n2298,n2299);
xor (n2298,n2221,n2222);
and (n2299,n122,n24);
and (n2300,n2301,n2302);
xor (n2301,n2298,n2299);
or (n2302,n2303,n2306);
and (n2303,n2304,n2305);
xor (n2304,n2227,n2228);
and (n2305,n116,n24);
and (n2306,n2307,n2308);
xor (n2307,n2304,n2305);
or (n2308,n2309,n2312);
and (n2309,n2310,n2311);
xor (n2310,n2233,n2234);
and (n2311,n335,n24);
and (n2312,n2313,n2314);
xor (n2313,n2310,n2311);
or (n2314,n2315,n2318);
and (n2315,n2316,n2317);
xor (n2316,n2238,n2239);
and (n2317,n329,n24);
and (n2318,n2319,n2320);
xor (n2319,n2316,n2317);
or (n2320,n2321,n2324);
and (n2321,n2322,n2323);
xor (n2322,n2244,n2245);
and (n2323,n360,n24);
and (n2324,n2325,n2326);
xor (n2325,n2322,n2323);
or (n2326,n2327,n2330);
and (n2327,n2328,n2329);
xor (n2328,n2249,n2250);
and (n2329,n476,n24);
and (n2330,n2331,n2332);
xor (n2331,n2328,n2329);
and (n2332,n2333,n905);
xor (n2333,n2255,n2256);
and (n2334,n59,n30);
or (n2335,n2336,n2339);
and (n2336,n2337,n2338);
xor (n2337,n2265,n2266);
and (n2338,n40,n30);
and (n2339,n2340,n2341);
xor (n2340,n2337,n2338);
or (n2341,n2342,n2345);
and (n2342,n2343,n2344);
xor (n2343,n2271,n2272);
and (n2344,n34,n30);
and (n2345,n2346,n2347);
xor (n2346,n2343,n2344);
or (n2347,n2348,n2351);
and (n2348,n2349,n2350);
xor (n2349,n2277,n2278);
and (n2350,n137,n30);
and (n2351,n2352,n2353);
xor (n2352,n2349,n2350);
or (n2353,n2354,n2357);
and (n2354,n2355,n2356);
xor (n2355,n2283,n2284);
and (n2356,n92,n30);
and (n2357,n2358,n2359);
xor (n2358,n2355,n2356);
or (n2359,n2360,n2363);
and (n2360,n2361,n2362);
xor (n2361,n2289,n2290);
and (n2362,n86,n30);
and (n2363,n2364,n2365);
xor (n2364,n2361,n2362);
or (n2365,n2366,n2369);
and (n2366,n2367,n2368);
xor (n2367,n2295,n2296);
and (n2368,n122,n30);
and (n2369,n2370,n2371);
xor (n2370,n2367,n2368);
or (n2371,n2372,n2375);
and (n2372,n2373,n2374);
xor (n2373,n2301,n2302);
and (n2374,n116,n30);
and (n2375,n2376,n2377);
xor (n2376,n2373,n2374);
or (n2377,n2378,n2381);
and (n2378,n2379,n2380);
xor (n2379,n2307,n2308);
and (n2380,n335,n30);
and (n2381,n2382,n2383);
xor (n2382,n2379,n2380);
or (n2383,n2384,n2387);
and (n2384,n2385,n2386);
xor (n2385,n2313,n2314);
and (n2386,n329,n30);
and (n2387,n2388,n2389);
xor (n2388,n2385,n2386);
or (n2389,n2390,n2393);
and (n2390,n2391,n2392);
xor (n2391,n2319,n2320);
and (n2392,n360,n30);
and (n2393,n2394,n2395);
xor (n2394,n2391,n2392);
or (n2395,n2396,n2399);
and (n2396,n2397,n2398);
xor (n2397,n2325,n2326);
and (n2398,n476,n30);
and (n2399,n2400,n2401);
xor (n2400,n2397,n2398);
and (n2401,n2402,n2403);
xor (n2402,n2331,n2332);
and (n2403,n408,n30);
and (n2404,n40,n77);
or (n2405,n2406,n2409);
and (n2406,n2407,n2408);
xor (n2407,n2340,n2341);
and (n2408,n34,n77);
and (n2409,n2410,n2411);
xor (n2410,n2407,n2408);
or (n2411,n2412,n2415);
and (n2412,n2413,n2414);
xor (n2413,n2346,n2347);
and (n2414,n137,n77);
and (n2415,n2416,n2417);
xor (n2416,n2413,n2414);
or (n2417,n2418,n2421);
and (n2418,n2419,n2420);
xor (n2419,n2352,n2353);
and (n2420,n92,n77);
and (n2421,n2422,n2423);
xor (n2422,n2419,n2420);
or (n2423,n2424,n2427);
and (n2424,n2425,n2426);
xor (n2425,n2358,n2359);
and (n2426,n86,n77);
and (n2427,n2428,n2429);
xor (n2428,n2425,n2426);
or (n2429,n2430,n2433);
and (n2430,n2431,n2432);
xor (n2431,n2364,n2365);
and (n2432,n122,n77);
and (n2433,n2434,n2435);
xor (n2434,n2431,n2432);
or (n2435,n2436,n2439);
and (n2436,n2437,n2438);
xor (n2437,n2370,n2371);
and (n2438,n116,n77);
and (n2439,n2440,n2441);
xor (n2440,n2437,n2438);
or (n2441,n2442,n2445);
and (n2442,n2443,n2444);
xor (n2443,n2376,n2377);
and (n2444,n335,n77);
and (n2445,n2446,n2447);
xor (n2446,n2443,n2444);
or (n2447,n2448,n2451);
and (n2448,n2449,n2450);
xor (n2449,n2382,n2383);
and (n2450,n329,n77);
and (n2451,n2452,n2453);
xor (n2452,n2449,n2450);
or (n2453,n2454,n2457);
and (n2454,n2455,n2456);
xor (n2455,n2388,n2389);
and (n2456,n360,n77);
and (n2457,n2458,n2459);
xor (n2458,n2455,n2456);
or (n2459,n2460,n2463);
and (n2460,n2461,n2462);
xor (n2461,n2394,n2395);
and (n2462,n476,n77);
and (n2463,n2464,n2465);
xor (n2464,n2461,n2462);
and (n2465,n2466,n2467);
xor (n2466,n2400,n2401);
not (n2467,n620);
and (n2468,n34,n78);
or (n2469,n2470,n2473);
and (n2470,n2471,n2472);
xor (n2471,n2410,n2411);
and (n2472,n137,n78);
and (n2473,n2474,n2475);
xor (n2474,n2471,n2472);
or (n2475,n2476,n2479);
and (n2476,n2477,n2478);
xor (n2477,n2416,n2417);
and (n2478,n92,n78);
and (n2479,n2480,n2481);
xor (n2480,n2477,n2478);
or (n2481,n2482,n2485);
and (n2482,n2483,n2484);
xor (n2483,n2422,n2423);
and (n2484,n86,n78);
and (n2485,n2486,n2487);
xor (n2486,n2483,n2484);
or (n2487,n2488,n2491);
and (n2488,n2489,n2490);
xor (n2489,n2428,n2429);
and (n2490,n122,n78);
and (n2491,n2492,n2493);
xor (n2492,n2489,n2490);
or (n2493,n2494,n2497);
and (n2494,n2495,n2496);
xor (n2495,n2434,n2435);
and (n2496,n116,n78);
and (n2497,n2498,n2499);
xor (n2498,n2495,n2496);
or (n2499,n2500,n2503);
and (n2500,n2501,n2502);
xor (n2501,n2440,n2441);
and (n2502,n335,n78);
and (n2503,n2504,n2505);
xor (n2504,n2501,n2502);
or (n2505,n2506,n2509);
and (n2506,n2507,n2508);
xor (n2507,n2446,n2447);
and (n2508,n329,n78);
and (n2509,n2510,n2511);
xor (n2510,n2507,n2508);
or (n2511,n2512,n2515);
and (n2512,n2513,n2514);
xor (n2513,n2452,n2453);
and (n2514,n360,n78);
and (n2515,n2516,n2517);
xor (n2516,n2513,n2514);
or (n2517,n2518,n2521);
and (n2518,n2519,n2520);
xor (n2519,n2458,n2459);
and (n2520,n476,n78);
and (n2521,n2522,n2523);
xor (n2522,n2519,n2520);
and (n2523,n2524,n2525);
xor (n2524,n2464,n2465);
and (n2525,n408,n78);
and (n2526,n137,n106);
or (n2527,n2528,n2531);
and (n2528,n2529,n2530);
xor (n2529,n2474,n2475);
and (n2530,n92,n106);
and (n2531,n2532,n2533);
xor (n2532,n2529,n2530);
or (n2533,n2534,n2537);
and (n2534,n2535,n2536);
xor (n2535,n2480,n2481);
and (n2536,n86,n106);
and (n2537,n2538,n2539);
xor (n2538,n2535,n2536);
or (n2539,n2540,n2543);
and (n2540,n2541,n2542);
xor (n2541,n2486,n2487);
and (n2542,n122,n106);
and (n2543,n2544,n2545);
xor (n2544,n2541,n2542);
or (n2545,n2546,n2549);
and (n2546,n2547,n2548);
xor (n2547,n2492,n2493);
and (n2548,n116,n106);
and (n2549,n2550,n2551);
xor (n2550,n2547,n2548);
or (n2551,n2552,n2555);
and (n2552,n2553,n2554);
xor (n2553,n2498,n2499);
and (n2554,n335,n106);
and (n2555,n2556,n2557);
xor (n2556,n2553,n2554);
or (n2557,n2558,n2561);
and (n2558,n2559,n2560);
xor (n2559,n2504,n2505);
and (n2560,n329,n106);
and (n2561,n2562,n2563);
xor (n2562,n2559,n2560);
or (n2563,n2564,n2567);
and (n2564,n2565,n2566);
xor (n2565,n2510,n2511);
and (n2566,n360,n106);
and (n2567,n2568,n2569);
xor (n2568,n2565,n2566);
or (n2569,n2570,n2573);
and (n2570,n2571,n2572);
xor (n2571,n2516,n2517);
and (n2572,n476,n106);
and (n2573,n2574,n2575);
xor (n2574,n2571,n2572);
and (n2575,n2576,n2577);
xor (n2576,n2522,n2523);
not (n2577,n407);
and (n2578,n92,n112);
or (n2579,n2580,n2583);
and (n2580,n2581,n2582);
xor (n2581,n2532,n2533);
and (n2582,n86,n112);
and (n2583,n2584,n2585);
xor (n2584,n2581,n2582);
or (n2585,n2586,n2589);
and (n2586,n2587,n2588);
xor (n2587,n2538,n2539);
and (n2588,n122,n112);
and (n2589,n2590,n2591);
xor (n2590,n2587,n2588);
or (n2591,n2592,n2595);
and (n2592,n2593,n2594);
xor (n2593,n2544,n2545);
and (n2594,n116,n112);
and (n2595,n2596,n2597);
xor (n2596,n2593,n2594);
or (n2597,n2598,n2601);
and (n2598,n2599,n2600);
xor (n2599,n2550,n2551);
and (n2600,n335,n112);
and (n2601,n2602,n2603);
xor (n2602,n2599,n2600);
or (n2603,n2604,n2607);
and (n2604,n2605,n2606);
xor (n2605,n2556,n2557);
and (n2606,n329,n112);
and (n2607,n2608,n2609);
xor (n2608,n2605,n2606);
or (n2609,n2610,n2613);
and (n2610,n2611,n2612);
xor (n2611,n2562,n2563);
and (n2612,n360,n112);
and (n2613,n2614,n2615);
xor (n2614,n2611,n2612);
or (n2615,n2616,n2619);
and (n2616,n2617,n2618);
xor (n2617,n2568,n2569);
and (n2618,n476,n112);
and (n2619,n2620,n2621);
xor (n2620,n2617,n2618);
and (n2621,n2622,n2623);
xor (n2622,n2574,n2575);
and (n2623,n408,n112);
or (n2624,n2625,n2627);
and (n2625,n2626,n2588);
xor (n2626,n2584,n2585);
and (n2627,n2628,n2629);
xor (n2628,n2626,n2588);
or (n2629,n2630,n2632);
and (n2630,n2631,n2594);
xor (n2631,n2590,n2591);
and (n2632,n2633,n2634);
xor (n2633,n2631,n2594);
or (n2634,n2635,n2637);
and (n2635,n2636,n2600);
xor (n2636,n2596,n2597);
and (n2637,n2638,n2639);
xor (n2638,n2636,n2600);
or (n2639,n2640,n2642);
and (n2640,n2641,n2606);
xor (n2641,n2602,n2603);
and (n2642,n2643,n2644);
xor (n2643,n2641,n2606);
or (n2644,n2645,n2647);
and (n2645,n2646,n2612);
xor (n2646,n2608,n2609);
and (n2647,n2648,n2649);
xor (n2648,n2646,n2612);
or (n2649,n2650,n2652);
and (n2650,n2651,n2618);
xor (n2651,n2614,n2615);
and (n2652,n2653,n2654);
xor (n2653,n2651,n2618);
and (n2654,n2655,n2623);
xor (n2655,n2620,n2621);
or (n2656,n2657,n2659);
and (n2657,n2658,n2594);
xor (n2658,n2628,n2629);
and (n2659,n2660,n2661);
xor (n2660,n2658,n2594);
or (n2661,n2662,n2664);
and (n2662,n2663,n2600);
xor (n2663,n2633,n2634);
and (n2664,n2665,n2666);
xor (n2665,n2663,n2600);
or (n2666,n2667,n2669);
and (n2667,n2668,n2606);
xor (n2668,n2638,n2639);
and (n2669,n2670,n2671);
xor (n2670,n2668,n2606);
or (n2671,n2672,n2674);
and (n2672,n2673,n2612);
xor (n2673,n2643,n2644);
and (n2674,n2675,n2676);
xor (n2675,n2673,n2612);
or (n2676,n2677,n2679);
and (n2677,n2678,n2618);
xor (n2678,n2648,n2649);
and (n2679,n2680,n2681);
xor (n2680,n2678,n2618);
and (n2681,n2682,n2623);
xor (n2682,n2653,n2654);
or (n2683,n2684,n2686);
and (n2684,n2685,n2600);
xor (n2685,n2660,n2661);
and (n2686,n2687,n2688);
xor (n2687,n2685,n2600);
or (n2688,n2689,n2691);
and (n2689,n2690,n2606);
xor (n2690,n2665,n2666);
and (n2691,n2692,n2693);
xor (n2692,n2690,n2606);
or (n2693,n2694,n2696);
and (n2694,n2695,n2612);
xor (n2695,n2670,n2671);
and (n2696,n2697,n2698);
xor (n2697,n2695,n2612);
or (n2698,n2699,n2701);
and (n2699,n2700,n2618);
xor (n2700,n2675,n2676);
and (n2701,n2702,n2703);
xor (n2702,n2700,n2618);
and (n2703,n2704,n2623);
xor (n2704,n2680,n2681);
or (n2705,n2706,n2708);
and (n2706,n2707,n2606);
xor (n2707,n2687,n2688);
and (n2708,n2709,n2710);
xor (n2709,n2707,n2606);
or (n2710,n2711,n2713);
and (n2711,n2712,n2612);
xor (n2712,n2692,n2693);
and (n2713,n2714,n2715);
xor (n2714,n2712,n2612);
or (n2715,n2716,n2718);
and (n2716,n2717,n2618);
xor (n2717,n2697,n2698);
and (n2718,n2719,n2720);
xor (n2719,n2717,n2618);
and (n2720,n2721,n2623);
xor (n2721,n2702,n2703);
or (n2722,n2723,n2725);
and (n2723,n2724,n2612);
xor (n2724,n2709,n2710);
and (n2725,n2726,n2727);
xor (n2726,n2724,n2612);
or (n2727,n2728,n2730);
and (n2728,n2729,n2618);
xor (n2729,n2714,n2715);
and (n2730,n2731,n2732);
xor (n2731,n2729,n2618);
and (n2732,n2733,n2623);
xor (n2733,n2719,n2720);
or (n2734,n2735,n2737);
and (n2735,n2736,n2618);
xor (n2736,n2726,n2727);
and (n2737,n2738,n2739);
xor (n2738,n2736,n2618);
and (n2739,n2740,n2623);
xor (n2740,n2731,n2732);
and (n2741,n2742,n2623);
xor (n2742,n2738,n2739);
endmodule
