module top (out,n9,n10,n12,n13,n16,n17,n24,n26,n27
        ,n31,n38,n42,n60,n65,n126,n128,n131,n139,n143
        ,n153,n171);
output out;
input n9;
input n10;
input n12;
input n13;
input n16;
input n17;
input n24;
input n26;
input n27;
input n31;
input n38;
input n42;
input n60;
input n65;
input n126;
input n128;
input n131;
input n139;
input n143;
input n153;
input n171;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n11;
wire n14;
wire n15;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n25;
wire n28;
wire n29;
wire n30;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n39;
wire n40;
wire n41;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n61;
wire n62;
wire n63;
wire n64;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n127;
wire n129;
wire n130;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n140;
wire n141;
wire n142;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
xor (out,n0,n265);
xor (n0,n1,n228);
xor (n1,n2,n119);
xor (n2,n3,n91);
xor (n3,n4,n66);
xor (n4,n5,n44);
xor (n5,n6,n19);
or (n6,n7,n14,n18);
and (n7,n8,n11);
and (n8,n9,n10);
and (n11,n12,n13);
and (n14,n11,n15);
and (n15,n16,n17);
and (n18,n8,n15);
or (n19,n20,n35,n43);
and (n20,n21,n33);
or (n21,n22,n28,n32);
and (n22,n23,n25);
and (n23,n16,n24);
and (n25,n26,n27);
and (n28,n29,n30);
and (n29,n26,n24);
and (n30,n31,n27);
and (n32,n22,n30);
xor (n33,n34,n15);
xor (n34,n8,n11);
and (n35,n33,n36);
xor (n36,n37,n39);
and (n37,n26,n38);
xor (n39,n40,n41);
and (n40,n31,n24);
and (n41,n42,n27);
and (n43,n21,n36);
xor (n44,n45,n61);
xor (n45,n46,n47);
and (n46,n37,n39);
xor (n47,n48,n55);
xor (n48,n49,n50);
and (n49,n40,n41);
xor (n50,n51,n54);
xor (n51,n52,n53);
and (n52,n12,n10);
and (n53,n16,n13);
and (n54,n26,n17);
xor (n55,n56,n59);
xor (n56,n57,n58);
and (n57,n31,n38);
and (n58,n42,n24);
and (n59,n60,n27);
nor (n61,n62,n63);
not (n62,n9);
and (n63,n64,n9);
not (n64,n65);
or (n66,n67,n87,n90);
and (n67,n68,n71);
and (n68,n69,n70);
and (n69,n12,n17);
and (n70,n16,n38);
or (n71,n72,n83,n86);
and (n72,n73,n82);
or (n73,n74,n79,n81);
and (n74,n75,n78);
and (n75,n76,n77);
and (n76,n12,n24);
and (n77,n16,n27);
and (n78,n12,n38);
and (n79,n78,n80);
xor (n80,n23,n25);
and (n81,n75,n80);
xor (n82,n69,n70);
and (n83,n82,n84);
xor (n84,n85,n30);
xor (n85,n22,n29);
and (n86,n73,n84);
and (n87,n71,n88);
xor (n88,n89,n36);
xor (n89,n21,n33);
and (n90,n68,n88);
or (n91,n92,n114);
and (n92,n93,n95);
xor (n93,n94,n88);
xor (n94,n68,n71);
and (n95,n96,n112);
or (n96,n97,n108,n111);
and (n97,n98,n107);
or (n98,n99,n104,n106);
and (n99,n100,n103);
and (n100,n101,n102);
and (n101,n9,n24);
and (n102,n12,n27);
and (n103,n9,n38);
and (n104,n103,n105);
xor (n105,n76,n77);
and (n106,n100,n105);
and (n107,n9,n17);
and (n108,n107,n109);
xor (n109,n110,n80);
xor (n110,n75,n78);
and (n111,n98,n109);
xor (n112,n113,n84);
xor (n113,n73,n82);
and (n114,n115,n116);
xor (n115,n93,n95);
and (n116,n117,n118);
and (n117,n9,n13);
xor (n118,n96,n112);
xor (n119,n120,n200);
xor (n120,n121,n175);
xor (n121,n122,n155);
xor (n122,n123,n133);
or (n123,n124,n129,n132);
and (n124,n125,n127);
and (n125,n126,n10);
and (n127,n128,n13);
and (n129,n127,n130);
and (n130,n131,n17);
and (n132,n125,n130);
or (n133,n134,n147,n154);
and (n134,n135,n145);
or (n135,n136,n140,n144);
and (n136,n137,n138);
and (n137,n131,n24);
and (n138,n139,n27);
and (n140,n141,n142);
and (n141,n139,n24);
and (n142,n143,n27);
and (n144,n136,n142);
xor (n145,n146,n130);
xor (n146,n125,n127);
and (n147,n145,n148);
xor (n148,n149,n150);
and (n149,n139,n38);
xor (n150,n151,n152);
and (n151,n143,n24);
and (n152,n153,n27);
and (n154,n135,n148);
xor (n155,n156,n172);
xor (n156,n157,n158);
and (n157,n149,n150);
xor (n158,n159,n166);
xor (n159,n160,n161);
and (n160,n151,n152);
xor (n161,n162,n165);
xor (n162,n163,n164);
and (n163,n128,n10);
and (n164,n131,n13);
and (n165,n139,n17);
xor (n166,n167,n170);
xor (n167,n168,n169);
and (n168,n143,n38);
and (n169,n153,n24);
and (n170,n171,n27);
nor (n172,n173,n174);
not (n173,n126);
and (n174,n64,n126);
or (n175,n176,n196,n199);
and (n176,n177,n180);
and (n177,n178,n179);
and (n178,n128,n17);
and (n179,n131,n38);
or (n180,n181,n192,n195);
and (n181,n182,n191);
or (n182,n183,n188,n190);
and (n183,n184,n187);
and (n184,n185,n186);
and (n185,n128,n24);
and (n186,n131,n27);
and (n187,n128,n38);
and (n188,n187,n189);
xor (n189,n137,n138);
and (n190,n184,n189);
xor (n191,n178,n179);
and (n192,n191,n193);
xor (n193,n194,n142);
xor (n194,n136,n141);
and (n195,n182,n193);
and (n196,n180,n197);
xor (n197,n198,n148);
xor (n198,n135,n145);
and (n199,n177,n197);
or (n200,n201,n223);
and (n201,n202,n204);
xor (n202,n203,n197);
xor (n203,n177,n180);
and (n204,n205,n221);
or (n205,n206,n217,n220);
and (n206,n207,n216);
or (n207,n208,n213,n215);
and (n208,n209,n212);
and (n209,n210,n211);
and (n210,n126,n24);
and (n211,n128,n27);
and (n212,n126,n38);
and (n213,n212,n214);
xor (n214,n185,n186);
and (n215,n209,n214);
and (n216,n126,n17);
and (n217,n216,n218);
xor (n218,n219,n189);
xor (n219,n184,n187);
and (n220,n207,n218);
xor (n221,n222,n193);
xor (n222,n182,n191);
and (n223,n224,n225);
xor (n224,n202,n204);
and (n225,n226,n227);
and (n226,n126,n13);
xor (n227,n205,n221);
or (n228,n229,n232,n264);
and (n229,n230,n231);
xor (n230,n115,n116);
xor (n231,n224,n225);
and (n232,n231,n233);
or (n233,n234,n237,n263);
and (n234,n235,n236);
xor (n235,n117,n118);
xor (n236,n226,n227);
and (n237,n236,n238);
or (n238,n239,n244,n262);
and (n239,n240,n242);
xor (n240,n241,n109);
xor (n241,n98,n107);
xor (n242,n243,n218);
xor (n243,n207,n216);
and (n244,n242,n245);
or (n245,n246,n251,n261);
and (n246,n247,n249);
xor (n247,n248,n105);
xor (n248,n100,n103);
xor (n249,n250,n214);
xor (n250,n209,n212);
and (n251,n249,n252);
or (n252,n253,n256,n260);
and (n253,n254,n255);
xor (n254,n101,n102);
xor (n255,n210,n211);
and (n256,n255,n257);
and (n257,n258,n259);
and (n258,n9,n27);
and (n259,n126,n27);
and (n260,n254,n257);
and (n261,n247,n252);
and (n262,n240,n245);
and (n263,n235,n238);
and (n264,n230,n233);
xor (n265,n266,n373);
xor (n266,n267,n348);
xor (n267,n268,n323);
xor (n268,n269,n286);
or (n269,n270,n277,n285);
and (n270,n271,n273);
and (n271,n272,n10);
xor (n272,n9,n126);
and (n273,n274,n13);
xor (n274,n275,n276);
xor (n275,n12,n128);
and (n276,n9,n126);
and (n277,n273,n278);
and (n278,n279,n17);
xor (n279,n280,n281);
xor (n280,n16,n131);
or (n281,n282,n283,n284);
and (n282,n12,n128);
and (n283,n128,n276);
and (n284,n12,n276);
and (n285,n271,n278);
or (n286,n287,n310,n322);
and (n287,n288,n308);
or (n288,n289,n298,n307);
and (n289,n290,n291);
and (n290,n279,n24);
and (n291,n292,n27);
xor (n292,n293,n294);
xor (n293,n26,n139);
or (n294,n295,n296,n297);
and (n295,n16,n131);
and (n296,n131,n281);
and (n297,n16,n281);
and (n298,n299,n300);
and (n299,n292,n24);
and (n300,n301,n27);
xor (n301,n302,n303);
xor (n302,n31,n143);
or (n303,n304,n305,n306);
and (n304,n26,n139);
and (n305,n139,n294);
and (n306,n26,n294);
and (n307,n289,n300);
xor (n308,n309,n278);
xor (n309,n271,n273);
and (n310,n308,n311);
xor (n311,n312,n313);
and (n312,n292,n38);
xor (n313,n314,n315);
and (n314,n301,n24);
and (n315,n316,n27);
xor (n316,n317,n318);
xor (n317,n42,n153);
or (n318,n319,n320,n321);
and (n319,n31,n143);
and (n320,n143,n303);
and (n321,n31,n303);
and (n322,n288,n311);
xor (n323,n324,n343);
xor (n324,n325,n326);
and (n325,n312,n313);
xor (n326,n327,n334);
xor (n327,n328,n329);
and (n328,n314,n315);
xor (n329,n330,n333);
xor (n330,n331,n332);
and (n331,n279,n13);
and (n332,n292,n17);
and (n333,n301,n38);
xor (n334,n335,n336);
and (n335,n316,n24);
and (n336,n337,n27);
xor (n337,n338,n339);
xor (n338,n60,n171);
or (n339,n340,n341,n342);
and (n340,n42,n153);
and (n341,n153,n318);
and (n342,n42,n318);
xor (n343,n344,n347);
nor (n344,n345,n346);
not (n345,n272);
and (n346,n64,n272);
and (n347,n274,n10);
or (n348,n349,n369,n372);
and (n349,n350,n353);
and (n350,n351,n352);
and (n351,n274,n17);
and (n352,n279,n38);
or (n353,n354,n365,n368);
and (n354,n355,n364);
or (n355,n356,n361,n363);
and (n356,n357,n360);
and (n357,n358,n359);
and (n358,n274,n24);
and (n359,n279,n27);
and (n360,n274,n38);
and (n361,n360,n362);
xor (n362,n290,n291);
and (n363,n357,n362);
xor (n364,n351,n352);
and (n365,n364,n366);
xor (n366,n367,n300);
xor (n367,n289,n299);
and (n368,n355,n366);
and (n369,n353,n370);
xor (n370,n371,n311);
xor (n371,n288,n308);
and (n372,n350,n370);
or (n373,n374,n396);
and (n374,n375,n377);
xor (n375,n376,n370);
xor (n376,n350,n353);
and (n377,n378,n394);
or (n378,n379,n390,n393);
and (n379,n380,n389);
or (n380,n381,n386,n388);
and (n381,n382,n385);
and (n382,n383,n384);
and (n383,n272,n24);
and (n384,n274,n27);
and (n385,n272,n38);
and (n386,n385,n387);
xor (n387,n358,n359);
and (n388,n382,n387);
and (n389,n272,n17);
and (n390,n389,n391);
xor (n391,n392,n362);
xor (n392,n357,n360);
and (n393,n380,n391);
xor (n394,n395,n366);
xor (n395,n355,n364);
and (n396,n397,n398);
xor (n397,n375,n377);
and (n398,n399,n400);
and (n399,n272,n13);
xor (n400,n378,n394);
endmodule
