module top (out,n20,n25,n26,n27,n29,n30,n41,n44,n47
        ,n50,n52,n55,n58,n69,n79,n84,n87,n90,n93
        ,n96,n99,n102,n105,n108,n110,n112,n120,n135,n140
        ,n143,n146,n149,n152,n156,n166,n196,n201,n253,n258
        ,n261,n270,n414,n428,n741,n754);
output out;
input n20;
input n25;
input n26;
input n27;
input n29;
input n30;
input n41;
input n44;
input n47;
input n50;
input n52;
input n55;
input n58;
input n69;
input n79;
input n84;
input n87;
input n90;
input n93;
input n96;
input n99;
input n102;
input n105;
input n108;
input n110;
input n112;
input n120;
input n135;
input n140;
input n143;
input n146;
input n149;
input n152;
input n156;
input n166;
input n196;
input n201;
input n253;
input n258;
input n261;
input n270;
input n414;
input n428;
input n741;
input n754;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n21;
wire n22;
wire n23;
wire n24;
wire n28;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n42;
wire n43;
wire n45;
wire n46;
wire n48;
wire n49;
wire n51;
wire n53;
wire n54;
wire n56;
wire n57;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n80;
wire n81;
wire n82;
wire n83;
wire n85;
wire n86;
wire n88;
wire n89;
wire n91;
wire n92;
wire n94;
wire n95;
wire n97;
wire n98;
wire n100;
wire n101;
wire n103;
wire n104;
wire n106;
wire n107;
wire n109;
wire n111;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n136;
wire n137;
wire n138;
wire n139;
wire n141;
wire n142;
wire n144;
wire n145;
wire n147;
wire n148;
wire n150;
wire n151;
wire n153;
wire n154;
wire n155;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n197;
wire n198;
wire n199;
wire n200;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n254;
wire n255;
wire n256;
wire n257;
wire n259;
wire n260;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
xor (out,n0,n1371);
nand (n0,n1,n1370);
or (n1,n2,n767);
not (n2,n3);
nor (n3,n4,n766);
and (n4,n5,n658);
or (n5,n6,n657);
and (n6,n7,n612);
xor (n7,n8,n434);
xor (n8,n9,n338);
xor (n9,n10,n226);
xor (n10,n11,n188);
xor (n11,n12,n126);
nand (n12,n13,n115);
or (n13,n14,n75);
nand (n14,n15,n65);
or (n15,n16,n62);
and (n16,n17,n56);
wire s0n17,s1n17,notn17;
or (n17,s0n17,s1n17);
not(notn17,n53);
and (s0n17,notn17,n18);
and (s1n17,n53,n37);
wire s0n18,s1n18,notn18;
or (n18,s0n18,s1n18);
not(notn18,n21);
and (s0n18,notn18,1'b0);
and (s1n18,n21,n20);
or (n21,n22,n33);
or (n22,n23,n31);
nor (n23,n24,n26,n27,n28,n30);
not (n24,n25);
not (n28,n29);
nor (n31,n25,n32,n27,n28,n30);
not (n32,n26);
or (n33,n34,n36);
and (n34,n24,n26,n27,n28,n35);
not (n35,n30);
nor (n36,n24,n32,n27,n28,n30);
xor (n37,n38,n39);
not (n38,n20);
and (n39,n40,n42);
not (n40,n41);
and (n42,n43,n45);
not (n43,n44);
and (n45,n46,n48);
not (n46,n47);
and (n48,n49,n51);
not (n49,n50);
not (n51,n52);
and (n53,n54,n55);
or (n54,n23,n34);
wire s0n56,s1n56,notn56;
or (n56,s0n56,s1n56);
not(notn56,n53);
and (s0n56,notn56,n57);
and (s1n56,n53,n59);
wire s0n57,s1n57,notn57;
or (n57,s0n57,s1n57);
not(notn57,n21);
and (s0n57,notn57,1'b0);
and (s1n57,n21,n58);
xor (n59,n60,n61);
not (n60,n58);
and (n61,n38,n39);
and (n62,n63,n64);
not (n63,n17);
not (n64,n56);
nor (n65,n66,n73);
and (n66,n67,n56);
wire s0n67,s1n67,notn67;
or (n67,s0n67,s1n67);
not(notn67,n53);
and (s0n67,notn67,n68);
and (s1n67,n53,n70);
wire s0n68,s1n68,notn68;
or (n68,s0n68,s1n68);
not(notn68,n21);
and (s0n68,notn68,1'b0);
and (s1n68,n21,n69);
xor (n70,n71,n72);
not (n71,n69);
and (n72,n60,n61);
and (n73,n74,n64);
not (n74,n67);
nor (n75,n76,n113);
and (n76,n77,n74);
wire s0n77,s1n77,notn77;
or (n77,s0n77,s1n77);
not(notn77,n111);
and (s0n77,notn77,n78);
and (s1n77,n111,n80);
wire s0n78,s1n78,notn78;
or (n78,s0n78,s1n78);
not(notn78,n21);
and (s0n78,notn78,1'b0);
and (s1n78,n21,n79);
xor (n80,n81,n82);
not (n81,n79);
and (n82,n83,n85);
not (n83,n84);
and (n85,n86,n88);
not (n86,n87);
and (n88,n89,n91);
not (n89,n90);
and (n91,n92,n94);
not (n92,n93);
and (n94,n95,n97);
not (n95,n96);
and (n97,n98,n100);
not (n98,n99);
and (n100,n101,n103);
not (n101,n102);
and (n103,n104,n106);
not (n104,n105);
and (n106,n107,n109);
not (n107,n108);
not (n109,n110);
and (n111,n54,n112);
and (n113,n114,n67);
not (n114,n77);
or (n115,n116,n15);
nor (n116,n117,n124);
and (n117,n118,n74);
wire s0n118,s1n118,notn118;
or (n118,s0n118,s1n118);
not(notn118,n111);
and (s0n118,notn118,n119);
and (s1n118,n111,n121);
wire s0n119,s1n119,notn119;
or (n119,s0n119,s1n119);
not(notn119,n21);
and (s0n119,notn119,1'b0);
and (s1n119,n21,n120);
xor (n121,n122,n123);
not (n122,n120);
and (n123,n81,n82);
and (n124,n125,n67);
not (n125,n118);
nand (n126,n127,n179);
or (n127,n128,n172);
not (n128,n129);
nor (n129,n130,n161);
nand (n130,n131,n160);
or (n131,n132,n154);
not (n132,n133);
wire s0n133,s1n133,notn133;
or (n133,s0n133,s1n133);
not(notn133,n53);
and (s0n133,notn133,n134);
and (s1n133,n53,n136);
wire s0n134,s1n134,notn134;
or (n134,s0n134,s1n134);
not(notn134,n21);
and (s0n134,notn134,1'b0);
and (s1n134,n21,n135);
xor (n136,n137,n138);
not (n137,n135);
and (n138,n139,n141);
not (n139,n140);
and (n141,n142,n144);
not (n142,n143);
and (n144,n145,n147);
not (n145,n146);
and (n147,n148,n150);
not (n148,n149);
and (n150,n151,n153);
not (n151,n152);
and (n153,n71,n72);
wire s0n154,s1n154,notn154;
or (n154,s0n154,s1n154);
not(notn154,n53);
and (s0n154,notn154,n155);
and (s1n154,n53,n157);
wire s0n155,s1n155,notn155;
or (n155,s0n155,s1n155);
not(notn155,n21);
and (s0n155,notn155,1'b0);
and (s1n155,n21,n156);
xor (n157,n158,n159);
not (n158,n156);
and (n159,n137,n138);
nand (n160,n132,n154);
nor (n161,n162,n170);
and (n162,n163,n154);
not (n163,n164);
wire s0n164,s1n164,notn164;
or (n164,s0n164,s1n164);
not(notn164,n53);
and (s0n164,notn164,n165);
and (s1n164,n53,n167);
wire s0n165,s1n165,notn165;
or (n165,s0n165,s1n165);
not(notn165,n21);
and (s0n165,notn165,1'b0);
and (s1n165,n21,n166);
xor (n167,n168,n169);
not (n168,n166);
and (n169,n158,n159);
and (n170,n171,n164);
not (n171,n154);
nor (n172,n173,n177);
and (n173,n174,n163);
wire s0n174,s1n174,notn174;
or (n174,s0n174,s1n174);
not(notn174,n111);
and (s0n174,notn174,n175);
and (s1n174,n111,n176);
wire s0n175,s1n175,notn175;
or (n175,s0n175,s1n175);
not(notn175,n21);
and (s0n175,notn175,1'b0);
and (s1n175,n21,n105);
xor (n176,n104,n106);
and (n177,n178,n164);
not (n178,n174);
or (n179,n180,n181);
not (n180,n130);
nor (n181,n182,n186);
and (n182,n183,n163);
wire s0n183,s1n183,notn183;
or (n183,s0n183,s1n183);
not(notn183,n111);
and (s0n183,notn183,n184);
and (s1n183,n111,n185);
wire s0n184,s1n184,notn184;
or (n184,s0n184,s1n184);
not(notn184,n21);
and (s0n184,notn184,1'b0);
and (s1n184,n21,n102);
xor (n185,n101,n103);
and (n186,n187,n164);
not (n187,n183);
nand (n188,n189,n218);
or (n189,n190,n206);
not (n190,n191);
nand (n191,n192,n204);
or (n192,n193,n203);
not (n193,n194);
wire s0n194,s1n194,notn194;
or (n194,s0n194,s1n194);
not(notn194,n53);
and (s0n194,notn194,n195);
and (s1n194,n53,n197);
wire s0n195,s1n195,notn195;
or (n195,s0n195,s1n195);
not(notn195,n21);
and (s0n195,notn195,1'b0);
and (s1n195,n21,n196);
xor (n197,n198,n199);
not (n198,n196);
and (n199,n200,n202);
not (n200,n201);
and (n202,n168,n169);
wire s0n203,s1n203,notn203;
or (n203,s0n203,s1n203);
not(notn203,n21);
and (s0n203,notn203,1'b0);
and (s1n203,n21,n110);
or (n204,n194,n205);
not (n205,n203);
not (n206,n207);
and (n207,n208,n215);
nor (n208,n209,n214);
and (n209,n164,n210);
not (n210,n211);
wire s0n211,s1n211,notn211;
or (n211,s0n211,s1n211);
not(notn211,n53);
and (s0n211,notn211,n212);
and (s1n211,n53,n213);
wire s0n212,s1n212,notn212;
or (n212,s0n212,s1n212);
not(notn212,n21);
and (s0n212,notn212,1'b0);
and (s1n212,n21,n201);
xor (n213,n200,n202);
and (n214,n163,n211);
nand (n215,n216,n217);
or (n216,n210,n194);
or (n217,n193,n211);
or (n218,n219,n208);
nor (n219,n220,n224);
and (n220,n221,n193);
wire s0n221,s1n221,notn221;
or (n221,s0n221,s1n221);
not(notn221,n111);
and (s0n221,notn221,n222);
and (s1n221,n111,n223);
wire s0n222,s1n222,notn222;
or (n222,s0n222,s1n222);
not(notn222,n21);
and (s0n222,notn222,1'b0);
and (s1n222,n21,n108);
xor (n223,n107,n109);
and (n224,n225,n194);
not (n225,n221);
xor (n226,n227,n309);
xor (n227,n228,n276);
nand (n228,n229,n265);
or (n229,n230,n249);
nand (n230,n231,n242);
nor (n231,n232,n240);
and (n232,n233,n237);
not (n233,n234);
wire s0n234,s1n234,notn234;
or (n234,s0n234,s1n234);
not(notn234,n53);
and (s0n234,notn234,n235);
and (s1n234,n53,n236);
wire s0n235,s1n235,notn235;
or (n235,s0n235,s1n235);
not(notn235,n21);
and (s0n235,notn235,1'b0);
and (s1n235,n21,n50);
xor (n236,n49,n51);
wire s0n237,s1n237,notn237;
or (n237,s0n237,s1n237);
not(notn237,n53);
and (s0n237,notn237,n238);
and (s1n237,n53,n239);
wire s0n238,s1n238,notn238;
or (n238,s0n238,s1n238);
not(notn238,n21);
and (s0n238,notn238,1'b0);
and (s1n238,n21,n47);
xor (n239,n46,n48);
and (n240,n234,n241);
not (n241,n237);
nand (n242,n243,n248);
or (n243,n244,n237);
not (n244,n245);
wire s0n245,s1n245,notn245;
or (n245,s0n245,s1n245);
not(notn245,n53);
and (s0n245,notn245,n246);
and (s1n245,n53,n247);
wire s0n246,s1n246,notn246;
or (n246,s0n246,s1n246);
not(notn246,n21);
and (s0n246,notn246,1'b0);
and (s1n246,n21,n44);
xor (n247,n43,n45);
nand (n248,n244,n237);
nor (n249,n250,n263);
and (n250,n244,n251);
wire s0n251,s1n251,notn251;
or (n251,s0n251,s1n251);
not(notn251,n111);
and (s0n251,notn251,n252);
and (s1n251,n111,n254);
wire s0n252,s1n252,notn252;
or (n252,s0n252,s1n252);
not(notn252,n21);
and (s0n252,notn252,1'b0);
and (s1n252,n21,n253);
xor (n254,n255,n256);
not (n255,n253);
and (n256,n257,n259);
not (n257,n258);
and (n259,n260,n262);
not (n260,n261);
and (n262,n122,n123);
and (n263,n264,n245);
not (n264,n251);
or (n265,n231,n266);
nor (n266,n267,n274);
and (n267,n244,n268);
wire s0n268,s1n268,notn268;
or (n268,s0n268,s1n268);
not(notn268,n111);
and (s0n268,notn268,n269);
and (s1n268,n111,n271);
wire s0n269,s1n269,notn269;
or (n269,s0n269,s1n269);
not(notn269,n21);
and (s0n269,notn269,1'b0);
and (s1n269,n21,n270);
xor (n271,n272,n273);
not (n272,n270);
and (n273,n255,n256);
and (n274,n275,n245);
not (n275,n268);
nand (n276,n277,n301);
or (n277,n278,n294);
nand (n278,n279,n290);
nor (n279,n280,n287);
and (n280,n281,n284);
wire s0n281,s1n281,notn281;
or (n281,s0n281,s1n281);
not(notn281,n53);
and (s0n281,notn281,n282);
and (s1n281,n53,n283);
wire s0n282,s1n282,notn282;
or (n282,s0n282,s1n282);
not(notn282,n21);
and (s0n282,notn282,1'b0);
and (s1n282,n21,n152);
xor (n283,n151,n153);
wire s0n284,s1n284,notn284;
or (n284,s0n284,s1n284);
not(notn284,n53);
and (s0n284,notn284,n285);
and (s1n284,n53,n286);
wire s0n285,s1n285,notn285;
or (n285,s0n285,s1n285);
not(notn285,n21);
and (s0n285,notn285,1'b0);
and (s1n285,n21,n149);
xor (n286,n148,n150);
and (n287,n288,n289);
not (n288,n281);
not (n289,n284);
not (n290,n291);
nor (n291,n292,n293);
and (n292,n67,n281);
and (n293,n74,n288);
nor (n294,n295,n299);
and (n295,n289,n296);
wire s0n296,s1n296,notn296;
or (n296,s0n296,s1n296);
not(notn296,n111);
and (s0n296,notn296,n297);
and (s1n296,n111,n298);
wire s0n297,s1n297,notn297;
or (n297,s0n297,s1n297);
not(notn297,n21);
and (s0n297,notn297,1'b0);
and (s1n297,n21,n87);
xor (n298,n86,n88);
and (n299,n284,n300);
not (n300,n296);
or (n301,n302,n290);
nor (n302,n303,n307);
and (n303,n289,n304);
wire s0n304,s1n304,notn304;
or (n304,s0n304,s1n304);
not(notn304,n111);
and (s0n304,notn304,n305);
and (s1n304,n111,n306);
wire s0n305,s1n305,notn305;
or (n305,s0n305,s1n305);
not(notn305,n21);
and (s0n305,notn305,1'b0);
and (s1n305,n21,n84);
xor (n306,n83,n85);
and (n307,n284,n308);
not (n308,n304);
nand (n309,n310,n330);
or (n310,n311,n318);
nor (n311,n312,n316);
and (n312,n313,n63);
wire s0n313,s1n313,notn313;
or (n313,s0n313,s1n313);
not(notn313,n111);
and (s0n313,notn313,n314);
and (s1n313,n111,n315);
wire s0n314,s1n314,notn314;
or (n314,s0n314,s1n314);
not(notn314,n21);
and (s0n314,notn314,1'b0);
and (s1n314,n21,n261);
xor (n315,n260,n262);
and (n316,n317,n17);
not (n317,n313);
nand (n318,n319,n326);
not (n319,n320);
nand (n320,n321,n325);
or (n321,n244,n322);
wire s0n322,s1n322,notn322;
or (n322,s0n322,s1n322);
not(notn322,n53);
and (s0n322,notn322,n323);
and (s1n322,n53,n324);
wire s0n323,s1n323,notn323;
or (n323,s0n323,s1n323);
not(notn323,n21);
and (s0n323,notn323,1'b0);
and (s1n323,n21,n41);
xor (n324,n40,n42);
nand (n325,n322,n244);
nor (n326,n327,n329);
and (n327,n63,n328);
not (n328,n322);
and (n329,n17,n322);
or (n330,n319,n331);
nor (n331,n332,n336);
and (n332,n333,n63);
wire s0n333,s1n333,notn333;
or (n333,s0n333,s1n333);
not(notn333,n111);
and (s0n333,notn333,n334);
and (s1n333,n111,n335);
wire s0n334,s1n334,notn334;
or (n334,s0n334,s1n334);
not(notn334,n21);
and (s0n334,notn334,1'b0);
and (s1n334,n21,n258);
xor (n335,n257,n259);
and (n336,n337,n17);
not (n337,n333);
xor (n338,n339,n401);
xor (n339,n340,n372);
nand (n340,n341,n364);
or (n341,n342,n357);
nand (n342,n343,n350);
or (n343,n344,n348);
and (n344,n345,n284);
wire s0n345,s1n345,notn345;
or (n345,s0n345,s1n345);
not(notn345,n53);
and (s0n345,notn345,n346);
and (s1n345,n53,n347);
wire s0n346,s1n346,notn346;
or (n346,s0n346,s1n346);
not(notn346,n21);
and (s0n346,notn346,1'b0);
and (s1n346,n21,n146);
xor (n347,n145,n147);
and (n348,n349,n289);
not (n349,n345);
nand (n350,n351,n355);
or (n351,n349,n352);
wire s0n352,s1n352,notn352;
or (n352,s0n352,s1n352);
not(notn352,n53);
and (s0n352,notn352,n353);
and (s1n352,n53,n354);
wire s0n353,s1n353,notn353;
or (n353,s0n353,s1n353);
not(notn353,n21);
and (s0n353,notn353,1'b0);
and (s1n353,n21,n143);
xor (n354,n142,n144);
or (n355,n356,n345);
not (n356,n352);
nor (n357,n358,n362);
and (n358,n356,n359);
wire s0n359,s1n359,notn359;
or (n359,s0n359,s1n359);
not(notn359,n111);
and (s0n359,notn359,n360);
and (s1n359,n111,n361);
wire s0n360,s1n360,notn360;
or (n360,s0n360,s1n360);
not(notn360,n21);
and (s0n360,notn360,1'b0);
and (s1n360,n21,n93);
xor (n361,n92,n94);
and (n362,n352,n363);
not (n363,n359);
or (n364,n365,n343);
nor (n365,n366,n370);
and (n366,n356,n367);
wire s0n367,s1n367,notn367;
or (n367,s0n367,s1n367);
not(notn367,n111);
and (s0n367,notn367,n368);
and (s1n367,n111,n369);
wire s0n368,s1n368,notn368;
or (n368,s0n368,s1n368);
not(notn368,n21);
and (s0n368,notn368,1'b0);
and (s1n368,n21,n90);
xor (n369,n89,n91);
and (n370,n352,n371);
not (n371,n367);
nand (n372,n373,n392);
or (n373,n374,n385);
or (n374,n375,n382);
nor (n375,n376,n380);
and (n376,n132,n377);
wire s0n377,s1n377,notn377;
or (n377,s0n377,s1n377);
not(notn377,n53);
and (s0n377,notn377,n378);
and (s1n377,n53,n379);
wire s0n378,s1n378,notn378;
or (n378,s0n378,s1n378);
not(notn378,n21);
and (s0n378,notn378,1'b0);
and (s1n378,n21,n140);
xor (n379,n139,n141);
and (n380,n381,n133);
not (n381,n377);
nor (n382,n383,n384);
and (n383,n377,n352);
and (n384,n381,n356);
nor (n385,n386,n390);
and (n386,n132,n387);
wire s0n387,s1n387,notn387;
or (n387,s0n387,s1n387);
not(notn387,n111);
and (s0n387,notn387,n388);
and (s1n387,n111,n389);
wire s0n388,s1n388,notn388;
or (n388,s0n388,s1n388);
not(notn388,n21);
and (s0n388,notn388,1'b0);
and (s1n388,n21,n99);
xor (n389,n98,n100);
and (n390,n391,n133);
not (n391,n387);
or (n392,n393,n394);
not (n393,n382);
nor (n394,n395,n399);
and (n395,n132,n396);
wire s0n396,s1n396,notn396;
or (n396,s0n396,s1n396);
not(notn396,n111);
and (s0n396,notn396,n397);
and (s1n396,n111,n398);
wire s0n397,s1n397,notn397;
or (n397,s0n397,s1n397);
not(notn397,n21);
and (s0n397,notn397,1'b0);
and (s1n397,n21,n96);
xor (n398,n95,n97);
and (n399,n133,n400);
not (n400,n396);
xor (n401,n402,n408);
nor (n402,n403,n193);
nor (n403,n404,n407);
and (n404,n163,n405);
not (n405,n406);
and (n406,n203,n211);
and (n407,n210,n205);
nand (n408,n409,n423);
or (n409,n410,n420);
nor (n410,n411,n418);
and (n411,n412,n233);
wire s0n412,s1n412,notn412;
or (n412,s0n412,s1n412);
not(notn412,n111);
and (s0n412,notn412,n413);
and (s1n412,n111,n415);
wire s0n413,s1n413,notn413;
or (n413,s0n413,s1n413);
not(notn413,n21);
and (s0n413,notn413,1'b0);
and (s1n413,n21,n414);
xor (n415,n416,n417);
not (n416,n414);
and (n417,n272,n273);
and (n418,n419,n234);
not (n419,n412);
nand (n420,n234,n421);
not (n421,n422);
wire s0n422,s1n422,notn422;
or (n422,s0n422,s1n422);
not(notn422,n21);
and (s0n422,notn422,1'b0);
and (s1n422,n21,n52);
or (n423,n424,n421);
nor (n424,n425,n432);
and (n425,n426,n233);
wire s0n426,s1n426,notn426;
or (n426,s0n426,s1n426);
not(notn426,n111);
and (s0n426,notn426,n427);
and (s1n426,n111,n429);
wire s0n427,s1n427,notn427;
or (n427,s0n427,s1n427);
not(notn427,n21);
and (s0n427,notn427,1'b0);
and (s1n427,n21,n428);
xor (n429,n430,n431);
not (n430,n428);
and (n431,n416,n417);
and (n432,n433,n234);
not (n433,n426);
or (n434,n435,n611);
and (n435,n436,n574);
xor (n436,n437,n486);
or (n437,n438,n485);
and (n438,n439,n465);
xor (n439,n440,n449);
nand (n440,n441,n445);
or (n441,n374,n442);
nor (n442,n443,n444);
and (n443,n174,n132);
and (n444,n178,n133);
or (n445,n446,n393);
nor (n446,n447,n448);
and (n447,n183,n132);
and (n448,n187,n133);
xor (n449,n450,n459);
nand (n450,n451,n455);
or (n451,n452,n420);
nor (n452,n453,n454);
and (n453,n251,n233);
and (n454,n264,n234);
or (n455,n456,n421);
nor (n456,n457,n458);
and (n457,n268,n233);
and (n458,n275,n234);
nor (n459,n460,n163);
nor (n460,n461,n464);
and (n461,n132,n462);
not (n462,n463);
and (n463,n203,n154);
and (n464,n171,n205);
or (n465,n466,n484);
and (n466,n467,n475);
xor (n467,n468,n469);
nor (n468,n180,n205);
nand (n469,n470,n474);
or (n470,n471,n420);
nor (n471,n472,n473);
and (n472,n233,n333);
and (n473,n337,n234);
or (n474,n452,n421);
nand (n475,n476,n480);
or (n476,n230,n477);
nor (n477,n478,n479);
and (n478,n244,n118);
and (n479,n125,n245);
or (n480,n231,n481);
nor (n481,n482,n483);
and (n482,n313,n244);
and (n483,n317,n245);
and (n484,n468,n469);
and (n485,n440,n449);
or (n486,n487,n573);
and (n487,n488,n552);
xor (n488,n489,n520);
or (n489,n490,n519);
and (n490,n491,n510);
xor (n491,n492,n501);
nand (n492,n493,n497);
or (n493,n14,n494);
nor (n494,n495,n496);
and (n495,n367,n74);
and (n496,n371,n67);
or (n497,n498,n15);
nor (n498,n499,n500);
and (n499,n296,n74);
and (n500,n300,n67);
nand (n501,n502,n506);
or (n502,n278,n503);
nor (n503,n504,n505);
and (n504,n289,n396);
and (n505,n284,n400);
or (n506,n507,n290);
nor (n507,n508,n509);
and (n508,n289,n359);
and (n509,n284,n363);
nand (n510,n511,n515);
or (n511,n319,n512);
nor (n512,n513,n514);
and (n513,n77,n63);
and (n514,n114,n17);
or (n515,n318,n516);
nor (n516,n517,n518);
and (n517,n304,n63);
and (n518,n308,n17);
and (n519,n492,n501);
or (n520,n521,n551);
and (n521,n522,n538);
xor (n522,n523,n532);
nand (n523,n524,n528);
or (n524,n342,n525);
nor (n525,n526,n527);
and (n526,n183,n356);
and (n527,n187,n352);
or (n528,n529,n343);
nor (n529,n530,n531);
and (n530,n356,n387);
and (n531,n352,n391);
nand (n532,n533,n537);
or (n533,n374,n534);
nor (n534,n535,n536);
and (n535,n221,n132);
and (n536,n225,n133);
or (n537,n442,n393);
and (n538,n539,n545);
nand (n539,n540,n544);
or (n540,n541,n420);
nor (n541,n542,n543);
and (n542,n233,n313);
and (n543,n317,n234);
or (n544,n471,n421);
nor (n545,n546,n132);
nor (n546,n547,n550);
and (n547,n356,n548);
not (n548,n549);
and (n549,n203,n377);
and (n550,n381,n205);
and (n551,n523,n532);
xor (n552,n553,n566);
xor (n553,n554,n560);
nand (n554,n555,n556);
or (n555,n278,n507);
or (n556,n557,n290);
nor (n557,n558,n559);
and (n558,n289,n367);
and (n559,n284,n371);
nand (n560,n561,n562);
or (n561,n318,n512);
or (n562,n319,n563);
nor (n563,n564,n565);
and (n564,n118,n63);
and (n565,n125,n17);
nand (n566,n567,n572);
or (n567,n343,n568);
not (n568,n569);
nand (n569,n570,n571);
or (n570,n400,n352);
or (n571,n356,n396);
or (n572,n342,n529);
and (n573,n489,n520);
xor (n574,n575,n589);
xor (n575,n576,n577);
and (n576,n450,n459);
xor (n577,n578,n583);
xor (n578,n579,n580);
nor (n579,n208,n205);
nand (n580,n581,n582);
or (n581,n456,n420);
or (n582,n410,n421);
nand (n583,n584,n588);
or (n584,n230,n585);
nor (n585,n586,n587);
and (n586,n244,n333);
and (n587,n337,n245);
or (n588,n231,n249);
or (n589,n590,n610);
and (n590,n591,n604);
xor (n591,n592,n595);
nand (n592,n593,n594);
or (n593,n230,n481);
or (n594,n231,n585);
nand (n595,n596,n600);
or (n596,n128,n597);
nor (n597,n598,n599);
and (n598,n164,n205);
and (n599,n163,n203);
or (n600,n601,n180);
nor (n601,n602,n603);
and (n602,n221,n163);
and (n603,n225,n164);
nand (n604,n605,n609);
or (n605,n606,n15);
nor (n606,n607,n608);
and (n607,n304,n74);
and (n608,n308,n67);
or (n609,n14,n498);
and (n610,n592,n595);
and (n611,n437,n486);
xor (n612,n613,n648);
xor (n613,n614,n617);
or (n614,n615,n616);
and (n615,n575,n589);
and (n616,n576,n577);
xor (n617,n618,n635);
xor (n618,n619,n622);
or (n619,n620,n621);
and (n620,n578,n583);
and (n621,n579,n580);
or (n622,n623,n634);
and (n623,n624,n631);
xor (n624,n625,n628);
nand (n625,n626,n627);
or (n626,n318,n563);
or (n627,n319,n311);
nand (n628,n629,n630);
or (n629,n568,n342);
or (n630,n357,n343);
nand (n631,n632,n633);
or (n632,n374,n446);
or (n633,n385,n393);
and (n634,n625,n628);
or (n635,n636,n647);
and (n636,n637,n644);
xor (n637,n638,n641);
nand (n638,n639,n640);
or (n639,n128,n601);
or (n640,n172,n180);
nand (n641,n642,n643);
or (n642,n14,n606);
or (n643,n75,n15);
nand (n644,n645,n646);
or (n645,n278,n557);
or (n646,n294,n290);
and (n647,n638,n641);
or (n648,n649,n656);
and (n649,n650,n655);
xor (n650,n651,n654);
or (n651,n652,n653);
and (n652,n553,n566);
and (n653,n554,n560);
xor (n654,n624,n631);
xor (n655,n637,n644);
and (n656,n651,n654);
and (n657,n8,n434);
xor (n658,n659,n700);
xor (n659,n660,n697);
xor (n660,n661,n685);
xor (n661,n662,n682);
xor (n662,n663,n676);
xor (n663,n664,n670);
nand (n664,n665,n666);
or (n665,n128,n181);
or (n666,n667,n180);
nor (n667,n668,n669);
and (n668,n163,n387);
and (n669,n391,n164);
nand (n670,n671,n672);
or (n671,n206,n219);
or (n672,n673,n208);
nor (n673,n674,n675);
and (n674,n174,n193);
and (n675,n178,n194);
nand (n676,n677,n678);
or (n677,n230,n266);
or (n678,n231,n679);
nor (n679,n680,n681);
and (n680,n244,n412);
and (n681,n419,n245);
or (n682,n683,n684);
and (n683,n339,n401);
and (n684,n340,n372);
xor (n685,n686,n694);
xor (n686,n687,n693);
nand (n687,n688,n689);
or (n688,n374,n394);
or (n689,n690,n393);
nor (n690,n691,n692);
and (n691,n132,n359);
and (n692,n133,n363);
and (n693,n402,n408);
or (n694,n695,n696);
and (n695,n11,n188);
and (n696,n12,n126);
or (n697,n698,n699);
and (n698,n613,n648);
and (n699,n614,n617);
xor (n700,n701,n708);
xor (n701,n702,n705);
or (n702,n703,n704);
and (n703,n618,n635);
and (n704,n619,n622);
or (n705,n706,n707);
and (n706,n9,n338);
and (n707,n10,n226);
xor (n708,n709,n733);
xor (n709,n710,n713);
or (n710,n711,n712);
and (n711,n227,n309);
and (n712,n228,n276);
xor (n713,n714,n727);
xor (n714,n715,n721);
nand (n715,n716,n717);
or (n716,n278,n302);
or (n717,n718,n290);
nor (n718,n719,n720);
and (n719,n289,n77);
and (n720,n284,n114);
nand (n721,n722,n723);
or (n722,n318,n331);
or (n723,n319,n724);
nor (n724,n725,n726);
and (n725,n251,n63);
and (n726,n264,n17);
nand (n727,n728,n729);
or (n728,n342,n365);
or (n729,n343,n730);
nor (n730,n731,n732);
and (n731,n356,n296);
and (n732,n352,n300);
xor (n733,n734,n760);
xor (n734,n735,n747);
nor (n735,n736,n205);
not (n736,n737);
nor (n737,n738,n745);
and (n738,n739,n194);
wire s0n739,s1n739,notn739;
or (n739,s0n739,s1n739);
not(notn739,n53);
and (s0n739,notn739,n740);
and (s1n739,n53,n742);
wire s0n740,s1n740,notn740;
or (n740,s0n740,s1n740);
not(notn740,n21);
and (s0n740,notn740,1'b0);
and (s1n740,n21,n741);
xor (n742,n743,n744);
not (n743,n741);
and (n744,n198,n199);
and (n745,n746,n193);
not (n746,n739);
nand (n747,n748,n749);
or (n748,n424,n420);
or (n749,n750,n421);
nor (n750,n751,n758);
and (n751,n752,n233);
wire s0n752,s1n752,notn752;
or (n752,s0n752,s1n752);
not(notn752,n111);
and (s0n752,notn752,n753);
and (s1n752,n111,n755);
wire s0n753,s1n753,notn753;
or (n753,s0n753,s1n753);
not(notn753,n21);
and (s0n753,notn753,1'b0);
and (s1n753,n21,n754);
xor (n755,n756,n757);
not (n756,n754);
and (n757,n430,n431);
and (n758,n759,n234);
not (n759,n752);
nand (n760,n761,n765);
or (n761,n762,n15);
nor (n762,n763,n764);
and (n763,n313,n74);
and (n764,n317,n67);
or (n765,n14,n116);
nor (n766,n5,n658);
not (n767,n768);
nor (n768,n769,n1366);
not (n769,n770);
nand (n770,n771,n1349);
or (n771,n772,n1348);
and (n772,n773,n938);
xor (n773,n774,n925);
or (n774,n775,n924);
and (n775,n776,n873);
xor (n776,n777,n825);
xor (n777,n778,n803);
xor (n778,n779,n780);
xor (n779,n467,n475);
or (n780,n781,n802);
and (n781,n782,n795);
xor (n782,n783,n789);
nand (n783,n784,n788);
or (n784,n230,n785);
nor (n785,n786,n787);
and (n786,n244,n77);
and (n787,n114,n245);
or (n788,n231,n477);
nand (n789,n790,n794);
or (n790,n14,n791);
nor (n791,n792,n793);
and (n792,n359,n74);
and (n793,n363,n67);
or (n794,n15,n494);
nand (n795,n796,n801);
or (n796,n797,n278);
not (n797,n798);
nand (n798,n799,n800);
or (n799,n284,n391);
or (n800,n289,n387);
or (n801,n503,n290);
and (n802,n783,n789);
or (n803,n804,n824);
and (n804,n805,n818);
xor (n805,n806,n812);
nand (n806,n807,n811);
or (n807,n318,n808);
nor (n808,n809,n810);
and (n809,n296,n63);
and (n810,n300,n17);
or (n811,n516,n319);
nand (n812,n813,n817);
or (n813,n342,n814);
nor (n814,n815,n816);
and (n815,n174,n356);
and (n816,n178,n352);
or (n817,n525,n343);
nand (n818,n819,n820);
or (n819,n393,n534);
or (n820,n374,n821);
nor (n821,n822,n823);
and (n822,n133,n205);
and (n823,n132,n203);
and (n824,n806,n812);
xor (n825,n826,n829);
xor (n826,n827,n828);
xor (n827,n522,n538);
xor (n828,n491,n510);
or (n829,n830,n872);
and (n830,n831,n850);
xor (n831,n832,n833);
xor (n832,n539,n545);
or (n833,n834,n849);
and (n834,n835,n843);
xor (n835,n836,n837);
nor (n836,n393,n205);
nand (n837,n838,n842);
or (n838,n839,n420);
nor (n839,n840,n841);
and (n840,n233,n118);
and (n841,n125,n234);
or (n842,n541,n421);
nand (n843,n844,n845);
or (n844,n231,n785);
or (n845,n230,n846);
nor (n846,n847,n848);
and (n847,n304,n244);
and (n848,n308,n245);
and (n849,n836,n837);
or (n850,n851,n871);
and (n851,n852,n865);
xor (n852,n853,n859);
nand (n853,n854,n858);
or (n854,n14,n855);
nor (n855,n856,n857);
and (n856,n396,n74);
and (n857,n400,n67);
or (n858,n791,n15);
nand (n859,n860,n861);
or (n860,n290,n797);
or (n861,n278,n862);
nor (n862,n863,n864);
and (n863,n289,n183);
and (n864,n284,n187);
nand (n865,n866,n867);
or (n866,n343,n814);
or (n867,n342,n868);
nor (n868,n869,n870);
and (n869,n221,n356);
and (n870,n225,n352);
and (n871,n853,n859);
and (n872,n832,n833);
or (n873,n874,n923);
and (n874,n875,n878);
xor (n875,n876,n877);
xor (n876,n805,n818);
xor (n877,n782,n795);
or (n878,n879,n922);
and (n879,n880,n900);
xor (n880,n881,n887);
nand (n881,n882,n886);
or (n882,n318,n883);
nor (n883,n884,n885);
and (n884,n367,n63);
and (n885,n371,n17);
or (n886,n319,n808);
and (n887,n888,n894);
nand (n888,n889,n893);
or (n889,n890,n420);
nor (n890,n891,n892);
and (n891,n77,n233);
and (n892,n114,n234);
or (n893,n839,n421);
nor (n894,n895,n356);
nor (n895,n896,n899);
and (n896,n289,n897);
not (n897,n898);
and (n898,n203,n345);
and (n899,n349,n205);
or (n900,n901,n921);
and (n901,n902,n915);
xor (n902,n903,n909);
nand (n903,n904,n908);
or (n904,n230,n905);
nor (n905,n906,n907);
and (n906,n296,n244);
and (n907,n300,n245);
or (n908,n231,n846);
nand (n909,n910,n914);
or (n910,n14,n911);
nor (n911,n912,n913);
and (n912,n387,n74);
and (n913,n391,n67);
or (n914,n855,n15);
nand (n915,n916,n920);
or (n916,n278,n917);
nor (n917,n918,n919);
and (n918,n174,n289);
and (n919,n178,n284);
or (n920,n862,n290);
and (n921,n903,n909);
and (n922,n881,n887);
and (n923,n876,n877);
and (n924,n777,n825);
xor (n925,n926,n931);
xor (n926,n927,n928);
xor (n927,n488,n552);
or (n928,n929,n930);
and (n929,n826,n829);
and (n930,n827,n828);
xor (n931,n932,n937);
xor (n932,n933,n934);
xor (n933,n591,n604);
or (n934,n935,n936);
and (n935,n778,n803);
and (n936,n779,n780);
xor (n937,n439,n465);
or (n938,n939,n1347);
and (n939,n940,n971);
xor (n940,n941,n970);
or (n941,n942,n969);
and (n942,n943,n968);
xor (n943,n944,n967);
or (n944,n945,n966);
and (n945,n946,n949);
xor (n946,n947,n948);
xor (n947,n835,n843);
xor (n948,n852,n865);
or (n949,n950,n965);
and (n950,n951,n964);
xor (n951,n952,n958);
nand (n952,n953,n957);
or (n953,n342,n954);
nor (n954,n955,n956);
and (n955,n352,n205);
and (n956,n356,n203);
or (n957,n868,n343);
nand (n958,n959,n963);
or (n959,n318,n960);
nor (n960,n961,n962);
and (n961,n359,n63);
and (n962,n363,n17);
or (n963,n883,n319);
xor (n964,n888,n894);
and (n965,n952,n958);
and (n966,n947,n948);
xor (n967,n831,n850);
xor (n968,n875,n878);
and (n969,n944,n967);
xor (n970,n776,n873);
nand (n971,n972,n1344,n1346);
or (n972,n973,n1339);
nand (n973,n974,n1328);
or (n974,n975,n1327);
and (n975,n976,n1097);
xor (n976,n977,n1082);
or (n977,n978,n1081);
and (n978,n979,n1047);
xor (n979,n980,n1002);
xor (n980,n981,n996);
xor (n981,n982,n989);
nand (n982,n983,n988);
or (n983,n14,n984);
not (n984,n985);
nor (n985,n986,n987);
and (n986,n74,n187);
and (n987,n183,n67);
or (n988,n911,n15);
nand (n989,n990,n995);
or (n990,n991,n278);
not (n991,n992);
nand (n992,n993,n994);
or (n993,n225,n284);
or (n994,n221,n289);
or (n995,n917,n290);
nand (n996,n997,n1001);
or (n997,n318,n998);
nor (n998,n999,n1000);
and (n999,n396,n63);
and (n1000,n400,n17);
or (n1001,n319,n960);
or (n1002,n1003,n1046);
and (n1003,n1004,n1026);
xor (n1004,n1005,n1011);
nand (n1005,n1006,n1010);
or (n1006,n318,n1007);
nor (n1007,n1008,n1009);
and (n1008,n387,n63);
and (n1009,n391,n17);
or (n1010,n998,n319);
xor (n1011,n1012,n1018);
nor (n1012,n1013,n289);
nor (n1013,n1014,n1017);
and (n1014,n1015,n74);
not (n1015,n1016);
and (n1016,n203,n281);
and (n1017,n288,n205);
nand (n1018,n1019,n1022);
or (n1019,n420,n1020);
not (n1020,n1021);
xnor (n1021,n296,n233);
or (n1022,n1023,n421);
nor (n1023,n1024,n1025);
and (n1024,n233,n304);
and (n1025,n308,n234);
or (n1026,n1027,n1045);
and (n1027,n1028,n1036);
xor (n1028,n1029,n1030);
nor (n1029,n290,n205);
nand (n1030,n1031,n1032);
or (n1031,n421,n1020);
or (n1032,n1033,n420);
nor (n1033,n1034,n1035);
and (n1034,n233,n367);
and (n1035,n371,n234);
nand (n1036,n1037,n1041);
or (n1037,n14,n1038);
nor (n1038,n1039,n1040);
and (n1039,n221,n74);
and (n1040,n225,n67);
or (n1041,n1042,n15);
nor (n1042,n1043,n1044);
and (n1043,n174,n74);
and (n1044,n178,n67);
and (n1045,n1029,n1030);
and (n1046,n1005,n1011);
xor (n1047,n1048,n1062);
xor (n1048,n1049,n1050);
and (n1049,n1012,n1018);
xor (n1050,n1051,n1056);
xor (n1051,n1052,n1053);
nor (n1052,n343,n205);
nand (n1053,n1054,n1055);
or (n1054,n1023,n420);
or (n1055,n890,n421);
nand (n1056,n1057,n1061);
or (n1057,n230,n1058);
nor (n1058,n1059,n1060);
and (n1059,n367,n244);
and (n1060,n371,n245);
or (n1061,n231,n905);
or (n1062,n1063,n1080);
and (n1063,n1064,n1074);
xor (n1064,n1065,n1071);
nand (n1065,n1066,n1070);
or (n1066,n230,n1067);
nor (n1067,n1068,n1069);
and (n1068,n244,n359);
and (n1069,n363,n245);
or (n1070,n1058,n231);
nand (n1071,n1072,n1073);
or (n1072,n15,n984);
or (n1073,n1042,n14);
nand (n1074,n1075,n1076);
or (n1075,n290,n991);
or (n1076,n278,n1077);
nor (n1077,n1078,n1079);
and (n1078,n284,n205);
and (n1079,n289,n203);
and (n1080,n1065,n1071);
and (n1081,n980,n1002);
xor (n1082,n1083,n1088);
xor (n1083,n1084,n1085);
xor (n1084,n902,n915);
or (n1085,n1086,n1087);
and (n1086,n1048,n1062);
and (n1087,n1049,n1050);
xor (n1088,n1089,n1096);
xor (n1089,n1090,n1093);
or (n1090,n1091,n1092);
and (n1091,n1051,n1056);
and (n1092,n1052,n1053);
or (n1093,n1094,n1095);
and (n1094,n981,n996);
and (n1095,n982,n989);
xor (n1096,n951,n964);
or (n1097,n1098,n1326);
and (n1098,n1099,n1136);
xor (n1099,n1100,n1135);
or (n1100,n1101,n1134);
and (n1101,n1102,n1133);
xor (n1102,n1103,n1132);
or (n1103,n1104,n1131);
and (n1104,n1105,n1118);
xor (n1105,n1106,n1112);
nand (n1106,n1107,n1111);
or (n1107,n230,n1108);
nor (n1108,n1109,n1110);
and (n1109,n396,n244);
and (n1110,n245,n400);
or (n1111,n1067,n231);
nand (n1112,n1113,n1117);
or (n1113,n318,n1114);
nor (n1114,n1115,n1116);
and (n1115,n183,n63);
and (n1116,n187,n17);
or (n1117,n1007,n319);
and (n1118,n1119,n1125);
nor (n1119,n1120,n74);
nor (n1120,n1121,n1124);
and (n1121,n1122,n63);
not (n1122,n1123);
and (n1123,n203,n56);
and (n1124,n64,n205);
nand (n1125,n1126,n1130);
or (n1126,n1127,n420);
nor (n1127,n1128,n1129);
and (n1128,n233,n359);
and (n1129,n363,n234);
or (n1130,n1033,n421);
and (n1131,n1106,n1112);
xor (n1132,n1064,n1074);
xor (n1133,n1004,n1026);
and (n1134,n1103,n1132);
xor (n1135,n979,n1047);
nand (n1136,n1137,n1323,n1325);
or (n1137,n1138,n1196);
nand (n1138,n1139,n1191);
not (n1139,n1140);
nor (n1140,n1141,n1167);
xor (n1141,n1142,n1166);
xor (n1142,n1143,n1165);
or (n1143,n1144,n1164);
and (n1144,n1145,n1158);
xor (n1145,n1146,n1152);
nand (n1146,n1147,n1151);
or (n1147,n14,n1148);
nor (n1148,n1149,n1150);
and (n1149,n67,n205);
and (n1150,n74,n203);
or (n1151,n1038,n15);
nand (n1152,n1153,n1157);
or (n1153,n1154,n230);
nor (n1154,n1155,n1156);
and (n1155,n245,n391);
and (n1156,n244,n387);
or (n1157,n1108,n231);
nand (n1158,n1159,n1163);
or (n1159,n318,n1160);
nor (n1160,n1161,n1162);
and (n1161,n174,n63);
and (n1162,n178,n17);
or (n1163,n1114,n319);
and (n1164,n1146,n1152);
xor (n1165,n1028,n1036);
xor (n1166,n1105,n1118);
or (n1167,n1168,n1190);
and (n1168,n1169,n1189);
xor (n1169,n1170,n1171);
xor (n1170,n1119,n1125);
or (n1171,n1172,n1188);
and (n1172,n1173,n1182);
xor (n1173,n1174,n1175);
nor (n1174,n15,n205);
nand (n1175,n1176,n1181);
or (n1176,n1177,n420);
not (n1177,n1178);
nand (n1178,n1179,n1180);
or (n1179,n234,n400);
nand (n1180,n400,n234);
or (n1181,n1127,n421);
nand (n1182,n1183,n1187);
or (n1183,n230,n1184);
nor (n1184,n1185,n1186);
and (n1185,n244,n183);
and (n1186,n245,n187);
or (n1187,n1154,n231);
and (n1188,n1174,n1175);
xor (n1189,n1145,n1158);
and (n1190,n1170,n1171);
or (n1191,n1192,n1193);
xor (n1192,n1102,n1133);
or (n1193,n1194,n1195);
and (n1194,n1142,n1166);
and (n1195,n1143,n1165);
nor (n1196,n1197,n1322);
and (n1197,n1198,n1317);
or (n1198,n1199,n1316);
and (n1199,n1200,n1241);
xor (n1200,n1201,n1234);
or (n1201,n1202,n1233);
and (n1202,n1203,n1219);
xor (n1203,n1204,n1210);
nand (n1204,n1205,n1209);
or (n1205,n230,n1206);
nor (n1206,n1207,n1208);
and (n1207,n245,n178);
and (n1208,n244,n174);
or (n1209,n1184,n231);
or (n1210,n1211,n1215);
nor (n1211,n1212,n319);
nor (n1212,n1213,n1214);
and (n1213,n63,n221);
and (n1214,n17,n225);
nor (n1215,n318,n1216);
nor (n1216,n1217,n1218);
and (n1217,n17,n205);
and (n1218,n63,n203);
xor (n1219,n1220,n1226);
nor (n1220,n1221,n63);
nor (n1221,n1222,n1225);
and (n1222,n1223,n244);
not (n1223,n1224);
and (n1224,n203,n322);
and (n1225,n328,n205);
nand (n1226,n1227,n1232);
or (n1227,n420,n1228);
not (n1228,n1229);
nand (n1229,n1230,n1231);
or (n1230,n233,n387);
nand (n1231,n387,n233);
nand (n1232,n1178,n422);
and (n1233,n1204,n1210);
xor (n1234,n1235,n1240);
xor (n1235,n1236,n1239);
nand (n1236,n1237,n1238);
or (n1237,n318,n1212);
or (n1238,n1160,n319);
and (n1239,n1220,n1226);
xor (n1240,n1173,n1182);
or (n1241,n1242,n1315);
and (n1242,n1243,n1263);
xor (n1243,n1244,n1262);
or (n1244,n1245,n1261);
and (n1245,n1246,n1255);
xor (n1246,n1247,n1248);
and (n1247,n320,n203);
nand (n1248,n1249,n1254);
or (n1249,n420,n1250);
not (n1250,n1251);
nand (n1251,n1252,n1253);
or (n1252,n234,n187);
nand (n1253,n187,n234);
nand (n1254,n1229,n422);
nand (n1255,n1256,n1260);
or (n1256,n230,n1257);
nor (n1257,n1258,n1259);
and (n1258,n244,n221);
and (n1259,n245,n225);
or (n1260,n1206,n231);
and (n1261,n1247,n1248);
xor (n1262,n1203,n1219);
or (n1263,n1264,n1314);
and (n1264,n1265,n1282);
xor (n1265,n1266,n1281);
and (n1266,n1267,n1273);
and (n1267,n1268,n245);
nand (n1268,n1269,n1272);
nand (n1269,n1270,n233);
not (n1270,n1271);
and (n1271,n203,n237);
nand (n1272,n241,n205);
nand (n1273,n1274,n1275);
or (n1274,n421,n1250);
nand (n1275,n1276,n1280);
not (n1276,n1277);
nor (n1277,n1278,n1279);
and (n1278,n178,n234);
and (n1279,n174,n233);
not (n1280,n420);
xor (n1281,n1246,n1255);
or (n1282,n1283,n1313);
and (n1283,n1284,n1292);
xor (n1284,n1285,n1291);
nand (n1285,n1286,n1290);
or (n1286,n230,n1287);
nor (n1287,n1288,n1289);
and (n1288,n245,n205);
and (n1289,n244,n203);
or (n1290,n1257,n231);
xor (n1291,n1267,n1273);
or (n1292,n1293,n1312);
and (n1293,n1294,n1302);
xor (n1294,n1295,n1296);
nor (n1295,n231,n205);
nand (n1296,n1297,n1301);
or (n1297,n1298,n420);
or (n1298,n1299,n1300);
and (n1299,n233,n225);
and (n1300,n221,n234);
or (n1301,n1277,n421);
nor (n1302,n1303,n1310);
nor (n1303,n1304,n1306);
and (n1304,n1305,n422);
not (n1305,n1298);
and (n1306,n1307,n1280);
nand (n1307,n1308,n1309);
or (n1308,n233,n203);
or (n1309,n234,n205);
or (n1310,n233,n1311);
and (n1311,n203,n422);
and (n1312,n1295,n1296);
and (n1313,n1285,n1291);
and (n1314,n1266,n1281);
and (n1315,n1244,n1262);
and (n1316,n1201,n1234);
or (n1317,n1318,n1319);
xor (n1318,n1169,n1189);
or (n1319,n1320,n1321);
and (n1320,n1235,n1240);
and (n1321,n1236,n1239);
and (n1322,n1318,n1319);
nand (n1323,n1191,n1324);
and (n1324,n1141,n1167);
nand (n1325,n1192,n1193);
and (n1326,n1100,n1135);
and (n1327,n977,n1082);
or (n1328,n1329,n1336);
xor (n1329,n1330,n1335);
xor (n1330,n1331,n1332);
xor (n1331,n880,n900);
or (n1332,n1333,n1334);
and (n1333,n1089,n1096);
and (n1334,n1090,n1093);
xor (n1335,n946,n949);
or (n1336,n1337,n1338);
and (n1337,n1083,n1088);
and (n1338,n1084,n1085);
nor (n1339,n1340,n1341);
xor (n1340,n943,n968);
or (n1341,n1342,n1343);
and (n1342,n1330,n1335);
and (n1343,n1331,n1332);
or (n1344,n1339,n1345);
nand (n1345,n1329,n1336);
nand (n1346,n1340,n1341);
and (n1347,n941,n970);
and (n1348,n774,n925);
nor (n1349,n1350,n1361);
nor (n1350,n1351,n1352);
xor (n1351,n7,n612);
or (n1352,n1353,n1360);
and (n1353,n1354,n1359);
xor (n1354,n1355,n1356);
xor (n1355,n650,n655);
or (n1356,n1357,n1358);
and (n1357,n932,n937);
and (n1358,n933,n934);
xor (n1359,n436,n574);
and (n1360,n1355,n1356);
nor (n1361,n1362,n1363);
xor (n1362,n1354,n1359);
or (n1363,n1364,n1365);
and (n1364,n926,n931);
and (n1365,n927,n928);
nand (n1366,n1367,n1369);
or (n1367,n1350,n1368);
nand (n1368,n1362,n1363);
nand (n1369,n1351,n1352);
or (n1370,n768,n3);
xor (n1371,n1372,n2281);
xor (n1372,n1373,n2278);
xor (n1373,n1374,n2277);
xor (n1374,n1375,n2269);
xor (n1375,n1376,n2268);
xor (n1376,n1377,n2253);
xor (n1377,n1378,n2252);
xor (n1378,n1379,n2232);
xor (n1379,n1380,n2231);
xor (n1380,n1381,n2204);
xor (n1381,n1382,n2203);
xor (n1382,n1383,n2171);
xor (n1383,n1384,n2170);
xor (n1384,n1385,n2131);
xor (n1385,n1386,n2130);
xor (n1386,n1387,n2086);
xor (n1387,n1388,n2085);
xor (n1388,n1389,n2034);
xor (n1389,n1390,n2033);
xor (n1390,n1391,n1977);
xor (n1391,n1392,n1976);
xor (n1392,n1393,n1914);
xor (n1393,n1394,n1913);
xor (n1394,n1395,n1845);
xor (n1395,n1396,n1844);
xor (n1396,n1397,n1769);
xor (n1397,n1398,n1768);
xor (n1398,n1399,n1688);
xor (n1399,n1400,n1687);
xor (n1400,n1401,n1600);
xor (n1401,n1402,n1599);
xor (n1402,n1403,n1507);
xor (n1403,n1404,n1506);
xor (n1404,n1405,n1408);
xor (n1405,n1406,n1407);
and (n1406,n752,n422);
and (n1407,n426,n234);
or (n1408,n1409,n1412);
and (n1409,n1410,n1411);
and (n1410,n426,n422);
and (n1411,n412,n234);
and (n1412,n1413,n1414);
xor (n1413,n1410,n1411);
or (n1414,n1415,n1418);
and (n1415,n1416,n1417);
and (n1416,n412,n422);
and (n1417,n268,n234);
and (n1418,n1419,n1420);
xor (n1419,n1416,n1417);
or (n1420,n1421,n1424);
and (n1421,n1422,n1423);
and (n1422,n268,n422);
and (n1423,n251,n234);
and (n1424,n1425,n1426);
xor (n1425,n1422,n1423);
or (n1426,n1427,n1430);
and (n1427,n1428,n1429);
and (n1428,n251,n422);
and (n1429,n333,n234);
and (n1430,n1431,n1432);
xor (n1431,n1428,n1429);
or (n1432,n1433,n1436);
and (n1433,n1434,n1435);
and (n1434,n333,n422);
and (n1435,n313,n234);
and (n1436,n1437,n1438);
xor (n1437,n1434,n1435);
or (n1438,n1439,n1442);
and (n1439,n1440,n1441);
and (n1440,n313,n422);
and (n1441,n118,n234);
and (n1442,n1443,n1444);
xor (n1443,n1440,n1441);
or (n1444,n1445,n1448);
and (n1445,n1446,n1447);
and (n1446,n118,n422);
and (n1447,n77,n234);
and (n1448,n1449,n1450);
xor (n1449,n1446,n1447);
or (n1450,n1451,n1454);
and (n1451,n1452,n1453);
and (n1452,n77,n422);
and (n1453,n304,n234);
and (n1454,n1455,n1456);
xor (n1455,n1452,n1453);
or (n1456,n1457,n1460);
and (n1457,n1458,n1459);
and (n1458,n304,n422);
and (n1459,n296,n234);
and (n1460,n1461,n1462);
xor (n1461,n1458,n1459);
or (n1462,n1463,n1466);
and (n1463,n1464,n1465);
and (n1464,n296,n422);
and (n1465,n367,n234);
and (n1466,n1467,n1468);
xor (n1467,n1464,n1465);
or (n1468,n1469,n1472);
and (n1469,n1470,n1471);
and (n1470,n367,n422);
and (n1471,n359,n234);
and (n1472,n1473,n1474);
xor (n1473,n1470,n1471);
or (n1474,n1475,n1478);
and (n1475,n1476,n1477);
and (n1476,n359,n422);
and (n1477,n396,n234);
and (n1478,n1479,n1480);
xor (n1479,n1476,n1477);
or (n1480,n1481,n1484);
and (n1481,n1482,n1483);
and (n1482,n396,n422);
and (n1483,n387,n234);
and (n1484,n1485,n1486);
xor (n1485,n1482,n1483);
or (n1486,n1487,n1490);
and (n1487,n1488,n1489);
and (n1488,n387,n422);
and (n1489,n183,n234);
and (n1490,n1491,n1492);
xor (n1491,n1488,n1489);
or (n1492,n1493,n1496);
and (n1493,n1494,n1495);
and (n1494,n183,n422);
and (n1495,n174,n234);
and (n1496,n1497,n1498);
xor (n1497,n1494,n1495);
or (n1498,n1499,n1501);
and (n1499,n1500,n1300);
and (n1500,n174,n422);
and (n1501,n1502,n1503);
xor (n1502,n1500,n1300);
and (n1503,n1504,n1505);
and (n1504,n221,n422);
and (n1505,n203,n234);
and (n1506,n412,n237);
or (n1507,n1508,n1511);
and (n1508,n1509,n1510);
xor (n1509,n1413,n1414);
and (n1510,n268,n237);
and (n1511,n1512,n1513);
xor (n1512,n1509,n1510);
or (n1513,n1514,n1517);
and (n1514,n1515,n1516);
xor (n1515,n1419,n1420);
and (n1516,n251,n237);
and (n1517,n1518,n1519);
xor (n1518,n1515,n1516);
or (n1519,n1520,n1523);
and (n1520,n1521,n1522);
xor (n1521,n1425,n1426);
and (n1522,n333,n237);
and (n1523,n1524,n1525);
xor (n1524,n1521,n1522);
or (n1525,n1526,n1529);
and (n1526,n1527,n1528);
xor (n1527,n1431,n1432);
and (n1528,n313,n237);
and (n1529,n1530,n1531);
xor (n1530,n1527,n1528);
or (n1531,n1532,n1535);
and (n1532,n1533,n1534);
xor (n1533,n1437,n1438);
and (n1534,n118,n237);
and (n1535,n1536,n1537);
xor (n1536,n1533,n1534);
or (n1537,n1538,n1541);
and (n1538,n1539,n1540);
xor (n1539,n1443,n1444);
and (n1540,n77,n237);
and (n1541,n1542,n1543);
xor (n1542,n1539,n1540);
or (n1543,n1544,n1547);
and (n1544,n1545,n1546);
xor (n1545,n1449,n1450);
and (n1546,n304,n237);
and (n1547,n1548,n1549);
xor (n1548,n1545,n1546);
or (n1549,n1550,n1553);
and (n1550,n1551,n1552);
xor (n1551,n1455,n1456);
and (n1552,n296,n237);
and (n1553,n1554,n1555);
xor (n1554,n1551,n1552);
or (n1555,n1556,n1559);
and (n1556,n1557,n1558);
xor (n1557,n1461,n1462);
and (n1558,n367,n237);
and (n1559,n1560,n1561);
xor (n1560,n1557,n1558);
or (n1561,n1562,n1565);
and (n1562,n1563,n1564);
xor (n1563,n1467,n1468);
and (n1564,n359,n237);
and (n1565,n1566,n1567);
xor (n1566,n1563,n1564);
or (n1567,n1568,n1571);
and (n1568,n1569,n1570);
xor (n1569,n1473,n1474);
and (n1570,n396,n237);
and (n1571,n1572,n1573);
xor (n1572,n1569,n1570);
or (n1573,n1574,n1577);
and (n1574,n1575,n1576);
xor (n1575,n1479,n1480);
and (n1576,n387,n237);
and (n1577,n1578,n1579);
xor (n1578,n1575,n1576);
or (n1579,n1580,n1583);
and (n1580,n1581,n1582);
xor (n1581,n1485,n1486);
and (n1582,n183,n237);
and (n1583,n1584,n1585);
xor (n1584,n1581,n1582);
or (n1585,n1586,n1589);
and (n1586,n1587,n1588);
xor (n1587,n1491,n1492);
and (n1588,n174,n237);
and (n1589,n1590,n1591);
xor (n1590,n1587,n1588);
or (n1591,n1592,n1595);
and (n1592,n1593,n1594);
xor (n1593,n1497,n1498);
and (n1594,n221,n237);
and (n1595,n1596,n1597);
xor (n1596,n1593,n1594);
and (n1597,n1598,n1271);
xor (n1598,n1502,n1503);
and (n1599,n268,n245);
or (n1600,n1601,n1604);
and (n1601,n1602,n1603);
xor (n1602,n1512,n1513);
and (n1603,n251,n245);
and (n1604,n1605,n1606);
xor (n1605,n1602,n1603);
or (n1606,n1607,n1610);
and (n1607,n1608,n1609);
xor (n1608,n1518,n1519);
and (n1609,n333,n245);
and (n1610,n1611,n1612);
xor (n1611,n1608,n1609);
or (n1612,n1613,n1616);
and (n1613,n1614,n1615);
xor (n1614,n1524,n1525);
and (n1615,n313,n245);
and (n1616,n1617,n1618);
xor (n1617,n1614,n1615);
or (n1618,n1619,n1622);
and (n1619,n1620,n1621);
xor (n1620,n1530,n1531);
and (n1621,n118,n245);
and (n1622,n1623,n1624);
xor (n1623,n1620,n1621);
or (n1624,n1625,n1628);
and (n1625,n1626,n1627);
xor (n1626,n1536,n1537);
and (n1627,n77,n245);
and (n1628,n1629,n1630);
xor (n1629,n1626,n1627);
or (n1630,n1631,n1634);
and (n1631,n1632,n1633);
xor (n1632,n1542,n1543);
and (n1633,n304,n245);
and (n1634,n1635,n1636);
xor (n1635,n1632,n1633);
or (n1636,n1637,n1640);
and (n1637,n1638,n1639);
xor (n1638,n1548,n1549);
and (n1639,n296,n245);
and (n1640,n1641,n1642);
xor (n1641,n1638,n1639);
or (n1642,n1643,n1646);
and (n1643,n1644,n1645);
xor (n1644,n1554,n1555);
and (n1645,n367,n245);
and (n1646,n1647,n1648);
xor (n1647,n1644,n1645);
or (n1648,n1649,n1652);
and (n1649,n1650,n1651);
xor (n1650,n1560,n1561);
and (n1651,n359,n245);
and (n1652,n1653,n1654);
xor (n1653,n1650,n1651);
or (n1654,n1655,n1658);
and (n1655,n1656,n1657);
xor (n1656,n1566,n1567);
and (n1657,n396,n245);
and (n1658,n1659,n1660);
xor (n1659,n1656,n1657);
or (n1660,n1661,n1664);
and (n1661,n1662,n1663);
xor (n1662,n1572,n1573);
and (n1663,n387,n245);
and (n1664,n1665,n1666);
xor (n1665,n1662,n1663);
or (n1666,n1667,n1670);
and (n1667,n1668,n1669);
xor (n1668,n1578,n1579);
and (n1669,n183,n245);
and (n1670,n1671,n1672);
xor (n1671,n1668,n1669);
or (n1672,n1673,n1676);
and (n1673,n1674,n1675);
xor (n1674,n1584,n1585);
and (n1675,n174,n245);
and (n1676,n1677,n1678);
xor (n1677,n1674,n1675);
or (n1678,n1679,n1682);
and (n1679,n1680,n1681);
xor (n1680,n1590,n1591);
and (n1681,n221,n245);
and (n1682,n1683,n1684);
xor (n1683,n1680,n1681);
and (n1684,n1685,n1686);
xor (n1685,n1596,n1597);
and (n1686,n203,n245);
and (n1687,n251,n322);
or (n1688,n1689,n1692);
and (n1689,n1690,n1691);
xor (n1690,n1605,n1606);
and (n1691,n333,n322);
and (n1692,n1693,n1694);
xor (n1693,n1690,n1691);
or (n1694,n1695,n1698);
and (n1695,n1696,n1697);
xor (n1696,n1611,n1612);
and (n1697,n313,n322);
and (n1698,n1699,n1700);
xor (n1699,n1696,n1697);
or (n1700,n1701,n1704);
and (n1701,n1702,n1703);
xor (n1702,n1617,n1618);
and (n1703,n118,n322);
and (n1704,n1705,n1706);
xor (n1705,n1702,n1703);
or (n1706,n1707,n1710);
and (n1707,n1708,n1709);
xor (n1708,n1623,n1624);
and (n1709,n77,n322);
and (n1710,n1711,n1712);
xor (n1711,n1708,n1709);
or (n1712,n1713,n1716);
and (n1713,n1714,n1715);
xor (n1714,n1629,n1630);
and (n1715,n304,n322);
and (n1716,n1717,n1718);
xor (n1717,n1714,n1715);
or (n1718,n1719,n1722);
and (n1719,n1720,n1721);
xor (n1720,n1635,n1636);
and (n1721,n296,n322);
and (n1722,n1723,n1724);
xor (n1723,n1720,n1721);
or (n1724,n1725,n1728);
and (n1725,n1726,n1727);
xor (n1726,n1641,n1642);
and (n1727,n367,n322);
and (n1728,n1729,n1730);
xor (n1729,n1726,n1727);
or (n1730,n1731,n1734);
and (n1731,n1732,n1733);
xor (n1732,n1647,n1648);
and (n1733,n359,n322);
and (n1734,n1735,n1736);
xor (n1735,n1732,n1733);
or (n1736,n1737,n1740);
and (n1737,n1738,n1739);
xor (n1738,n1653,n1654);
and (n1739,n396,n322);
and (n1740,n1741,n1742);
xor (n1741,n1738,n1739);
or (n1742,n1743,n1746);
and (n1743,n1744,n1745);
xor (n1744,n1659,n1660);
and (n1745,n387,n322);
and (n1746,n1747,n1748);
xor (n1747,n1744,n1745);
or (n1748,n1749,n1752);
and (n1749,n1750,n1751);
xor (n1750,n1665,n1666);
and (n1751,n183,n322);
and (n1752,n1753,n1754);
xor (n1753,n1750,n1751);
or (n1754,n1755,n1758);
and (n1755,n1756,n1757);
xor (n1756,n1671,n1672);
and (n1757,n174,n322);
and (n1758,n1759,n1760);
xor (n1759,n1756,n1757);
or (n1760,n1761,n1764);
and (n1761,n1762,n1763);
xor (n1762,n1677,n1678);
and (n1763,n221,n322);
and (n1764,n1765,n1766);
xor (n1765,n1762,n1763);
and (n1766,n1767,n1224);
xor (n1767,n1683,n1684);
and (n1768,n333,n17);
or (n1769,n1770,n1773);
and (n1770,n1771,n1772);
xor (n1771,n1693,n1694);
and (n1772,n313,n17);
and (n1773,n1774,n1775);
xor (n1774,n1771,n1772);
or (n1775,n1776,n1779);
and (n1776,n1777,n1778);
xor (n1777,n1699,n1700);
and (n1778,n118,n17);
and (n1779,n1780,n1781);
xor (n1780,n1777,n1778);
or (n1781,n1782,n1785);
and (n1782,n1783,n1784);
xor (n1783,n1705,n1706);
and (n1784,n77,n17);
and (n1785,n1786,n1787);
xor (n1786,n1783,n1784);
or (n1787,n1788,n1791);
and (n1788,n1789,n1790);
xor (n1789,n1711,n1712);
and (n1790,n304,n17);
and (n1791,n1792,n1793);
xor (n1792,n1789,n1790);
or (n1793,n1794,n1797);
and (n1794,n1795,n1796);
xor (n1795,n1717,n1718);
and (n1796,n296,n17);
and (n1797,n1798,n1799);
xor (n1798,n1795,n1796);
or (n1799,n1800,n1803);
and (n1800,n1801,n1802);
xor (n1801,n1723,n1724);
and (n1802,n367,n17);
and (n1803,n1804,n1805);
xor (n1804,n1801,n1802);
or (n1805,n1806,n1809);
and (n1806,n1807,n1808);
xor (n1807,n1729,n1730);
and (n1808,n359,n17);
and (n1809,n1810,n1811);
xor (n1810,n1807,n1808);
or (n1811,n1812,n1815);
and (n1812,n1813,n1814);
xor (n1813,n1735,n1736);
and (n1814,n396,n17);
and (n1815,n1816,n1817);
xor (n1816,n1813,n1814);
or (n1817,n1818,n1821);
and (n1818,n1819,n1820);
xor (n1819,n1741,n1742);
and (n1820,n387,n17);
and (n1821,n1822,n1823);
xor (n1822,n1819,n1820);
or (n1823,n1824,n1827);
and (n1824,n1825,n1826);
xor (n1825,n1747,n1748);
and (n1826,n183,n17);
and (n1827,n1828,n1829);
xor (n1828,n1825,n1826);
or (n1829,n1830,n1833);
and (n1830,n1831,n1832);
xor (n1831,n1753,n1754);
and (n1832,n174,n17);
and (n1833,n1834,n1835);
xor (n1834,n1831,n1832);
or (n1835,n1836,n1839);
and (n1836,n1837,n1838);
xor (n1837,n1759,n1760);
and (n1838,n221,n17);
and (n1839,n1840,n1841);
xor (n1840,n1837,n1838);
and (n1841,n1842,n1843);
xor (n1842,n1765,n1766);
and (n1843,n203,n17);
and (n1844,n313,n56);
or (n1845,n1846,n1849);
and (n1846,n1847,n1848);
xor (n1847,n1774,n1775);
and (n1848,n118,n56);
and (n1849,n1850,n1851);
xor (n1850,n1847,n1848);
or (n1851,n1852,n1855);
and (n1852,n1853,n1854);
xor (n1853,n1780,n1781);
and (n1854,n77,n56);
and (n1855,n1856,n1857);
xor (n1856,n1853,n1854);
or (n1857,n1858,n1861);
and (n1858,n1859,n1860);
xor (n1859,n1786,n1787);
and (n1860,n304,n56);
and (n1861,n1862,n1863);
xor (n1862,n1859,n1860);
or (n1863,n1864,n1867);
and (n1864,n1865,n1866);
xor (n1865,n1792,n1793);
and (n1866,n296,n56);
and (n1867,n1868,n1869);
xor (n1868,n1865,n1866);
or (n1869,n1870,n1873);
and (n1870,n1871,n1872);
xor (n1871,n1798,n1799);
and (n1872,n367,n56);
and (n1873,n1874,n1875);
xor (n1874,n1871,n1872);
or (n1875,n1876,n1879);
and (n1876,n1877,n1878);
xor (n1877,n1804,n1805);
and (n1878,n359,n56);
and (n1879,n1880,n1881);
xor (n1880,n1877,n1878);
or (n1881,n1882,n1885);
and (n1882,n1883,n1884);
xor (n1883,n1810,n1811);
and (n1884,n396,n56);
and (n1885,n1886,n1887);
xor (n1886,n1883,n1884);
or (n1887,n1888,n1891);
and (n1888,n1889,n1890);
xor (n1889,n1816,n1817);
and (n1890,n387,n56);
and (n1891,n1892,n1893);
xor (n1892,n1889,n1890);
or (n1893,n1894,n1897);
and (n1894,n1895,n1896);
xor (n1895,n1822,n1823);
and (n1896,n183,n56);
and (n1897,n1898,n1899);
xor (n1898,n1895,n1896);
or (n1899,n1900,n1903);
and (n1900,n1901,n1902);
xor (n1901,n1828,n1829);
and (n1902,n174,n56);
and (n1903,n1904,n1905);
xor (n1904,n1901,n1902);
or (n1905,n1906,n1909);
and (n1906,n1907,n1908);
xor (n1907,n1834,n1835);
and (n1908,n221,n56);
and (n1909,n1910,n1911);
xor (n1910,n1907,n1908);
and (n1911,n1912,n1123);
xor (n1912,n1840,n1841);
and (n1913,n118,n67);
or (n1914,n1915,n1918);
and (n1915,n1916,n1917);
xor (n1916,n1850,n1851);
and (n1917,n77,n67);
and (n1918,n1919,n1920);
xor (n1919,n1916,n1917);
or (n1920,n1921,n1924);
and (n1921,n1922,n1923);
xor (n1922,n1856,n1857);
and (n1923,n304,n67);
and (n1924,n1925,n1926);
xor (n1925,n1922,n1923);
or (n1926,n1927,n1930);
and (n1927,n1928,n1929);
xor (n1928,n1862,n1863);
and (n1929,n296,n67);
and (n1930,n1931,n1932);
xor (n1931,n1928,n1929);
or (n1932,n1933,n1936);
and (n1933,n1934,n1935);
xor (n1934,n1868,n1869);
and (n1935,n367,n67);
and (n1936,n1937,n1938);
xor (n1937,n1934,n1935);
or (n1938,n1939,n1942);
and (n1939,n1940,n1941);
xor (n1940,n1874,n1875);
and (n1941,n359,n67);
and (n1942,n1943,n1944);
xor (n1943,n1940,n1941);
or (n1944,n1945,n1948);
and (n1945,n1946,n1947);
xor (n1946,n1880,n1881);
and (n1947,n396,n67);
and (n1948,n1949,n1950);
xor (n1949,n1946,n1947);
or (n1950,n1951,n1954);
and (n1951,n1952,n1953);
xor (n1952,n1886,n1887);
and (n1953,n387,n67);
and (n1954,n1955,n1956);
xor (n1955,n1952,n1953);
or (n1956,n1957,n1959);
and (n1957,n1958,n987);
xor (n1958,n1892,n1893);
and (n1959,n1960,n1961);
xor (n1960,n1958,n987);
or (n1961,n1962,n1965);
and (n1962,n1963,n1964);
xor (n1963,n1898,n1899);
and (n1964,n174,n67);
and (n1965,n1966,n1967);
xor (n1966,n1963,n1964);
or (n1967,n1968,n1971);
and (n1968,n1969,n1970);
xor (n1969,n1904,n1905);
and (n1970,n221,n67);
and (n1971,n1972,n1973);
xor (n1972,n1969,n1970);
and (n1973,n1974,n1975);
xor (n1974,n1910,n1911);
and (n1975,n203,n67);
and (n1976,n77,n281);
or (n1977,n1978,n1981);
and (n1978,n1979,n1980);
xor (n1979,n1919,n1920);
and (n1980,n304,n281);
and (n1981,n1982,n1983);
xor (n1982,n1979,n1980);
or (n1983,n1984,n1987);
and (n1984,n1985,n1986);
xor (n1985,n1925,n1926);
and (n1986,n296,n281);
and (n1987,n1988,n1989);
xor (n1988,n1985,n1986);
or (n1989,n1990,n1993);
and (n1990,n1991,n1992);
xor (n1991,n1931,n1932);
and (n1992,n367,n281);
and (n1993,n1994,n1995);
xor (n1994,n1991,n1992);
or (n1995,n1996,n1999);
and (n1996,n1997,n1998);
xor (n1997,n1937,n1938);
and (n1998,n359,n281);
and (n1999,n2000,n2001);
xor (n2000,n1997,n1998);
or (n2001,n2002,n2005);
and (n2002,n2003,n2004);
xor (n2003,n1943,n1944);
and (n2004,n396,n281);
and (n2005,n2006,n2007);
xor (n2006,n2003,n2004);
or (n2007,n2008,n2011);
and (n2008,n2009,n2010);
xor (n2009,n1949,n1950);
and (n2010,n387,n281);
and (n2011,n2012,n2013);
xor (n2012,n2009,n2010);
or (n2013,n2014,n2017);
and (n2014,n2015,n2016);
xor (n2015,n1955,n1956);
and (n2016,n183,n281);
and (n2017,n2018,n2019);
xor (n2018,n2015,n2016);
or (n2019,n2020,n2023);
and (n2020,n2021,n2022);
xor (n2021,n1960,n1961);
and (n2022,n174,n281);
and (n2023,n2024,n2025);
xor (n2024,n2021,n2022);
or (n2025,n2026,n2029);
and (n2026,n2027,n2028);
xor (n2027,n1966,n1967);
and (n2028,n221,n281);
and (n2029,n2030,n2031);
xor (n2030,n2027,n2028);
and (n2031,n2032,n1016);
xor (n2032,n1972,n1973);
and (n2033,n304,n284);
or (n2034,n2035,n2038);
and (n2035,n2036,n2037);
xor (n2036,n1982,n1983);
and (n2037,n296,n284);
and (n2038,n2039,n2040);
xor (n2039,n2036,n2037);
or (n2040,n2041,n2044);
and (n2041,n2042,n2043);
xor (n2042,n1988,n1989);
and (n2043,n367,n284);
and (n2044,n2045,n2046);
xor (n2045,n2042,n2043);
or (n2046,n2047,n2050);
and (n2047,n2048,n2049);
xor (n2048,n1994,n1995);
and (n2049,n359,n284);
and (n2050,n2051,n2052);
xor (n2051,n2048,n2049);
or (n2052,n2053,n2056);
and (n2053,n2054,n2055);
xor (n2054,n2000,n2001);
and (n2055,n396,n284);
and (n2056,n2057,n2058);
xor (n2057,n2054,n2055);
or (n2058,n2059,n2062);
and (n2059,n2060,n2061);
xor (n2060,n2006,n2007);
and (n2061,n387,n284);
and (n2062,n2063,n2064);
xor (n2063,n2060,n2061);
or (n2064,n2065,n2068);
and (n2065,n2066,n2067);
xor (n2066,n2012,n2013);
and (n2067,n183,n284);
and (n2068,n2069,n2070);
xor (n2069,n2066,n2067);
or (n2070,n2071,n2074);
and (n2071,n2072,n2073);
xor (n2072,n2018,n2019);
and (n2073,n174,n284);
and (n2074,n2075,n2076);
xor (n2075,n2072,n2073);
or (n2076,n2077,n2080);
and (n2077,n2078,n2079);
xor (n2078,n2024,n2025);
and (n2079,n221,n284);
and (n2080,n2081,n2082);
xor (n2081,n2078,n2079);
and (n2082,n2083,n2084);
xor (n2083,n2030,n2031);
and (n2084,n203,n284);
and (n2085,n296,n345);
or (n2086,n2087,n2090);
and (n2087,n2088,n2089);
xor (n2088,n2039,n2040);
and (n2089,n367,n345);
and (n2090,n2091,n2092);
xor (n2091,n2088,n2089);
or (n2092,n2093,n2096);
and (n2093,n2094,n2095);
xor (n2094,n2045,n2046);
and (n2095,n359,n345);
and (n2096,n2097,n2098);
xor (n2097,n2094,n2095);
or (n2098,n2099,n2102);
and (n2099,n2100,n2101);
xor (n2100,n2051,n2052);
and (n2101,n396,n345);
and (n2102,n2103,n2104);
xor (n2103,n2100,n2101);
or (n2104,n2105,n2108);
and (n2105,n2106,n2107);
xor (n2106,n2057,n2058);
and (n2107,n387,n345);
and (n2108,n2109,n2110);
xor (n2109,n2106,n2107);
or (n2110,n2111,n2114);
and (n2111,n2112,n2113);
xor (n2112,n2063,n2064);
and (n2113,n183,n345);
and (n2114,n2115,n2116);
xor (n2115,n2112,n2113);
or (n2116,n2117,n2120);
and (n2117,n2118,n2119);
xor (n2118,n2069,n2070);
and (n2119,n174,n345);
and (n2120,n2121,n2122);
xor (n2121,n2118,n2119);
or (n2122,n2123,n2126);
and (n2123,n2124,n2125);
xor (n2124,n2075,n2076);
and (n2125,n221,n345);
and (n2126,n2127,n2128);
xor (n2127,n2124,n2125);
and (n2128,n2129,n898);
xor (n2129,n2081,n2082);
and (n2130,n367,n352);
or (n2131,n2132,n2135);
and (n2132,n2133,n2134);
xor (n2133,n2091,n2092);
and (n2134,n359,n352);
and (n2135,n2136,n2137);
xor (n2136,n2133,n2134);
or (n2137,n2138,n2141);
and (n2138,n2139,n2140);
xor (n2139,n2097,n2098);
and (n2140,n396,n352);
and (n2141,n2142,n2143);
xor (n2142,n2139,n2140);
or (n2143,n2144,n2147);
and (n2144,n2145,n2146);
xor (n2145,n2103,n2104);
and (n2146,n387,n352);
and (n2147,n2148,n2149);
xor (n2148,n2145,n2146);
or (n2149,n2150,n2153);
and (n2150,n2151,n2152);
xor (n2151,n2109,n2110);
and (n2152,n183,n352);
and (n2153,n2154,n2155);
xor (n2154,n2151,n2152);
or (n2155,n2156,n2159);
and (n2156,n2157,n2158);
xor (n2157,n2115,n2116);
and (n2158,n174,n352);
and (n2159,n2160,n2161);
xor (n2160,n2157,n2158);
or (n2161,n2162,n2165);
and (n2162,n2163,n2164);
xor (n2163,n2121,n2122);
and (n2164,n221,n352);
and (n2165,n2166,n2167);
xor (n2166,n2163,n2164);
and (n2167,n2168,n2169);
xor (n2168,n2127,n2128);
and (n2169,n203,n352);
and (n2170,n359,n377);
or (n2171,n2172,n2175);
and (n2172,n2173,n2174);
xor (n2173,n2136,n2137);
and (n2174,n396,n377);
and (n2175,n2176,n2177);
xor (n2176,n2173,n2174);
or (n2177,n2178,n2181);
and (n2178,n2179,n2180);
xor (n2179,n2142,n2143);
and (n2180,n387,n377);
and (n2181,n2182,n2183);
xor (n2182,n2179,n2180);
or (n2183,n2184,n2187);
and (n2184,n2185,n2186);
xor (n2185,n2148,n2149);
and (n2186,n183,n377);
and (n2187,n2188,n2189);
xor (n2188,n2185,n2186);
or (n2189,n2190,n2193);
and (n2190,n2191,n2192);
xor (n2191,n2154,n2155);
and (n2192,n174,n377);
and (n2193,n2194,n2195);
xor (n2194,n2191,n2192);
or (n2195,n2196,n2199);
and (n2196,n2197,n2198);
xor (n2197,n2160,n2161);
and (n2198,n221,n377);
and (n2199,n2200,n2201);
xor (n2200,n2197,n2198);
and (n2201,n2202,n549);
xor (n2202,n2166,n2167);
and (n2203,n396,n133);
or (n2204,n2205,n2208);
and (n2205,n2206,n2207);
xor (n2206,n2176,n2177);
and (n2207,n387,n133);
and (n2208,n2209,n2210);
xor (n2209,n2206,n2207);
or (n2210,n2211,n2214);
and (n2211,n2212,n2213);
xor (n2212,n2182,n2183);
and (n2213,n183,n133);
and (n2214,n2215,n2216);
xor (n2215,n2212,n2213);
or (n2216,n2217,n2220);
and (n2217,n2218,n2219);
xor (n2218,n2188,n2189);
and (n2219,n174,n133);
and (n2220,n2221,n2222);
xor (n2221,n2218,n2219);
or (n2222,n2223,n2226);
and (n2223,n2224,n2225);
xor (n2224,n2194,n2195);
and (n2225,n221,n133);
and (n2226,n2227,n2228);
xor (n2227,n2224,n2225);
and (n2228,n2229,n2230);
xor (n2229,n2200,n2201);
and (n2230,n203,n133);
and (n2231,n387,n154);
or (n2232,n2233,n2236);
and (n2233,n2234,n2235);
xor (n2234,n2209,n2210);
and (n2235,n183,n154);
and (n2236,n2237,n2238);
xor (n2237,n2234,n2235);
or (n2238,n2239,n2242);
and (n2239,n2240,n2241);
xor (n2240,n2215,n2216);
and (n2241,n174,n154);
and (n2242,n2243,n2244);
xor (n2243,n2240,n2241);
or (n2244,n2245,n2248);
and (n2245,n2246,n2247);
xor (n2246,n2221,n2222);
and (n2247,n221,n154);
and (n2248,n2249,n2250);
xor (n2249,n2246,n2247);
and (n2250,n2251,n463);
xor (n2251,n2227,n2228);
and (n2252,n183,n164);
or (n2253,n2254,n2257);
and (n2254,n2255,n2256);
xor (n2255,n2237,n2238);
and (n2256,n174,n164);
and (n2257,n2258,n2259);
xor (n2258,n2255,n2256);
or (n2259,n2260,n2263);
and (n2260,n2261,n2262);
xor (n2261,n2243,n2244);
and (n2262,n221,n164);
and (n2263,n2264,n2265);
xor (n2264,n2261,n2262);
and (n2265,n2266,n2267);
xor (n2266,n2249,n2250);
and (n2267,n203,n164);
and (n2268,n174,n211);
or (n2269,n2270,n2273);
and (n2270,n2271,n2272);
xor (n2271,n2258,n2259);
and (n2272,n221,n211);
and (n2273,n2274,n2275);
xor (n2274,n2271,n2272);
and (n2275,n2276,n406);
xor (n2276,n2264,n2265);
and (n2277,n221,n194);
and (n2278,n2279,n2280);
xor (n2279,n2274,n2275);
and (n2280,n203,n194);
and (n2281,n203,n739);
endmodule
