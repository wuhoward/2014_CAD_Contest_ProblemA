module top (out,n3,n7,n9,n10,n33,n34,n41,n45,n51
        ,n59,n65,n69,n75,n85,n86,n92,n97,n103,n115
        ,n117,n121,n126,n132,n141,n143,n151,n158,n168,n169
        ,n175,n179,n185,n195,n209,n215,n226,n241,n242,n250
        ,n257,n270,n272,n281,n289,n300,n308,n315,n324,n329
        ,n345,n351,n360,n372,n483,n513,n515,n545,n619,n621
        ,n719,n837,n906,n908,n1141,n1147,n1175,n1187,n1193);
output out;
input n3;
input n7;
input n9;
input n10;
input n33;
input n34;
input n41;
input n45;
input n51;
input n59;
input n65;
input n69;
input n75;
input n85;
input n86;
input n92;
input n97;
input n103;
input n115;
input n117;
input n121;
input n126;
input n132;
input n141;
input n143;
input n151;
input n158;
input n168;
input n169;
input n175;
input n179;
input n185;
input n195;
input n209;
input n215;
input n226;
input n241;
input n242;
input n250;
input n257;
input n270;
input n272;
input n281;
input n289;
input n300;
input n308;
input n315;
input n324;
input n329;
input n345;
input n351;
input n360;
input n372;
input n483;
input n513;
input n515;
input n545;
input n619;
input n621;
input n719;
input n837;
input n906;
input n908;
input n1141;
input n1147;
input n1175;
input n1187;
input n1193;
wire n0;
wire n1;
wire n2;
wire n4;
wire n5;
wire n6;
wire n8;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n24;
wire n25;
wire n26;
wire n27;
wire n28;
wire n29;
wire n30;
wire n31;
wire n32;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n42;
wire n43;
wire n44;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n66;
wire n67;
wire n68;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n93;
wire n94;
wire n95;
wire n96;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n116;
wire n118;
wire n119;
wire n120;
wire n122;
wire n123;
wire n124;
wire n125;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n142;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n176;
wire n177;
wire n178;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n271;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n325;
wire n326;
wire n327;
wire n328;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n514;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n620;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n907;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2988;
wire n2989;
wire n2990;
wire n2991;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2996;
wire n2997;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3003;
wire n3004;
wire n3005;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3010;
wire n3011;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3038;
wire n3039;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
wire n3056;
wire n3057;
wire n3058;
wire n3059;
wire n3060;
wire n3061;
wire n3062;
wire n3063;
wire n3064;
wire n3065;
wire n3066;
wire n3067;
wire n3068;
wire n3069;
wire n3070;
wire n3071;
wire n3072;
wire n3073;
wire n3074;
wire n3075;
wire n3076;
wire n3077;
wire n3078;
wire n3079;
wire n3080;
wire n3081;
wire n3082;
wire n3083;
wire n3084;
wire n3085;
wire n3086;
wire n3087;
wire n3088;
wire n3089;
wire n3090;
wire n3091;
wire n3092;
wire n3093;
wire n3094;
wire n3095;
wire n3096;
wire n3097;
wire n3098;
wire n3099;
wire n3100;
wire n3101;
wire n3102;
wire n3103;
wire n3104;
wire n3105;
wire n3106;
wire n3107;
wire n3108;
wire n3109;
wire n3110;
wire n3111;
wire n3112;
wire n3113;
wire n3114;
wire n3115;
wire n3116;
wire n3117;
wire n3118;
wire n3119;
wire n3120;
wire n3121;
wire n3122;
wire n3123;
wire n3124;
wire n3125;
wire n3126;
wire n3127;
wire n3128;
wire n3129;
wire n3130;
wire n3131;
wire n3132;
wire n3133;
wire n3134;
wire n3135;
wire n3136;
wire n3137;
wire n3138;
wire n3139;
wire n3140;
wire n3141;
wire n3142;
wire n3143;
wire n3144;
wire n3145;
wire n3146;
wire n3147;
wire n3148;
wire n3149;
wire n3150;
wire n3151;
wire n3152;
wire n3153;
wire n3154;
wire n3155;
wire n3156;
wire n3157;
wire n3158;
wire n3159;
wire n3160;
wire n3161;
wire n3162;
wire n3163;
wire n3164;
wire n3165;
wire n3166;
wire n3167;
wire n3168;
wire n3169;
wire n3170;
wire n3171;
wire n3172;
wire n3173;
wire n3174;
wire n3175;
wire n3176;
wire n3177;
wire n3178;
wire n3179;
wire n3180;
wire n3181;
wire n3182;
wire n3183;
wire n3184;
wire n3185;
wire n3186;
wire n3187;
wire n3188;
wire n3189;
wire n3190;
wire n3191;
wire n3192;
wire n3193;
wire n3194;
wire n3195;
wire n3196;
wire n3197;
wire n3198;
wire n3199;
wire n3200;
wire n3201;
wire n3202;
wire n3203;
wire n3204;
wire n3205;
wire n3206;
wire n3207;
wire n3208;
wire n3209;
wire n3210;
wire n3211;
wire n3212;
wire n3213;
wire n3214;
wire n3215;
wire n3216;
wire n3217;
wire n3218;
wire n3219;
wire n3220;
wire n3221;
wire n3222;
wire n3223;
wire n3224;
wire n3225;
wire n3226;
wire n3227;
wire n3228;
wire n3229;
wire n3230;
wire n3231;
wire n3232;
wire n3233;
wire n3234;
wire n3235;
wire n3236;
wire n3237;
wire n3238;
wire n3239;
wire n3240;
wire n3241;
wire n3242;
wire n3243;
wire n3244;
wire n3245;
wire n3246;
wire n3247;
wire n3248;
wire n3249;
wire n3250;
wire n3251;
wire n3252;
wire n3253;
wire n3254;
wire n3255;
wire n3256;
wire n3257;
wire n3258;
wire n3259;
wire n3260;
wire n3261;
wire n3262;
wire n3263;
wire n3264;
wire n3265;
wire n3266;
wire n3267;
wire n3268;
wire n3269;
wire n3270;
wire n3271;
wire n3272;
wire n3273;
wire n3274;
wire n3275;
wire n3276;
wire n3277;
wire n3278;
wire n3279;
wire n3280;
wire n3281;
wire n3282;
wire n3283;
wire n3284;
wire n3285;
wire n3286;
wire n3287;
wire n3288;
wire n3289;
wire n3290;
wire n3291;
wire n3292;
wire n3293;
wire n3294;
wire n3295;
wire n3296;
wire n3297;
wire n3298;
wire n3299;
wire n3300;
wire n3301;
wire n3302;
wire n3303;
wire n3304;
wire n3305;
wire n3306;
wire n3307;
wire n3308;
wire n3309;
wire n3310;
wire n3311;
wire n3312;
wire n3313;
wire n3314;
wire n3315;
wire n3316;
wire n3317;
wire n3318;
wire n3319;
wire n3320;
wire n3321;
wire n3322;
wire n3323;
wire n3324;
wire n3325;
wire n3326;
wire n3327;
wire n3328;
wire n3329;
wire n3330;
wire n3331;
wire n3332;
wire n3333;
wire n3334;
wire n3335;
wire n3336;
wire n3337;
wire n3338;
wire n3339;
wire n3340;
wire n3341;
wire n3342;
wire n3343;
wire n3344;
wire n3345;
wire n3346;
wire n3347;
wire n3348;
wire n3349;
wire n3350;
wire n3351;
wire n3352;
wire n3353;
wire n3354;
wire n3355;
wire n3356;
wire n3357;
wire n3358;
wire n3359;
wire n3360;
wire n3361;
wire n3362;
wire n3363;
wire n3364;
wire n3365;
wire n3366;
wire n3367;
wire n3368;
wire n3369;
wire n3370;
wire n3371;
wire n3372;
wire n3373;
wire n3374;
wire n3375;
wire n3376;
wire n3377;
wire n3378;
wire n3379;
wire n3380;
wire n3381;
wire n3382;
wire n3383;
wire n3384;
wire n3385;
wire n3386;
wire n3387;
wire n3388;
wire n3389;
wire n3390;
wire n3391;
wire n3392;
wire n3393;
wire n3394;
wire n3395;
wire n3396;
wire n3397;
wire n3398;
wire n3399;
wire n3400;
wire n3401;
wire n3402;
wire n3403;
wire n3404;
wire n3405;
wire n3406;
wire n3407;
wire n3408;
wire n3409;
wire n3410;
wire n3411;
wire n3412;
wire n3413;
wire n3414;
wire n3415;
wire n3416;
wire n3417;
wire n3418;
wire n3419;
wire n3420;
wire n3421;
wire n3422;
wire n3423;
wire n3424;
wire n3425;
wire n3426;
wire n3427;
wire n3428;
wire n3429;
wire n3430;
wire n3431;
wire n3432;
wire n3433;
wire n3434;
wire n3435;
wire n3436;
wire n3437;
wire n3438;
wire n3439;
wire n3440;
wire n3441;
wire n3442;
wire n3443;
wire n3444;
wire n3445;
wire n3446;
wire n3447;
wire n3448;
wire n3449;
wire n3450;
wire n3451;
wire n3452;
wire n3453;
wire n3454;
wire n3455;
wire n3456;
wire n3457;
wire n3458;
wire n3459;
wire n3460;
wire n3461;
wire n3462;
wire n3463;
wire n3464;
wire n3465;
wire n3466;
wire n3467;
wire n3468;
wire n3469;
wire n3470;
wire n3471;
wire n3472;
wire n3473;
wire n3474;
wire n3475;
wire n3476;
wire n3477;
wire n3478;
wire n3479;
wire n3480;
wire n3481;
wire n3482;
wire n3483;
wire n3484;
wire n3485;
wire n3486;
wire n3487;
wire n3488;
wire n3489;
wire n3490;
wire n3491;
wire n3492;
wire n3493;
wire n3494;
wire n3495;
wire n3496;
wire n3497;
wire n3498;
wire n3499;
wire n3500;
wire n3501;
wire n3502;
wire n3503;
wire n3504;
wire n3505;
wire n3506;
wire n3507;
wire n3508;
wire n3509;
wire n3510;
wire n3511;
wire n3512;
wire n3513;
wire n3514;
wire n3515;
wire n3516;
wire n3517;
wire n3518;
wire n3519;
wire n3520;
wire n3521;
wire n3522;
wire n3523;
wire n3524;
wire n3525;
wire n3526;
wire n3527;
wire n3528;
wire n3529;
wire n3530;
wire n3531;
wire n3532;
wire n3533;
wire n3534;
wire n3535;
wire n3536;
wire n3537;
wire n3538;
wire n3539;
wire n3540;
wire n3541;
wire n3542;
wire n3543;
wire n3544;
wire n3545;
wire n3546;
wire n3547;
wire n3548;
wire n3549;
wire n3550;
wire n3551;
wire n3552;
wire n3553;
wire n3554;
wire n3555;
wire n3556;
wire n3557;
wire n3558;
wire n3559;
wire n3560;
wire n3561;
wire n3562;
wire n3563;
wire n3564;
wire n3565;
wire n3566;
wire n3567;
wire n3568;
wire n3569;
wire n3570;
wire n3571;
wire n3572;
wire n3573;
wire n3574;
wire n3575;
wire n3576;
wire n3577;
wire n3578;
wire n3579;
wire n3580;
wire n3581;
wire n3582;
wire n3583;
wire n3584;
wire n3585;
wire n3586;
wire n3587;
wire n3588;
wire n3589;
wire n3590;
wire n3591;
wire n3592;
wire n3593;
wire n3594;
wire n3595;
wire n3596;
wire n3597;
wire n3598;
wire n3599;
wire n3600;
wire n3601;
wire n3602;
wire n3603;
wire n3604;
wire n3605;
wire n3606;
wire n3607;
wire n3608;
wire n3609;
wire n3610;
wire n3611;
wire n3612;
wire n3613;
wire n3614;
wire n3615;
wire n3616;
wire n3617;
wire n3618;
wire n3619;
wire n3620;
wire n3621;
wire n3622;
wire n3623;
wire n3624;
wire n3625;
wire n3626;
wire n3627;
wire n3628;
wire n3629;
wire n3630;
wire n3631;
wire n3632;
wire n3633;
wire n3634;
wire n3635;
wire n3636;
wire n3637;
wire n3638;
wire n3639;
wire n3640;
wire n3641;
wire n3642;
wire n3643;
wire n3644;
wire n3645;
wire n3646;
wire n3647;
wire n3648;
wire n3649;
wire n3650;
wire n3651;
wire n3652;
wire n3653;
wire n3654;
wire n3655;
wire n3656;
wire n3657;
wire n3658;
wire n3659;
wire n3660;
wire n3661;
wire n3662;
wire n3663;
wire n3664;
wire n3665;
wire n3666;
wire n3667;
wire n3668;
wire n3669;
wire n3670;
wire n3671;
wire n3672;
wire n3673;
wire n3674;
wire n3675;
wire n3676;
wire n3677;
wire n3678;
wire n3679;
wire n3680;
wire n3681;
wire n3682;
wire n3683;
wire n3684;
wire n3685;
wire n3686;
wire n3687;
wire n3688;
wire n3689;
wire n3690;
wire n3691;
wire n3692;
wire n3693;
wire n3694;
wire n3695;
wire n3696;
wire n3697;
wire n3698;
wire n3699;
wire n3700;
wire n3701;
wire n3702;
wire n3703;
wire n3704;
wire n3705;
wire n3706;
wire n3707;
wire n3708;
wire n3709;
wire n3710;
wire n3711;
wire n3712;
wire n3713;
wire n3714;
wire n3715;
wire n3716;
wire n3717;
wire n3718;
wire n3719;
wire n3720;
wire n3721;
wire n3722;
wire n3723;
wire n3724;
wire n3725;
wire n3726;
wire n3727;
wire n3728;
wire n3729;
wire n3730;
wire n3731;
wire n3732;
wire n3733;
wire n3734;
wire n3735;
wire n3736;
wire n3737;
wire n3738;
wire n3739;
wire n3740;
wire n3741;
wire n3742;
wire n3743;
wire n3744;
wire n3745;
wire n3746;
wire n3747;
wire n3748;
wire n3749;
wire n3750;
wire n3751;
wire n3752;
wire n3753;
wire n3754;
wire n3755;
wire n3756;
wire n3757;
wire n3758;
wire n3759;
wire n3760;
wire n3761;
wire n3762;
wire n3763;
wire n3764;
wire n3765;
wire n3766;
wire n3767;
wire n3768;
wire n3769;
wire n3770;
wire n3771;
wire n3772;
wire n3773;
wire n3774;
wire n3775;
wire n3776;
wire n3777;
wire n3778;
wire n3779;
wire n3780;
wire n3781;
wire n3782;
wire n3783;
wire n3784;
wire n3785;
wire n3786;
wire n3787;
wire n3788;
wire n3789;
wire n3790;
wire n3791;
wire n3792;
wire n3793;
wire n3794;
wire n3795;
wire n3796;
wire n3797;
wire n3798;
wire n3799;
wire n3800;
wire n3801;
wire n3802;
wire n3803;
wire n3804;
wire n3805;
wire n3806;
wire n3807;
wire n3808;
wire n3809;
wire n3810;
wire n3811;
wire n3812;
wire n3813;
wire n3814;
wire n3815;
wire n3816;
wire n3817;
wire n3818;
wire n3819;
wire n3820;
wire n3821;
wire n3822;
wire n3823;
wire n3824;
wire n3825;
wire n3826;
wire n3827;
wire n3828;
wire n3829;
wire n3830;
wire n3831;
wire n3832;
wire n3833;
wire n3834;
wire n3835;
wire n3836;
wire n3837;
wire n3838;
wire n3839;
wire n3840;
wire n3841;
wire n3842;
wire n3843;
wire n3844;
wire n3845;
wire n3846;
wire n3847;
wire n3848;
wire n3849;
wire n3850;
wire n3851;
wire n3852;
wire n3853;
wire n3854;
wire n3855;
wire n3856;
wire n3857;
wire n3858;
wire n3859;
wire n3860;
wire n3861;
wire n3862;
wire n3863;
wire n3864;
wire n3865;
wire n3866;
wire n3867;
wire n3868;
wire n3869;
wire n3870;
wire n3871;
wire n3872;
wire n3873;
wire n3874;
wire n3875;
wire n3876;
wire n3877;
wire n3878;
wire n3879;
wire n3880;
wire n3881;
wire n3882;
wire n3883;
wire n3884;
wire n3885;
wire n3886;
wire n3887;
wire n3888;
wire n3889;
wire n3890;
wire n3891;
wire n3892;
wire n3893;
wire n3894;
wire n3895;
wire n3896;
wire n3897;
wire n3898;
wire n3899;
wire n3900;
wire n3901;
wire n3902;
wire n3903;
wire n3904;
wire n3905;
wire n3906;
wire n3907;
wire n3908;
wire n3909;
wire n3910;
wire n3911;
wire n3912;
wire n3913;
wire n3914;
wire n3915;
wire n3916;
wire n3917;
wire n3918;
wire n3919;
wire n3920;
wire n3921;
wire n3922;
wire n3923;
wire n3924;
wire n3925;
wire n3926;
wire n3927;
wire n3928;
wire n3929;
wire n3930;
wire n3931;
wire n3932;
wire n3933;
wire n3934;
wire n3935;
wire n3936;
wire n3937;
wire n3938;
wire n3939;
wire n3940;
wire n3941;
wire n3942;
wire n3943;
wire n3944;
wire n3945;
wire n3946;
wire n3947;
wire n3948;
wire n3949;
wire n3950;
wire n3951;
wire n3952;
wire n3953;
wire n3954;
wire n3955;
wire n3956;
wire n3957;
wire n3958;
wire n3959;
wire n3960;
wire n3961;
wire n3962;
wire n3963;
wire n3964;
wire n3965;
wire n3966;
wire n3967;
wire n3968;
wire n3969;
wire n3970;
wire n3971;
wire n3972;
wire n3973;
wire n3974;
wire n3975;
wire n3976;
wire n3977;
wire n3978;
wire n3979;
wire n3980;
wire n3981;
wire n3982;
wire n3983;
wire n3984;
wire n3985;
wire n3986;
wire n3987;
wire n3988;
wire n3989;
wire n3990;
wire n3991;
wire n3992;
wire n3993;
wire n3994;
wire n3995;
wire n3996;
wire n3997;
wire n3998;
wire n3999;
wire n4000;
wire n4001;
wire n4002;
wire n4003;
wire n4004;
wire n4005;
wire n4006;
wire n4007;
wire n4008;
wire n4009;
wire n4010;
wire n4011;
wire n4012;
wire n4013;
wire n4014;
wire n4015;
wire n4016;
wire n4017;
wire n4018;
wire n4019;
wire n4020;
wire n4021;
wire n4022;
wire n4023;
wire n4024;
wire n4025;
wire n4026;
wire n4027;
wire n4028;
wire n4029;
wire n4030;
wire n4031;
wire n4032;
wire n4033;
wire n4034;
wire n4035;
wire n4036;
wire n4037;
wire n4038;
wire n4039;
wire n4040;
wire n4041;
wire n4042;
wire n4043;
wire n4044;
wire n4045;
wire n4046;
wire n4047;
wire n4048;
wire n4049;
wire n4050;
wire n4051;
wire n4052;
wire n4053;
wire n4054;
wire n4055;
wire n4056;
wire n4057;
wire n4058;
wire n4059;
wire n4060;
wire n4061;
wire n4062;
wire n4063;
wire n4064;
wire n4065;
wire n4066;
wire n4067;
wire n4068;
wire n4069;
wire n4070;
wire n4071;
wire n4072;
wire n4073;
wire n4074;
wire n4075;
wire n4076;
wire n4077;
wire n4078;
wire n4079;
wire n4080;
wire n4081;
wire n4082;
wire n4083;
wire n4084;
wire n4085;
wire n4086;
wire n4087;
wire n4088;
wire n4089;
wire n4090;
wire n4091;
wire n4092;
wire n4093;
wire n4094;
wire n4095;
wire n4096;
wire n4097;
wire n4098;
wire n4099;
wire n4100;
wire n4101;
wire n4102;
wire n4103;
wire n4104;
wire n4105;
wire n4106;
wire n4107;
wire n4108;
wire n4109;
wire n4110;
wire n4111;
wire n4112;
wire n4113;
wire n4114;
wire n4115;
wire n4116;
wire n4117;
wire n4118;
wire n4119;
wire n4120;
wire n4121;
wire n4122;
wire n4123;
wire n4124;
wire n4125;
wire n4126;
wire n4127;
wire n4128;
wire n4129;
wire n4130;
wire n4131;
wire n4132;
wire n4133;
wire n4134;
wire n4135;
wire n4136;
wire n4137;
wire n4138;
wire n4139;
wire n4140;
wire n4141;
wire n4142;
wire n4143;
wire n4144;
wire n4145;
wire n4146;
wire n4147;
wire n4148;
wire n4149;
wire n4150;
wire n4151;
wire n4152;
wire n4153;
wire n4154;
wire n4155;
wire n4156;
wire n4157;
wire n4158;
wire n4159;
wire n4160;
wire n4161;
wire n4162;
wire n4163;
wire n4164;
wire n4165;
wire n4166;
wire n4167;
wire n4168;
wire n4169;
wire n4170;
wire n4171;
wire n4172;
wire n4173;
wire n4174;
wire n4175;
wire n4176;
wire n4177;
wire n4178;
wire n4179;
wire n4180;
wire n4181;
wire n4182;
wire n4183;
wire n4184;
wire n4185;
wire n4186;
wire n4187;
wire n4188;
wire n4189;
wire n4190;
wire n4191;
wire n4192;
wire n4193;
wire n4194;
wire n4195;
wire n4196;
wire n4197;
wire n4198;
wire n4199;
wire n4200;
wire n4201;
wire n4202;
wire n4203;
wire n4204;
wire n4205;
wire n4206;
wire n4207;
wire n4208;
wire n4209;
wire n4210;
wire n4211;
wire n4212;
wire n4213;
wire n4214;
wire n4215;
wire n4216;
wire n4217;
wire n4218;
wire n4219;
wire n4220;
wire n4221;
wire n4222;
wire n4223;
wire n4224;
wire n4225;
wire n4226;
wire n4227;
wire n4228;
wire n4229;
wire n4230;
wire n4231;
wire n4232;
wire n4233;
wire n4234;
wire n4235;
wire n4236;
wire n4237;
wire n4238;
wire n4239;
wire n4240;
wire n4241;
wire n4242;
wire n4243;
wire n4244;
wire n4245;
wire n4246;
wire n4247;
wire n4248;
wire n4249;
wire n4250;
wire n4251;
wire n4252;
wire n4253;
wire n4254;
wire n4255;
wire n4256;
wire n4257;
wire n4258;
wire n4259;
wire n4260;
wire n4261;
wire n4262;
wire n4263;
wire n4264;
wire n4265;
wire n4266;
wire n4267;
wire n4268;
wire n4269;
wire n4270;
wire n4271;
wire n4272;
wire n4273;
wire n4274;
wire n4275;
wire n4276;
wire n4277;
wire n4278;
wire n4279;
wire n4280;
wire n4281;
wire n4282;
wire n4283;
wire n4284;
wire n4285;
wire n4286;
wire n4287;
wire n4288;
wire n4289;
wire n4290;
wire n4291;
wire n4292;
wire n4293;
wire n4294;
wire n4295;
wire n4296;
wire n4297;
wire n4298;
wire n4299;
wire n4300;
wire n4301;
wire n4302;
wire n4303;
wire n4304;
wire n4305;
wire n4306;
wire n4307;
wire n4308;
wire n4309;
wire n4310;
wire n4311;
wire n4312;
wire n4313;
wire n4314;
wire n4315;
wire n4316;
wire n4317;
wire n4318;
wire n4319;
wire n4320;
wire n4321;
wire n4322;
wire n4323;
wire n4324;
wire n4325;
wire n4326;
wire n4327;
wire n4328;
wire n4329;
wire n4330;
wire n4331;
wire n4332;
wire n4333;
wire n4334;
wire n4335;
wire n4336;
wire n4337;
wire n4338;
wire n4339;
wire n4340;
wire n4341;
wire n4342;
wire n4343;
wire n4344;
wire n4345;
wire n4346;
wire n4347;
wire n4348;
wire n4349;
wire n4350;
wire n4351;
wire n4352;
wire n4353;
wire n4354;
wire n4355;
wire n4356;
wire n4357;
wire n4358;
wire n4359;
wire n4360;
wire n4361;
wire n4362;
wire n4363;
wire n4364;
wire n4365;
wire n4366;
wire n4367;
wire n4368;
wire n4369;
wire n4370;
wire n4371;
wire n4372;
wire n4373;
wire n4374;
wire n4375;
wire n4376;
wire n4377;
wire n4378;
wire n4379;
wire n4380;
wire n4381;
wire n4382;
wire n4383;
wire n4384;
wire n4385;
wire n4386;
wire n4387;
wire n4388;
wire n4389;
wire n4390;
wire n4391;
wire n4392;
wire n4393;
wire n4394;
wire n4395;
wire n4396;
wire n4397;
wire n4398;
wire n4399;
wire n4400;
wire n4401;
wire n4402;
wire n4403;
wire n4404;
wire n4405;
wire n4406;
wire n4407;
wire n4408;
wire n4409;
wire n4410;
wire n4411;
wire n4412;
wire n4413;
wire n4414;
wire n4415;
wire n4416;
wire n4417;
wire n4418;
wire n4419;
wire n4420;
wire n4421;
wire n4422;
wire n4423;
wire n4424;
wire n4425;
wire n4426;
wire n4427;
wire n4428;
wire n4429;
wire n4430;
wire n4431;
wire n4432;
wire n4433;
wire n4434;
wire n4435;
wire n4436;
wire n4437;
wire n4438;
wire n4439;
wire n4440;
wire n4441;
wire n4442;
wire n4443;
wire n4444;
wire n4445;
wire n4446;
wire n4447;
wire n4448;
wire n4449;
wire n4450;
wire n4451;
wire n4452;
wire n4453;
wire n4454;
wire n4455;
wire n4456;
wire n4457;
wire n4458;
wire n4459;
wire n4460;
wire n4461;
wire n4462;
wire n4463;
wire n4464;
wire n4465;
wire n4466;
wire n4467;
wire n4468;
wire n4469;
wire n4470;
wire n4471;
wire n4472;
wire n4473;
wire n4474;
wire n4475;
wire n4476;
wire n4477;
wire n4478;
wire n4479;
wire n4480;
wire n4481;
wire n4482;
wire n4483;
wire n4484;
wire n4485;
wire n4486;
wire n4487;
wire n4488;
wire n4489;
wire n4490;
wire n4491;
wire n4492;
wire n4493;
wire n4494;
wire n4495;
wire n4496;
wire n4497;
wire n4498;
wire n4499;
wire n4500;
wire n4501;
wire n4502;
wire n4503;
wire n4504;
wire n4505;
wire n4506;
wire n4507;
wire n4508;
wire n4509;
wire n4510;
wire n4511;
wire n4512;
wire n4513;
wire n4514;
wire n4515;
wire n4516;
wire n4517;
wire n4518;
wire n4519;
wire n4520;
wire n4521;
wire n4522;
wire n4523;
wire n4524;
wire n4525;
wire n4526;
wire n4527;
wire n4528;
wire n4529;
wire n4530;
wire n4531;
wire n4532;
wire n4533;
wire n4534;
wire n4535;
wire n4536;
wire n4537;
wire n4538;
wire n4539;
wire n4540;
wire n4541;
wire n4542;
wire n4543;
wire n4544;
wire n4545;
wire n4546;
wire n4547;
wire n4548;
wire n4549;
wire n4550;
wire n4551;
wire n4552;
wire n4553;
wire n4554;
wire n4555;
wire n4556;
wire n4557;
wire n4558;
wire n4559;
wire n4560;
wire n4561;
wire n4562;
wire n4563;
wire n4564;
wire n4565;
wire n4566;
wire n4567;
wire n4568;
wire n4569;
wire n4570;
wire n4571;
wire n4572;
wire n4573;
wire n4574;
wire n4575;
wire n4576;
wire n4577;
wire n4578;
wire n4579;
wire n4580;
wire n4581;
wire n4582;
wire n4583;
wire n4584;
wire n4585;
wire n4586;
wire n4587;
wire n4588;
wire n4589;
wire n4590;
wire n4591;
wire n4592;
wire n4593;
wire n4594;
wire n4595;
wire n4596;
wire n4597;
wire n4598;
wire n4599;
wire n4600;
wire n4601;
wire n4602;
wire n4603;
wire n4604;
wire n4605;
wire n4606;
wire n4607;
wire n4608;
wire n4609;
wire n4610;
wire n4611;
wire n4612;
wire n4613;
wire n4614;
wire n4615;
wire n4616;
wire n4617;
wire n4618;
wire n4619;
wire n4620;
wire n4621;
wire n4622;
wire n4623;
wire n4624;
wire n4625;
wire n4626;
wire n4627;
wire n4628;
wire n4629;
wire n4630;
wire n4631;
wire n4632;
wire n4633;
wire n4634;
wire n4635;
wire n4636;
wire n4637;
wire n4638;
wire n4639;
wire n4640;
wire n4641;
wire n4642;
wire n4643;
wire n4644;
wire n4645;
wire n4646;
wire n4647;
wire n4648;
wire n4649;
wire n4650;
wire n4651;
wire n4652;
wire n4653;
wire n4654;
wire n4655;
wire n4656;
wire n4657;
wire n4658;
wire n4659;
wire n4660;
wire n4661;
wire n4662;
wire n4663;
wire n4664;
wire n4665;
wire n4666;
wire n4667;
wire n4668;
wire n4669;
wire n4670;
wire n4671;
wire n4672;
wire n4673;
wire n4674;
wire n4675;
wire n4676;
wire n4677;
wire n4678;
wire n4679;
wire n4680;
wire n4681;
wire n4682;
wire n4683;
wire n4684;
wire n4685;
wire n4686;
wire n4687;
wire n4688;
wire n4689;
wire n4690;
wire n4691;
wire n4692;
wire n4693;
wire n4694;
wire n4695;
wire n4696;
wire n4697;
wire n4698;
wire n4699;
wire n4700;
wire n4701;
wire n4702;
wire n4703;
wire n4704;
wire n4705;
wire n4706;
wire n4707;
wire n4708;
wire n4709;
wire n4710;
wire n4711;
wire n4712;
wire n4713;
wire n4714;
wire n4715;
wire n4716;
wire n4717;
wire n4718;
wire n4719;
wire n4720;
wire n4721;
wire n4722;
wire n4723;
wire n4724;
wire n4725;
wire n4726;
wire n4727;
wire n4728;
wire n4729;
wire n4730;
wire n4731;
wire n4732;
wire n4733;
wire n4734;
wire n4735;
wire n4736;
wire n4737;
wire n4738;
wire n4739;
wire n4740;
wire n4741;
wire n4742;
wire n4743;
wire n4744;
wire n4745;
wire n4746;
wire n4747;
wire n4748;
wire n4749;
wire n4750;
wire n4751;
wire n4752;
wire n4753;
wire n4754;
wire n4755;
wire n4756;
wire n4757;
wire n4758;
wire n4759;
wire n4760;
wire n4761;
wire n4762;
wire n4763;
wire n4764;
wire n4765;
wire n4766;
wire n4767;
wire n4768;
wire n4769;
wire n4770;
wire n4771;
wire n4772;
wire n4773;
wire n4774;
wire n4775;
wire n4776;
wire n4777;
wire n4778;
wire n4779;
wire n4780;
wire n4781;
wire n4782;
wire n4783;
wire n4784;
wire n4785;
wire n4786;
wire n4787;
wire n4788;
wire n4789;
wire n4790;
wire n4791;
wire n4792;
wire n4793;
wire n4794;
wire n4795;
wire n4796;
wire n4797;
wire n4798;
wire n4799;
wire n4800;
wire n4801;
wire n4802;
wire n4803;
wire n4804;
wire n4805;
wire n4806;
wire n4807;
wire n4808;
wire n4809;
wire n4810;
wire n4811;
wire n4812;
wire n4813;
wire n4814;
wire n4815;
wire n4816;
wire n4817;
wire n4818;
wire n4819;
wire n4820;
wire n4821;
wire n4822;
wire n4823;
wire n4824;
wire n4825;
wire n4826;
wire n4827;
wire n4828;
wire n4829;
wire n4830;
wire n4831;
wire n4832;
wire n4833;
wire n4834;
wire n4835;
wire n4836;
wire n4837;
wire n4838;
wire n4839;
wire n4840;
wire n4841;
wire n4842;
wire n4843;
wire n4844;
wire n4845;
wire n4846;
wire n4847;
wire n4848;
wire n4849;
wire n4850;
wire n4851;
wire n4852;
wire n4853;
wire n4854;
wire n4855;
wire n4856;
wire n4857;
wire n4858;
wire n4859;
wire n4860;
wire n4861;
wire n4862;
wire n4863;
wire n4864;
wire n4865;
wire n4866;
wire n4867;
wire n4868;
wire n4869;
wire n4870;
wire n4871;
wire n4872;
wire n4873;
wire n4874;
wire n4875;
wire n4876;
wire n4877;
wire n4878;
wire n4879;
wire n4880;
wire n4881;
wire n4882;
wire n4883;
wire n4884;
wire n4885;
wire n4886;
wire n4887;
wire n4888;
wire n4889;
wire n4890;
wire n4891;
wire n4892;
wire n4893;
wire n4894;
wire n4895;
wire n4896;
wire n4897;
wire n4898;
wire n4899;
wire n4900;
wire n4901;
wire n4902;
wire n4903;
wire n4904;
wire n4905;
wire n4906;
wire n4907;
wire n4908;
wire n4909;
wire n4910;
wire n4911;
wire n4912;
wire n4913;
wire n4914;
wire n4915;
wire n4916;
wire n4917;
wire n4918;
wire n4919;
wire n4920;
wire n4921;
wire n4922;
wire n4923;
wire n4924;
wire n4925;
wire n4926;
wire n4927;
wire n4928;
wire n4929;
wire n4930;
wire n4931;
wire n4932;
wire n4933;
wire n4934;
wire n4935;
wire n4936;
wire n4937;
wire n4938;
wire n4939;
wire n4940;
wire n4941;
wire n4942;
wire n4943;
wire n4944;
wire n4945;
wire n4946;
wire n4947;
wire n4948;
wire n4949;
wire n4950;
wire n4951;
wire n4952;
wire n4953;
wire n4954;
wire n4955;
wire n4956;
wire n4957;
wire n4958;
wire n4959;
wire n4960;
wire n4961;
wire n4962;
wire n4963;
wire n4964;
wire n4965;
wire n4966;
wire n4967;
wire n4968;
wire n4969;
wire n4970;
wire n4971;
wire n4972;
wire n4973;
wire n4974;
wire n4975;
wire n4976;
wire n4977;
wire n4978;
wire n4979;
wire n4980;
wire n4981;
wire n4982;
wire n4983;
wire n4984;
wire n4985;
wire n4986;
wire n4987;
wire n4988;
wire n4989;
wire n4990;
wire n4991;
wire n4992;
wire n4993;
wire n4994;
wire n4995;
wire n4996;
wire n4997;
wire n4998;
wire n4999;
wire n5000;
wire n5001;
wire n5002;
wire n5003;
wire n5004;
wire n5005;
wire n5006;
wire n5007;
wire n5008;
wire n5009;
wire n5010;
wire n5011;
wire n5012;
wire n5013;
wire n5014;
wire n5015;
wire n5016;
wire n5017;
wire n5018;
wire n5019;
wire n5020;
wire n5021;
wire n5022;
wire n5023;
wire n5024;
wire n5025;
wire n5026;
wire n5027;
wire n5028;
wire n5029;
wire n5030;
wire n5031;
wire n5032;
wire n5033;
wire n5034;
wire n5035;
wire n5036;
wire n5037;
wire n5038;
wire n5039;
wire n5040;
wire n5041;
wire n5042;
wire n5043;
wire n5044;
wire n5045;
wire n5046;
wire n5047;
wire n5048;
wire n5049;
wire n5050;
wire n5051;
wire n5052;
wire n5053;
wire n5054;
wire n5055;
wire n5056;
wire n5057;
wire n5058;
wire n5059;
wire n5060;
wire n5061;
wire n5062;
wire n5063;
wire n5064;
wire n5065;
wire n5066;
wire n5067;
wire n5068;
wire n5069;
wire n5070;
wire n5071;
wire n5072;
wire n5073;
wire n5074;
wire n5075;
wire n5076;
wire n5077;
wire n5078;
wire n5079;
wire n5080;
wire n5081;
wire n5082;
wire n5083;
wire n5084;
wire n5085;
wire n5086;
wire n5087;
wire n5088;
wire n5089;
wire n5090;
wire n5091;
wire n5092;
wire n5093;
wire n5094;
wire n5095;
wire n5096;
wire n5097;
wire n5098;
wire n5099;
wire n5100;
wire n5101;
wire n5102;
wire n5103;
wire n5104;
wire n5105;
wire n5106;
wire n5107;
wire n5108;
wire n5109;
wire n5110;
wire n5111;
wire n5112;
wire n5113;
wire n5114;
wire n5115;
wire n5116;
wire n5117;
wire n5118;
wire n5119;
wire n5120;
wire n5121;
wire n5122;
wire n5123;
wire n5124;
wire n5125;
wire n5126;
wire n5127;
wire n5128;
wire n5129;
wire n5130;
wire n5131;
wire n5132;
wire n5133;
wire n5134;
wire n5135;
wire n5136;
wire n5137;
wire n5138;
wire n5139;
wire n5140;
wire n5141;
wire n5142;
wire n5143;
wire n5144;
wire n5145;
wire n5146;
wire n5147;
wire n5148;
wire n5149;
wire n5150;
wire n5151;
wire n5152;
wire n5153;
wire n5154;
wire n5155;
wire n5156;
wire n5157;
wire n5158;
wire n5159;
wire n5160;
wire n5161;
wire n5162;
wire n5163;
wire n5164;
wire n5165;
wire n5166;
wire n5167;
wire n5168;
wire n5169;
wire n5170;
wire n5171;
wire n5172;
wire n5173;
wire n5174;
wire n5175;
wire n5176;
wire n5177;
wire n5178;
wire n5179;
wire n5180;
wire n5181;
wire n5182;
wire n5183;
wire n5184;
wire n5185;
wire n5186;
wire n5187;
wire n5188;
wire n5189;
wire n5190;
wire n5191;
wire n5192;
wire n5193;
wire n5194;
wire n5195;
wire n5196;
wire n5197;
wire n5198;
wire n5199;
wire n5200;
wire n5201;
wire n5202;
wire n5203;
wire n5204;
wire n5205;
wire n5206;
wire n5207;
wire n5208;
wire n5209;
wire n5210;
wire n5211;
wire n5212;
wire n5213;
wire n5214;
wire n5215;
wire n5216;
wire n5217;
wire n5218;
wire n5219;
wire n5220;
wire n5221;
wire n5222;
wire n5223;
wire n5224;
wire n5225;
wire n5226;
wire n5227;
wire n5228;
wire n5229;
wire n5230;
wire n5231;
wire n5232;
wire n5233;
wire n5234;
wire n5235;
wire n5236;
wire n5237;
wire n5238;
wire n5239;
wire n5240;
wire n5241;
wire n5242;
wire n5243;
wire n5244;
wire n5245;
wire n5246;
wire n5247;
wire n5248;
wire n5249;
wire n5250;
wire n5251;
wire n5252;
wire n5253;
wire n5254;
wire n5255;
wire n5256;
wire n5257;
wire n5258;
wire n5259;
wire n5260;
wire n5261;
wire n5262;
wire n5263;
wire n5264;
wire n5265;
wire n5266;
wire n5267;
wire n5268;
wire n5269;
wire n5270;
wire n5271;
wire n5272;
wire n5273;
wire n5274;
wire n5275;
wire n5276;
wire n5277;
wire n5278;
wire n5279;
wire n5280;
wire n5281;
wire n5282;
wire n5283;
wire n5284;
wire n5285;
wire n5286;
wire n5287;
wire n5288;
wire n5289;
wire n5290;
wire n5291;
wire n5292;
wire n5293;
wire n5294;
wire n5295;
wire n5296;
wire n5297;
wire n5298;
wire n5299;
wire n5300;
wire n5301;
wire n5302;
wire n5303;
wire n5304;
wire n5305;
wire n5306;
wire n5307;
wire n5308;
wire n5309;
wire n5310;
wire n5311;
wire n5312;
wire n5313;
wire n5314;
wire n5315;
wire n5316;
wire n5317;
wire n5318;
wire n5319;
wire n5320;
wire n5321;
wire n5322;
wire n5323;
wire n5324;
wire n5325;
wire n5326;
wire n5327;
wire n5328;
wire n5329;
wire n5330;
wire n5331;
wire n5332;
wire n5333;
wire n5334;
wire n5335;
wire n5336;
wire n5337;
wire n5338;
wire n5339;
wire n5340;
wire n5341;
wire n5342;
wire n5343;
wire n5344;
wire n5345;
wire n5346;
wire n5347;
wire n5348;
wire n5349;
wire n5350;
wire n5351;
wire n5352;
wire n5353;
wire n5354;
wire n5355;
wire n5356;
wire n5357;
wire n5358;
wire n5359;
wire n5360;
wire n5361;
wire n5362;
wire n5363;
wire n5364;
wire n5365;
wire n5366;
wire n5367;
wire n5368;
wire n5369;
wire n5370;
wire n5371;
wire n5372;
wire n5373;
wire n5374;
wire n5375;
wire n5376;
wire n5377;
wire n5378;
wire n5379;
wire n5380;
wire n5381;
wire n5382;
wire n5383;
wire n5384;
wire n5385;
wire n5386;
wire n5387;
wire n5388;
wire n5389;
wire n5390;
wire n5391;
wire n5392;
wire n5393;
wire n5394;
wire n5395;
wire n5396;
wire n5397;
wire n5398;
wire n5399;
wire n5400;
wire n5401;
wire n5402;
wire n5403;
wire n5404;
wire n5405;
wire n5406;
wire n5407;
wire n5408;
wire n5409;
wire n5410;
wire n5411;
wire n5412;
wire n5413;
wire n5414;
wire n5415;
wire n5416;
wire n5417;
wire n5418;
wire n5419;
wire n5420;
wire n5421;
wire n5422;
wire n5423;
wire n5424;
wire n5425;
wire n5426;
wire n5427;
wire n5428;
wire n5429;
wire n5430;
wire n5431;
wire n5432;
wire n5433;
wire n5434;
wire n5435;
wire n5436;
wire n5437;
wire n5438;
wire n5439;
wire n5440;
wire n5441;
wire n5442;
wire n5443;
wire n5444;
wire n5445;
wire n5446;
wire n5447;
wire n5448;
wire n5449;
wire n5450;
wire n5451;
wire n5452;
wire n5453;
wire n5454;
wire n5455;
wire n5456;
wire n5457;
wire n5458;
wire n5459;
wire n5460;
wire n5461;
wire n5462;
wire n5463;
wire n5464;
wire n5465;
wire n5466;
wire n5467;
wire n5468;
wire n5469;
wire n5470;
wire n5471;
wire n5472;
wire n5473;
wire n5474;
wire n5475;
wire n5476;
wire n5477;
wire n5478;
wire n5479;
wire n5480;
wire n5481;
wire n5482;
wire n5483;
wire n5484;
wire n5485;
wire n5486;
wire n5487;
wire n5488;
wire n5489;
wire n5490;
wire n5491;
wire n5492;
wire n5493;
wire n5494;
wire n5495;
wire n5496;
wire n5497;
wire n5498;
wire n5499;
wire n5500;
wire n5501;
wire n5502;
wire n5503;
wire n5504;
wire n5505;
wire n5506;
wire n5507;
wire n5508;
wire n5509;
wire n5510;
wire n5511;
wire n5512;
wire n5513;
wire n5514;
wire n5515;
wire n5516;
wire n5517;
wire n5518;
wire n5519;
wire n5520;
wire n5521;
wire n5522;
wire n5523;
wire n5524;
wire n5525;
wire n5526;
wire n5527;
wire n5528;
wire n5529;
wire n5530;
wire n5531;
wire n5532;
wire n5533;
wire n5534;
wire n5535;
wire n5536;
wire n5537;
wire n5538;
wire n5539;
wire n5540;
wire n5541;
wire n5542;
wire n5543;
wire n5544;
wire n5545;
wire n5546;
wire n5547;
wire n5548;
wire n5549;
wire n5550;
wire n5551;
wire n5552;
wire n5553;
wire n5554;
wire n5555;
wire n5556;
wire n5557;
wire n5558;
wire n5559;
wire n5560;
wire n5561;
wire n5562;
wire n5563;
wire n5564;
wire n5565;
wire n5566;
wire n5567;
wire n5568;
wire n5569;
wire n5570;
wire n5571;
wire n5572;
wire n5573;
wire n5574;
wire n5575;
wire n5576;
wire n5577;
wire n5578;
wire n5579;
wire n5580;
wire n5581;
wire n5582;
wire n5583;
wire n5584;
wire n5585;
wire n5586;
wire n5587;
wire n5588;
wire n5589;
wire n5590;
wire n5591;
wire n5592;
wire n5593;
wire n5594;
wire n5595;
wire n5596;
wire n5597;
wire n5598;
wire n5599;
wire n5600;
wire n5601;
wire n5602;
wire n5603;
wire n5604;
wire n5605;
wire n5606;
wire n5607;
wire n5608;
wire n5609;
wire n5610;
wire n5611;
wire n5612;
wire n5613;
wire n5614;
wire n5615;
wire n5616;
wire n5617;
wire n5618;
wire n5619;
wire n5620;
wire n5621;
wire n5622;
wire n5623;
wire n5624;
wire n5625;
wire n5626;
wire n5627;
wire n5628;
wire n5629;
wire n5630;
wire n5631;
wire n5632;
wire n5633;
wire n5634;
wire n5635;
wire n5636;
wire n5637;
wire n5638;
wire n5639;
wire n5640;
wire n5641;
wire n5642;
wire n5643;
wire n5644;
wire n5645;
wire n5646;
wire n5647;
wire n5648;
wire n5649;
wire n5650;
wire n5651;
wire n5652;
wire n5653;
wire n5654;
wire n5655;
wire n5656;
wire n5657;
wire n5658;
wire n5659;
wire n5660;
wire n5661;
wire n5662;
wire n5663;
wire n5664;
wire n5665;
wire n5666;
wire n5667;
wire n5668;
wire n5669;
wire n5670;
wire n5671;
wire n5672;
wire n5673;
wire n5674;
wire n5675;
wire n5676;
wire n5677;
wire n5678;
wire n5679;
wire n5680;
wire n5681;
wire n5682;
wire n5683;
wire n5684;
wire n5685;
wire n5686;
wire n5687;
wire n5688;
wire n5689;
wire n5690;
wire n5691;
wire n5692;
wire n5693;
wire n5694;
wire n5695;
wire n5696;
wire n5697;
wire n5698;
wire n5699;
wire n5700;
wire n5701;
wire n5702;
wire n5703;
wire n5704;
wire n5705;
wire n5706;
wire n5707;
wire n5708;
wire n5709;
wire n5710;
wire n5711;
wire n5712;
wire n5713;
wire n5714;
wire n5715;
wire n5716;
wire n5717;
wire n5718;
wire n5719;
wire n5720;
wire n5721;
wire n5722;
wire n5723;
wire n5724;
wire n5725;
wire n5726;
wire n5727;
wire n5728;
wire n5729;
wire n5730;
wire n5731;
wire n5732;
wire n5733;
wire n5734;
wire n5735;
wire n5736;
wire n5737;
wire n5738;
wire n5739;
wire n5740;
wire n5741;
wire n5742;
wire n5743;
wire n5744;
wire n5745;
wire n5746;
wire n5747;
wire n5748;
wire n5749;
wire n5750;
wire n5751;
wire n5752;
wire n5753;
wire n5754;
wire n5755;
wire n5756;
wire n5757;
wire n5758;
wire n5759;
wire n5760;
wire n5761;
wire n5762;
wire n5763;
wire n5764;
wire n5765;
wire n5766;
wire n5767;
wire n5768;
wire n5769;
wire n5770;
wire n5771;
wire n5772;
wire n5773;
wire n5774;
wire n5775;
wire n5776;
wire n5777;
wire n5778;
wire n5779;
wire n5780;
wire n5781;
wire n5782;
wire n5783;
wire n5784;
wire n5785;
wire n5786;
wire n5787;
wire n5788;
wire n5789;
wire n5790;
wire n5791;
wire n5792;
wire n5793;
wire n5794;
wire n5795;
wire n5796;
wire n5797;
wire n5798;
wire n5799;
wire n5800;
wire n5801;
wire n5802;
wire n5803;
wire n5804;
wire n5805;
wire n5806;
wire n5807;
wire n5808;
wire n5809;
wire n5810;
wire n5811;
wire n5812;
wire n5813;
wire n5814;
wire n5815;
wire n5816;
wire n5817;
wire n5818;
wire n5819;
wire n5820;
wire n5821;
wire n5822;
wire n5823;
wire n5824;
wire n5825;
wire n5826;
wire n5827;
wire n5828;
wire n5829;
wire n5830;
wire n5831;
wire n5832;
wire n5833;
wire n5834;
wire n5835;
wire n5836;
wire n5837;
wire n5838;
wire n5839;
wire n5840;
wire n5841;
wire n5842;
wire n5843;
wire n5844;
wire n5845;
wire n5846;
wire n5847;
wire n5848;
wire n5849;
wire n5850;
wire n5851;
wire n5852;
wire n5853;
wire n5854;
wire n5855;
wire n5856;
wire n5857;
wire n5858;
wire n5859;
wire n5860;
wire n5861;
wire n5862;
wire n5863;
wire n5864;
wire n5865;
wire n5866;
wire n5867;
wire n5868;
wire n5869;
wire n5870;
wire n5871;
wire n5872;
wire n5873;
wire n5874;
wire n5875;
wire n5876;
wire n5877;
wire n5878;
wire n5879;
wire n5880;
wire n5881;
wire n5882;
wire n5883;
wire n5884;
wire n5885;
wire n5886;
wire n5887;
wire n5888;
wire n5889;
wire n5890;
wire n5891;
wire n5892;
wire n5893;
wire n5894;
wire n5895;
wire n5896;
wire n5897;
wire n5898;
wire n5899;
wire n5900;
wire n5901;
wire n5902;
wire n5903;
wire n5904;
wire n5905;
wire n5906;
wire n5907;
wire n5908;
wire n5909;
wire n5910;
wire n5911;
wire n5912;
wire n5913;
wire n5914;
wire n5915;
wire n5916;
wire n5917;
wire n5918;
wire n5919;
wire n5920;
wire n5921;
wire n5922;
wire n5923;
wire n5924;
wire n5925;
wire n5926;
wire n5927;
wire n5928;
wire n5929;
wire n5930;
wire n5931;
wire n5932;
wire n5933;
wire n5934;
wire n5935;
wire n5936;
wire n5937;
wire n5938;
wire n5939;
wire n5940;
wire n5941;
wire n5942;
wire n5943;
wire n5944;
wire n5945;
wire n5946;
wire n5947;
wire n5948;
wire n5949;
wire n5950;
wire n5951;
wire n5952;
wire n5953;
wire n5954;
wire n5955;
wire n5956;
wire n5957;
wire n5958;
wire n5959;
wire n5960;
wire n5961;
wire n5962;
wire n5963;
wire n5964;
wire n5965;
wire n5966;
wire n5967;
wire n5968;
wire n5969;
wire n5970;
wire n5971;
wire n5972;
wire n5973;
wire n5974;
wire n5975;
wire n5976;
wire n5977;
wire n5978;
wire n5979;
wire n5980;
wire n5981;
wire n5982;
wire n5983;
wire n5984;
wire n5985;
wire n5986;
wire n5987;
wire n5988;
wire n5989;
wire n5990;
wire n5991;
wire n5992;
wire n5993;
wire n5994;
wire n5995;
wire n5996;
wire n5997;
wire n5998;
wire n5999;
wire n6000;
wire n6001;
wire n6002;
wire n6003;
wire n6004;
wire n6005;
wire n6006;
wire n6007;
wire n6008;
wire n6009;
wire n6010;
wire n6011;
wire n6012;
wire n6013;
wire n6014;
wire n6015;
wire n6016;
wire n6017;
wire n6018;
wire n6019;
wire n6020;
wire n6021;
wire n6022;
wire n6023;
wire n6024;
wire n6025;
wire n6026;
wire n6027;
wire n6028;
wire n6029;
wire n6030;
wire n6031;
wire n6032;
wire n6033;
wire n6034;
wire n6035;
wire n6036;
wire n6037;
wire n6038;
wire n6039;
wire n6040;
wire n6041;
wire n6042;
wire n6043;
wire n6044;
wire n6045;
wire n6046;
wire n6047;
wire n6048;
wire n6049;
wire n6050;
wire n6051;
wire n6052;
wire n6053;
wire n6054;
wire n6055;
wire n6056;
wire n6057;
wire n6058;
wire n6059;
wire n6060;
wire n6061;
wire n6062;
wire n6063;
wire n6064;
wire n6065;
wire n6066;
wire n6067;
wire n6068;
wire n6069;
wire n6070;
wire n6071;
wire n6072;
wire n6073;
wire n6074;
wire n6075;
wire n6076;
wire n6077;
wire n6078;
wire n6079;
wire n6080;
wire n6081;
wire n6082;
wire n6083;
wire n6084;
wire n6085;
wire n6086;
wire n6087;
wire n6088;
wire n6089;
wire n6090;
wire n6091;
wire n6092;
wire n6093;
wire n6094;
wire n6095;
wire n6096;
wire n6097;
wire n6098;
wire n6099;
wire n6100;
wire n6101;
wire n6102;
wire n6103;
wire n6104;
wire n6105;
wire n6106;
wire n6107;
wire n6108;
wire n6109;
wire n6110;
wire n6111;
wire n6112;
wire n6113;
wire n6114;
wire n6115;
wire n6116;
wire n6117;
wire n6118;
wire n6119;
wire n6120;
wire n6121;
wire n6122;
wire n6123;
wire n6124;
wire n6125;
wire n6126;
wire n6127;
wire n6128;
wire n6129;
wire n6130;
wire n6131;
wire n6132;
wire n6133;
wire n6134;
wire n6135;
wire n6136;
wire n6137;
wire n6138;
wire n6139;
wire n6140;
wire n6141;
wire n6142;
wire n6143;
wire n6144;
wire n6145;
wire n6146;
wire n6147;
wire n6148;
wire n6149;
wire n6150;
wire n6151;
wire n6152;
wire n6153;
wire n6154;
wire n6155;
wire n6156;
wire n6157;
wire n6158;
wire n6159;
wire n6160;
wire n6161;
wire n6162;
wire n6163;
wire n6164;
wire n6165;
wire n6166;
wire n6167;
wire n6168;
wire n6169;
wire n6170;
wire n6171;
wire n6172;
wire n6173;
wire n6174;
wire n6175;
wire n6176;
wire n6177;
wire n6178;
wire n6179;
wire n6180;
wire n6181;
wire n6182;
wire n6183;
wire n6184;
wire n6185;
wire n6186;
wire n6187;
wire n6188;
wire n6189;
wire n6190;
wire n6191;
wire n6192;
wire n6193;
wire n6194;
wire n6195;
wire n6196;
wire n6197;
wire n6198;
wire n6199;
wire n6200;
wire n6201;
wire n6202;
wire n6203;
wire n6204;
wire n6205;
wire n6206;
wire n6207;
wire n6208;
wire n6209;
wire n6210;
wire n6211;
wire n6212;
wire n6213;
wire n6214;
wire n6215;
wire n6216;
wire n6217;
wire n6218;
wire n6219;
wire n6220;
wire n6221;
wire n6222;
wire n6223;
wire n6224;
wire n6225;
wire n6226;
wire n6227;
wire n6228;
wire n6229;
wire n6230;
wire n6231;
wire n6232;
wire n6233;
wire n6234;
wire n6235;
wire n6236;
wire n6237;
wire n6238;
wire n6239;
wire n6240;
wire n6241;
wire n6242;
wire n6243;
wire n6244;
wire n6245;
wire n6246;
wire n6247;
wire n6248;
wire n6249;
wire n6250;
wire n6251;
wire n6252;
wire n6253;
wire n6254;
wire n6255;
wire n6256;
wire n6257;
wire n6258;
wire n6259;
wire n6260;
wire n6261;
wire n6262;
wire n6263;
wire n6264;
wire n6265;
wire n6266;
wire n6267;
wire n6268;
wire n6269;
wire n6270;
wire n6271;
wire n6272;
wire n6273;
wire n6274;
wire n6275;
wire n6276;
wire n6277;
wire n6278;
wire n6279;
wire n6280;
wire n6281;
wire n6282;
wire n6283;
wire n6284;
wire n6285;
wire n6286;
wire n6287;
wire n6288;
wire n6289;
wire n6290;
wire n6291;
wire n6292;
wire n6293;
wire n6294;
wire n6295;
wire n6296;
wire n6297;
wire n6298;
wire n6299;
wire n6300;
wire n6301;
wire n6302;
wire n6303;
wire n6304;
wire n6305;
wire n6306;
wire n6307;
wire n6308;
wire n6309;
wire n6310;
wire n6311;
wire n6312;
wire n6313;
wire n6314;
wire n6315;
wire n6316;
wire n6317;
wire n6318;
wire n6319;
wire n6320;
wire n6321;
wire n6322;
wire n6323;
wire n6324;
wire n6325;
wire n6326;
wire n6327;
wire n6328;
wire n6329;
wire n6330;
wire n6331;
wire n6332;
wire n6333;
wire n6334;
wire n6335;
wire n6336;
wire n6337;
wire n6338;
wire n6339;
wire n6340;
wire n6341;
wire n6342;
wire n6343;
wire n6344;
wire n6345;
wire n6346;
wire n6347;
wire n6348;
wire n6349;
wire n6350;
wire n6351;
wire n6352;
wire n6353;
wire n6354;
wire n6355;
wire n6356;
wire n6357;
wire n6358;
wire n6359;
wire n6360;
wire n6361;
wire n6362;
wire n6363;
wire n6364;
wire n6365;
wire n6366;
wire n6367;
wire n6368;
wire n6369;
wire n6370;
wire n6371;
wire n6372;
wire n6373;
wire n6374;
wire n6375;
wire n6376;
wire n6377;
wire n6378;
wire n6379;
wire n6380;
wire n6381;
wire n6382;
wire n6383;
wire n6384;
wire n6385;
wire n6386;
wire n6387;
wire n6388;
wire n6389;
wire n6390;
wire n6391;
wire n6392;
wire n6393;
wire n6394;
wire n6395;
wire n6396;
wire n6397;
wire n6398;
wire n6399;
wire n6400;
wire n6401;
wire n6402;
wire n6403;
wire n6404;
wire n6405;
wire n6406;
wire n6407;
wire n6408;
wire n6409;
wire n6410;
wire n6411;
wire n6412;
wire n6413;
wire n6414;
wire n6415;
wire n6416;
wire n6417;
wire n6418;
wire n6419;
wire n6420;
wire n6421;
wire n6422;
wire n6423;
wire n6424;
wire n6425;
wire n6426;
wire n6427;
wire n6428;
wire n6429;
wire n6430;
wire n6431;
wire n6432;
wire n6433;
wire n6434;
wire n6435;
wire n6436;
wire n6437;
wire n6438;
wire n6439;
wire n6440;
wire n6441;
wire n6442;
wire n6443;
wire n6444;
wire n6445;
wire n6446;
wire n6447;
wire n6448;
wire n6449;
wire n6450;
wire n6451;
wire n6452;
wire n6453;
wire n6454;
wire n6455;
wire n6456;
wire n6457;
wire n6458;
wire n6459;
wire n6460;
wire n6461;
wire n6462;
wire n6463;
wire n6464;
wire n6465;
wire n6466;
wire n6467;
wire n6468;
wire n6469;
wire n6470;
wire n6471;
wire n6472;
wire n6473;
wire n6474;
wire n6475;
wire n6476;
wire n6477;
wire n6478;
wire n6479;
wire n6480;
wire n6481;
wire n6482;
wire n6483;
wire n6484;
wire n6485;
wire n6486;
wire n6487;
wire n6488;
wire n6489;
wire n6490;
wire n6491;
wire n6492;
wire n6493;
wire n6494;
wire n6495;
wire n6496;
wire n6497;
wire n6498;
wire n6499;
wire n6500;
wire n6501;
wire n6502;
wire n6503;
wire n6504;
wire n6505;
wire n6506;
wire n6507;
wire n6508;
wire n6509;
wire n6510;
wire n6511;
wire n6512;
wire n6513;
wire n6514;
wire n6515;
wire n6516;
wire n6517;
wire n6518;
wire n6519;
wire n6520;
wire n6521;
wire n6522;
wire n6523;
wire n6524;
wire n6525;
wire n6526;
wire n6527;
wire n6528;
wire n6529;
wire n6530;
wire n6531;
wire n6532;
wire n6533;
wire n6534;
wire n6535;
wire n6536;
wire n6537;
wire n6538;
wire n6539;
wire n6540;
wire n6541;
wire n6542;
wire n6543;
wire n6544;
wire n6545;
wire n6546;
wire n6547;
wire n6548;
wire n6549;
wire n6550;
wire n6551;
wire n6552;
wire n6553;
wire n6554;
wire n6555;
wire n6556;
wire n6557;
wire n6558;
wire n6559;
wire n6560;
wire n6561;
wire n6562;
wire n6563;
wire n6564;
wire n6565;
wire n6566;
wire n6567;
wire n6568;
wire n6569;
wire n6570;
wire n6571;
wire n6572;
wire n6573;
wire n6574;
wire n6575;
wire n6576;
wire n6577;
wire n6578;
wire n6579;
wire n6580;
wire n6581;
wire n6582;
wire n6583;
wire n6584;
wire n6585;
wire n6586;
wire n6587;
wire n6588;
wire n6589;
wire n6590;
wire n6591;
wire n6592;
wire n6593;
wire n6594;
wire n6595;
wire n6596;
wire n6597;
wire n6598;
wire n6599;
wire n6600;
wire n6601;
wire n6602;
wire n6603;
wire n6604;
wire n6605;
wire n6606;
wire n6607;
wire n6608;
wire n6609;
wire n6610;
wire n6611;
wire n6612;
wire n6613;
wire n6614;
wire n6615;
wire n6616;
wire n6617;
wire n6618;
wire n6619;
wire n6620;
wire n6621;
wire n6622;
wire n6623;
wire n6624;
wire n6625;
wire n6626;
wire n6627;
wire n6628;
wire n6629;
wire n6630;
wire n6631;
wire n6632;
wire n6633;
wire n6634;
wire n6635;
wire n6636;
wire n6637;
wire n6638;
wire n6639;
wire n6640;
wire n6641;
wire n6642;
wire n6643;
wire n6644;
wire n6645;
wire n6646;
wire n6647;
wire n6648;
wire n6649;
wire n6650;
wire n6651;
wire n6652;
wire n6653;
wire n6654;
wire n6655;
wire n6656;
wire n6657;
wire n6658;
wire n6659;
wire n6660;
wire n6661;
wire n6662;
wire n6663;
wire n6664;
wire n6665;
wire n6666;
wire n6667;
wire n6668;
wire n6669;
wire n6670;
wire n6671;
wire n6672;
wire n6673;
wire n6674;
wire n6675;
wire n6676;
wire n6677;
wire n6678;
wire n6679;
wire n6680;
wire n6681;
wire n6682;
wire n6683;
wire n6684;
wire n6685;
wire n6686;
wire n6687;
wire n6688;
wire n6689;
wire n6690;
wire n6691;
wire n6692;
wire n6693;
wire n6694;
wire n6695;
wire n6696;
wire n6697;
wire n6698;
wire n6699;
wire n6700;
wire n6701;
wire n6702;
wire n6703;
wire n6704;
wire n6705;
wire n6706;
wire n6707;
wire n6708;
wire n6709;
wire n6710;
wire n6711;
wire n6712;
wire n6713;
wire n6714;
wire n6715;
wire n6716;
wire n6717;
wire n6718;
wire n6719;
wire n6720;
wire n6721;
wire n6722;
wire n6723;
wire n6724;
wire n6725;
wire n6726;
wire n6727;
wire n6728;
wire n6729;
wire n6730;
wire n6731;
wire n6732;
wire n6733;
wire n6734;
wire n6735;
wire n6736;
wire n6737;
wire n6738;
wire n6739;
wire n6740;
wire n6741;
wire n6742;
wire n6743;
wire n6744;
wire n6745;
wire n6746;
wire n6747;
wire n6748;
wire n6749;
wire n6750;
wire n6751;
wire n6752;
wire n6753;
wire n6754;
wire n6755;
wire n6756;
wire n6757;
wire n6758;
wire n6759;
wire n6760;
wire n6761;
wire n6762;
wire n6763;
wire n6764;
wire n6765;
wire n6766;
wire n6767;
wire n6768;
wire n6769;
wire n6770;
wire n6771;
wire n6772;
wire n6773;
wire n6774;
wire n6775;
wire n6776;
wire n6777;
wire n6778;
wire n6779;
wire n6780;
wire n6781;
wire n6782;
wire n6783;
wire n6784;
wire n6785;
wire n6786;
wire n6787;
wire n6788;
wire n6789;
wire n6790;
wire n6791;
wire n6792;
wire n6793;
wire n6794;
wire n6795;
wire n6796;
wire n6797;
wire n6798;
wire n6799;
wire n6800;
wire n6801;
wire n6802;
wire n6803;
wire n6804;
wire n6805;
wire n6806;
wire n6807;
wire n6808;
wire n6809;
wire n6810;
wire n6811;
wire n6812;
wire n6813;
wire n6814;
wire n6815;
wire n6816;
wire n6817;
wire n6818;
wire n6819;
wire n6820;
wire n6821;
wire n6822;
wire n6823;
wire n6824;
wire n6825;
wire n6826;
wire n6827;
wire n6828;
wire n6829;
wire n6830;
wire n6831;
wire n6832;
wire n6833;
wire n6834;
wire n6835;
wire n6836;
wire n6837;
wire n6838;
wire n6839;
wire n6840;
wire n6841;
wire n6842;
wire n6843;
wire n6844;
wire n6845;
wire n6846;
wire n6847;
wire n6848;
wire n6849;
wire n6850;
wire n6851;
wire n6852;
wire n6853;
wire n6854;
wire n6855;
wire n6856;
wire n6857;
wire n6858;
wire n6859;
wire n6860;
wire n6861;
wire n6862;
wire n6863;
wire n6864;
wire n6865;
wire n6866;
wire n6867;
wire n6868;
wire n6869;
wire n6870;
wire n6871;
wire n6872;
wire n6873;
wire n6874;
wire n6875;
wire n6876;
wire n6877;
wire n6878;
wire n6879;
wire n6880;
wire n6881;
wire n6882;
wire n6883;
wire n6884;
wire n6885;
wire n6886;
wire n6887;
wire n6888;
wire n6889;
wire n6890;
wire n6891;
wire n6892;
wire n6893;
wire n6894;
wire n6895;
wire n6896;
wire n6897;
wire n6898;
wire n6899;
wire n6900;
wire n6901;
wire n6902;
wire n6903;
wire n6904;
wire n6905;
wire n6906;
wire n6907;
wire n6908;
wire n6909;
wire n6910;
wire n6911;
wire n6912;
wire n6913;
wire n6914;
wire n6915;
wire n6916;
wire n6917;
wire n6918;
wire n6919;
wire n6920;
wire n6921;
wire n6922;
wire n6923;
wire n6924;
wire n6925;
wire n6926;
wire n6927;
wire n6928;
wire n6929;
wire n6930;
wire n6931;
wire n6932;
wire n6933;
wire n6934;
wire n6935;
wire n6936;
wire n6937;
wire n6938;
wire n6939;
wire n6940;
wire n6941;
wire n6942;
wire n6943;
wire n6944;
wire n6945;
wire n6946;
wire n6947;
wire n6948;
wire n6949;
wire n6950;
wire n6951;
wire n6952;
wire n6953;
wire n6954;
wire n6955;
wire n6956;
wire n6957;
wire n6958;
wire n6959;
wire n6960;
wire n6961;
wire n6962;
wire n6963;
wire n6964;
wire n6965;
wire n6966;
wire n6967;
wire n6968;
wire n6969;
wire n6970;
wire n6971;
wire n6972;
wire n6973;
wire n6974;
wire n6975;
wire n6976;
wire n6977;
wire n6978;
wire n6979;
wire n6980;
wire n6981;
wire n6982;
wire n6983;
wire n6984;
wire n6985;
wire n6986;
wire n6987;
wire n6988;
wire n6989;
wire n6990;
wire n6991;
wire n6992;
wire n6993;
wire n6994;
wire n6995;
wire n6996;
wire n6997;
wire n6998;
wire n6999;
wire n7000;
wire n7001;
wire n7002;
wire n7003;
wire n7004;
wire n7005;
wire n7006;
wire n7007;
wire n7008;
wire n7009;
wire n7010;
wire n7011;
wire n7012;
wire n7013;
wire n7014;
wire n7015;
wire n7016;
wire n7017;
wire n7018;
wire n7019;
wire n7020;
wire n7021;
wire n7022;
wire n7023;
wire n7024;
wire n7025;
wire n7026;
wire n7027;
wire n7028;
wire n7029;
wire n7030;
wire n7031;
wire n7032;
wire n7033;
wire n7034;
wire n7035;
wire n7036;
wire n7037;
wire n7038;
wire n7039;
wire n7040;
wire n7041;
wire n7042;
wire n7043;
wire n7044;
wire n7045;
wire n7046;
wire n7047;
wire n7048;
wire n7049;
wire n7050;
wire n7051;
wire n7052;
wire n7053;
wire n7054;
wire n7055;
wire n7056;
wire n7057;
wire n7058;
wire n7059;
wire n7060;
wire n7061;
wire n7062;
wire n7063;
wire n7064;
wire n7065;
wire n7066;
wire n7067;
wire n7068;
wire n7069;
wire n7070;
wire n7071;
wire n7072;
wire n7073;
wire n7074;
wire n7075;
wire n7076;
wire n7077;
wire n7078;
wire n7079;
wire n7080;
wire n7081;
wire n7082;
wire n7083;
wire n7084;
wire n7085;
wire n7086;
wire n7087;
wire n7088;
wire n7089;
wire n7090;
wire n7091;
wire n7092;
wire n7093;
wire n7094;
wire n7095;
wire n7096;
wire n7097;
wire n7098;
wire n7099;
wire n7100;
wire n7101;
wire n7102;
wire n7103;
wire n7104;
wire n7105;
wire n7106;
wire n7107;
wire n7108;
wire n7109;
wire n7110;
wire n7111;
wire n7112;
wire n7113;
wire n7114;
wire n7115;
wire n7116;
wire n7117;
wire n7118;
wire n7119;
wire n7120;
wire n7121;
wire n7122;
wire n7123;
wire n7124;
wire n7125;
wire n7126;
wire n7127;
wire n7128;
wire n7129;
wire n7130;
wire n7131;
wire n7132;
wire n7133;
wire n7134;
wire n7135;
wire n7136;
wire n7137;
wire n7138;
wire n7139;
wire n7140;
wire n7141;
wire n7142;
wire n7143;
wire n7144;
wire n7145;
wire n7146;
wire n7147;
wire n7148;
wire n7149;
wire n7150;
wire n7151;
wire n7152;
wire n7153;
wire n7154;
wire n7155;
wire n7156;
wire n7157;
wire n7158;
wire n7159;
wire n7160;
wire n7161;
wire n7162;
wire n7163;
wire n7164;
wire n7165;
wire n7166;
wire n7167;
wire n7168;
wire n7169;
wire n7170;
wire n7171;
wire n7172;
wire n7173;
wire n7174;
wire n7175;
wire n7176;
wire n7177;
wire n7178;
wire n7179;
wire n7180;
wire n7181;
wire n7182;
wire n7183;
wire n7184;
wire n7185;
wire n7186;
wire n7187;
wire n7188;
wire n7189;
wire n7190;
wire n7191;
wire n7192;
wire n7193;
wire n7194;
wire n7195;
wire n7196;
wire n7197;
wire n7198;
wire n7199;
wire n7200;
wire n7201;
wire n7202;
wire n7203;
wire n7204;
wire n7205;
wire n7206;
wire n7207;
wire n7208;
wire n7209;
wire n7210;
wire n7211;
wire n7212;
wire n7213;
wire n7214;
wire n7215;
wire n7216;
wire n7217;
wire n7218;
wire n7219;
wire n7220;
wire n7221;
wire n7222;
wire n7223;
wire n7224;
wire n7225;
wire n7226;
wire n7227;
wire n7228;
wire n7229;
wire n7230;
wire n7231;
wire n7232;
wire n7233;
wire n7234;
wire n7235;
wire n7236;
wire n7237;
wire n7238;
wire n7239;
wire n7240;
wire n7241;
wire n7242;
wire n7243;
wire n7244;
wire n7245;
wire n7246;
wire n7247;
wire n7248;
wire n7249;
wire n7250;
wire n7251;
wire n7252;
wire n7253;
wire n7254;
wire n7255;
wire n7256;
wire n7257;
wire n7258;
wire n7259;
wire n7260;
wire n7261;
wire n7262;
wire n7263;
wire n7264;
wire n7265;
wire n7266;
wire n7267;
wire n7268;
wire n7269;
wire n7270;
wire n7271;
wire n7272;
wire n7273;
wire n7274;
wire n7275;
wire n7276;
wire n7277;
wire n7278;
wire n7279;
wire n7280;
wire n7281;
wire n7282;
wire n7283;
wire n7284;
wire n7285;
wire n7286;
wire n7287;
wire n7288;
wire n7289;
wire n7290;
wire n7291;
wire n7292;
wire n7293;
wire n7294;
wire n7295;
wire n7296;
wire n7297;
wire n7298;
wire n7299;
wire n7300;
wire n7301;
wire n7302;
wire n7303;
wire n7304;
wire n7305;
wire n7306;
wire n7307;
wire n7308;
wire n7309;
wire n7310;
wire n7311;
wire n7312;
wire n7313;
wire n7314;
wire n7315;
wire n7316;
wire n7317;
wire n7318;
wire n7319;
wire n7320;
wire n7321;
wire n7322;
wire n7323;
wire n7324;
wire n7325;
wire n7326;
wire n7327;
wire n7328;
wire n7329;
wire n7330;
wire n7331;
wire n7332;
wire n7333;
wire n7334;
wire n7335;
wire n7336;
wire n7337;
wire n7338;
wire n7339;
wire n7340;
wire n7341;
wire n7342;
wire n7343;
wire n7344;
wire n7345;
wire n7346;
wire n7347;
wire n7348;
wire n7349;
wire n7350;
wire n7351;
wire n7352;
wire n7353;
wire n7354;
wire n7355;
wire n7356;
wire n7357;
wire n7358;
wire n7359;
wire n7360;
wire n7361;
wire n7362;
wire n7363;
wire n7364;
wire n7365;
wire n7366;
wire n7367;
wire n7368;
wire n7369;
wire n7370;
wire n7371;
wire n7372;
wire n7373;
wire n7374;
wire n7375;
wire n7376;
wire n7377;
wire n7378;
wire n7379;
wire n7380;
wire n7381;
wire n7382;
wire n7383;
wire n7384;
wire n7385;
wire n7386;
wire n7387;
wire n7388;
wire n7389;
wire n7390;
wire n7391;
wire n7392;
wire n7393;
wire n7394;
wire n7395;
wire n7396;
wire n7397;
wire n7398;
wire n7399;
wire n7400;
wire n7401;
wire n7402;
wire n7403;
wire n7404;
wire n7405;
wire n7406;
wire n7407;
wire n7408;
wire n7409;
wire n7410;
wire n7411;
wire n7412;
wire n7413;
wire n7414;
wire n7415;
wire n7416;
wire n7417;
wire n7418;
wire n7419;
wire n7420;
wire n7421;
wire n7422;
wire n7423;
wire n7424;
wire n7425;
wire n7426;
wire n7427;
wire n7428;
wire n7429;
wire n7430;
wire n7431;
wire n7432;
wire n7433;
wire n7434;
wire n7435;
wire n7436;
wire n7437;
wire n7438;
wire n7439;
wire n7440;
wire n7441;
wire n7442;
wire n7443;
wire n7444;
wire n7445;
wire n7446;
wire n7447;
wire n7448;
wire n7449;
wire n7450;
wire n7451;
wire n7452;
wire n7453;
wire n7454;
wire n7455;
wire n7456;
wire n7457;
wire n7458;
wire n7459;
wire n7460;
wire n7461;
wire n7462;
wire n7463;
wire n7464;
wire n7465;
wire n7466;
wire n7467;
wire n7468;
wire n7469;
wire n7470;
wire n7471;
wire n7472;
wire n7473;
wire n7474;
wire n7475;
wire n7476;
wire n7477;
wire n7478;
wire n7479;
wire n7480;
wire n7481;
wire n7482;
wire n7483;
wire n7484;
wire n7485;
wire n7486;
wire n7487;
wire n7488;
wire n7489;
wire n7490;
wire n7491;
wire n7492;
wire n7493;
wire n7494;
wire n7495;
wire n7496;
wire n7497;
wire n7498;
wire n7499;
wire n7500;
wire n7501;
wire n7502;
wire n7503;
wire n7504;
wire n7505;
wire n7506;
wire n7507;
wire n7508;
wire n7509;
wire n7510;
wire n7511;
wire n7512;
wire n7513;
wire n7514;
wire n7515;
wire n7516;
wire n7517;
wire n7518;
wire n7519;
wire n7520;
wire n7521;
wire n7522;
wire n7523;
wire n7524;
wire n7525;
wire n7526;
wire n7527;
wire n7528;
wire n7529;
wire n7530;
wire n7531;
wire n7532;
wire n7533;
wire n7534;
wire n7535;
wire n7536;
wire n7537;
wire n7538;
wire n7539;
wire n7540;
wire n7541;
wire n7542;
wire n7543;
wire n7544;
wire n7545;
wire n7546;
wire n7547;
wire n7548;
wire n7549;
wire n7550;
wire n7551;
wire n7552;
wire n7553;
wire n7554;
wire n7555;
wire n7556;
wire n7557;
wire n7558;
wire n7559;
wire n7560;
wire n7561;
wire n7562;
wire n7563;
wire n7564;
wire n7565;
wire n7566;
wire n7567;
wire n7568;
wire n7569;
wire n7570;
wire n7571;
wire n7572;
wire n7573;
wire n7574;
wire n7575;
wire n7576;
wire n7577;
wire n7578;
wire n7579;
wire n7580;
wire n7581;
wire n7582;
wire n7583;
wire n7584;
wire n7585;
wire n7586;
wire n7587;
wire n7588;
wire n7589;
wire n7590;
wire n7591;
wire n7592;
wire n7593;
wire n7594;
wire n7595;
wire n7596;
wire n7597;
wire n7598;
wire n7599;
wire n7600;
wire n7601;
wire n7602;
wire n7603;
wire n7604;
wire n7605;
wire n7606;
wire n7607;
wire n7608;
wire n7609;
wire n7610;
wire n7611;
wire n7612;
wire n7613;
wire n7614;
wire n7615;
wire n7616;
wire n7617;
wire n7618;
wire n7619;
wire n7620;
wire n7621;
wire n7622;
wire n7623;
wire n7624;
wire n7625;
wire n7626;
wire n7627;
wire n7628;
wire n7629;
wire n7630;
wire n7631;
wire n7632;
wire n7633;
wire n7634;
wire n7635;
wire n7636;
wire n7637;
wire n7638;
wire n7639;
wire n7640;
wire n7641;
wire n7642;
wire n7643;
wire n7644;
wire n7645;
wire n7646;
wire n7647;
wire n7648;
wire n7649;
wire n7650;
wire n7651;
wire n7652;
wire n7653;
wire n7654;
wire n7655;
wire n7656;
wire n7657;
wire n7658;
wire n7659;
wire n7660;
wire n7661;
wire n7662;
wire n7663;
wire n7664;
wire n7665;
wire n7666;
wire n7667;
wire n7668;
wire n7669;
wire n7670;
wire n7671;
wire n7672;
wire n7673;
wire n7674;
wire n7675;
wire n7676;
wire n7677;
wire n7678;
wire n7679;
wire n7680;
wire n7681;
wire n7682;
wire n7683;
wire n7684;
wire n7685;
wire n7686;
wire n7687;
wire n7688;
wire n7689;
wire n7690;
wire n7691;
wire n7692;
wire n7693;
wire n7694;
wire n7695;
wire n7696;
wire n7697;
wire n7698;
wire n7699;
wire n7700;
wire n7701;
wire n7702;
wire n7703;
wire n7704;
wire n7705;
wire n7706;
wire n7707;
wire n7708;
wire n7709;
wire n7710;
wire n7711;
wire n7712;
wire n7713;
wire n7714;
wire n7715;
wire n7716;
wire n7717;
wire n7718;
wire n7719;
wire n7720;
wire n7721;
wire n7722;
wire n7723;
wire n7724;
wire n7725;
wire n7726;
wire n7727;
wire n7728;
wire n7729;
wire n7730;
wire n7731;
wire n7732;
wire n7733;
wire n7734;
wire n7735;
wire n7736;
wire n7737;
wire n7738;
wire n7739;
wire n7740;
wire n7741;
wire n7742;
wire n7743;
wire n7744;
wire n7745;
wire n7746;
wire n7747;
wire n7748;
wire n7749;
wire n7750;
wire n7751;
wire n7752;
wire n7753;
wire n7754;
wire n7755;
wire n7756;
wire n7757;
wire n7758;
wire n7759;
wire n7760;
wire n7761;
wire n7762;
wire n7763;
wire n7764;
wire n7765;
wire n7766;
wire n7767;
wire n7768;
wire n7769;
wire n7770;
wire n7771;
wire n7772;
wire n7773;
wire n7774;
wire n7775;
wire n7776;
wire n7777;
wire n7778;
wire n7779;
wire n7780;
wire n7781;
wire n7782;
wire n7783;
wire n7784;
wire n7785;
wire n7786;
wire n7787;
wire n7788;
wire n7789;
wire n7790;
wire n7791;
wire n7792;
wire n7793;
wire n7794;
wire n7795;
wire n7796;
wire n7797;
wire n7798;
wire n7799;
wire n7800;
wire n7801;
wire n7802;
wire n7803;
wire n7804;
wire n7805;
wire n7806;
wire n7807;
wire n7808;
wire n7809;
wire n7810;
wire n7811;
wire n7812;
wire n7813;
wire n7814;
wire n7815;
wire n7816;
wire n7817;
wire n7818;
wire n7819;
wire n7820;
wire n7821;
wire n7822;
wire n7823;
wire n7824;
wire n7825;
wire n7826;
wire n7827;
wire n7828;
wire n7829;
wire n7830;
wire n7831;
wire n7832;
wire n7833;
wire n7834;
wire n7835;
wire n7836;
wire n7837;
wire n7838;
wire n7839;
wire n7840;
wire n7841;
wire n7842;
wire n7843;
wire n7844;
wire n7845;
wire n7846;
wire n7847;
wire n7848;
wire n7849;
wire n7850;
wire n7851;
wire n7852;
wire n7853;
wire n7854;
wire n7855;
wire n7856;
wire n7857;
wire n7858;
wire n7859;
wire n7860;
wire n7861;
wire n7862;
wire n7863;
wire n7864;
wire n7865;
wire n7866;
wire n7867;
wire n7868;
wire n7869;
wire n7870;
wire n7871;
wire n7872;
wire n7873;
wire n7874;
wire n7875;
wire n7876;
wire n7877;
wire n7878;
wire n7879;
wire n7880;
wire n7881;
wire n7882;
wire n7883;
wire n7884;
wire n7885;
wire n7886;
wire n7887;
wire n7888;
wire n7889;
wire n7890;
wire n7891;
wire n7892;
wire n7893;
wire n7894;
wire n7895;
wire n7896;
wire n7897;
wire n7898;
wire n7899;
wire n7900;
wire n7901;
wire n7902;
wire n7903;
wire n7904;
wire n7905;
wire n7906;
wire n7907;
wire n7908;
wire n7909;
wire n7910;
wire n7911;
wire n7912;
wire n7913;
wire n7914;
wire n7915;
wire n7916;
wire n7917;
wire n7918;
wire n7919;
wire n7920;
wire n7921;
wire n7922;
wire n7923;
wire n7924;
wire n7925;
wire n7926;
wire n7927;
wire n7928;
wire n7929;
wire n7930;
wire n7931;
wire n7932;
wire n7933;
wire n7934;
wire n7935;
wire n7936;
wire n7937;
wire n7938;
wire n7939;
wire n7940;
wire n7941;
wire n7942;
wire n7943;
wire n7944;
wire n7945;
wire n7946;
wire n7947;
wire n7948;
wire n7949;
wire n7950;
wire n7951;
wire n7952;
wire n7953;
wire n7954;
wire n7955;
wire n7956;
wire n7957;
wire n7958;
wire n7959;
wire n7960;
wire n7961;
wire n7962;
wire n7963;
wire n7964;
wire n7965;
wire n7966;
wire n7967;
wire n7968;
wire n7969;
wire n7970;
wire n7971;
wire n7972;
wire n7973;
wire n7974;
wire n7975;
wire n7976;
wire n7977;
wire n7978;
wire n7979;
wire n7980;
wire n7981;
wire n7982;
wire n7983;
wire n7984;
wire n7985;
wire n7986;
wire n7987;
wire n7988;
wire n7989;
wire n7990;
wire n7991;
wire n7992;
wire n7993;
wire n7994;
wire n7995;
wire n7996;
wire n7997;
wire n7998;
wire n7999;
wire n8000;
wire n8001;
wire n8002;
wire n8003;
wire n8004;
wire n8005;
wire n8006;
wire n8007;
wire n8008;
wire n8009;
wire n8010;
wire n8011;
wire n8012;
wire n8013;
wire n8014;
wire n8015;
wire n8016;
wire n8017;
wire n8018;
wire n8019;
wire n8020;
wire n8021;
wire n8022;
wire n8023;
wire n8024;
wire n8025;
wire n8026;
wire n8027;
wire n8028;
wire n8029;
wire n8030;
wire n8031;
wire n8032;
wire n8033;
wire n8034;
wire n8035;
wire n8036;
wire n8037;
wire n8038;
wire n8039;
wire n8040;
wire n8041;
wire n8042;
wire n8043;
wire n8044;
wire n8045;
wire n8046;
wire n8047;
wire n8048;
wire n8049;
wire n8050;
wire n8051;
wire n8052;
wire n8053;
wire n8054;
wire n8055;
wire n8056;
wire n8057;
wire n8058;
wire n8059;
wire n8060;
wire n8061;
wire n8062;
wire n8063;
wire n8064;
wire n8065;
wire n8066;
wire n8067;
wire n8068;
wire n8069;
wire n8070;
wire n8071;
wire n8072;
wire n8073;
wire n8074;
wire n8075;
wire n8076;
wire n8077;
wire n8078;
wire n8079;
wire n8080;
wire n8081;
wire n8082;
wire n8083;
wire n8084;
wire n8085;
wire n8086;
wire n8087;
wire n8088;
wire n8089;
wire n8090;
wire n8091;
wire n8092;
wire n8093;
wire n8094;
wire n8095;
wire n8096;
wire n8097;
wire n8098;
wire n8099;
wire n8100;
wire n8101;
wire n8102;
wire n8103;
wire n8104;
wire n8105;
wire n8106;
wire n8107;
wire n8108;
wire n8109;
wire n8110;
wire n8111;
wire n8112;
wire n8113;
wire n8114;
wire n8115;
wire n8116;
wire n8117;
wire n8118;
wire n8119;
wire n8120;
wire n8121;
wire n8122;
wire n8123;
wire n8124;
wire n8125;
wire n8126;
wire n8127;
wire n8128;
wire n8129;
wire n8130;
wire n8131;
wire n8132;
wire n8133;
wire n8134;
wire n8135;
wire n8136;
wire n8137;
wire n8138;
wire n8139;
wire n8140;
wire n8141;
wire n8142;
wire n8143;
wire n8144;
wire n8145;
wire n8146;
wire n8147;
wire n8148;
wire n8149;
wire n8150;
wire n8151;
wire n8152;
wire n8153;
wire n8154;
wire n8155;
wire n8156;
wire n8157;
wire n8158;
wire n8159;
wire n8160;
wire n8161;
wire n8162;
wire n8163;
wire n8164;
wire n8165;
wire n8166;
wire n8167;
wire n8168;
wire n8169;
wire n8170;
wire n8171;
wire n8172;
wire n8173;
wire n8174;
wire n8175;
wire n8176;
wire n8177;
wire n8178;
wire n8179;
wire n8180;
wire n8181;
wire n8182;
wire n8183;
wire n8184;
wire n8185;
wire n8186;
wire n8187;
wire n8188;
wire n8189;
wire n8190;
wire n8191;
wire n8192;
wire n8193;
wire n8194;
wire n8195;
wire n8196;
wire n8197;
wire n8198;
wire n8199;
wire n8200;
wire n8201;
wire n8202;
wire n8203;
wire n8204;
wire n8205;
wire n8206;
wire n8207;
wire n8208;
wire n8209;
wire n8210;
wire n8211;
wire n8212;
wire n8213;
wire n8214;
wire n8215;
wire n8216;
wire n8217;
wire n8218;
wire n8219;
wire n8220;
wire n8221;
wire n8222;
wire n8223;
wire n8224;
wire n8225;
wire n8226;
wire n8227;
wire n8228;
wire n8229;
wire n8230;
wire n8231;
wire n8232;
wire n8233;
wire n8234;
wire n8235;
wire n8236;
wire n8237;
wire n8238;
wire n8239;
wire n8240;
wire n8241;
wire n8242;
wire n8243;
wire n8244;
wire n8245;
wire n8246;
wire n8247;
wire n8248;
wire n8249;
wire n8250;
wire n8251;
wire n8252;
wire n8253;
wire n8254;
wire n8255;
wire n8256;
wire n8257;
wire n8258;
wire n8259;
wire n8260;
wire n8261;
wire n8262;
wire n8263;
wire n8264;
wire n8265;
wire n8266;
wire n8267;
wire n8268;
wire n8269;
wire n8270;
wire n8271;
wire n8272;
wire n8273;
wire n8274;
wire n8275;
wire n8276;
wire n8277;
wire n8278;
wire n8279;
wire n8280;
wire n8281;
wire n8282;
wire n8283;
wire n8284;
wire n8285;
wire n8286;
wire n8287;
wire n8288;
wire n8289;
wire n8290;
wire n8291;
wire n8292;
wire n8293;
wire n8294;
wire n8295;
wire n8296;
wire n8297;
wire n8298;
wire n8299;
wire n8300;
wire n8301;
wire n8302;
wire n8303;
wire n8304;
wire n8305;
wire n8306;
wire n8307;
wire n8308;
wire n8309;
wire n8310;
wire n8311;
wire n8312;
wire n8313;
wire n8314;
wire n8315;
wire n8316;
wire n8317;
wire n8318;
wire n8319;
wire n8320;
wire n8321;
wire n8322;
wire n8323;
wire n8324;
wire n8325;
wire n8326;
wire n8327;
wire n8328;
wire n8329;
wire n8330;
wire n8331;
wire n8332;
wire n8333;
wire n8334;
wire n8335;
wire n8336;
wire n8337;
wire n8338;
wire n8339;
wire n8340;
wire n8341;
wire n8342;
wire n8343;
wire n8344;
wire n8345;
wire n8346;
wire n8347;
wire n8348;
wire n8349;
wire n8350;
wire n8351;
wire n8352;
wire n8353;
wire n8354;
wire n8355;
wire n8356;
wire n8357;
wire n8358;
wire n8359;
wire n8360;
wire n8361;
wire n8362;
wire n8363;
wire n8364;
wire n8365;
wire n8366;
wire n8367;
wire n8368;
wire n8369;
wire n8370;
wire n8371;
wire n8372;
wire n8373;
wire n8374;
wire n8375;
wire n8376;
wire n8377;
wire n8378;
wire n8379;
wire n8380;
wire n8381;
wire n8382;
wire n8383;
wire n8384;
wire n8385;
wire n8386;
wire n8387;
wire n8388;
wire n8389;
wire n8390;
wire n8391;
wire n8392;
wire n8393;
wire n8394;
wire n8395;
wire n8396;
wire n8397;
wire n8398;
wire n8399;
wire n8400;
wire n8401;
wire n8402;
wire n8403;
wire n8404;
wire n8405;
wire n8406;
wire n8407;
wire n8408;
wire n8409;
wire n8410;
wire n8411;
wire n8412;
wire n8413;
wire n8414;
wire n8415;
wire n8416;
wire n8417;
wire n8418;
wire n8419;
wire n8420;
wire n8421;
wire n8422;
wire n8423;
wire n8424;
wire n8425;
wire n8426;
wire n8427;
wire n8428;
wire n8429;
wire n8430;
wire n8431;
wire n8432;
wire n8433;
wire n8434;
wire n8435;
wire n8436;
wire n8437;
wire n8438;
wire n8439;
wire n8440;
wire n8441;
wire n8442;
wire n8443;
wire n8444;
wire n8445;
wire n8446;
wire n8447;
wire n8448;
wire n8449;
wire n8450;
wire n8451;
wire n8452;
wire n8453;
wire n8454;
wire n8455;
wire n8456;
wire n8457;
wire n8458;
wire n8459;
wire n8460;
wire n8461;
wire n8462;
wire n8463;
wire n8464;
wire n8465;
wire n8466;
wire n8467;
wire n8468;
wire n8469;
wire n8470;
wire n8471;
wire n8472;
wire n8473;
wire n8474;
wire n8475;
wire n8476;
wire n8477;
wire n8478;
wire n8479;
wire n8480;
wire n8481;
wire n8482;
wire n8483;
wire n8484;
wire n8485;
wire n8486;
wire n8487;
wire n8488;
wire n8489;
wire n8490;
wire n8491;
wire n8492;
wire n8493;
wire n8494;
wire n8495;
wire n8496;
wire n8497;
wire n8498;
wire n8499;
wire n8500;
wire n8501;
wire n8502;
wire n8503;
wire n8504;
wire n8505;
wire n8506;
wire n8507;
wire n8508;
wire n8509;
wire n8510;
wire n8511;
wire n8512;
wire n8513;
wire n8514;
wire n8515;
wire n8516;
wire n8517;
wire n8518;
wire n8519;
wire n8520;
wire n8521;
wire n8522;
wire n8523;
wire n8524;
wire n8525;
wire n8526;
wire n8527;
wire n8528;
wire n8529;
wire n8530;
wire n8531;
wire n8532;
wire n8533;
wire n8534;
wire n8535;
wire n8536;
wire n8537;
wire n8538;
wire n8539;
wire n8540;
wire n8541;
wire n8542;
wire n8543;
wire n8544;
wire n8545;
wire n8546;
wire n8547;
wire n8548;
wire n8549;
wire n8550;
wire n8551;
wire n8552;
wire n8553;
wire n8554;
wire n8555;
wire n8556;
wire n8557;
wire n8558;
wire n8559;
wire n8560;
wire n8561;
wire n8562;
wire n8563;
wire n8564;
wire n8565;
wire n8566;
wire n8567;
wire n8568;
wire n8569;
wire n8570;
wire n8571;
wire n8572;
wire n8573;
wire n8574;
wire n8575;
wire n8576;
wire n8577;
wire n8578;
wire n8579;
wire n8580;
wire n8581;
wire n8582;
wire n8583;
wire n8584;
wire n8585;
wire n8586;
wire n8587;
wire n8588;
wire n8589;
wire n8590;
wire n8591;
wire n8592;
wire n8593;
wire n8594;
wire n8595;
wire n8596;
wire n8597;
wire n8598;
wire n8599;
wire n8600;
wire n8601;
wire n8602;
wire n8603;
wire n8604;
wire n8605;
wire n8606;
wire n8607;
wire n8608;
wire n8609;
wire n8610;
wire n8611;
wire n8612;
wire n8613;
wire n8614;
wire n8615;
wire n8616;
wire n8617;
wire n8618;
wire n8619;
wire n8620;
wire n8621;
wire n8622;
wire n8623;
wire n8624;
wire n8625;
wire n8626;
wire n8627;
wire n8628;
wire n8629;
wire n8630;
wire n8631;
wire n8632;
wire n8633;
wire n8634;
wire n8635;
wire n8636;
wire n8637;
wire n8638;
wire n8639;
wire n8640;
wire n8641;
wire n8642;
wire n8643;
wire n8644;
wire n8645;
wire n8646;
wire n8647;
wire n8648;
wire n8649;
wire n8650;
wire n8651;
wire n8652;
wire n8653;
wire n8654;
wire n8655;
wire n8656;
wire n8657;
wire n8658;
wire n8659;
wire n8660;
wire n8661;
wire n8662;
wire n8663;
wire n8664;
wire n8665;
wire n8666;
wire n8667;
wire n8668;
wire n8669;
wire n8670;
wire n8671;
wire n8672;
wire n8673;
wire n8674;
wire n8675;
wire n8676;
wire n8677;
wire n8678;
wire n8679;
wire n8680;
wire n8681;
wire n8682;
wire n8683;
wire n8684;
wire n8685;
wire n8686;
wire n8687;
wire n8688;
wire n8689;
wire n8690;
wire n8691;
wire n8692;
wire n8693;
wire n8694;
wire n8695;
wire n8696;
wire n8697;
wire n8698;
wire n8699;
wire n8700;
wire n8701;
wire n8702;
wire n8703;
wire n8704;
wire n8705;
wire n8706;
wire n8707;
wire n8708;
wire n8709;
wire n8710;
wire n8711;
wire n8712;
wire n8713;
wire n8714;
wire n8715;
wire n8716;
wire n8717;
wire n8718;
wire n8719;
wire n8720;
wire n8721;
wire n8722;
wire n8723;
wire n8724;
wire n8725;
wire n8726;
wire n8727;
wire n8728;
wire n8729;
wire n8730;
wire n8731;
wire n8732;
wire n8733;
wire n8734;
wire n8735;
wire n8736;
wire n8737;
wire n8738;
wire n8739;
wire n8740;
wire n8741;
wire n8742;
wire n8743;
wire n8744;
wire n8745;
wire n8746;
wire n8747;
wire n8748;
wire n8749;
wire n8750;
wire n8751;
wire n8752;
wire n8753;
wire n8754;
wire n8755;
wire n8756;
wire n8757;
wire n8758;
wire n8759;
wire n8760;
wire n8761;
wire n8762;
wire n8763;
wire n8764;
wire n8765;
wire n8766;
wire n8767;
wire n8768;
wire n8769;
wire n8770;
wire n8771;
wire n8772;
wire n8773;
wire n8774;
wire n8775;
wire n8776;
wire n8777;
wire n8778;
wire n8779;
wire n8780;
wire n8781;
wire n8782;
wire n8783;
wire n8784;
wire n8785;
wire n8786;
wire n8787;
wire n8788;
wire n8789;
wire n8790;
wire n8791;
wire n8792;
wire n8793;
wire n8794;
wire n8795;
wire n8796;
wire n8797;
wire n8798;
wire n8799;
wire n8800;
wire n8801;
wire n8802;
wire n8803;
wire n8804;
wire n8805;
wire n8806;
wire n8807;
wire n8808;
wire n8809;
wire n8810;
wire n8811;
wire n8812;
wire n8813;
wire n8814;
wire n8815;
wire n8816;
wire n8817;
wire n8818;
wire n8819;
wire n8820;
wire n8821;
wire n8822;
wire n8823;
wire n8824;
wire n8825;
wire n8826;
wire n8827;
wire n8828;
wire n8829;
wire n8830;
wire n8831;
wire n8832;
wire n8833;
wire n8834;
wire n8835;
wire n8836;
wire n8837;
wire n8838;
wire n8839;
wire n8840;
wire n8841;
wire n8842;
wire n8843;
wire n8844;
wire n8845;
wire n8846;
wire n8847;
wire n8848;
wire n8849;
wire n8850;
wire n8851;
wire n8852;
wire n8853;
wire n8854;
wire n8855;
wire n8856;
wire n8857;
wire n8858;
wire n8859;
wire n8860;
wire n8861;
wire n8862;
wire n8863;
wire n8864;
wire n8865;
wire n8866;
wire n8867;
wire n8868;
wire n8869;
wire n8870;
wire n8871;
wire n8872;
wire n8873;
wire n8874;
wire n8875;
wire n8876;
wire n8877;
wire n8878;
wire n8879;
wire n8880;
wire n8881;
wire n8882;
wire n8883;
wire n8884;
wire n8885;
wire n8886;
wire n8887;
wire n8888;
wire n8889;
wire n8890;
wire n8891;
wire n8892;
wire n8893;
wire n8894;
wire n8895;
wire n8896;
wire n8897;
wire n8898;
wire n8899;
wire n8900;
wire n8901;
wire n8902;
wire n8903;
wire n8904;
wire n8905;
wire n8906;
wire n8907;
wire n8908;
wire n8909;
wire n8910;
wire n8911;
wire n8912;
wire n8913;
wire n8914;
wire n8915;
wire n8916;
wire n8917;
wire n8918;
wire n8919;
wire n8920;
wire n8921;
wire n8922;
wire n8923;
wire n8924;
wire n8925;
wire n8926;
wire n8927;
wire n8928;
wire n8929;
wire n8930;
wire n8931;
wire n8932;
wire n8933;
wire n8934;
wire n8935;
wire n8936;
wire n8937;
wire n8938;
wire n8939;
wire n8940;
wire n8941;
wire n8942;
wire n8943;
wire n8944;
wire n8945;
wire n8946;
wire n8947;
wire n8948;
wire n8949;
wire n8950;
wire n8951;
wire n8952;
wire n8953;
wire n8954;
wire n8955;
wire n8956;
wire n8957;
wire n8958;
wire n8959;
wire n8960;
wire n8961;
wire n8962;
wire n8963;
wire n8964;
wire n8965;
wire n8966;
wire n8967;
wire n8968;
wire n8969;
wire n8970;
wire n8971;
wire n8972;
wire n8973;
wire n8974;
wire n8975;
wire n8976;
wire n8977;
wire n8978;
wire n8979;
wire n8980;
wire n8981;
wire n8982;
wire n8983;
wire n8984;
wire n8985;
wire n8986;
wire n8987;
wire n8988;
wire n8989;
wire n8990;
wire n8991;
wire n8992;
wire n8993;
wire n8994;
wire n8995;
wire n8996;
wire n8997;
wire n8998;
wire n8999;
wire n9000;
wire n9001;
wire n9002;
wire n9003;
wire n9004;
wire n9005;
wire n9006;
wire n9007;
wire n9008;
wire n9009;
wire n9010;
wire n9011;
wire n9012;
wire n9013;
wire n9014;
wire n9015;
wire n9016;
wire n9017;
wire n9018;
wire n9019;
wire n9020;
wire n9021;
wire n9022;
wire n9023;
wire n9024;
wire n9025;
wire n9026;
wire n9027;
wire n9028;
wire n9029;
wire n9030;
wire n9031;
wire n9032;
wire n9033;
wire n9034;
wire n9035;
wire n9036;
wire n9037;
wire n9038;
wire n9039;
wire n9040;
wire n9041;
wire n9042;
xor (out,n0,n4650);
nand (n0,n1,n11);
or (n1,n2,n4);
not (n2,n3);
not (n4,n5);
nand (n5,n6,n8,n10);
not (n6,n7);
not (n8,n9);
nand (n11,n12,n4);
xor (n12,n13,n1109);
and (n13,n14,n1108);
not (n14,n15);
nor (n15,n16,n986);
or (n16,n17,n985);
and (n17,n18,n807);
xor (n18,n19,n579);
xor (n19,n20,n438);
xor (n20,n21,n229);
xor (n21,n22,n188);
xor (n22,n23,n107);
or (n23,n24,n106);
and (n24,n25,n78);
xor (n25,n26,n54);
nand (n26,n27,n48);
or (n27,n28,n43);
nand (n28,n29,n37);
not (n29,n30);
nor (n30,n31,n35);
and (n31,n32,n34);
not (n32,n33);
and (n35,n33,n36);
not (n36,n34);
not (n37,n38);
nand (n38,n39,n42);
nand (n39,n40,n33);
not (n40,n41);
nand (n42,n32,n41);
nor (n43,n44,n46);
and (n44,n36,n45);
and (n46,n34,n47);
not (n47,n45);
or (n48,n37,n49);
nor (n49,n50,n52);
and (n50,n36,n51);
and (n52,n34,n53);
not (n53,n51);
nand (n54,n55,n72);
or (n55,n56,n67);
nand (n56,n57,n62);
nor (n57,n58,n60);
and (n58,n36,n59);
and (n60,n34,n61);
not (n61,n59);
nand (n62,n63,n66);
or (n63,n59,n64);
not (n64,n65);
nand (n66,n64,n59);
nor (n67,n68,n70);
and (n68,n64,n69);
and (n70,n65,n71);
not (n71,n69);
or (n72,n57,n73);
nor (n73,n74,n76);
and (n74,n64,n75);
and (n76,n65,n77);
not (n77,n75);
nand (n78,n79,n100);
or (n79,n80,n95);
nand (n80,n81,n88);
not (n81,n82);
nand (n82,n83,n87);
or (n83,n84,n86);
not (n84,n85);
nand (n87,n84,n86);
not (n88,n89);
nor (n89,n90,n93);
and (n90,n91,n92);
not (n91,n86);
and (n93,n86,n94);
not (n94,n92);
nor (n95,n96,n98);
and (n96,n94,n97);
and (n98,n92,n99);
not (n99,n97);
or (n100,n81,n101);
nor (n101,n102,n104);
and (n102,n94,n103);
and (n104,n92,n105);
not (n105,n103);
and (n106,n26,n54);
xor (n107,n108,n161);
xor (n108,n109,n135);
nand (n109,n110,n129);
or (n110,n111,n123);
nand (n111,n112,n119);
not (n112,n113);
nand (n113,n114,n118);
or (n114,n115,n116);
not (n116,n117);
nand (n118,n115,n116);
nand (n119,n120,n122);
or (n120,n121,n116);
nand (n122,n121,n116);
nor (n123,n124,n127);
and (n124,n125,n126);
not (n125,n121);
and (n127,n121,n128);
not (n128,n126);
or (n129,n112,n130);
nor (n130,n131,n133);
and (n131,n125,n132);
and (n133,n121,n134);
not (n134,n132);
nand (n135,n136,n154);
or (n136,n137,n149);
not (n137,n138);
nor (n138,n139,n145);
nand (n139,n140,n144);
or (n140,n141,n142);
not (n142,n143);
nand (n144,n141,n142);
nor (n145,n146,n147);
and (n146,n84,n141);
and (n147,n85,n148);
not (n148,n141);
nor (n149,n150,n152);
and (n150,n84,n151);
and (n152,n85,n153);
not (n153,n151);
or (n154,n155,n156);
not (n155,n139);
nor (n156,n157,n159);
and (n157,n84,n158);
and (n159,n85,n160);
not (n160,n158);
nand (n161,n162,n182);
or (n162,n163,n177);
not (n163,n164);
and (n164,n165,n172);
nor (n165,n166,n170);
and (n166,n167,n169);
not (n167,n168);
and (n170,n168,n171);
not (n171,n169);
nor (n172,n173,n176);
and (n173,n174,n171);
not (n174,n175);
and (n176,n175,n169);
nor (n177,n178,n180);
and (n178,n179,n174);
and (n180,n181,n175);
not (n181,n179);
or (n182,n165,n183);
nor (n183,n184,n186);
and (n184,n185,n174);
and (n186,n187,n175);
not (n187,n185);
xor (n188,n189,n204);
xor (n189,n190,n198);
nand (n190,n191,n192);
or (n191,n80,n101);
or (n192,n81,n193);
nor (n193,n194,n196);
and (n194,n94,n195);
and (n196,n92,n197);
not (n197,n195);
nand (n198,n199,n200);
or (n199,n56,n73);
or (n200,n57,n201);
nor (n201,n202,n203);
and (n202,n64,n45);
and (n203,n65,n47);
nand (n204,n205,n217);
or (n205,n206,n212);
not (n206,n207);
nand (n207,n208,n210);
or (n208,n71,n209);
or (n210,n211,n69);
not (n211,n209);
not (n212,n213);
nand (n213,n214,n216);
or (n214,n64,n215);
nand (n216,n215,n64);
or (n217,n218,n224);
not (n218,n219);
nor (n219,n220,n213);
nor (n220,n221,n223);
and (n221,n209,n222);
not (n222,n215);
and (n223,n211,n215);
nor (n224,n225,n227);
and (n225,n211,n226);
and (n227,n209,n228);
not (n228,n226);
or (n229,n230,n437);
and (n230,n231,n376);
xor (n231,n232,n292);
xor (n232,n233,n284);
xor (n233,n234,n260);
nand (n234,n235,n253);
or (n235,n236,n248);
not (n236,n237);
nor (n237,n238,n245);
nor (n238,n239,n243);
and (n239,n240,n242);
not (n240,n241);
and (n243,n241,n244);
not (n244,n242);
nand (n245,n246,n247);
or (n246,n244,n92);
or (n247,n94,n242);
nor (n248,n249,n251);
and (n249,n240,n250);
and (n251,n241,n252);
not (n252,n250);
or (n253,n254,n255);
not (n254,n245);
nor (n255,n256,n258);
and (n256,n240,n257);
and (n258,n241,n259);
not (n259,n257);
nand (n260,n261,n278);
or (n261,n262,n266);
not (n262,n263);
nand (n263,n264,n265);
or (n264,n187,n168);
or (n265,n167,n185);
nand (n266,n267,n274);
not (n267,n268);
nand (n268,n269,n273);
or (n269,n270,n271);
not (n271,n272);
nand (n273,n270,n271);
nor (n274,n275,n277);
and (n275,n276,n167);
not (n276,n270);
and (n277,n270,n168);
or (n278,n267,n279);
nor (n279,n280,n282);
and (n280,n281,n167);
and (n282,n283,n168);
not (n283,n281);
nand (n284,n285,n286);
or (n285,n177,n165);
or (n286,n163,n287);
nor (n287,n288,n290);
and (n288,n289,n174);
and (n290,n291,n175);
not (n291,n289);
xor (n292,n293,n332);
xor (n293,n294,n318);
nand (n294,n295,n311);
or (n295,n296,n306);
not (n296,n297);
nor (n297,n298,n302);
nand (n298,n299,n301);
or (n299,n300,n240);
nand (n301,n300,n240);
nor (n302,n303,n304);
and (n303,n40,n300);
and (n304,n41,n305);
not (n305,n300);
nor (n306,n307,n309);
and (n307,n40,n308);
and (n309,n41,n310);
not (n310,n308);
or (n311,n312,n313);
not (n312,n298);
nor (n313,n314,n316);
and (n314,n40,n315);
and (n316,n41,n317);
not (n317,n315);
nand (n318,n319,n326);
or (n319,n320,n111);
not (n320,n321);
nand (n321,n322,n325);
or (n322,n121,n323);
not (n323,n324);
or (n325,n125,n324);
or (n326,n112,n327);
nor (n327,n328,n330);
and (n328,n125,n329);
and (n330,n121,n331);
not (n331,n329);
or (n332,n333,n375);
and (n333,n334,n354);
xor (n334,n335,n341);
nand (n335,n336,n340);
or (n336,n80,n337);
nor (n337,n338,n339);
and (n338,n259,n92);
and (n339,n257,n94);
or (n340,n81,n95);
nand (n341,n342,n348);
or (n342,n218,n343);
nor (n343,n344,n346);
and (n344,n211,n345);
and (n346,n209,n347);
not (n347,n345);
or (n348,n349,n212);
nor (n349,n350,n352);
and (n350,n211,n351);
and (n352,n209,n353);
not (n353,n351);
nand (n354,n355,n369);
or (n355,n356,n366);
not (n356,n357);
and (n357,n358,n363);
nor (n358,n359,n361);
and (n359,n211,n360);
and (n361,n209,n362);
not (n362,n360);
nor (n363,n364,n365);
and (n364,n271,n362);
and (n365,n272,n360);
nor (n366,n367,n368);
and (n367,n271,n281);
and (n368,n272,n283);
or (n369,n358,n370);
nor (n370,n371,n373);
and (n371,n271,n372);
and (n373,n272,n374);
not (n374,n372);
and (n375,n335,n341);
or (n376,n377,n436);
and (n377,n378,n411);
xor (n378,n379,n380);
not (n379,n318);
or (n380,n381,n410);
and (n381,n382,n401);
xor (n382,n383,n392);
nand (n383,n384,n388);
or (n384,n296,n385);
nor (n385,n386,n387);
and (n386,n40,n45);
and (n387,n41,n47);
or (n388,n312,n389);
nor (n389,n390,n391);
and (n390,n40,n51);
and (n391,n41,n53);
nand (n392,n393,n397);
or (n393,n28,n394);
nor (n394,n395,n396);
and (n395,n36,n69);
and (n396,n34,n71);
or (n397,n37,n398);
nor (n398,n399,n400);
and (n399,n36,n75);
and (n400,n34,n77);
nand (n401,n402,n406);
or (n402,n137,n403);
nor (n403,n404,n405);
and (n404,n84,n97);
and (n405,n85,n99);
or (n406,n155,n407);
nor (n407,n408,n409);
and (n408,n84,n103);
and (n409,n85,n105);
and (n410,n383,n392);
or (n411,n412,n435);
and (n412,n413,n429);
xor (n413,n414,n423);
nand (n414,n415,n419);
or (n415,n56,n416);
nor (n416,n417,n418);
and (n417,n64,n351);
and (n418,n65,n353);
or (n419,n57,n420);
nor (n420,n421,n422);
and (n421,n64,n226);
and (n422,n65,n228);
nand (n423,n424,n428);
or (n424,n218,n425);
nor (n425,n426,n427);
and (n426,n211,n372);
and (n427,n209,n374);
or (n428,n212,n343);
nand (n429,n430,n431);
or (n430,n320,n112);
or (n431,n111,n432);
nor (n432,n433,n434);
and (n433,n125,n158);
and (n434,n121,n160);
and (n435,n414,n423);
and (n436,n379,n380);
and (n437,n232,n292);
xor (n438,n439,n496);
xor (n439,n440,n463);
xor (n440,n441,n457);
xor (n441,n442,n448);
nand (n442,n443,n444);
or (n443,n236,n255);
or (n444,n254,n445);
nor (n445,n446,n447);
and (n446,n240,n97);
and (n447,n241,n99);
nand (n448,n449,n453);
or (n449,n356,n450);
nor (n450,n451,n452);
and (n451,n271,n345);
and (n452,n272,n347);
or (n453,n358,n454);
nor (n454,n455,n456);
and (n455,n271,n351);
and (n456,n272,n353);
nand (n457,n458,n459);
or (n458,n266,n279);
or (n459,n267,n460);
nor (n460,n461,n462);
and (n461,n167,n372);
and (n462,n374,n168);
xor (n463,n464,n477);
xor (n464,n465,n471);
nand (n465,n466,n467);
or (n466,n296,n313);
or (n467,n312,n468);
nor (n468,n469,n470);
and (n469,n40,n250);
and (n470,n41,n252);
nand (n471,n472,n473);
or (n472,n28,n49);
or (n473,n37,n474);
nor (n474,n475,n476);
and (n475,n36,n308);
and (n476,n34,n310);
not (n477,n478);
nand (n478,n479,n492);
or (n479,n480,n489);
nand (n480,n481,n486);
nor (n481,n482,n484);
and (n482,n125,n483);
and (n484,n121,n485);
not (n485,n483);
nand (n486,n487,n488);
or (n487,n483,n142);
nand (n488,n142,n483);
nor (n489,n490,n491);
and (n490,n142,n324);
and (n491,n143,n323);
or (n492,n481,n493);
nor (n493,n494,n495);
and (n494,n142,n329);
and (n495,n143,n331);
or (n496,n497,n578);
and (n497,n498,n562);
xor (n498,n499,n538);
or (n499,n500,n537);
and (n500,n501,n531);
xor (n501,n502,n525);
nand (n502,n503,n521);
or (n503,n504,n509);
not (n504,n505);
nand (n505,n506,n507);
or (n506,n115,n128);
or (n507,n508,n126);
not (n508,n115);
not (n509,n510);
nor (n510,n511,n517);
nand (n511,n512,n516);
or (n512,n513,n514);
not (n514,n515);
nand (n516,n513,n514);
nor (n517,n518,n519);
and (n518,n513,n508);
and (n519,n115,n520);
not (n520,n513);
nand (n521,n511,n522);
nand (n522,n523,n524);
or (n523,n115,n134);
or (n524,n508,n132);
nand (n525,n526,n530);
or (n526,n236,n527);
nor (n527,n528,n529);
and (n528,n240,n315);
and (n529,n241,n317);
or (n530,n254,n248);
nand (n531,n532,n536);
or (n532,n266,n533);
nor (n533,n534,n535);
and (n534,n179,n167);
and (n535,n181,n168);
or (n536,n267,n262);
and (n537,n502,n525);
or (n538,n539,n561);
and (n539,n540,n558);
xor (n540,n541,n549);
nand (n541,n542,n548);
or (n542,n163,n543);
nor (n543,n544,n546);
and (n544,n545,n174);
and (n546,n547,n175);
not (n547,n545);
or (n548,n165,n287);
nand (n549,n550,n554);
or (n550,n480,n551);
nor (n551,n552,n553);
and (n552,n142,n151);
and (n553,n143,n153);
or (n554,n481,n555);
nor (n555,n556,n557);
and (n556,n142,n158);
and (n557,n143,n160);
nand (n558,n559,n560);
or (n559,n296,n389);
or (n560,n312,n306);
and (n561,n541,n549);
or (n562,n563,n577);
and (n563,n564,n574);
xor (n564,n565,n571);
nand (n565,n566,n567);
or (n566,n137,n407);
or (n567,n155,n568);
nor (n568,n569,n570);
and (n569,n84,n195);
and (n570,n85,n197);
nand (n571,n572,n573);
or (n572,n28,n398);
or (n573,n37,n43);
nand (n574,n575,n576);
or (n575,n56,n420);
or (n576,n57,n67);
and (n577,n565,n571);
and (n578,n499,n538);
xor (n579,n580,n699);
xor (n580,n581,n657);
or (n581,n582,n656);
and (n582,n583,n649);
xor (n583,n584,n585);
xor (n584,n498,n562);
or (n585,n586,n648);
and (n586,n587,n647);
xor (n587,n588,n611);
or (n588,n589,n610);
and (n589,n590,n604);
xor (n590,n591,n598);
nand (n591,n592,n596);
or (n592,n593,n80);
nor (n593,n594,n595);
and (n594,n94,n250);
and (n595,n92,n252);
nand (n596,n597,n82);
not (n597,n337);
nand (n598,n599,n603);
or (n599,n356,n600);
nor (n600,n601,n602);
and (n601,n271,n185);
and (n602,n272,n187);
or (n603,n358,n366);
nand (n604,n605,n609);
or (n605,n266,n606);
nor (n606,n607,n608);
and (n607,n289,n167);
and (n608,n168,n291);
or (n609,n267,n533);
and (n610,n591,n598);
or (n611,n612,n646);
and (n612,n613,n640);
xor (n613,n614,n633);
nand (n614,n615,n629);
or (n615,n616,n624);
not (n616,n617);
nor (n617,n618,n622);
and (n618,n619,n620);
not (n620,n621);
and (n622,n623,n621);
not (n623,n619);
not (n624,n625);
nand (n625,n617,n626);
nand (n626,n627,n628);
or (n627,n619,n514);
nand (n628,n619,n514);
not (n629,n630);
nor (n630,n631,n632);
and (n631,n514,n132);
and (n632,n515,n134);
nand (n633,n634,n638);
or (n634,n509,n635);
nor (n635,n636,n637);
and (n636,n508,n329);
and (n637,n115,n331);
or (n638,n639,n504);
not (n639,n511);
nand (n640,n641,n645);
or (n641,n480,n642);
nor (n642,n643,n644);
and (n643,n142,n195);
and (n644,n143,n197);
or (n645,n481,n551);
and (n646,n614,n633);
xor (n647,n540,n558);
and (n648,n588,n611);
or (n649,n650,n655);
and (n650,n651,n654);
xor (n651,n652,n653);
xor (n652,n564,n574);
xor (n653,n501,n531);
xor (n654,n334,n354);
and (n655,n652,n653);
and (n656,n584,n585);
xor (n657,n658,n692);
xor (n658,n659,n662);
or (n659,n660,n661);
and (n660,n293,n332);
and (n661,n294,n318);
xor (n662,n663,n680);
xor (n663,n664,n677);
or (n664,n665,n676);
and (n665,n666,n673);
xor (n666,n667,n670);
nand (n667,n668,n669);
or (n668,n218,n349);
or (n669,n224,n212);
nand (n670,n671,n672);
or (n671,n356,n370);
or (n672,n358,n450);
nand (n673,n674,n675);
or (n674,n480,n555);
or (n675,n481,n489);
and (n676,n667,n670);
or (n677,n678,n679);
and (n678,n233,n284);
and (n679,n234,n260);
or (n680,n681,n691);
and (n681,n682,n688);
xor (n682,n683,n685);
nand (n683,n684,n522);
or (n684,n510,n511);
nand (n685,n686,n687);
or (n686,n111,n327);
or (n687,n112,n123);
nand (n688,n689,n690);
or (n689,n137,n568);
or (n690,n155,n149);
and (n691,n683,n685);
or (n692,n693,n698);
and (n693,n694,n697);
xor (n694,n695,n696);
xor (n695,n682,n688);
xor (n696,n666,n673);
xor (n697,n25,n78);
and (n698,n695,n696);
or (n699,n700,n806);
and (n700,n701,n805);
xor (n701,n702,n703);
xor (n702,n694,n697);
or (n703,n704,n804);
and (n704,n705,n803);
xor (n705,n706,n730);
or (n706,n707,n729);
and (n707,n708,n723);
xor (n708,n709,n715);
nand (n709,n710,n714);
or (n710,n236,n711);
nor (n711,n712,n713);
and (n712,n240,n308);
and (n713,n241,n310);
or (n714,n254,n527);
nand (n715,n716,n722);
or (n716,n163,n717);
nor (n717,n718,n720);
and (n718,n174,n719);
and (n720,n721,n175);
not (n721,n719);
or (n722,n165,n543);
nand (n723,n724,n728);
or (n724,n509,n725);
nor (n725,n726,n727);
and (n726,n508,n324);
and (n727,n115,n323);
or (n728,n639,n635);
and (n729,n709,n715);
or (n730,n731,n802);
and (n731,n732,n780);
xor (n732,n733,n757);
or (n733,n734,n756);
and (n734,n735,n750);
xor (n735,n736,n742);
nand (n736,n737,n741);
or (n737,n480,n738);
nor (n738,n739,n740);
and (n739,n142,n103);
and (n740,n143,n105);
or (n741,n481,n642);
nand (n742,n743,n748);
or (n743,n744,n296);
not (n744,n745);
nand (n745,n746,n747);
or (n746,n41,n77);
or (n747,n40,n75);
nand (n748,n749,n298);
not (n749,n385);
nand (n750,n751,n755);
or (n751,n28,n752);
nor (n752,n753,n754);
and (n753,n36,n226);
and (n754,n34,n228);
or (n755,n37,n394);
and (n756,n736,n742);
or (n757,n758,n779);
and (n758,n759,n772);
xor (n759,n760,n766);
nand (n760,n761,n765);
or (n761,n137,n762);
nor (n762,n763,n764);
and (n763,n259,n85);
and (n764,n257,n84);
or (n765,n155,n403);
nand (n766,n767,n771);
or (n767,n56,n768);
nor (n768,n769,n770);
and (n769,n64,n345);
and (n770,n65,n347);
or (n771,n57,n416);
nand (n772,n773,n778);
or (n773,n218,n774);
not (n774,n775);
nor (n775,n776,n777);
and (n776,n283,n211);
and (n777,n281,n209);
or (n778,n425,n212);
and (n779,n760,n766);
or (n780,n781,n801);
and (n781,n782,n795);
xor (n782,n783,n789);
nand (n783,n784,n788);
or (n784,n625,n785);
nor (n785,n786,n787);
and (n786,n128,n515);
and (n787,n126,n514);
or (n788,n617,n630);
nand (n789,n790,n794);
or (n790,n80,n791);
nor (n791,n792,n793);
and (n792,n94,n315);
and (n793,n92,n317);
or (n794,n81,n593);
nand (n795,n796,n800);
or (n796,n356,n797);
nor (n797,n798,n799);
and (n798,n271,n179);
and (n799,n272,n181);
or (n800,n358,n600);
and (n801,n783,n789);
and (n802,n733,n757);
xor (n803,n378,n411);
and (n804,n706,n730);
xor (n805,n231,n376);
and (n806,n702,n703);
or (n807,n808,n984);
and (n808,n809,n854);
xor (n809,n810,n853);
or (n810,n811,n852);
and (n811,n812,n845);
xor (n812,n813,n814);
xor (n813,n587,n647);
or (n814,n815,n844);
and (n815,n816,n843);
xor (n816,n817,n842);
or (n817,n818,n841);
and (n818,n819,n833);
xor (n819,n820,n826);
nand (n820,n821,n825);
or (n821,n266,n822);
nor (n822,n823,n824);
and (n823,n545,n167);
and (n824,n168,n547);
or (n825,n267,n606);
nand (n826,n827,n831);
or (n827,n828,n111);
nor (n828,n829,n830);
and (n829,n125,n151);
and (n830,n121,n153);
nand (n831,n832,n113);
not (n832,n432);
nand (n833,n834,n840);
or (n834,n163,n835);
nor (n835,n836,n838);
and (n836,n174,n837);
and (n838,n839,n175);
not (n839,n837);
or (n840,n165,n717);
and (n841,n820,n826);
xor (n842,n382,n401);
xor (n843,n613,n640);
and (n844,n817,n842);
or (n845,n846,n851);
and (n846,n847,n850);
xor (n847,n848,n849);
xor (n848,n590,n604);
xor (n849,n413,n429);
xor (n850,n708,n723);
and (n851,n848,n849);
and (n852,n813,n814);
xor (n853,n583,n649);
or (n854,n855,n983);
and (n855,n856,n982);
xor (n856,n857,n858);
xor (n857,n651,n654);
or (n858,n859,n981);
and (n859,n860,n980);
xor (n860,n861,n896);
or (n861,n862,n895);
and (n862,n863,n871);
xor (n863,n864,n870);
nand (n864,n865,n869);
or (n865,n236,n866);
nor (n866,n867,n868);
and (n867,n240,n51);
and (n868,n241,n53);
or (n869,n254,n711);
not (n870,n723);
or (n871,n872,n894);
and (n872,n873,n887);
xor (n873,n874,n880);
nand (n874,n875,n879);
or (n875,n137,n876);
nor (n876,n877,n878);
and (n877,n250,n84);
and (n878,n85,n252);
or (n879,n155,n762);
nand (n880,n881,n886);
or (n881,n882,n218);
not (n882,n883);
nor (n883,n884,n885);
and (n884,n187,n211);
and (n885,n185,n209);
nand (n886,n775,n213);
nand (n887,n888,n893);
or (n888,n356,n889);
not (n889,n890);
nand (n890,n891,n892);
or (n891,n291,n272);
or (n892,n271,n289);
or (n893,n358,n797);
and (n894,n874,n880);
and (n895,n864,n870);
or (n896,n897,n979);
and (n897,n898,n957);
xor (n898,n899,n933);
or (n899,n900,n932);
and (n900,n901,n926);
xor (n901,n902,n918);
nand (n902,n903,n915);
or (n903,n904,n910);
nand (n904,n905,n909);
or (n905,n906,n907);
not (n907,n908);
nand (n909,n907,n906);
nor (n910,n904,n911);
nor (n911,n912,n913);
and (n912,n620,n906);
and (n913,n621,n914);
not (n914,n906);
nor (n915,n916,n917);
and (n916,n132,n621);
and (n917,n134,n620);
nand (n918,n919,n924);
or (n919,n920,n625);
not (n920,n921);
nor (n921,n922,n923);
and (n922,n329,n515);
and (n923,n331,n514);
nand (n924,n925,n616);
not (n925,n785);
nand (n926,n927,n931);
or (n927,n111,n928);
nor (n928,n929,n930);
and (n929,n125,n195);
and (n930,n121,n197);
or (n931,n112,n828);
and (n932,n902,n918);
or (n933,n934,n956);
and (n934,n935,n950);
xor (n935,n936,n943);
nand (n936,n937,n938);
or (n937,n254,n866);
nand (n938,n939,n237);
not (n939,n940);
nor (n940,n941,n942);
and (n941,n240,n45);
and (n942,n241,n47);
nand (n943,n944,n949);
or (n944,n945,n296);
not (n945,n946);
nand (n946,n947,n948);
or (n947,n41,n71);
or (n948,n40,n69);
nand (n949,n298,n745);
nand (n950,n951,n955);
or (n951,n480,n952);
nor (n952,n953,n954);
and (n953,n142,n97);
and (n954,n143,n99);
or (n955,n481,n738);
and (n956,n936,n943);
or (n957,n958,n978);
and (n958,n959,n972);
xor (n959,n960,n966);
nand (n960,n961,n965);
or (n961,n28,n962);
nor (n962,n963,n964);
and (n963,n36,n351);
and (n964,n34,n353);
or (n965,n37,n752);
nand (n966,n967,n971);
or (n967,n56,n968);
nor (n968,n969,n970);
and (n969,n372,n64);
and (n970,n65,n374);
or (n971,n57,n768);
nand (n972,n973,n977);
or (n973,n509,n974);
nor (n974,n975,n976);
and (n975,n508,n158);
and (n976,n115,n160);
or (n977,n639,n725);
and (n978,n960,n966);
and (n979,n899,n933);
xor (n980,n732,n780);
and (n981,n861,n896);
xor (n982,n705,n803);
and (n983,n857,n858);
and (n984,n810,n853);
and (n985,n19,n579);
xor (n986,n987,n1105);
xor (n987,n988,n1081);
xor (n988,n989,n1078);
xor (n989,n990,n1035);
xor (n990,n991,n1015);
xor (n991,n992,n995);
or (n992,n993,n994);
and (n993,n441,n457);
and (n994,n442,n448);
xor (n995,n996,n1009);
xor (n996,n997,n1003);
nand (n997,n998,n999);
or (n998,n356,n454);
or (n999,n358,n1000);
nor (n1000,n1001,n1002);
and (n1001,n271,n226);
and (n1002,n228,n272);
nand (n1003,n1004,n1005);
or (n1004,n266,n460);
or (n1005,n267,n1006);
nor (n1006,n1007,n1008);
and (n1007,n167,n345);
and (n1008,n347,n168);
nand (n1009,n1010,n1011);
or (n1010,n137,n156);
or (n1011,n155,n1012);
nor (n1012,n1013,n1014);
and (n1013,n84,n324);
and (n1014,n85,n323);
xor (n1015,n1016,n1029);
xor (n1016,n1017,n1023);
nand (n1017,n1018,n1019);
or (n1018,n296,n468);
or (n1019,n312,n1020);
nor (n1020,n1021,n1022);
and (n1021,n40,n257);
and (n1022,n41,n259);
nand (n1023,n1024,n1025);
or (n1024,n163,n183);
or (n1025,n165,n1026);
nor (n1026,n1027,n1028);
and (n1027,n281,n174);
and (n1028,n283,n175);
nand (n1029,n1030,n1031);
or (n1030,n474,n28);
or (n1031,n37,n1032);
nor (n1032,n1033,n1034);
and (n1033,n36,n315);
and (n1034,n34,n317);
xor (n1035,n1036,n1075);
xor (n1036,n1037,n1055);
xor (n1037,n1038,n1049);
xor (n1038,n1039,n1043);
nand (n1039,n1040,n1042);
or (n1040,n1041,n113);
not (n1041,n111);
not (n1042,n130);
nand (n1043,n1044,n1045);
or (n1044,n480,n493);
or (n1045,n481,n1046);
nor (n1046,n1047,n1048);
and (n1047,n142,n126);
and (n1048,n143,n128);
nand (n1049,n1050,n1051);
or (n1050,n80,n193);
or (n1051,n81,n1052);
nor (n1052,n1053,n1054);
and (n1053,n94,n151);
and (n1054,n92,n153);
xor (n1055,n1056,n1069);
xor (n1056,n1057,n1063);
nand (n1057,n1058,n1059);
or (n1058,n56,n201);
or (n1059,n57,n1060);
nor (n1060,n1061,n1062);
and (n1061,n64,n51);
and (n1062,n65,n53);
nand (n1063,n1064,n1065);
or (n1064,n206,n218);
or (n1065,n212,n1066);
nor (n1066,n1067,n1068);
and (n1067,n211,n75);
and (n1068,n209,n77);
nand (n1069,n1070,n1074);
or (n1070,n1071,n254);
nor (n1071,n1072,n1073);
and (n1072,n240,n103);
and (n1073,n241,n105);
or (n1074,n236,n445);
or (n1075,n1076,n1077);
and (n1076,n464,n477);
and (n1077,n465,n471);
or (n1078,n1079,n1080);
and (n1079,n439,n496);
and (n1080,n440,n463);
xor (n1081,n1082,n1102);
xor (n1082,n1083,n1086);
or (n1083,n1084,n1085);
and (n1084,n658,n692);
and (n1085,n659,n662);
xor (n1086,n1087,n1094);
xor (n1087,n1088,n1091);
or (n1088,n1089,n1090);
and (n1089,n663,n680);
and (n1090,n664,n677);
or (n1091,n1092,n1093);
and (n1092,n22,n188);
and (n1093,n23,n107);
xor (n1094,n1095,n1099);
xor (n1095,n478,n1096);
or (n1096,n1097,n1098);
and (n1097,n108,n161);
and (n1098,n109,n135);
or (n1099,n1100,n1101);
and (n1100,n189,n204);
and (n1101,n190,n198);
or (n1102,n1103,n1104);
and (n1103,n20,n438);
and (n1104,n21,n229);
or (n1105,n1106,n1107);
and (n1106,n580,n699);
and (n1107,n581,n657);
nand (n1108,n16,n986);
nand (n1109,n1110,n2504);
not (n1110,n1111);
nand (n1111,n1112,n2492,n2503);
nand (n1112,n1113,n2421);
nand (n1113,n1114,n2415);
or (n1114,n1115,n2284);
not (n1115,n1116);
nand (n1116,n1117,n2283);
or (n1117,n1118,n2146);
nor (n1118,n1119,n1856);
xor (n1119,n1120,n1849);
xor (n1120,n1121,n1576);
xor (n1121,n1122,n1475);
xor (n1122,n1123,n1307);
or (n1123,n1124,n1306);
and (n1124,n1125,n1204);
xor (n1125,n1126,n1159);
xor (n1126,n1127,n1150);
xor (n1127,n1128,n1137);
nand (n1128,n1129,n1133);
or (n1129,n509,n1130);
nor (n1130,n1131,n1132);
and (n1131,n197,n115);
and (n1132,n195,n508);
or (n1133,n639,n1134);
nor (n1134,n1135,n1136);
and (n1135,n153,n115);
and (n1136,n151,n508);
nand (n1137,n1138,n1144);
or (n1138,n163,n1139);
nor (n1139,n1140,n1142);
and (n1140,n1141,n174);
and (n1142,n175,n1143);
not (n1143,n1141);
or (n1144,n1145,n165);
nor (n1145,n1146,n1148);
and (n1146,n1147,n174);
and (n1148,n175,n1149);
not (n1149,n1147);
nand (n1150,n1151,n1155);
or (n1151,n80,n1152);
nor (n1152,n1153,n1154);
and (n1153,n94,n45);
and (n1154,n92,n47);
or (n1155,n81,n1156);
nor (n1156,n1157,n1158);
and (n1157,n94,n51);
and (n1158,n92,n53);
xor (n1159,n1160,n1182);
xor (n1160,n1161,n1171);
nand (n1161,n1162,n1166);
or (n1162,n356,n1163);
nor (n1163,n1164,n1165);
and (n1164,n271,n719);
and (n1165,n272,n721);
or (n1166,n358,n1167);
not (n1167,n1168);
nand (n1168,n1169,n1170);
or (n1169,n547,n272);
or (n1170,n271,n545);
nand (n1171,n1172,n1178);
or (n1172,n266,n1173);
nor (n1173,n1174,n1176);
and (n1174,n1175,n167);
and (n1176,n1177,n168);
not (n1177,n1175);
or (n1178,n267,n1179);
nor (n1179,n1180,n1181);
and (n1180,n837,n167);
and (n1181,n839,n168);
and (n1182,n1183,n1190);
nor (n1183,n1184,n174);
nor (n1184,n1185,n1188);
and (n1185,n1186,n167);
nand (n1186,n1187,n169);
and (n1188,n1189,n171);
not (n1189,n1187);
nand (n1190,n1191,n1198);
or (n1191,n1192,n1194);
not (n1192,n1193);
not (n1194,n1195);
nor (n1195,n1196,n1197);
and (n1196,n132,n908);
and (n1197,n134,n907);
or (n1198,n1199,n1200);
nand (n1199,n908,n1192);
not (n1200,n1201);
nand (n1201,n1202,n1203);
or (n1202,n126,n907);
nand (n1203,n907,n126);
or (n1204,n1205,n1305);
and (n1205,n1206,n1272);
xor (n1206,n1207,n1240);
or (n1207,n1208,n1239);
and (n1208,n1209,n1230);
xor (n1209,n1210,n1221);
nand (n1210,n1211,n1216);
or (n1211,n1212,n111);
not (n1212,n1213);
nor (n1213,n1214,n1215);
and (n1214,n250,n121);
and (n1215,n252,n125);
nand (n1216,n1217,n113);
not (n1217,n1218);
nor (n1218,n1219,n1220);
and (n1219,n259,n121);
and (n1220,n257,n125);
nand (n1221,n1222,n1226);
or (n1222,n296,n1223);
nor (n1223,n1224,n1225);
and (n1224,n40,n372);
and (n1225,n41,n374);
or (n1226,n312,n1227);
nor (n1227,n1228,n1229);
and (n1228,n347,n41);
and (n1229,n345,n40);
nand (n1230,n1231,n1235);
or (n1231,n28,n1232);
nor (n1232,n1233,n1234);
and (n1233,n36,n185);
and (n1234,n34,n187);
or (n1235,n37,n1236);
nor (n1236,n1237,n1238);
and (n1237,n36,n281);
and (n1238,n34,n283);
and (n1239,n1210,n1221);
or (n1240,n1241,n1271);
and (n1241,n1242,n1262);
xor (n1242,n1243,n1253);
nand (n1243,n1244,n1248);
or (n1244,n1245,n625);
nor (n1245,n1246,n1247);
and (n1246,n197,n515);
and (n1247,n195,n514);
nand (n1248,n1249,n616);
not (n1249,n1250);
nor (n1250,n1251,n1252);
and (n1251,n514,n151);
and (n1252,n515,n153);
nand (n1253,n1254,n1258);
or (n1254,n480,n1255);
nor (n1255,n1256,n1257);
and (n1256,n142,n308);
and (n1257,n143,n310);
or (n1258,n481,n1259);
nor (n1259,n1260,n1261);
and (n1260,n317,n143);
and (n1261,n315,n142);
nand (n1262,n1263,n1267);
or (n1263,n56,n1264);
nor (n1264,n1265,n1266);
and (n1265,n64,n289);
and (n1266,n65,n291);
or (n1267,n57,n1268);
nor (n1268,n1269,n1270);
and (n1269,n64,n179);
and (n1270,n65,n181);
and (n1271,n1243,n1253);
or (n1272,n1273,n1304);
and (n1273,n1274,n1295);
xor (n1274,n1275,n1285);
nand (n1275,n1276,n1281);
or (n1276,n1277,n218);
not (n1277,n1278);
nand (n1278,n1279,n1280);
or (n1279,n209,n721);
or (n1280,n211,n719);
or (n1281,n212,n1282);
nor (n1282,n1283,n1284);
and (n1283,n211,n545);
and (n1284,n209,n547);
nand (n1285,n1286,n1291);
or (n1286,n1287,n137);
not (n1287,n1288);
nand (n1288,n1289,n1290);
or (n1289,n85,n47);
or (n1290,n84,n45);
nand (n1291,n139,n1292);
nand (n1292,n1293,n1294);
or (n1293,n85,n53);
or (n1294,n84,n51);
nand (n1295,n1296,n1300);
or (n1296,n356,n1297);
nor (n1297,n1298,n1299);
and (n1298,n271,n1175);
and (n1299,n272,n1177);
or (n1300,n358,n1301);
nor (n1301,n1302,n1303);
and (n1302,n271,n837);
and (n1303,n272,n839);
and (n1304,n1275,n1285);
and (n1305,n1207,n1240);
and (n1306,n1126,n1159);
or (n1307,n1308,n1474);
and (n1308,n1309,n1430);
xor (n1309,n1310,n1370);
or (n1310,n1311,n1369);
and (n1311,n1312,n1337);
xor (n1312,n1313,n1314);
xor (n1313,n1183,n1190);
or (n1314,n1315,n1336);
and (n1315,n1316,n1325);
xor (n1316,n1317,n1318);
nor (n1317,n165,n1189);
nand (n1318,n1319,n1324);
or (n1319,n1199,n1320);
not (n1320,n1321);
nor (n1321,n1322,n1323);
and (n1322,n331,n907);
and (n1323,n329,n908);
nand (n1324,n1201,n1193);
nand (n1325,n1326,n1332);
or (n1326,n1327,n1331);
not (n1327,n1328);
nand (n1328,n1329,n1330);
or (n1329,n621,n160);
or (n1330,n620,n158);
not (n1331,n910);
nand (n1332,n904,n1333);
nor (n1333,n1334,n1335);
and (n1334,n324,n621);
and (n1335,n323,n620);
and (n1336,n1317,n1318);
or (n1337,n1338,n1368);
and (n1338,n1339,n1359);
xor (n1339,n1340,n1350);
nand (n1340,n1341,n1346);
or (n1341,n1342,n509);
not (n1342,n1343);
nand (n1343,n1344,n1345);
or (n1344,n115,n99);
or (n1345,n508,n97);
nand (n1346,n511,n1347);
nand (n1347,n1348,n1349);
or (n1348,n115,n105);
or (n1349,n508,n103);
nand (n1350,n1351,n1355);
or (n1351,n80,n1352);
nor (n1352,n1353,n1354);
and (n1353,n94,n69);
and (n1354,n92,n71);
or (n1355,n81,n1356);
nor (n1356,n1357,n1358);
and (n1357,n75,n94);
and (n1358,n77,n92);
nand (n1359,n1360,n1364);
or (n1360,n236,n1361);
nor (n1361,n1362,n1363);
and (n1362,n240,n351);
and (n1363,n241,n353);
or (n1364,n254,n1365);
nor (n1365,n1366,n1367);
and (n1366,n240,n226);
and (n1367,n241,n228);
and (n1368,n1340,n1350);
and (n1369,n1313,n1314);
or (n1370,n1371,n1429);
and (n1371,n1372,n1412);
xor (n1372,n1373,n1391);
xor (n1373,n1374,n1385);
xor (n1374,n1375,n1382);
nand (n1375,n1376,n1378);
or (n1376,n1377,n137);
not (n1377,n1292);
or (n1378,n1379,n155);
nor (n1379,n1380,n1381);
and (n1380,n84,n308);
and (n1381,n85,n310);
nand (n1382,n1383,n1384);
or (n1383,n1301,n356);
or (n1384,n358,n1163);
nand (n1385,n1386,n1390);
or (n1386,n266,n1387);
nor (n1387,n1388,n1389);
and (n1388,n1147,n167);
and (n1389,n1149,n168);
or (n1390,n267,n1173);
xor (n1391,n1392,n1406);
xor (n1392,n1393,n1401);
nand (n1393,n1394,n1396);
or (n1394,n1395,n1331);
not (n1395,n1333);
nand (n1396,n1397,n904);
not (n1397,n1398);
nor (n1398,n1399,n1400);
and (n1399,n331,n621);
and (n1400,n329,n620);
nand (n1401,n1402,n1404);
or (n1402,n1403,n509);
not (n1403,n1347);
nand (n1404,n1405,n511);
not (n1405,n1130);
nand (n1406,n1407,n1411);
or (n1407,n163,n1408);
nor (n1408,n1409,n1410);
and (n1409,n1189,n175);
and (n1410,n1187,n174);
or (n1411,n165,n1139);
xor (n1412,n1413,n1423);
xor (n1413,n1414,n1417);
nand (n1414,n1415,n1416);
or (n1415,n80,n1356);
or (n1416,n81,n1152);
nand (n1417,n1418,n1419);
or (n1418,n236,n1365);
or (n1419,n254,n1420);
nor (n1420,n1421,n1422);
and (n1421,n240,n69);
and (n1422,n241,n71);
nand (n1423,n1424,n1425);
or (n1424,n111,n1218);
or (n1425,n112,n1426);
nor (n1426,n1427,n1428);
and (n1427,n125,n97);
and (n1428,n121,n99);
and (n1429,n1373,n1391);
xor (n1430,n1431,n1459);
xor (n1431,n1432,n1456);
or (n1432,n1433,n1455);
and (n1433,n1434,n1449);
xor (n1434,n1435,n1443);
nand (n1435,n1436,n1437);
or (n1436,n1259,n480);
nand (n1437,n1438,n1442);
not (n1438,n1439);
nor (n1439,n1440,n1441);
and (n1440,n142,n250);
and (n1441,n143,n252);
not (n1442,n481);
nand (n1443,n1444,n1445);
or (n1444,n56,n1268);
or (n1445,n57,n1446);
nor (n1446,n1447,n1448);
and (n1447,n64,n185);
and (n1448,n65,n187);
nand (n1449,n1450,n1451);
or (n1450,n218,n1282);
or (n1451,n212,n1452);
nor (n1452,n1453,n1454);
and (n1453,n211,n289);
and (n1454,n209,n291);
and (n1455,n1435,n1443);
or (n1456,n1457,n1458);
and (n1457,n1374,n1385);
and (n1458,n1375,n1382);
nand (n1459,n1460,n1473);
or (n1460,n1461,n1465);
not (n1461,n1462);
nand (n1462,n1463,n1195);
or (n1463,n1464,n1193);
not (n1464,n1199);
not (n1465,n1466);
nand (n1466,n1467,n1468);
or (n1467,n1331,n1398);
or (n1468,n1469,n1470);
not (n1469,n904);
nor (n1470,n1471,n1472);
and (n1471,n620,n126);
and (n1472,n621,n128);
or (n1473,n1466,n1462);
and (n1474,n1310,n1370);
xor (n1475,n1476,n1512);
xor (n1476,n1477,n1480);
or (n1477,n1478,n1479);
and (n1478,n1431,n1459);
and (n1479,n1432,n1456);
xor (n1480,n1481,n1485);
xor (n1481,n1473,n1482);
or (n1482,n1483,n1484);
and (n1483,n1127,n1150);
and (n1484,n1128,n1137);
or (n1485,n1486,n1511);
and (n1486,n1487,n1502);
xor (n1487,n1488,n1494);
nand (n1488,n1489,n1490);
or (n1489,n236,n1420);
or (n1490,n254,n1491);
nor (n1491,n1492,n1493);
and (n1492,n240,n75);
and (n1493,n241,n77);
nand (n1494,n1495,n1500);
or (n1495,n1496,n112);
not (n1496,n1497);
nand (n1497,n1498,n1499);
or (n1498,n121,n105);
or (n1499,n125,n103);
nand (n1500,n1501,n1041);
not (n1501,n1426);
nand (n1502,n1503,n1507);
or (n1503,n296,n1504);
nor (n1504,n1505,n1506);
and (n1505,n40,n351);
and (n1506,n41,n353);
or (n1507,n312,n1508);
nor (n1508,n1509,n1510);
and (n1509,n40,n226);
and (n1510,n41,n228);
and (n1511,n1488,n1494);
xor (n1512,n1513,n1564);
xor (n1513,n1514,n1542);
or (n1514,n1515,n1541);
and (n1515,n1516,n1535);
xor (n1516,n1517,n1526);
nand (n1517,n1518,n1522);
or (n1518,n1519,n28);
nor (n1519,n1520,n1521);
and (n1520,n374,n34);
and (n1521,n372,n36);
or (n1522,n37,n1523);
nor (n1523,n1524,n1525);
and (n1524,n36,n345);
and (n1525,n34,n347);
nand (n1526,n1527,n1531);
or (n1527,n1528,n625);
nor (n1528,n1529,n1530);
and (n1529,n514,n158);
and (n1530,n515,n160);
nand (n1531,n616,n1532);
nand (n1532,n1533,n1534);
or (n1533,n515,n323);
or (n1534,n514,n324);
nand (n1535,n1536,n1537);
or (n1536,n480,n1439);
or (n1537,n481,n1538);
nor (n1538,n1539,n1540);
and (n1539,n142,n257);
and (n1540,n143,n259);
and (n1541,n1517,n1526);
or (n1542,n1543,n1563);
and (n1543,n1544,n1557);
xor (n1544,n1545,n1551);
nand (n1545,n1546,n1547);
or (n1546,n56,n1446);
or (n1547,n57,n1548);
nor (n1548,n1549,n1550);
and (n1549,n281,n64);
and (n1550,n65,n283);
nand (n1551,n1552,n1553);
or (n1552,n218,n1452);
or (n1553,n212,n1554);
nor (n1554,n1555,n1556);
and (n1555,n211,n179);
and (n1556,n209,n181);
nand (n1557,n1558,n1562);
or (n1558,n1559,n155);
nor (n1559,n1560,n1561);
and (n1560,n84,n315);
and (n1561,n85,n317);
or (n1562,n137,n1379);
and (n1563,n1545,n1551);
xor (n1564,n1565,n1573);
xor (n1565,n1566,n1570);
nand (n1566,n1567,n1569);
or (n1567,n1568,n625);
not (n1568,n1532);
nand (n1569,n616,n921);
nand (n1570,n1571,n1572);
or (n1571,n1496,n111);
or (n1572,n112,n928);
nand (n1573,n1574,n1575);
or (n1574,n236,n1491);
or (n1575,n254,n940);
xor (n1576,n1577,n1759);
xor (n1577,n1578,n1673);
xor (n1578,n1579,n1627);
xor (n1579,n1580,n1587);
or (n1580,n1581,n1586);
and (n1581,n1582,n1585);
xor (n1582,n1583,n1584);
xor (n1583,n1487,n1502);
xor (n1584,n1516,n1535);
xor (n1585,n1544,n1557);
and (n1586,n1583,n1584);
xor (n1587,n1588,n1615);
xor (n1588,n1589,n1604);
xor (n1589,n1590,n1598);
xor (n1590,n1591,n1594);
nand (n1591,n1592,n1593);
or (n1592,n212,n882);
or (n1593,n218,n1554);
nand (n1594,n1595,n1596);
or (n1595,n1167,n356);
nand (n1596,n890,n1597);
not (n1597,n358);
nand (n1598,n1599,n1600);
or (n1599,n80,n1156);
or (n1600,n81,n1601);
nor (n1601,n1602,n1603);
and (n1602,n94,n308);
and (n1603,n92,n310);
xor (n1604,n1605,n1612);
xor (n1605,n1606,n1609);
nand (n1606,n1607,n1608);
or (n1607,n1508,n296);
nand (n1608,n298,n946);
nand (n1609,n1610,n1611);
or (n1610,n480,n1538);
or (n1611,n481,n952);
nand (n1612,n1613,n1614);
or (n1613,n28,n1523);
or (n1614,n37,n962);
xor (n1615,n1616,n1624);
xor (n1616,n1617,n1620);
nand (n1617,n1618,n1619);
or (n1618,n56,n1548);
or (n1619,n968,n57);
nand (n1620,n1621,n1622);
or (n1621,n1134,n509);
nand (n1622,n1623,n511);
not (n1623,n974);
nand (n1624,n1625,n1626);
or (n1625,n137,n1559);
or (n1626,n155,n876);
xor (n1627,n1628,n1650);
xor (n1628,n1629,n1647);
xor (n1629,n1630,n1643);
xor (n1630,n1631,n1637);
nand (n1631,n1632,n1633);
or (n1632,n266,n1179);
or (n1633,n267,n1634);
nor (n1634,n1635,n1636);
and (n1635,n719,n167);
and (n1636,n168,n721);
nand (n1637,n1638,n1639);
or (n1638,n163,n1145);
or (n1639,n165,n1640);
nor (n1640,n1641,n1642);
and (n1641,n1175,n174);
and (n1642,n1177,n175);
nor (n1643,n1644,n1646);
and (n1644,n910,n1645);
not (n1645,n1470);
and (n1646,n904,n915);
or (n1647,n1648,n1649);
and (n1648,n1160,n1182);
and (n1649,n1161,n1171);
or (n1650,n1651,n1672);
and (n1651,n1652,n1659);
xor (n1652,n1653,n1656);
or (n1653,n1654,n1655);
and (n1654,n1392,n1406);
and (n1655,n1393,n1401);
or (n1656,n1657,n1658);
and (n1657,n1413,n1423);
and (n1658,n1414,n1417);
or (n1659,n1660,n1671);
and (n1660,n1661,n1668);
xor (n1661,n1662,n1665);
nand (n1662,n1663,n1664);
or (n1663,n296,n1227);
or (n1664,n312,n1504);
nand (n1665,n1666,n1667);
or (n1666,n28,n1236);
or (n1667,n37,n1519);
nand (n1668,n1669,n1670);
or (n1669,n625,n1250);
or (n1670,n617,n1528);
and (n1671,n1662,n1665);
and (n1672,n1653,n1656);
or (n1673,n1674,n1758);
and (n1674,n1675,n1678);
xor (n1675,n1676,n1677);
xor (n1676,n1652,n1659);
xor (n1677,n1582,n1585);
or (n1678,n1679,n1757);
and (n1679,n1680,n1683);
xor (n1680,n1681,n1682);
xor (n1681,n1661,n1668);
xor (n1682,n1434,n1449);
or (n1683,n1684,n1756);
and (n1684,n1685,n1733);
xor (n1685,n1686,n1709);
or (n1686,n1687,n1708);
and (n1687,n1688,n1701);
xor (n1688,n1689,n1695);
nand (n1689,n1690,n1694);
or (n1690,n236,n1691);
nor (n1691,n1692,n1693);
and (n1692,n240,n345);
and (n1693,n241,n347);
or (n1694,n254,n1361);
nand (n1695,n1696,n1700);
or (n1696,n111,n1697);
nor (n1697,n1698,n1699);
and (n1698,n125,n315);
and (n1699,n121,n317);
or (n1700,n112,n1212);
nand (n1701,n1702,n1707);
or (n1702,n296,n1703);
not (n1703,n1704);
nor (n1704,n1705,n1706);
and (n1705,n281,n41);
and (n1706,n283,n40);
or (n1707,n312,n1223);
and (n1708,n1689,n1695);
or (n1709,n1710,n1732);
and (n1710,n1711,n1726);
xor (n1711,n1712,n1720);
nand (n1712,n1713,n1718);
or (n1713,n1714,n28);
not (n1714,n1715);
nand (n1715,n1716,n1717);
or (n1716,n34,n181);
or (n1717,n36,n179);
nand (n1718,n1719,n38);
not (n1719,n1232);
nand (n1720,n1721,n1725);
or (n1721,n625,n1722);
nor (n1722,n1723,n1724);
and (n1723,n514,n103);
and (n1724,n515,n105);
or (n1725,n617,n1245);
nand (n1726,n1727,n1731);
or (n1727,n480,n1728);
nor (n1728,n1729,n1730);
and (n1729,n142,n51);
and (n1730,n143,n53);
or (n1731,n481,n1255);
and (n1732,n1712,n1720);
or (n1733,n1734,n1755);
and (n1734,n1735,n1749);
xor (n1735,n1736,n1742);
nand (n1736,n1737,n1741);
or (n1737,n56,n1738);
nor (n1738,n1739,n1740);
and (n1739,n64,n545);
and (n1740,n65,n547);
or (n1741,n57,n1264);
nand (n1742,n1743,n1744);
or (n1743,n1277,n212);
nand (n1744,n1745,n219);
not (n1745,n1746);
nor (n1746,n1747,n1748);
and (n1747,n211,n837);
and (n1748,n839,n209);
nand (n1749,n1750,n1754);
or (n1750,n1751,n137);
nor (n1751,n1752,n1753);
and (n1752,n84,n75);
and (n1753,n85,n77);
or (n1754,n155,n1287);
and (n1755,n1736,n1742);
and (n1756,n1686,n1709);
and (n1757,n1681,n1682);
and (n1758,n1676,n1677);
or (n1759,n1760,n1848);
and (n1760,n1761,n1813);
xor (n1761,n1762,n1763);
xor (n1762,n1125,n1204);
or (n1763,n1764,n1812);
and (n1764,n1765,n1811);
xor (n1765,n1766,n1810);
or (n1766,n1767,n1809);
and (n1767,n1768,n1787);
xor (n1768,n1769,n1775);
nand (n1769,n1770,n1774);
or (n1770,n266,n1771);
nor (n1771,n1772,n1773);
and (n1772,n167,n1141);
and (n1773,n1143,n168);
or (n1774,n267,n1387);
and (n1775,n1776,n1781);
nor (n1776,n1777,n167);
nor (n1777,n1778,n1780);
and (n1778,n1779,n271);
nand (n1779,n1187,n270);
and (n1780,n1189,n276);
nand (n1781,n1782,n1783);
or (n1782,n1192,n1320);
or (n1783,n1199,n1784);
nor (n1784,n1785,n1786);
and (n1785,n907,n324);
and (n1786,n908,n323);
or (n1787,n1788,n1808);
and (n1788,n1789,n1802);
xor (n1789,n1790,n1796);
nand (n1790,n1791,n1792);
or (n1791,n1327,n1469);
or (n1792,n1331,n1793);
nor (n1793,n1794,n1795);
and (n1794,n153,n621);
and (n1795,n151,n620);
nand (n1796,n1797,n1798);
or (n1797,n1342,n639);
or (n1798,n509,n1799);
nor (n1799,n1800,n1801);
and (n1800,n508,n257);
and (n1801,n115,n259);
nand (n1802,n1803,n1807);
or (n1803,n80,n1804);
nor (n1804,n1805,n1806);
and (n1805,n94,n226);
and (n1806,n92,n228);
or (n1807,n81,n1352);
and (n1808,n1790,n1796);
and (n1809,n1769,n1775);
xor (n1810,n1206,n1272);
xor (n1811,n1312,n1337);
and (n1812,n1766,n1810);
or (n1813,n1814,n1847);
and (n1814,n1815,n1846);
xor (n1815,n1816,n1823);
or (n1816,n1817,n1822);
and (n1817,n1818,n1821);
xor (n1818,n1819,n1820);
xor (n1819,n1316,n1325);
xor (n1820,n1274,n1295);
xor (n1821,n1242,n1262);
and (n1822,n1819,n1820);
or (n1823,n1824,n1845);
and (n1824,n1825,n1828);
xor (n1825,n1826,n1827);
xor (n1826,n1209,n1230);
xor (n1827,n1339,n1359);
or (n1828,n1829,n1844);
and (n1829,n1830,n1843);
xor (n1830,n1831,n1837);
nand (n1831,n1832,n1836);
or (n1832,n356,n1833);
nor (n1833,n1834,n1835);
and (n1834,n271,n1147);
and (n1835,n272,n1149);
or (n1836,n358,n1297);
nand (n1837,n1838,n1842);
or (n1838,n266,n1839);
nor (n1839,n1840,n1841);
and (n1840,n1189,n168);
and (n1841,n1187,n167);
or (n1842,n267,n1771);
xor (n1843,n1776,n1781);
and (n1844,n1831,n1837);
and (n1845,n1826,n1827);
xor (n1846,n1372,n1412);
and (n1847,n1816,n1823);
and (n1848,n1762,n1763);
or (n1849,n1850,n1855);
and (n1850,n1851,n1854);
xor (n1851,n1852,n1853);
xor (n1852,n1309,n1430);
xor (n1853,n1675,n1678);
xor (n1854,n1761,n1813);
and (n1855,n1852,n1853);
or (n1856,n1857,n2145);
and (n1857,n1858,n2144);
xor (n1858,n1859,n2001);
or (n1859,n1860,n2000);
and (n1860,n1861,n1944);
xor (n1861,n1862,n1863);
xor (n1862,n1680,n1683);
or (n1863,n1864,n1943);
and (n1864,n1865,n1936);
xor (n1865,n1866,n1867);
xor (n1866,n1768,n1787);
or (n1867,n1868,n1935);
and (n1868,n1869,n1912);
xor (n1869,n1870,n1893);
or (n1870,n1871,n1892);
and (n1871,n1872,n1886);
xor (n1872,n1873,n1880);
nand (n1873,n1874,n1879);
or (n1874,n1875,n296);
not (n1875,n1876);
nor (n1876,n1877,n1878);
and (n1877,n185,n41);
and (n1878,n187,n40);
nand (n1879,n1704,n298);
nand (n1880,n1881,n1885);
or (n1881,n1882,n28);
nor (n1882,n1883,n1884);
and (n1883,n291,n34);
and (n1884,n289,n36);
nand (n1885,n1715,n38);
nand (n1886,n1887,n1891);
or (n1887,n1199,n1888);
nor (n1888,n1889,n1890);
and (n1889,n907,n158);
and (n1890,n908,n160);
or (n1891,n1784,n1192);
and (n1892,n1873,n1880);
or (n1893,n1894,n1911);
and (n1894,n1895,n1905);
xor (n1895,n1896,n1897);
nor (n1896,n267,n1189);
nand (n1897,n1898,n1903);
or (n1898,n1899,n1331);
not (n1899,n1900);
nand (n1900,n1901,n1902);
or (n1901,n621,n197);
or (n1902,n620,n195);
nand (n1903,n1904,n904);
not (n1904,n1793);
nand (n1905,n1906,n1910);
or (n1906,n509,n1907);
nor (n1907,n1908,n1909);
and (n1908,n508,n250);
and (n1909,n115,n252);
or (n1910,n639,n1799);
and (n1911,n1896,n1897);
or (n1912,n1913,n1934);
and (n1913,n1914,n1928);
xor (n1914,n1915,n1922);
nand (n1915,n1916,n1920);
or (n1916,n1917,n80);
nor (n1917,n1918,n1919);
and (n1918,n351,n94);
and (n1919,n353,n92);
nand (n1920,n1921,n82);
not (n1921,n1804);
nand (n1922,n1923,n1927);
or (n1923,n236,n1924);
nor (n1924,n1925,n1926);
and (n1925,n240,n372);
and (n1926,n241,n374);
or (n1927,n254,n1691);
nand (n1928,n1929,n1933);
or (n1929,n111,n1930);
nor (n1930,n1931,n1932);
and (n1931,n125,n308);
and (n1932,n121,n310);
or (n1933,n112,n1697);
and (n1934,n1915,n1922);
and (n1935,n1870,n1893);
or (n1936,n1937,n1942);
and (n1937,n1938,n1941);
xor (n1938,n1939,n1940);
xor (n1939,n1735,n1749);
xor (n1940,n1688,n1701);
xor (n1941,n1711,n1726);
and (n1942,n1939,n1940);
and (n1943,n1866,n1867);
or (n1944,n1945,n1999);
and (n1945,n1946,n1998);
xor (n1946,n1947,n1948);
xor (n1947,n1685,n1733);
or (n1948,n1949,n1997);
and (n1949,n1950,n1996);
xor (n1950,n1951,n1974);
or (n1951,n1952,n1973);
and (n1952,n1953,n1967);
xor (n1953,n1954,n1961);
nand (n1954,n1955,n1960);
or (n1955,n1956,n480);
not (n1956,n1957);
nor (n1957,n1958,n1959);
and (n1958,n45,n143);
and (n1959,n47,n142);
or (n1960,n481,n1728);
nand (n1961,n1962,n1966);
or (n1962,n56,n1963);
nor (n1963,n1964,n1965);
and (n1964,n64,n719);
and (n1965,n65,n721);
or (n1966,n57,n1738);
nand (n1967,n1968,n1972);
or (n1968,n218,n1969);
nor (n1969,n1970,n1971);
and (n1970,n1175,n211);
and (n1971,n209,n1177);
or (n1972,n1746,n212);
and (n1973,n1954,n1961);
or (n1974,n1975,n1995);
and (n1975,n1976,n1989);
xor (n1976,n1977,n1983);
nand (n1977,n1978,n1982);
or (n1978,n625,n1979);
nor (n1979,n1980,n1981);
and (n1980,n99,n515);
and (n1981,n97,n514);
or (n1982,n617,n1722);
nand (n1983,n1984,n1988);
or (n1984,n356,n1985);
nor (n1985,n1986,n1987);
and (n1986,n1141,n271);
and (n1987,n272,n1143);
or (n1988,n358,n1833);
nand (n1989,n1990,n1994);
or (n1990,n137,n1991);
nor (n1991,n1992,n1993);
and (n1992,n84,n69);
and (n1993,n85,n71);
or (n1994,n155,n1751);
and (n1995,n1977,n1983);
xor (n1996,n1789,n1802);
and (n1997,n1951,n1974);
xor (n1998,n1825,n1828);
and (n1999,n1947,n1948);
and (n2000,n1862,n1863);
or (n2001,n2002,n2143);
and (n2002,n2003,n2006);
xor (n2003,n2004,n2005);
xor (n2004,n1765,n1811);
xor (n2005,n1815,n1846);
or (n2006,n2007,n2142);
and (n2007,n2008,n2065);
xor (n2008,n2009,n2010);
xor (n2009,n1818,n1821);
or (n2010,n2011,n2064);
and (n2011,n2012,n2063);
xor (n2012,n2013,n2014);
xor (n2013,n1869,n1912);
or (n2014,n2015,n2062);
and (n2015,n2016,n2061);
xor (n2016,n2017,n2039);
or (n2017,n2018,n2038);
and (n2018,n2019,n2032);
xor (n2019,n2020,n2026);
nand (n2020,n2021,n2025);
or (n2021,n218,n2022);
nor (n2022,n2023,n2024);
and (n2023,n1149,n209);
and (n2024,n1147,n211);
or (n2025,n1969,n212);
nand (n2026,n2027,n2031);
or (n2027,n625,n2028);
nor (n2028,n2029,n2030);
and (n2029,n514,n257);
and (n2030,n515,n259);
or (n2031,n617,n1979);
nand (n2032,n2033,n2037);
or (n2033,n356,n2034);
nor (n2034,n2035,n2036);
and (n2035,n1189,n272);
and (n2036,n1187,n271);
or (n2037,n1985,n358);
and (n2038,n2020,n2026);
or (n2039,n2040,n2060);
and (n2040,n2041,n2054);
xor (n2041,n2042,n2048);
nand (n2042,n2043,n2047);
or (n2043,n1199,n2044);
nor (n2044,n2045,n2046);
and (n2045,n153,n908);
and (n2046,n151,n907);
or (n2047,n1888,n1192);
nand (n2048,n2049,n2053);
or (n2049,n2050,n480);
nor (n2050,n2051,n2052);
and (n2051,n142,n75);
and (n2052,n143,n77);
nand (n2053,n1442,n1957);
nand (n2054,n2055,n2059);
or (n2055,n56,n2056);
nor (n2056,n2057,n2058);
and (n2057,n64,n837);
and (n2058,n65,n839);
or (n2059,n57,n1963);
and (n2060,n2042,n2048);
xor (n2061,n1914,n1928);
and (n2062,n2017,n2039);
xor (n2063,n1950,n1996);
and (n2064,n2013,n2014);
or (n2065,n2066,n2141);
and (n2066,n2067,n2134);
xor (n2067,n2068,n2069);
xor (n2068,n1830,n1843);
or (n2069,n2070,n2133);
and (n2070,n2071,n2109);
xor (n2071,n2072,n2086);
and (n2072,n2073,n2079);
nand (n2073,n2074,n2078);
or (n2074,n2075,n1331);
nor (n2075,n2076,n2077);
and (n2076,n620,n103);
and (n2077,n621,n105);
nand (n2078,n904,n1900);
not (n2079,n2080);
nand (n2080,n2081,n272);
nand (n2081,n2082,n2083);
or (n2082,n1187,n360);
nand (n2083,n2084,n211);
not (n2084,n2085);
and (n2085,n1187,n360);
or (n2086,n2087,n2108);
and (n2087,n2088,n2102);
xor (n2088,n2089,n2096);
nand (n2089,n2090,n2094);
or (n2090,n2091,n509);
nor (n2091,n2092,n2093);
and (n2092,n508,n315);
and (n2093,n115,n317);
nand (n2094,n2095,n511);
not (n2095,n1907);
nand (n2096,n2097,n2101);
or (n2097,n80,n2098);
nor (n2098,n2099,n2100);
and (n2099,n94,n345);
and (n2100,n92,n347);
or (n2101,n81,n1917);
nand (n2102,n2103,n2107);
or (n2103,n236,n2104);
nor (n2104,n2105,n2106);
and (n2105,n281,n240);
and (n2106,n241,n283);
or (n2107,n254,n1924);
and (n2108,n2089,n2096);
or (n2109,n2110,n2132);
and (n2110,n2111,n2126);
xor (n2111,n2112,n2119);
nand (n2112,n2113,n2117);
or (n2113,n2114,n111);
nor (n2114,n2115,n2116);
and (n2115,n125,n51);
and (n2116,n121,n53);
nand (n2117,n2118,n113);
not (n2118,n1930);
nand (n2119,n2120,n2125);
or (n2120,n2121,n296);
not (n2121,n2122);
nand (n2122,n2123,n2124);
or (n2123,n41,n181);
or (n2124,n40,n179);
nand (n2125,n298,n1876);
nand (n2126,n2127,n2131);
or (n2127,n28,n2128);
nor (n2128,n2129,n2130);
and (n2129,n36,n545);
and (n2130,n34,n547);
or (n2131,n37,n1882);
and (n2132,n2112,n2119);
and (n2133,n2072,n2086);
or (n2134,n2135,n2140);
and (n2135,n2136,n2139);
xor (n2136,n2137,n2138);
xor (n2137,n1976,n1989);
xor (n2138,n1895,n1905);
xor (n2139,n1872,n1886);
and (n2140,n2137,n2138);
and (n2141,n2068,n2069);
and (n2142,n2009,n2010);
and (n2143,n2004,n2005);
xor (n2144,n1851,n1854);
and (n2145,n1859,n2001);
nand (n2146,n2147,n2282);
or (n2147,n2148,n2281);
and (n2148,n2149,n2152);
xor (n2149,n2150,n2151);
xor (n2150,n1861,n1944);
xor (n2151,n2003,n2006);
or (n2152,n2153,n2280);
and (n2153,n2154,n2157);
xor (n2154,n2155,n2156);
xor (n2155,n1865,n1936);
xor (n2156,n1946,n1998);
or (n2157,n2158,n2279);
and (n2158,n2159,n2266);
xor (n2159,n2160,n2161);
xor (n2160,n1938,n1941);
or (n2161,n2162,n2265);
and (n2162,n2163,n2235);
xor (n2163,n2164,n2165);
xor (n2164,n1953,n1967);
or (n2165,n2166,n2234);
and (n2166,n2167,n2212);
xor (n2167,n2168,n2190);
or (n2168,n2169,n2189);
and (n2169,n2170,n2183);
xor (n2170,n2171,n2177);
nand (n2171,n2172,n2176);
or (n2172,n80,n2173);
nor (n2173,n2174,n2175);
and (n2174,n374,n92);
and (n2175,n372,n94);
or (n2176,n2098,n81);
nand (n2177,n2178,n2182);
or (n2178,n236,n2179);
nor (n2179,n2180,n2181);
and (n2180,n185,n240);
and (n2181,n241,n187);
or (n2182,n254,n2104);
nand (n2183,n2184,n2188);
or (n2184,n111,n2185);
nor (n2185,n2186,n2187);
and (n2186,n125,n45);
and (n2187,n121,n47);
or (n2188,n112,n2114);
and (n2189,n2171,n2177);
or (n2190,n2191,n2211);
and (n2191,n2192,n2205);
xor (n2192,n2193,n2199);
nand (n2193,n2194,n2195);
or (n2194,n312,n2121);
nand (n2195,n297,n2196);
nand (n2196,n2197,n2198);
or (n2197,n41,n291);
or (n2198,n40,n289);
nand (n2199,n2200,n2204);
or (n2200,n28,n2201);
nor (n2201,n2202,n2203);
and (n2202,n36,n719);
and (n2203,n34,n721);
or (n2204,n37,n2128);
nand (n2205,n2206,n2210);
or (n2206,n1199,n2207);
nor (n2207,n2208,n2209);
and (n2208,n907,n195);
and (n2209,n908,n197);
or (n2210,n2044,n1192);
and (n2211,n2193,n2199);
or (n2212,n2213,n2233);
and (n2213,n2214,n2227);
xor (n2214,n2215,n2221);
nand (n2215,n2216,n2220);
or (n2216,n480,n2217);
nor (n2217,n2218,n2219);
and (n2218,n142,n69);
and (n2219,n143,n71);
or (n2220,n481,n2050);
nand (n2221,n2222,n2226);
or (n2222,n56,n2223);
nor (n2223,n2224,n2225);
and (n2224,n64,n1175);
and (n2225,n65,n1177);
or (n2226,n57,n2056);
nand (n2227,n2228,n2232);
or (n2228,n218,n2229);
nor (n2229,n2230,n2231);
and (n2230,n211,n1141);
and (n2231,n209,n1143);
or (n2232,n212,n2022);
and (n2233,n2215,n2221);
and (n2234,n2168,n2190);
or (n2235,n2236,n2264);
and (n2236,n2237,n2247);
xor (n2237,n2238,n2244);
nand (n2238,n2239,n2243);
or (n2239,n137,n2240);
nor (n2240,n2241,n2242);
and (n2241,n84,n226);
and (n2242,n85,n228);
or (n2243,n155,n1991);
nor (n2244,n2072,n2245);
and (n2245,n2246,n2080);
not (n2246,n2073);
or (n2247,n2248,n2263);
and (n2248,n2249,n2257);
xor (n2249,n2250,n2251);
nor (n2250,n358,n1189);
nand (n2251,n2252,n2256);
or (n2252,n1331,n2253);
nor (n2253,n2254,n2255);
and (n2254,n620,n97);
and (n2255,n621,n99);
or (n2256,n1469,n2075);
nand (n2257,n2258,n2262);
or (n2258,n509,n2259);
nor (n2259,n2260,n2261);
and (n2260,n508,n308);
and (n2261,n115,n310);
or (n2262,n639,n2091);
and (n2263,n2250,n2251);
and (n2264,n2238,n2244);
and (n2265,n2164,n2165);
or (n2266,n2267,n2278);
and (n2267,n2268,n2271);
xor (n2268,n2269,n2270);
xor (n2269,n2071,n2109);
xor (n2270,n2016,n2061);
or (n2271,n2272,n2277);
and (n2272,n2273,n2276);
xor (n2273,n2274,n2275);
xor (n2274,n2019,n2032);
xor (n2275,n2088,n2102);
xor (n2276,n2041,n2054);
and (n2277,n2274,n2275);
and (n2278,n2269,n2270);
and (n2279,n2160,n2161);
and (n2280,n2155,n2156);
and (n2281,n2150,n2151);
xor (n2282,n1858,n2144);
nand (n2283,n1119,n1856);
not (n2284,n2285);
nor (n2285,n2286,n2410);
nor (n2286,n2287,n2401);
xor (n2287,n2288,n2390);
xor (n2288,n2289,n2322);
or (n2289,n2290,n2321);
and (n2290,n2291,n2298);
xor (n2291,n2292,n2295);
or (n2292,n2293,n2294);
and (n2293,n1628,n1650);
and (n2294,n1629,n1647);
or (n2295,n2296,n2297);
and (n2296,n1476,n1512);
and (n2297,n1477,n1480);
xor (n2298,n2299,n2318);
xor (n2299,n2300,n2309);
xor (n2300,n2301,n2306);
xor (n2301,n2302,n2303);
not (n2302,n1643);
or (n2303,n2304,n2305);
and (n2304,n1565,n1573);
and (n2305,n1566,n1570);
or (n2306,n2307,n2308);
and (n2307,n1605,n1612);
and (n2308,n1606,n1609);
xor (n2309,n2310,n2317);
xor (n2310,n2311,n2314);
or (n2311,n2312,n2313);
and (n2312,n1616,n1624);
and (n2313,n1617,n1620);
or (n2314,n2315,n2316);
and (n2315,n1590,n1598);
and (n2316,n1591,n1594);
xor (n2317,n935,n950);
or (n2318,n2319,n2320);
and (n2319,n1513,n1564);
and (n2320,n1514,n1542);
and (n2321,n2292,n2295);
xor (n2322,n2323,n2371);
xor (n2323,n2324,n2362);
xor (n2324,n2325,n2351);
xor (n2325,n2326,n2344);
or (n2326,n2327,n2343);
and (n2327,n2328,n2342);
xor (n2328,n2329,n2341);
xor (n2329,n2330,n2338);
xor (n2330,n2331,n2335);
nand (n2331,n2332,n2333);
or (n2332,n1601,n80);
nand (n2333,n2334,n82);
not (n2334,n791);
nand (n2335,n2336,n2337);
or (n2336,n266,n1634);
or (n2337,n267,n822);
nand (n2338,n2339,n2340);
or (n2339,n163,n1640);
or (n2340,n165,n835);
xor (n2341,n901,n926);
xor (n2342,n873,n887);
and (n2343,n2329,n2341);
xor (n2344,n2345,n2350);
xor (n2345,n2346,n2349);
or (n2346,n2347,n2348);
and (n2347,n2330,n2338);
and (n2348,n2331,n2335);
xor (n2349,n819,n833);
xor (n2350,n735,n750);
or (n2351,n2352,n2361);
and (n2352,n2353,n2358);
xor (n2353,n2354,n2355);
xor (n2354,n959,n972);
or (n2355,n2356,n2357);
and (n2356,n1630,n1643);
and (n2357,n1631,n1637);
or (n2358,n2359,n2360);
and (n2359,n1481,n1485);
and (n2360,n1473,n1482);
and (n2361,n2354,n2355);
or (n2362,n2363,n2370);
and (n2363,n2364,n2369);
xor (n2364,n2365,n2368);
or (n2365,n2366,n2367);
and (n2366,n1588,n1615);
and (n2367,n1589,n1604);
xor (n2368,n2328,n2342);
xor (n2369,n2353,n2358);
and (n2370,n2365,n2368);
xor (n2371,n2372,n2381);
xor (n2372,n2373,n2378);
xor (n2373,n2374,n2377);
xor (n2374,n2375,n2376);
xor (n2375,n782,n795);
xor (n2376,n759,n772);
xor (n2377,n863,n871);
or (n2378,n2379,n2380);
and (n2379,n2299,n2318);
and (n2380,n2300,n2309);
xor (n2381,n2382,n2387);
xor (n2382,n2383,n2386);
or (n2383,n2384,n2385);
and (n2384,n2301,n2306);
and (n2385,n2302,n2303);
xor (n2386,n898,n957);
or (n2387,n2388,n2389);
and (n2388,n2310,n2317);
and (n2389,n2311,n2314);
or (n2390,n2391,n2400);
and (n2391,n2392,n2397);
xor (n2392,n2393,n2394);
xor (n2393,n2364,n2369);
or (n2394,n2395,n2396);
and (n2395,n1579,n1627);
and (n2396,n1580,n1587);
or (n2397,n2398,n2399);
and (n2398,n1122,n1475);
and (n2399,n1123,n1307);
and (n2400,n2393,n2394);
or (n2401,n2402,n2409);
and (n2402,n2403,n2406);
xor (n2403,n2404,n2405);
xor (n2404,n2291,n2298);
xor (n2405,n2392,n2397);
or (n2406,n2407,n2408);
and (n2407,n1577,n1759);
and (n2408,n1578,n1673);
and (n2409,n2404,n2405);
nor (n2410,n2411,n2414);
or (n2411,n2412,n2413);
and (n2412,n1120,n1849);
and (n2413,n1121,n1576);
xor (n2414,n2403,n2406);
nor (n2415,n2416,n2420);
and (n2416,n2417,n2418);
not (n2417,n2286);
not (n2418,n2419);
nand (n2419,n2411,n2414);
and (n2420,n2287,n2401);
nor (n2421,n2422,n2487);
nand (n2422,n2423,n2476);
nor (n2423,n2424,n2457);
nor (n2424,n2425,n2454);
xor (n2425,n2426,n2451);
xor (n2426,n2427,n2430);
or (n2427,n2428,n2429);
and (n2428,n2372,n2381);
and (n2429,n2373,n2378);
xor (n2430,n2431,n2442);
xor (n2431,n2432,n2435);
or (n2432,n2433,n2434);
and (n2433,n2325,n2351);
and (n2434,n2326,n2344);
xor (n2435,n2436,n2441);
xor (n2436,n2437,n2440);
or (n2437,n2438,n2439);
and (n2438,n2345,n2350);
and (n2439,n2346,n2349);
xor (n2440,n816,n843);
xor (n2441,n847,n850);
xor (n2442,n2443,n2448);
xor (n2443,n2444,n2447);
or (n2444,n2445,n2446);
and (n2445,n2374,n2377);
and (n2446,n2375,n2376);
xor (n2447,n860,n980);
or (n2448,n2449,n2450);
and (n2449,n2382,n2387);
and (n2450,n2383,n2386);
or (n2451,n2452,n2453);
and (n2452,n2323,n2371);
and (n2453,n2324,n2362);
or (n2454,n2455,n2456);
and (n2455,n2288,n2390);
and (n2456,n2289,n2322);
nor (n2457,n2458,n2473);
xor (n2458,n2459,n2470);
xor (n2459,n2460,n2461);
xor (n2460,n856,n982);
xor (n2461,n2462,n2467);
xor (n2462,n2463,n2464);
xor (n2463,n812,n845);
or (n2464,n2465,n2466);
and (n2465,n2436,n2441);
and (n2466,n2437,n2440);
or (n2467,n2468,n2469);
and (n2468,n2443,n2448);
and (n2469,n2444,n2447);
or (n2470,n2471,n2472);
and (n2471,n2431,n2442);
and (n2472,n2432,n2435);
or (n2473,n2474,n2475);
and (n2474,n2426,n2451);
and (n2475,n2427,n2430);
or (n2476,n2477,n2484);
xor (n2477,n2478,n2481);
xor (n2478,n2479,n2480);
xor (n2479,n701,n805);
xor (n2480,n809,n854);
or (n2481,n2482,n2483);
and (n2482,n2462,n2467);
and (n2483,n2463,n2464);
or (n2484,n2485,n2486);
and (n2485,n2459,n2470);
and (n2486,n2460,n2461);
nor (n2487,n2488,n2491);
or (n2488,n2489,n2490);
and (n2489,n2478,n2481);
and (n2490,n2479,n2480);
xor (n2491,n18,n807);
nand (n2492,n2493,n2502);
nand (n2493,n2494,n2501);
or (n2494,n2495,n2496);
not (n2495,n2476);
not (n2496,n2497);
nand (n2497,n2498,n2500);
or (n2498,n2457,n2499);
nand (n2499,n2425,n2454);
nand (n2500,n2458,n2473);
nand (n2501,n2477,n2484);
not (n2502,n2487);
nand (n2503,n2488,n2491);
nand (n2504,n2505,n4645);
nand (n2505,n2506,n4622,n4635);
nand (n2506,n2507,n2693,n4401,n4605);
nor (n2507,n2508,n2523);
nor (n2508,n2509,n2510);
xor (n2509,n2149,n2152);
or (n2510,n2511,n2522);
and (n2511,n2512,n2515);
xor (n2512,n2513,n2514);
xor (n2513,n2008,n2065);
xor (n2514,n2154,n2157);
or (n2515,n2516,n2521);
and (n2516,n2517,n2520);
xor (n2517,n2518,n2519);
xor (n2518,n2067,n2134);
xor (n2519,n2012,n2063);
xor (n2520,n2159,n2266);
and (n2521,n2518,n2519);
and (n2522,n2513,n2514);
nor (n2523,n2524,n2525);
xor (n2524,n2512,n2515);
or (n2525,n2526,n2692);
and (n2526,n2527,n2691);
xor (n2527,n2528,n2672);
or (n2528,n2529,n2671);
and (n2529,n2530,n2566);
xor (n2530,n2531,n2532);
xor (n2531,n2136,n2139);
or (n2532,n2533,n2565);
and (n2533,n2534,n2564);
xor (n2534,n2535,n2536);
xor (n2535,n2111,n2126);
or (n2536,n2537,n2563);
and (n2537,n2538,n2551);
xor (n2538,n2539,n2545);
nand (n2539,n2540,n2544);
or (n2540,n625,n2541);
nor (n2541,n2542,n2543);
and (n2542,n514,n250);
and (n2543,n515,n252);
or (n2544,n617,n2028);
nand (n2545,n2546,n2550);
or (n2546,n137,n2547);
nor (n2547,n2548,n2549);
and (n2548,n84,n351);
and (n2549,n85,n353);
or (n2550,n155,n2240);
and (n2551,n2552,n2557);
nor (n2552,n2553,n211);
nor (n2553,n2554,n2556);
and (n2554,n2555,n64);
nand (n2555,n1187,n215);
and (n2556,n1189,n222);
nand (n2557,n2558,n2562);
or (n2558,n1331,n2559);
nor (n2559,n2560,n2561);
and (n2560,n620,n257);
and (n2561,n621,n259);
or (n2562,n1469,n2253);
and (n2563,n2539,n2545);
xor (n2564,n2237,n2247);
and (n2565,n2535,n2536);
or (n2566,n2567,n2670);
and (n2567,n2568,n2669);
xor (n2568,n2569,n2641);
or (n2569,n2570,n2640);
and (n2570,n2571,n2618);
xor (n2571,n2572,n2595);
or (n2572,n2573,n2594);
and (n2573,n2574,n2588);
xor (n2574,n2575,n2582);
nand (n2575,n2576,n2580);
or (n2576,n2577,n509);
nor (n2577,n2578,n2579);
and (n2578,n508,n51);
and (n2579,n115,n53);
nand (n2580,n2581,n511);
not (n2581,n2259);
nand (n2582,n2583,n2587);
or (n2583,n80,n2584);
nor (n2584,n2585,n2586);
and (n2585,n94,n281);
and (n2586,n92,n283);
or (n2587,n81,n2173);
nand (n2588,n2589,n2593);
or (n2589,n236,n2590);
nor (n2590,n2591,n2592);
and (n2591,n240,n179);
and (n2592,n241,n181);
or (n2593,n254,n2179);
and (n2594,n2575,n2582);
or (n2595,n2596,n2617);
and (n2596,n2597,n2611);
xor (n2597,n2598,n2604);
nand (n2598,n2599,n2603);
or (n2599,n111,n2600);
nor (n2600,n2601,n2602);
and (n2601,n125,n75);
and (n2602,n121,n77);
or (n2603,n112,n2185);
nand (n2604,n2605,n2609);
or (n2605,n296,n2606);
nor (n2606,n2607,n2608);
and (n2607,n40,n545);
and (n2608,n41,n547);
or (n2609,n312,n2610);
not (n2610,n2196);
nand (n2611,n2612,n2616);
or (n2612,n28,n2613);
nor (n2613,n2614,n2615);
and (n2614,n36,n837);
and (n2615,n34,n839);
or (n2616,n37,n2201);
and (n2617,n2598,n2604);
or (n2618,n2619,n2639);
and (n2619,n2620,n2633);
xor (n2620,n2621,n2627);
nand (n2621,n2622,n2626);
or (n2622,n1199,n2623);
nor (n2623,n2624,n2625);
and (n2624,n907,n103);
and (n2625,n908,n105);
or (n2626,n2207,n1192);
nand (n2627,n2628,n2632);
or (n2628,n480,n2629);
nor (n2629,n2630,n2631);
and (n2630,n142,n226);
and (n2631,n143,n228);
or (n2632,n481,n2217);
nand (n2633,n2634,n2635);
or (n2634,n2223,n57);
or (n2635,n56,n2636);
nor (n2636,n2637,n2638);
and (n2637,n1147,n64);
and (n2638,n65,n1149);
and (n2639,n2621,n2627);
and (n2640,n2572,n2595);
or (n2641,n2642,n2668);
and (n2642,n2643,n2667);
xor (n2643,n2644,n2666);
or (n2644,n2645,n2665);
and (n2645,n2646,n2659);
xor (n2646,n2647,n2653);
nand (n2647,n2648,n2652);
or (n2648,n218,n2649);
nor (n2649,n2650,n2651);
and (n2650,n1189,n209);
and (n2651,n1187,n211);
or (n2652,n2229,n212);
nand (n2653,n2654,n2658);
or (n2654,n625,n2655);
nor (n2655,n2656,n2657);
and (n2656,n514,n315);
and (n2657,n515,n317);
or (n2658,n617,n2541);
nand (n2659,n2660,n2664);
or (n2660,n137,n2661);
nor (n2661,n2662,n2663);
and (n2662,n84,n345);
and (n2663,n85,n347);
or (n2664,n155,n2547);
and (n2665,n2647,n2653);
xor (n2666,n2249,n2257);
xor (n2667,n2192,n2205);
and (n2668,n2644,n2666);
xor (n2669,n2167,n2212);
and (n2670,n2569,n2641);
and (n2671,n2531,n2532);
or (n2672,n2673,n2690);
and (n2673,n2674,n2677);
xor (n2674,n2675,n2676);
xor (n2675,n2163,n2235);
xor (n2676,n2268,n2271);
or (n2677,n2678,n2689);
and (n2678,n2679,n2688);
xor (n2679,n2680,n2687);
or (n2680,n2681,n2686);
and (n2681,n2682,n2685);
xor (n2682,n2683,n2684);
xor (n2683,n2170,n2183);
xor (n2684,n2214,n2227);
xor (n2685,n2538,n2551);
and (n2686,n2683,n2684);
xor (n2687,n2273,n2276);
xor (n2688,n2534,n2564);
and (n2689,n2680,n2687);
and (n2690,n2675,n2676);
xor (n2691,n2517,n2520);
and (n2692,n2528,n2672);
nand (n2693,n2694,n3882);
nor (n2694,n2695,n3868);
and (n2695,n2696,n3282,n3602);
nor (n2696,n2697,n3197);
nor (n2697,n2698,n3085);
xor (n2698,n2699,n3078);
xor (n2699,n2700,n2871);
or (n2700,n2701,n2870);
and (n2701,n2702,n2795);
xor (n2702,n2703,n2738);
xor (n2703,n2704,n2723);
xor (n2704,n2705,n2714);
nand (n2705,n2706,n2710);
or (n2706,n480,n2707);
nor (n2707,n2708,n2709);
and (n2708,n142,n185);
and (n2709,n143,n187);
or (n2710,n481,n2711);
nor (n2711,n2712,n2713);
and (n2712,n142,n281);
and (n2713,n143,n283);
nand (n2714,n2715,n2719);
or (n2715,n137,n2716);
nor (n2716,n2717,n2718);
and (n2717,n289,n84);
and (n2718,n85,n291);
or (n2719,n155,n2720);
nor (n2720,n2721,n2722);
and (n2721,n84,n179);
and (n2722,n85,n181);
and (n2723,n2724,n2729);
nor (n2724,n2725,n40);
nor (n2725,n2726,n2728);
and (n2726,n2727,n240);
nand (n2727,n1187,n300);
and (n2728,n1189,n305);
nand (n2729,n2730,n2734);
or (n2730,n1199,n2731);
nor (n2731,n2732,n2733);
and (n2732,n907,n51);
and (n2733,n908,n53);
or (n2734,n2735,n1192);
nor (n2735,n2736,n2737);
and (n2736,n907,n308);
and (n2737,n908,n310);
or (n2738,n2739,n2794);
and (n2739,n2740,n2763);
xor (n2740,n2741,n2742);
xor (n2741,n2724,n2729);
or (n2742,n2743,n2762);
and (n2743,n2744,n2752);
xor (n2744,n2745,n2746);
and (n2745,n298,n1187);
nand (n2746,n2747,n2751);
or (n2747,n1199,n2748);
nor (n2748,n2749,n2750);
and (n2749,n907,n45);
and (n2750,n908,n47);
or (n2751,n2731,n1192);
nand (n2752,n2753,n2757);
or (n2753,n509,n2754);
nor (n2754,n2755,n2756);
and (n2755,n508,n372);
and (n2756,n115,n374);
or (n2757,n639,n2758);
not (n2758,n2759);
nor (n2759,n2760,n2761);
and (n2760,n345,n115);
and (n2761,n347,n508);
and (n2762,n2745,n2746);
or (n2763,n2764,n2793);
and (n2764,n2765,n2784);
xor (n2765,n2766,n2775);
nand (n2766,n2767,n2771);
or (n2767,n80,n2768);
nor (n2768,n2769,n2770);
and (n2769,n94,n1175);
and (n2770,n92,n1177);
or (n2771,n81,n2772);
nor (n2772,n2773,n2774);
and (n2773,n837,n94);
and (n2774,n839,n92);
nand (n2775,n2776,n2780);
or (n2776,n236,n2777);
nor (n2777,n2778,n2779);
and (n2778,n240,n1141);
and (n2779,n241,n1143);
or (n2780,n254,n2781);
nor (n2781,n2782,n2783);
and (n2782,n240,n1147);
and (n2783,n241,n1149);
nand (n2784,n2785,n2789);
or (n2785,n1331,n2786);
nor (n2786,n2787,n2788);
and (n2787,n620,n69);
and (n2788,n621,n71);
or (n2789,n1469,n2790);
nor (n2790,n2791,n2792);
and (n2791,n75,n620);
and (n2792,n77,n621);
and (n2793,n2766,n2775);
and (n2794,n2741,n2742);
or (n2795,n2796,n2869);
and (n2796,n2797,n2849);
xor (n2797,n2798,n2830);
or (n2798,n2799,n2829);
and (n2799,n2800,n2820);
xor (n2800,n2801,n2811);
nand (n2801,n2802,n2807);
or (n2802,n2803,n111);
not (n2803,n2804);
nand (n2804,n2805,n2806);
or (n2805,n121,n187);
or (n2806,n125,n185);
nand (n2807,n113,n2808);
nor (n2808,n2809,n2810);
and (n2809,n283,n125);
and (n2810,n281,n121);
nand (n2811,n2812,n2816);
or (n2812,n2813,n625);
nor (n2813,n2814,n2815);
and (n2814,n514,n351);
and (n2815,n515,n353);
nand (n2816,n616,n2817);
nand (n2817,n2818,n2819);
or (n2818,n515,n228);
or (n2819,n514,n226);
nand (n2820,n2821,n2825);
or (n2821,n480,n2822);
nor (n2822,n2823,n2824);
and (n2823,n142,n289);
and (n2824,n143,n291);
or (n2825,n481,n2826);
nor (n2826,n2827,n2828);
and (n2827,n179,n142);
and (n2828,n143,n181);
and (n2829,n2801,n2811);
xor (n2830,n2831,n2843);
xor (n2831,n2832,n2840);
nand (n2832,n2833,n2835);
or (n2833,n2834,n625);
not (n2834,n2817);
nand (n2835,n2836,n616);
not (n2836,n2837);
nor (n2837,n2838,n2839);
and (n2838,n71,n515);
and (n2839,n69,n514);
nand (n2840,n2841,n2842);
or (n2841,n480,n2826);
or (n2842,n2707,n481);
nand (n2843,n2844,n2848);
or (n2844,n137,n2845);
nor (n2845,n2846,n2847);
and (n2846,n545,n84);
and (n2847,n85,n547);
or (n2848,n155,n2716);
xor (n2849,n2850,n2863);
xor (n2850,n2851,n2857);
nand (n2851,n2852,n2853);
or (n2852,n2758,n509);
nand (n2853,n2854,n511);
nor (n2854,n2855,n2856);
and (n2855,n353,n508);
and (n2856,n351,n115);
nand (n2857,n2858,n2859);
or (n2858,n2772,n80);
nand (n2859,n2860,n82);
nor (n2860,n2861,n2862);
and (n2861,n721,n94);
and (n2862,n719,n92);
nand (n2863,n2864,n2865);
or (n2864,n236,n2781);
or (n2865,n2866,n254);
nor (n2866,n2867,n2868);
and (n2867,n240,n1175);
and (n2868,n241,n1177);
and (n2869,n2798,n2830);
and (n2870,n2703,n2738);
xor (n2871,n2872,n2996);
xor (n2872,n2873,n2947);
or (n2873,n2874,n2946);
and (n2874,n2875,n2917);
xor (n2875,n2876,n2893);
xor (n2876,n2877,n2885);
xor (n2877,n2878,n2879);
and (n2878,n38,n1187);
nand (n2879,n2880,n2881);
or (n2880,n1199,n2735);
or (n2881,n2882,n1192);
nor (n2882,n2883,n2884);
and (n2883,n317,n908);
and (n2884,n315,n907);
nand (n2885,n2886,n2888);
or (n2886,n509,n2887);
not (n2887,n2854);
or (n2888,n639,n2889);
not (n2889,n2890);
nor (n2890,n2891,n2892);
and (n2891,n226,n115);
and (n2892,n228,n508);
xor (n2893,n2894,n2908);
xor (n2894,n2895,n2902);
nand (n2895,n2896,n2898);
or (n2896,n2897,n80);
not (n2897,n2860);
or (n2898,n81,n2899);
nor (n2899,n2900,n2901);
and (n2900,n547,n92);
and (n2901,n545,n94);
nand (n2902,n2903,n2904);
or (n2903,n236,n2866);
or (n2904,n254,n2905);
nor (n2905,n2906,n2907);
and (n2906,n240,n837);
and (n2907,n241,n839);
nand (n2908,n2909,n2913);
or (n2909,n1331,n2910);
nor (n2910,n2911,n2912);
and (n2911,n620,n45);
and (n2912,n621,n47);
or (n2913,n1469,n2914);
nor (n2914,n2915,n2916);
and (n2915,n620,n51);
and (n2916,n621,n53);
xor (n2917,n2918,n2940);
xor (n2918,n2919,n2929);
nand (n2919,n2920,n2925);
or (n2920,n2921,n296);
not (n2921,n2922);
nand (n2922,n2923,n2924);
or (n2923,n41,n1143);
or (n2924,n40,n1141);
or (n2925,n312,n2926);
nor (n2926,n2927,n2928);
and (n2927,n1149,n41);
and (n2928,n1147,n40);
nand (n2929,n2930,n2935);
or (n2930,n2931,n112);
not (n2931,n2932);
nand (n2932,n2933,n2934);
or (n2933,n121,n347);
or (n2934,n125,n345);
nand (n2935,n2936,n1041);
not (n2936,n2937);
nor (n2937,n2938,n2939);
and (n2938,n125,n372);
and (n2939,n121,n374);
nand (n2940,n2941,n2942);
or (n2941,n625,n2837);
or (n2942,n617,n2943);
nor (n2943,n2944,n2945);
and (n2944,n514,n75);
and (n2945,n515,n77);
and (n2946,n2876,n2893);
xor (n2947,n2948,n2993);
xor (n2948,n2949,n2969);
xor (n2949,n2950,n2963);
xor (n2950,n2951,n2957);
nand (n2951,n2952,n2953);
or (n2952,n2889,n509);
nand (n2953,n511,n2954);
nor (n2954,n2955,n2956);
and (n2955,n69,n115);
and (n2956,n71,n508);
nand (n2957,n2958,n2959);
or (n2958,n2899,n80);
nand (n2959,n82,n2960);
nand (n2960,n2961,n2962);
or (n2961,n92,n291);
or (n2962,n94,n289);
nand (n2963,n2964,n2965);
or (n2964,n236,n2905);
or (n2965,n254,n2966);
nor (n2966,n2967,n2968);
and (n2967,n240,n719);
and (n2968,n241,n721);
xor (n2969,n2970,n2984);
xor (n2970,n2971,n2978);
nand (n2971,n2972,n2973);
or (n2972,n2931,n111);
nand (n2973,n2974,n113);
not (n2974,n2975);
nor (n2975,n2976,n2977);
and (n2976,n353,n121);
and (n2977,n351,n125);
nand (n2978,n2979,n2980);
or (n2979,n296,n2926);
nand (n2980,n298,n2981);
nor (n2981,n2982,n2983);
and (n2982,n1177,n40);
and (n2983,n1175,n41);
nand (n2984,n2985,n2989);
or (n2985,n28,n2986);
nor (n2986,n2987,n2988);
and (n2987,n1189,n34);
and (n2988,n36,n1187);
or (n2989,n37,n2990);
nor (n2990,n2991,n2992);
and (n2991,n36,n1141);
and (n2992,n34,n1143);
or (n2993,n2994,n2995);
and (n2994,n2704,n2723);
and (n2995,n2705,n2714);
xor (n2996,n2997,n3050);
xor (n2997,n2998,n3026);
or (n2998,n2999,n3025);
and (n2999,n3000,n3007);
xor (n3000,n3001,n3004);
or (n3001,n3002,n3003);
and (n3002,n2850,n2863);
and (n3003,n2851,n2857);
or (n3004,n3005,n3006);
and (n3005,n2831,n2843);
and (n3006,n2832,n2840);
or (n3007,n3008,n3024);
and (n3008,n3009,n3020);
xor (n3009,n3010,n3014);
nand (n3010,n3011,n3012);
or (n3011,n2790,n1331);
nand (n3012,n3013,n904);
not (n3013,n2910);
nand (n3014,n3015,n3016);
or (n3015,n2921,n312);
or (n3016,n296,n3017);
nor (n3017,n3018,n3019);
and (n3018,n41,n1189);
and (n3019,n40,n1187);
nand (n3020,n3021,n3023);
or (n3021,n111,n3022);
not (n3022,n2808);
or (n3023,n112,n2937);
and (n3024,n3010,n3014);
and (n3025,n3001,n3004);
xor (n3026,n3027,n3047);
xor (n3027,n3028,n3034);
nand (n3028,n3029,n3030);
or (n3029,n137,n2720);
or (n3030,n155,n3031);
nor (n3031,n3032,n3033);
and (n3032,n84,n185);
and (n3033,n85,n187);
xor (n3034,n3035,n3041);
and (n3035,n3036,n34);
nand (n3036,n3037,n3038);
or (n3037,n1187,n33);
nand (n3038,n3039,n40);
not (n3039,n3040);
and (n3040,n1187,n33);
nand (n3041,n3042,n3043);
or (n3042,n2914,n1331);
nand (n3043,n904,n3044);
nor (n3044,n3045,n3046);
and (n3045,n308,n621);
and (n3046,n310,n620);
or (n3047,n3048,n3049);
and (n3048,n2894,n2908);
and (n3049,n2895,n2902);
xor (n3050,n3051,n3058);
xor (n3051,n3052,n3055);
or (n3052,n3053,n3054);
and (n3053,n2877,n2885);
and (n3054,n2878,n2879);
or (n3055,n3056,n3057);
and (n3056,n2918,n2940);
and (n3057,n2919,n2929);
xor (n3058,n3059,n3072);
xor (n3059,n3060,n3066);
nand (n3060,n3061,n3062);
or (n3061,n1199,n2882);
or (n3062,n3063,n1192);
nor (n3063,n3064,n3065);
and (n3064,n907,n250);
and (n3065,n908,n252);
nand (n3066,n3067,n3068);
or (n3067,n625,n2943);
nand (n3068,n616,n3069);
nor (n3069,n3070,n3071);
and (n3070,n45,n515);
and (n3071,n47,n514);
nand (n3072,n3073,n3074);
or (n3073,n480,n2711);
or (n3074,n481,n3075);
nor (n3075,n3076,n3077);
and (n3076,n142,n372);
and (n3077,n143,n374);
or (n3078,n3079,n3084);
and (n3079,n3080,n3083);
xor (n3080,n3081,n3082);
xor (n3081,n3000,n3007);
xor (n3082,n2875,n2917);
xor (n3083,n2702,n2795);
and (n3084,n3081,n3082);
or (n3085,n3086,n3196);
and (n3086,n3087,n3195);
xor (n3087,n3088,n3139);
or (n3088,n3089,n3138);
and (n3089,n3090,n3137);
xor (n3090,n3091,n3092);
xor (n3091,n3009,n3020);
or (n3092,n3093,n3136);
and (n3093,n3094,n3113);
xor (n3094,n3095,n3101);
nand (n3095,n3096,n3100);
or (n3096,n137,n3097);
nor (n3097,n3098,n3099);
and (n3098,n84,n719);
and (n3099,n85,n721);
or (n3100,n155,n2845);
and (n3101,n3102,n3107);
nor (n3102,n3103,n240);
nor (n3103,n3104,n3106);
and (n3104,n3105,n94);
nand (n3105,n1187,n242);
and (n3106,n1189,n244);
nand (n3107,n3108,n3112);
or (n3108,n1199,n3109);
nor (n3109,n3110,n3111);
and (n3110,n907,n75);
and (n3111,n908,n77);
or (n3112,n2748,n1192);
or (n3113,n3114,n3135);
and (n3114,n3115,n3129);
xor (n3115,n3116,n3123);
nand (n3116,n3117,n3121);
or (n3117,n3118,n509);
nor (n3118,n3119,n3120);
and (n3119,n508,n281);
and (n3120,n115,n283);
nand (n3121,n3122,n511);
not (n3122,n2754);
nand (n3123,n3124,n3128);
or (n3124,n80,n3125);
nor (n3125,n3126,n3127);
and (n3126,n94,n1147);
and (n3127,n92,n1149);
or (n3128,n81,n2768);
nand (n3129,n3130,n3134);
or (n3130,n236,n3131);
nor (n3131,n3132,n3133);
and (n3132,n1189,n241);
and (n3133,n240,n1187);
or (n3134,n254,n2777);
and (n3135,n3116,n3123);
and (n3136,n3095,n3101);
xor (n3137,n2740,n2763);
and (n3138,n3091,n3092);
or (n3139,n3140,n3194);
and (n3140,n3141,n3171);
xor (n3141,n3142,n3170);
or (n3142,n3143,n3169);
and (n3143,n3144,n3168);
xor (n3144,n3145,n3167);
or (n3145,n3146,n3166);
and (n3146,n3147,n3160);
xor (n3147,n3148,n3154);
nand (n3148,n3149,n3153);
or (n3149,n1331,n3150);
nor (n3150,n3151,n3152);
and (n3151,n620,n226);
and (n3152,n621,n228);
or (n3153,n1469,n2786);
nand (n3154,n3155,n3159);
or (n3155,n111,n3156);
nor (n3156,n3157,n3158);
and (n3157,n125,n179);
and (n3158,n121,n181);
or (n3159,n112,n2803);
nand (n3160,n3161,n3165);
or (n3161,n625,n3162);
nor (n3162,n3163,n3164);
and (n3163,n514,n345);
and (n3164,n515,n347);
or (n3165,n617,n2813);
and (n3166,n3148,n3154);
xor (n3167,n2800,n2820);
xor (n3168,n2744,n2752);
and (n3169,n3145,n3167);
xor (n3170,n2797,n2849);
or (n3171,n3172,n3193);
and (n3172,n3173,n3192);
xor (n3173,n3174,n3175);
xor (n3174,n2765,n2784);
or (n3175,n3176,n3191);
and (n3176,n3177,n3190);
xor (n3177,n3178,n3184);
nand (n3178,n3179,n3183);
or (n3179,n480,n3180);
nor (n3180,n3181,n3182);
and (n3181,n142,n545);
and (n3182,n143,n547);
or (n3183,n481,n2822);
nand (n3184,n3185,n3189);
or (n3185,n137,n3186);
nor (n3186,n3187,n3188);
and (n3187,n84,n837);
and (n3188,n85,n839);
or (n3189,n155,n3097);
xor (n3190,n3102,n3107);
and (n3191,n3178,n3184);
xor (n3192,n3094,n3113);
and (n3193,n3174,n3175);
and (n3194,n3142,n3170);
xor (n3195,n3080,n3083);
and (n3196,n3088,n3139);
nor (n3197,n3198,n3199);
xor (n3198,n3087,n3195);
or (n3199,n3200,n3281);
and (n3200,n3201,n3280);
xor (n3201,n3202,n3203);
xor (n3202,n3090,n3137);
or (n3203,n3204,n3279);
and (n3204,n3205,n3278);
xor (n3205,n3206,n3271);
or (n3206,n3207,n3270);
and (n3207,n3208,n3248);
xor (n3208,n3209,n3226);
or (n3209,n3210,n3225);
and (n3210,n3211,n3219);
xor (n3211,n3212,n3213);
and (n3212,n245,n1187);
nand (n3213,n3214,n3218);
or (n3214,n1199,n3215);
nor (n3215,n3216,n3217);
and (n3216,n907,n69);
and (n3217,n908,n71);
or (n3218,n3109,n1192);
nand (n3219,n3220,n3224);
or (n3220,n1331,n3221);
nor (n3221,n3222,n3223);
and (n3222,n620,n351);
and (n3223,n621,n353);
or (n3224,n1469,n3150);
and (n3225,n3212,n3213);
or (n3226,n3227,n3247);
and (n3227,n3228,n3241);
xor (n3228,n3229,n3235);
nand (n3229,n3230,n3234);
or (n3230,n625,n3231);
nor (n3231,n3232,n3233);
and (n3232,n514,n372);
and (n3233,n515,n374);
or (n3234,n617,n3162);
nand (n3235,n3236,n3240);
or (n3236,n480,n3237);
nor (n3237,n3238,n3239);
and (n3238,n142,n719);
and (n3239,n143,n721);
or (n3240,n481,n3180);
nand (n3241,n3242,n3246);
or (n3242,n137,n3243);
nor (n3243,n3244,n3245);
and (n3244,n84,n1175);
and (n3245,n85,n1177);
or (n3246,n155,n3186);
and (n3247,n3229,n3235);
or (n3248,n3249,n3269);
and (n3249,n3250,n3263);
xor (n3250,n3251,n3257);
nand (n3251,n3252,n3256);
or (n3252,n80,n3253);
nor (n3253,n3254,n3255);
and (n3254,n94,n1141);
and (n3255,n92,n1143);
or (n3256,n81,n3125);
nand (n3257,n3258,n3262);
or (n3258,n509,n3259);
nor (n3259,n3260,n3261);
and (n3260,n508,n185);
and (n3261,n115,n187);
or (n3262,n639,n3118);
nand (n3263,n3264,n3268);
or (n3264,n111,n3265);
nor (n3265,n3266,n3267);
and (n3266,n289,n125);
and (n3267,n121,n291);
or (n3268,n112,n3156);
and (n3269,n3251,n3257);
and (n3270,n3209,n3226);
or (n3271,n3272,n3277);
and (n3272,n3273,n3276);
xor (n3273,n3274,n3275);
xor (n3274,n3115,n3129);
xor (n3275,n3147,n3160);
xor (n3276,n3177,n3190);
and (n3277,n3274,n3275);
xor (n3278,n3144,n3168);
and (n3279,n3206,n3271);
xor (n3280,n3141,n3171);
and (n3281,n3202,n3203);
nand (n3282,n3283,n3601);
or (n3283,n3284,n3596);
nor (n3284,n3285,n3595);
and (n3285,n3286,n3583);
not (n3286,n3287);
nand (n3287,n3288,n3580);
or (n3288,n3289,n3560);
not (n3289,n3290);
nand (n3290,n3291,n3502);
xor (n3291,n3292,n3433);
xor (n3292,n3293,n3298);
xor (n3293,n3294,n3297);
xor (n3294,n3295,n3296);
xor (n3295,n3228,n3241);
xor (n3296,n3211,n3219);
xor (n3297,n3250,n3263);
or (n3298,n3299,n3432);
and (n3299,n3300,n3373);
xor (n3300,n3301,n3339);
or (n3301,n3302,n3338);
and (n3302,n3303,n3323);
xor (n3303,n3304,n3313);
nand (n3304,n3305,n3309);
or (n3305,n480,n3306);
nor (n3306,n3307,n3308);
and (n3307,n142,n1175);
and (n3308,n143,n1177);
or (n3309,n481,n3310);
nor (n3310,n3311,n3312);
and (n3311,n142,n837);
and (n3312,n143,n839);
nand (n3313,n3314,n3319);
or (n3314,n3315,n137);
not (n3315,n3316);
nand (n3316,n3317,n3318);
or (n3317,n1143,n85);
or (n3318,n84,n1141);
or (n3319,n155,n3320);
nor (n3320,n3321,n3322);
and (n3321,n84,n1147);
and (n3322,n85,n1149);
and (n3323,n3324,n3329);
nor (n3324,n3325,n84);
nor (n3325,n3326,n3328);
and (n3326,n3327,n142);
nand (n3327,n1187,n141);
and (n3328,n1189,n148);
nand (n3329,n3330,n3334);
or (n3330,n3331,n1199);
nor (n3331,n3332,n3333);
and (n3332,n907,n345);
and (n3333,n908,n347);
or (n3334,n3335,n1192);
nor (n3335,n3336,n3337);
and (n3336,n907,n351);
and (n3337,n908,n353);
and (n3338,n3304,n3313);
xor (n3339,n3340,n3356);
xor (n3340,n3341,n3344);
nand (n3341,n3342,n3343);
or (n3342,n137,n3320);
or (n3343,n155,n3243);
xor (n3344,n3345,n3350);
nor (n3345,n3346,n94);
nor (n3346,n3347,n3349);
and (n3347,n3348,n84);
nand (n3348,n1187,n86);
and (n3349,n1189,n91);
nand (n3350,n3351,n3355);
or (n3351,n1199,n3352);
nor (n3352,n3353,n3354);
and (n3353,n907,n226);
and (n3354,n908,n228);
or (n3355,n3215,n1192);
or (n3356,n3357,n3372);
and (n3357,n3358,n3363);
xor (n3358,n3359,n3360);
nor (n3359,n81,n1189);
nand (n3360,n3361,n3362);
or (n3361,n1199,n3335);
or (n3362,n3352,n1192);
nand (n3363,n3364,n3368);
or (n3364,n1331,n3365);
nor (n3365,n3366,n3367);
and (n3366,n620,n372);
and (n3367,n621,n374);
or (n3368,n1469,n3369);
nor (n3369,n3370,n3371);
and (n3370,n620,n345);
and (n3371,n621,n347);
and (n3372,n3359,n3360);
or (n3373,n3374,n3431);
and (n3374,n3375,n3430);
xor (n3375,n3376,n3405);
or (n3376,n3377,n3404);
and (n3377,n3378,n3395);
xor (n3378,n3379,n3385);
nand (n3379,n3380,n3384);
or (n3380,n1331,n3381);
nor (n3381,n3382,n3383);
and (n3382,n620,n281);
and (n3383,n621,n283);
or (n3384,n1469,n3365);
nand (n3385,n3386,n3390);
or (n3386,n509,n3387);
nor (n3387,n3388,n3389);
and (n3388,n508,n545);
and (n3389,n115,n547);
or (n3390,n639,n3391);
not (n3391,n3392);
nor (n3392,n3393,n3394);
and (n3393,n289,n115);
and (n3394,n291,n508);
nand (n3395,n3396,n3400);
or (n3396,n111,n3397);
nor (n3397,n3398,n3399);
and (n3398,n125,n837);
and (n3399,n121,n839);
or (n3400,n112,n3401);
nor (n3401,n3402,n3403);
and (n3402,n125,n719);
and (n3403,n121,n721);
and (n3404,n3379,n3385);
or (n3405,n3406,n3429);
and (n3406,n3407,n3423);
xor (n3407,n3408,n3417);
nand (n3408,n3409,n3413);
or (n3409,n625,n3410);
nor (n3410,n3411,n3412);
and (n3411,n514,n179);
and (n3412,n515,n181);
or (n3413,n617,n3414);
nor (n3414,n3415,n3416);
and (n3415,n514,n185);
and (n3416,n515,n187);
nand (n3417,n3418,n3422);
or (n3418,n480,n3419);
nor (n3419,n3420,n3421);
and (n3420,n142,n1147);
and (n3421,n143,n1149);
or (n3422,n481,n3306);
nand (n3423,n3424,n3425);
or (n3424,n3315,n155);
or (n3425,n137,n3426);
nor (n3426,n3427,n3428);
and (n3427,n1189,n85);
and (n3428,n1187,n84);
and (n3429,n3408,n3417);
xor (n3430,n3358,n3363);
and (n3431,n3376,n3405);
and (n3432,n3301,n3339);
xor (n3433,n3434,n3482);
xor (n3434,n3435,n3438);
or (n3435,n3436,n3437);
and (n3436,n3340,n3356);
and (n3437,n3341,n3344);
xor (n3438,n3439,n3461);
xor (n3439,n3440,n3441);
and (n3440,n3345,n3350);
or (n3441,n3442,n3460);
and (n3442,n3443,n3454);
xor (n3443,n3444,n3448);
nand (n3444,n3445,n3446);
or (n3445,n3221,n1469);
nand (n3446,n3447,n910);
not (n3447,n3369);
nand (n3448,n3449,n3453);
or (n3449,n80,n3450);
nor (n3450,n3451,n3452);
and (n3451,n92,n1189);
and (n3452,n94,n1187);
or (n3453,n81,n3253);
nand (n3454,n3455,n3459);
or (n3455,n509,n3456);
nor (n3456,n3457,n3458);
and (n3457,n508,n179);
and (n3458,n115,n181);
or (n3459,n639,n3259);
and (n3460,n3444,n3448);
or (n3461,n3462,n3481);
and (n3462,n3463,n3478);
xor (n3463,n3464,n3471);
nand (n3464,n3465,n3469);
or (n3465,n3466,n111);
nor (n3466,n3467,n3468);
and (n3467,n547,n121);
and (n3468,n545,n125);
nand (n3469,n3470,n113);
not (n3470,n3265);
nand (n3471,n3472,n3476);
or (n3472,n3473,n625);
nor (n3473,n3474,n3475);
and (n3474,n514,n281);
and (n3475,n515,n283);
nand (n3476,n3477,n616);
not (n3477,n3231);
nand (n3478,n3479,n3480);
or (n3479,n480,n3310);
or (n3480,n481,n3237);
and (n3481,n3464,n3471);
or (n3482,n3483,n3501);
and (n3483,n3484,n3500);
xor (n3484,n3485,n3499);
or (n3485,n3486,n3498);
and (n3486,n3487,n3495);
xor (n3487,n3488,n3492);
nand (n3488,n3489,n3490);
or (n3489,n3391,n509);
nand (n3490,n3491,n511);
not (n3491,n3456);
nand (n3492,n3493,n3494);
or (n3493,n111,n3401);
or (n3494,n112,n3466);
nand (n3495,n3496,n3497);
or (n3496,n625,n3414);
or (n3497,n617,n3473);
and (n3498,n3488,n3492);
xor (n3499,n3463,n3478);
xor (n3500,n3443,n3454);
and (n3501,n3485,n3499);
or (n3502,n3503,n3559);
and (n3503,n3504,n3558);
xor (n3504,n3505,n3506);
xor (n3505,n3484,n3500);
or (n3506,n3507,n3557);
and (n3507,n3508,n3511);
xor (n3508,n3509,n3510);
xor (n3509,n3487,n3495);
xor (n3510,n3303,n3323);
or (n3511,n3512,n3556);
and (n3512,n3513,n3533);
xor (n3513,n3514,n3515);
xor (n3514,n3324,n3329);
or (n3515,n3516,n3532);
and (n3516,n3517,n3526);
xor (n3517,n3518,n3519);
nor (n3518,n155,n1189);
nand (n3519,n3520,n3525);
or (n3520,n3521,n1331);
not (n3521,n3522);
nand (n3522,n3523,n3524);
or (n3523,n621,n187);
or (n3524,n620,n185);
or (n3525,n1469,n3381);
nand (n3526,n3527,n3531);
or (n3527,n509,n3528);
nor (n3528,n3529,n3530);
and (n3529,n508,n719);
and (n3530,n115,n721);
or (n3531,n639,n3387);
and (n3532,n3518,n3519);
or (n3533,n3534,n3555);
and (n3534,n3535,n3549);
xor (n3535,n3536,n3542);
nand (n3536,n3537,n3541);
or (n3537,n111,n3538);
nor (n3538,n3539,n3540);
and (n3539,n125,n1175);
and (n3540,n121,n1177);
or (n3541,n112,n3397);
nand (n3542,n3543,n3548);
or (n3543,n1199,n3544);
not (n3544,n3545);
nor (n3545,n3546,n3547);
and (n3546,n372,n908);
and (n3547,n374,n907);
or (n3548,n3331,n1192);
nand (n3549,n3550,n3554);
or (n3550,n480,n3551);
nor (n3551,n3552,n3553);
and (n3552,n142,n1141);
and (n3553,n143,n1143);
or (n3554,n481,n3419);
and (n3555,n3536,n3542);
and (n3556,n3514,n3515);
and (n3557,n3509,n3510);
xor (n3558,n3300,n3373);
and (n3559,n3505,n3506);
not (n3560,n3561);
nand (n3561,n3562,n3577);
xor (n3562,n3563,n3568);
xor (n3563,n3564,n3565);
xor (n3564,n3273,n3276);
or (n3565,n3566,n3567);
and (n3566,n3434,n3482);
and (n3567,n3435,n3438);
xor (n3568,n3569,n3574);
xor (n3569,n3570,n3573);
or (n3570,n3571,n3572);
and (n3571,n3439,n3461);
and (n3572,n3440,n3441);
xor (n3573,n3208,n3248);
or (n3574,n3575,n3576);
and (n3575,n3294,n3297);
and (n3576,n3295,n3296);
or (n3577,n3578,n3579);
and (n3578,n3292,n3433);
and (n3579,n3293,n3298);
nand (n3580,n3581,n3582);
not (n3581,n3562);
not (n3582,n3577);
not (n3583,n3584);
nor (n3584,n3585,n3592);
xor (n3585,n3586,n3591);
xor (n3586,n3587,n3588);
xor (n3587,n3173,n3192);
or (n3588,n3589,n3590);
and (n3589,n3569,n3574);
and (n3590,n3570,n3573);
xor (n3591,n3205,n3278);
or (n3592,n3593,n3594);
and (n3593,n3563,n3568);
and (n3594,n3564,n3565);
and (n3595,n3585,n3592);
nor (n3596,n3597,n3598);
xor (n3597,n3201,n3280);
or (n3598,n3599,n3600);
and (n3599,n3586,n3591);
and (n3600,n3587,n3588);
nand (n3601,n3597,n3598);
nor (n3602,n3603,n3729);
nor (n3603,n3604,n3726);
xor (n3604,n3605,n3723);
xor (n3605,n3606,n3623);
xor (n3606,n3607,n3620);
xor (n3607,n3608,n3611);
or (n3608,n3609,n3610);
and (n3609,n3051,n3058);
and (n3610,n3052,n3055);
xor (n3611,n3612,n3617);
xor (n3612,n3613,n3614);
and (n3613,n3035,n3041);
or (n3614,n3615,n3616);
and (n3615,n3059,n3072);
and (n3616,n3060,n3066);
or (n3617,n3618,n3619);
and (n3618,n2970,n2984);
and (n3619,n2971,n2978);
or (n3620,n3621,n3622);
and (n3621,n2948,n2993);
and (n3622,n2949,n2969);
xor (n3623,n3624,n3720);
xor (n3624,n3625,n3673);
xor (n3625,n3626,n3651);
xor (n3626,n3627,n3630);
or (n3627,n3628,n3629);
and (n3628,n2950,n2963);
and (n3629,n2951,n2957);
xor (n3630,n3631,n3645);
xor (n3631,n3632,n3639);
nand (n3632,n3633,n3635);
or (n3633,n3634,n625);
not (n3634,n3069);
nand (n3635,n616,n3636);
nor (n3636,n3637,n3638);
and (n3637,n51,n515);
and (n3638,n53,n514);
nand (n3639,n3640,n3641);
or (n3640,n480,n3075);
or (n3641,n3642,n481);
nor (n3642,n3643,n3644);
and (n3643,n142,n345);
and (n3644,n143,n347);
nand (n3645,n3646,n3647);
or (n3646,n137,n3031);
or (n3647,n155,n3648);
nor (n3648,n3649,n3650);
and (n3649,n84,n281);
and (n3650,n85,n283);
xor (n3651,n3652,n3666);
xor (n3652,n3653,n3660);
nand (n3653,n3654,n3656);
or (n3654,n3655,n80);
not (n3655,n2960);
nand (n3656,n3657,n82);
nor (n3657,n3658,n3659);
and (n3658,n179,n92);
and (n3659,n181,n94);
nand (n3660,n3661,n3662);
or (n3661,n236,n2966);
or (n3662,n254,n3663);
nor (n3663,n3664,n3665);
and (n3664,n240,n545);
and (n3665,n241,n547);
nand (n3666,n3667,n3668);
or (n3667,n111,n2975);
or (n3668,n112,n3669);
not (n3669,n3670);
nand (n3670,n3671,n3672);
or (n3671,n121,n228);
or (n3672,n125,n226);
xor (n3673,n3674,n3717);
xor (n3674,n3675,n3699);
xor (n3675,n3676,n3693);
xor (n3676,n3677,n3684);
nand (n3677,n3678,n3680);
or (n3678,n3679,n296);
not (n3679,n2981);
nand (n3680,n3681,n298);
nor (n3681,n3682,n3683);
and (n3682,n839,n40);
and (n3683,n837,n41);
nand (n3684,n3685,n3690);
or (n3685,n3686,n37);
not (n3686,n3687);
nand (n3687,n3688,n3689);
or (n3688,n34,n1149);
or (n3689,n36,n1147);
nand (n3690,n3691,n3692);
not (n3691,n2990);
not (n3692,n28);
nand (n3693,n3694,n3695);
or (n3694,n1199,n3063);
or (n3695,n3696,n1192);
nor (n3696,n3697,n3698);
and (n3697,n259,n908);
and (n3698,n257,n907);
xor (n3699,n3700,n3710);
xor (n3700,n3701,n3702);
nor (n3701,n57,n1189);
nand (n3702,n3703,n3705);
or (n3703,n3704,n1331);
not (n3704,n3044);
nand (n3705,n3706,n904);
not (n3706,n3707);
nor (n3707,n3708,n3709);
and (n3708,n317,n621);
and (n3709,n315,n620);
nand (n3710,n3711,n3713);
or (n3711,n3712,n509);
not (n3712,n2954);
nand (n3713,n511,n3714);
nand (n3714,n3715,n3716);
or (n3715,n115,n77);
or (n3716,n508,n75);
or (n3717,n3718,n3719);
and (n3718,n3027,n3047);
and (n3719,n3028,n3034);
or (n3720,n3721,n3722);
and (n3721,n2997,n3050);
and (n3722,n2998,n3026);
or (n3723,n3724,n3725);
and (n3724,n2872,n2996);
and (n3725,n2873,n2947);
or (n3726,n3727,n3728);
and (n3727,n2699,n3078);
and (n3728,n2700,n2871);
nor (n3729,n3730,n3733);
or (n3730,n3731,n3732);
and (n3731,n3605,n3723);
and (n3732,n3606,n3623);
xor (n3733,n3734,n3741);
xor (n3734,n3735,n3738);
or (n3735,n3736,n3737);
and (n3736,n3607,n3620);
and (n3737,n3608,n3611);
or (n3738,n3739,n3740);
and (n3739,n3624,n3720);
and (n3740,n3625,n3673);
xor (n3741,n3742,n3801);
xor (n3742,n3743,n3798);
xor (n3743,n3744,n3795);
xor (n3744,n3745,n3768);
xor (n3745,n3746,n3762);
xor (n3746,n3747,n3755);
nand (n3747,n3748,n3750);
or (n3748,n3749,n509);
not (n3749,n3714);
nand (n3750,n3751,n511);
not (n3751,n3752);
nor (n3752,n3753,n3754);
and (n3753,n508,n45);
and (n3754,n115,n47);
nand (n3755,n3756,n3758);
or (n3756,n80,n3757);
not (n3757,n3657);
or (n3758,n81,n3759);
nor (n3759,n3760,n3761);
and (n3760,n94,n185);
and (n3761,n92,n187);
nand (n3762,n3763,n3764);
or (n3763,n236,n3663);
or (n3764,n254,n3765);
nor (n3765,n3766,n3767);
and (n3766,n240,n289);
and (n3767,n241,n291);
xor (n3768,n3769,n3782);
xor (n3769,n3770,n3776);
nand (n3770,n3771,n3772);
or (n3771,n480,n3642);
or (n3772,n481,n3773);
nor (n3773,n3774,n3775);
and (n3774,n142,n351);
and (n3775,n143,n353);
nand (n3776,n3777,n3778);
or (n3777,n137,n3648);
or (n3778,n155,n3779);
nor (n3779,n3780,n3781);
and (n3780,n84,n372);
and (n3781,n85,n374);
xor (n3782,n3783,n3788);
nor (n3783,n3784,n64);
nor (n3784,n3785,n3787);
and (n3785,n3786,n36);
nand (n3786,n1187,n59);
and (n3787,n1189,n61);
nand (n3788,n3789,n3794);
or (n3789,n3790,n1469);
not (n3790,n3791);
nand (n3791,n3792,n3793);
or (n3792,n621,n252);
or (n3793,n620,n250);
or (n3794,n1331,n3707);
or (n3795,n3796,n3797);
and (n3796,n3612,n3617);
and (n3797,n3613,n3614);
or (n3798,n3799,n3800);
and (n3799,n3674,n3717);
and (n3800,n3675,n3699);
xor (n3801,n3802,n3817);
xor (n3802,n3803,n3814);
xor (n3803,n3804,n3811);
xor (n3804,n3805,n3808);
or (n3805,n3806,n3807);
and (n3806,n3676,n3693);
and (n3807,n3677,n3684);
or (n3808,n3809,n3810);
and (n3809,n3631,n3645);
and (n3810,n3632,n3639);
or (n3811,n3812,n3813);
and (n3812,n3700,n3710);
and (n3813,n3701,n3702);
or (n3814,n3815,n3816);
and (n3815,n3626,n3651);
and (n3816,n3627,n3630);
xor (n3817,n3818,n3846);
xor (n3818,n3819,n3822);
or (n3819,n3820,n3821);
and (n3820,n3652,n3666);
and (n3821,n3653,n3660);
xor (n3822,n3823,n3837);
xor (n3823,n3824,n3830);
nand (n3824,n3825,n3826);
or (n3825,n1199,n3696);
or (n3826,n3827,n1192);
nor (n3827,n3828,n3829);
and (n3828,n97,n907);
and (n3829,n99,n908);
nand (n3830,n3831,n3833);
or (n3831,n3832,n625);
not (n3832,n3636);
nand (n3833,n616,n3834);
nand (n3834,n3835,n3836);
or (n3835,n515,n310);
or (n3836,n514,n308);
nand (n3837,n3838,n3842);
or (n3838,n56,n3839);
nor (n3839,n3840,n3841);
and (n3840,n1189,n65);
and (n3841,n1187,n64);
or (n3842,n57,n3843);
nor (n3843,n3844,n3845);
and (n3844,n1141,n64);
and (n3845,n65,n1143);
xor (n3846,n3847,n3862);
xor (n3847,n3848,n3855);
nand (n3848,n3849,n3854);
or (n3849,n3850,n112);
not (n3850,n3851);
nand (n3851,n3852,n3853);
or (n3852,n121,n71);
or (n3853,n125,n69);
nand (n3854,n1041,n3670);
nand (n3855,n3856,n3858);
or (n3856,n296,n3857);
not (n3857,n3681);
or (n3858,n312,n3859);
nor (n3859,n3860,n3861);
and (n3860,n40,n719);
and (n3861,n41,n721);
nand (n3862,n3863,n3864);
or (n3863,n28,n3686);
or (n3864,n37,n3865);
nor (n3865,n3866,n3867);
and (n3866,n36,n1175);
and (n3867,n34,n1177);
nand (n3868,n3869,n3876);
or (n3869,n3870,n3871);
not (n3870,n3602);
not (n3871,n3872);
nand (n3872,n3873,n3875);
or (n3873,n2697,n3874);
nand (n3874,n3198,n3199);
nand (n3875,n2698,n3085);
nor (n3876,n3877,n3881);
and (n3877,n3878,n3880);
not (n3878,n3879);
nand (n3879,n3604,n3726);
not (n3880,n3729);
and (n3881,n3730,n3733);
nand (n3882,n2696,n3602,n3883,n3887);
and (n3883,n3884,n3885,n3583);
not (n3884,n3596);
and (n3885,n3580,n3886);
or (n3886,n3502,n3291);
nand (n3887,n3888,n4391,n4400);
nand (n3888,n3889,n4325,n4384);
or (n3889,n3890,n4324);
and (n3890,n3891,n4067);
xor (n3891,n3892,n4015);
or (n3892,n3893,n4014);
and (n3893,n3894,n3975);
xor (n3894,n3895,n3924);
xor (n3895,n3896,n3915);
xor (n3896,n3897,n3906);
nand (n3897,n3898,n3902);
or (n3898,n111,n3899);
nor (n3899,n3900,n3901);
and (n3900,n125,n1141);
and (n3901,n121,n1143);
or (n3902,n112,n3903);
nor (n3903,n3904,n3905);
and (n3904,n125,n1147);
and (n3905,n121,n1149);
nand (n3906,n3907,n3911);
or (n3907,n3908,n1199);
nor (n3908,n3909,n3910);
and (n3909,n907,n185);
and (n3910,n908,n187);
or (n3911,n3912,n1192);
nor (n3912,n3913,n3914);
and (n3913,n907,n281);
and (n3914,n908,n283);
nand (n3915,n3916,n3920);
or (n3916,n625,n3917);
nor (n3917,n3918,n3919);
and (n3918,n514,n719);
and (n3919,n515,n721);
or (n3920,n617,n3921);
nor (n3921,n3922,n3923);
and (n3922,n514,n545);
and (n3923,n515,n547);
or (n3924,n3925,n3974);
and (n3925,n3926,n3949);
xor (n3926,n3927,n3933);
nand (n3927,n3928,n3932);
or (n3928,n625,n3929);
nor (n3929,n3930,n3931);
and (n3930,n514,n837);
and (n3931,n515,n839);
or (n3932,n617,n3917);
xor (n3933,n3934,n3940);
and (n3934,n3935,n121);
nand (n3935,n3936,n3937);
or (n3936,n1187,n117);
nand (n3937,n3938,n508);
not (n3938,n3939);
and (n3939,n1187,n117);
nand (n3940,n3941,n3945);
or (n3941,n1331,n3942);
nor (n3942,n3943,n3944);
and (n3943,n620,n545);
and (n3944,n621,n547);
or (n3945,n1469,n3946);
nor (n3946,n3947,n3948);
and (n3947,n620,n289);
and (n3948,n621,n291);
or (n3949,n3950,n3973);
and (n3950,n3951,n3962);
xor (n3951,n3952,n3953);
and (n3952,n113,n1187);
nand (n3953,n3954,n3958);
or (n3954,n1199,n3955);
nor (n3955,n3956,n3957);
and (n3956,n907,n289);
and (n3957,n908,n291);
or (n3958,n3959,n1192);
nor (n3959,n3960,n3961);
and (n3960,n907,n179);
and (n3961,n908,n181);
nand (n3962,n3963,n3968);
or (n3963,n3964,n509);
not (n3964,n3965);
nor (n3965,n3966,n3967);
and (n3966,n1141,n115);
and (n3967,n1143,n508);
nand (n3968,n3969,n511);
not (n3969,n3970);
nor (n3970,n3971,n3972);
and (n3971,n508,n1147);
and (n3972,n115,n1149);
and (n3973,n3952,n3953);
and (n3974,n3927,n3933);
xor (n3975,n3976,n3999);
xor (n3976,n3977,n3978);
and (n3977,n3934,n3940);
or (n3978,n3979,n3998);
and (n3979,n3980,n3995);
xor (n3980,n3981,n3987);
nand (n3981,n3982,n3983);
or (n3982,n509,n3970);
or (n3983,n639,n3984);
nor (n3984,n3985,n3986);
and (n3985,n508,n1175);
and (n3986,n115,n1177);
nand (n3987,n3988,n3993);
or (n3988,n3989,n111);
not (n3989,n3990);
nand (n3990,n3991,n3992);
or (n3991,n125,n1187);
or (n3992,n1189,n121);
nand (n3993,n3994,n113);
not (n3994,n3899);
nand (n3995,n3996,n3997);
or (n3996,n1199,n3959);
or (n3997,n3908,n1192);
and (n3998,n3981,n3987);
xor (n3999,n4000,n4008);
xor (n4000,n4001,n4002);
nor (n4001,n481,n1189);
nand (n4002,n4003,n4004);
or (n4003,n1331,n3946);
or (n4004,n1469,n4005);
nor (n4005,n4006,n4007);
and (n4006,n620,n179);
and (n4007,n621,n181);
nand (n4008,n4009,n4010);
or (n4009,n509,n3984);
or (n4010,n639,n4011);
nor (n4011,n4012,n4013);
and (n4012,n508,n837);
and (n4013,n115,n839);
and (n4014,n3895,n3924);
xor (n4015,n4016,n4064);
xor (n4016,n4017,n4045);
xor (n4017,n4018,n4031);
xor (n4018,n4019,n4025);
nand (n4019,n4020,n4024);
or (n4020,n480,n4021);
nor (n4021,n4022,n4023);
and (n4022,n1189,n143);
and (n4023,n142,n1187);
or (n4024,n481,n3551);
nand (n4025,n4026,n4027);
or (n4026,n625,n3921);
or (n4027,n617,n4028);
nor (n4028,n4029,n4030);
and (n4029,n514,n289);
and (n4030,n515,n291);
nand (n4031,n4032,n4044);
or (n4032,n4033,n4040);
not (n4033,n4034);
nand (n4034,n4035,n143);
nand (n4035,n4036,n4037);
or (n4036,n1187,n483);
nand (n4037,n4038,n125);
not (n4038,n4039);
and (n4039,n1187,n483);
not (n4040,n4041);
nand (n4041,n4042,n4043);
or (n4042,n1331,n4005);
or (n4043,n1469,n3521);
or (n4044,n4041,n4034);
xor (n4045,n4046,n4053);
xor (n4046,n4047,n4050);
or (n4047,n4048,n4049);
and (n4048,n4000,n4008);
and (n4049,n4001,n4002);
or (n4050,n4051,n4052);
and (n4051,n3896,n3915);
and (n4052,n3897,n3906);
xor (n4053,n4054,n4061);
xor (n4054,n4055,n4058);
nand (n4055,n4056,n4057);
or (n4056,n509,n4011);
or (n4057,n639,n3528);
nand (n4058,n4059,n4060);
or (n4059,n111,n3903);
or (n4060,n112,n3538);
nand (n4061,n4062,n4063);
or (n4062,n1192,n3544);
or (n4063,n3912,n1199);
or (n4064,n4065,n4066);
and (n4065,n3976,n3999);
and (n4066,n3977,n3978);
or (n4067,n4068,n4323);
and (n4068,n4069,n4109);
xor (n4069,n4070,n4108);
or (n4070,n4071,n4107);
and (n4071,n4072,n4106);
xor (n4072,n4073,n4074);
xor (n4073,n3980,n3995);
or (n4074,n4075,n4105);
and (n4075,n4076,n4091);
xor (n4076,n4077,n4083);
nand (n4077,n4078,n4082);
or (n4078,n1331,n4079);
nor (n4079,n4080,n4081);
and (n4080,n721,n621);
and (n4081,n719,n620);
or (n4082,n1469,n3942);
nand (n4083,n4084,n4089);
or (n4084,n4085,n625);
not (n4085,n4086);
nand (n4086,n4087,n4088);
or (n4087,n515,n1177);
or (n4088,n514,n1175);
nand (n4089,n4090,n616);
not (n4090,n3929);
and (n4091,n4092,n4098);
nor (n4092,n4093,n508);
nor (n4093,n4094,n4097);
and (n4094,n4095,n514);
not (n4095,n4096);
and (n4096,n1187,n513);
and (n4097,n1189,n520);
nand (n4098,n4099,n4104);
or (n4099,n1199,n4100);
not (n4100,n4101);
nor (n4101,n4102,n4103);
and (n4102,n547,n907);
and (n4103,n545,n908);
or (n4104,n3955,n1192);
and (n4105,n4077,n4083);
xor (n4106,n3926,n3949);
and (n4107,n4073,n4074);
xor (n4108,n3894,n3975);
or (n4109,n4110,n4322);
and (n4110,n4111,n4145);
xor (n4111,n4112,n4144);
or (n4112,n4113,n4143);
and (n4113,n4114,n4142);
xor (n4114,n4115,n4141);
or (n4115,n4116,n4140);
and (n4116,n4117,n4133);
xor (n4117,n4118,n4125);
nand (n4118,n4119,n4124);
or (n4119,n4120,n509);
not (n4120,n4121);
nand (n4121,n4122,n4123);
or (n4122,n508,n1187);
or (n4123,n1189,n115);
nand (n4124,n511,n3965);
nand (n4125,n4126,n4131);
or (n4126,n4127,n1331);
not (n4127,n4128);
nor (n4128,n4129,n4130);
and (n4129,n839,n620);
and (n4130,n837,n621);
nand (n4131,n4132,n904);
not (n4132,n4079);
nand (n4133,n4134,n4139);
or (n4134,n4135,n625);
not (n4135,n4136);
nor (n4136,n4137,n4138);
and (n4137,n1147,n515);
and (n4138,n1149,n514);
nand (n4139,n616,n4086);
and (n4140,n4118,n4125);
xor (n4141,n3951,n3962);
xor (n4142,n4076,n4091);
and (n4143,n4115,n4141);
xor (n4144,n4072,n4106);
nand (n4145,n4146,n4321);
or (n4146,n4147,n4177);
not (n4147,n4148);
nand (n4148,n4149,n4151);
not (n4149,n4150);
xor (n4150,n4114,n4142);
not (n4151,n4152);
or (n4152,n4153,n4176);
and (n4153,n4154,n4175);
xor (n4154,n4155,n4156);
xor (n4155,n4092,n4098);
or (n4156,n4157,n4174);
and (n4157,n4158,n4167);
xor (n4158,n4159,n4160);
and (n4159,n511,n1187);
nand (n4160,n4161,n4166);
or (n4161,n1199,n4162);
not (n4162,n4163);
nor (n4163,n4164,n4165);
and (n4164,n719,n908);
and (n4165,n721,n907);
nand (n4166,n4101,n1193);
nand (n4167,n4168,n4173);
or (n4168,n4169,n1331);
not (n4169,n4170);
nor (n4170,n4171,n4172);
and (n4171,n1177,n620);
and (n4172,n1175,n621);
nand (n4173,n904,n4128);
and (n4174,n4159,n4160);
xor (n4175,n4117,n4133);
and (n4176,n4155,n4156);
not (n4177,n4178);
nand (n4178,n4179,n4320);
or (n4179,n4180,n4210);
not (n4180,n4181);
nand (n4181,n4182,n4184);
not (n4182,n4183);
xor (n4183,n4154,n4175);
not (n4184,n4185);
or (n4185,n4186,n4209);
and (n4186,n4187,n4208);
xor (n4187,n4188,n4195);
nand (n4188,n4189,n4194);
or (n4189,n4190,n625);
not (n4190,n4191);
nor (n4191,n4192,n4193);
and (n4192,n1141,n515);
and (n4193,n1143,n514);
nand (n4194,n616,n4136);
and (n4195,n4196,n4201);
and (n4196,n4197,n515);
nand (n4197,n4198,n4200);
or (n4198,n4199,n621);
and (n4199,n1187,n619);
or (n4200,n1187,n619);
nand (n4201,n4202,n4203);
or (n4202,n1192,n4162);
nand (n4203,n4204,n1464);
not (n4204,n4205);
nor (n4205,n4206,n4207);
and (n4206,n837,n907);
and (n4207,n839,n908);
xor (n4208,n4158,n4167);
and (n4209,n4188,n4195);
not (n4210,n4211);
nand (n4211,n4212,n4319);
or (n4212,n4213,n4237);
not (n4213,n4214);
nand (n4214,n4215,n4217);
not (n4215,n4216);
xor (n4216,n4187,n4208);
not (n4217,n4218);
or (n4218,n4219,n4236);
and (n4219,n4220,n4235);
xor (n4220,n4221,n4228);
nand (n4221,n4222,n4227);
or (n4222,n4223,n1331);
not (n4223,n4224);
nor (n4224,n4225,n4226);
and (n4225,n1149,n620);
and (n4226,n1147,n621);
nand (n4227,n904,n4170);
nand (n4228,n4229,n4234);
or (n4229,n4230,n625);
not (n4230,n4231);
nand (n4231,n4232,n4233);
or (n4232,n514,n1187);
or (n4233,n515,n1189);
nand (n4234,n616,n4191);
xor (n4235,n4196,n4201);
and (n4236,n4221,n4228);
not (n4237,n4238);
nand (n4238,n4239,n4318);
or (n4239,n4240,n4264);
not (n4240,n4241);
nand (n4241,n4242,n4244);
not (n4242,n4243);
xor (n4243,n4220,n4235);
not (n4244,n4245);
or (n4245,n4246,n4263);
and (n4246,n4247,n4256);
xor (n4247,n4248,n4249);
and (n4248,n616,n1187);
nand (n4249,n4250,n4255);
or (n4250,n4251,n1331);
not (n4251,n4252);
nor (n4252,n4253,n4254);
and (n4253,n1141,n621);
and (n4254,n1143,n620);
nand (n4255,n904,n4224);
nand (n4256,n4257,n4262);
or (n4257,n1199,n4258);
not (n4258,n4259);
nor (n4259,n4260,n4261);
and (n4260,n1177,n907);
and (n4261,n1175,n908);
or (n4262,n4205,n1192);
and (n4263,n4248,n4249);
not (n4264,n4265);
nand (n4265,n4266,n4317);
or (n4266,n4267,n4283);
nor (n4267,n4268,n4269);
xor (n4268,n4247,n4256);
and (n4269,n4270,n4276);
nor (n4270,n4271,n620);
nor (n4271,n4272,n4273);
and (n4272,n914,n1189);
and (n4273,n4274,n907);
not (n4274,n4275);
and (n4275,n1187,n906);
nand (n4276,n4277,n4278);
or (n4277,n1192,n4258);
nand (n4278,n4279,n1464);
not (n4279,n4280);
nor (n4280,n4281,n4282);
and (n4281,n907,n1147);
and (n4282,n908,n1149);
not (n4283,n4284);
or (n4284,n4285,n4316);
and (n4285,n4286,n4295);
xor (n4286,n4287,n4294);
nand (n4287,n4288,n4293);
or (n4288,n4289,n1331);
not (n4289,n4290);
nand (n4290,n4291,n4292);
or (n4291,n620,n1187);
or (n4292,n621,n1189);
nand (n4293,n904,n4252);
xor (n4294,n4270,n4276);
or (n4295,n4296,n4315);
and (n4296,n4297,n4305);
xor (n4297,n4298,n4299);
nor (n4298,n1469,n1189);
nand (n4299,n4300,n4304);
or (n4300,n4301,n1199);
nor (n4301,n4302,n4303);
and (n4302,n907,n1141);
and (n4303,n908,n1143);
or (n4304,n4280,n1192);
nor (n4305,n4306,n4313);
nor (n4306,n4307,n4309);
and (n4307,n4308,n1193);
not (n4308,n4301);
nor (n4309,n4310,n1199);
nor (n4310,n4311,n4312);
and (n4311,n1187,n907);
and (n4312,n1189,n908);
or (n4313,n4314,n907);
and (n4314,n1187,n1193);
and (n4315,n4298,n4299);
and (n4316,n4287,n4294);
nand (n4317,n4268,n4269);
nand (n4318,n4243,n4245);
nand (n4319,n4216,n4218);
nand (n4320,n4183,n4185);
nand (n4321,n4150,n4152);
and (n4322,n4112,n4144);
and (n4323,n4070,n4108);
and (n4324,n3892,n4015);
nor (n4325,n4326,n4366);
not (n4326,n4327);
nand (n4327,n4328,n4350);
not (n4328,n4329);
xor (n4329,n4330,n4333);
xor (n4330,n4331,n4332);
xor (n4331,n3375,n3430);
xor (n4332,n3508,n3511);
or (n4333,n4334,n4349);
and (n4334,n4335,n4338);
xor (n4335,n4336,n4337);
xor (n4336,n3407,n3423);
xor (n4337,n3378,n3395);
or (n4338,n4339,n4348);
and (n4339,n4340,n4345);
xor (n4340,n4341,n4344);
nand (n4341,n4342,n4343);
or (n4342,n625,n4028);
or (n4343,n617,n3410);
and (n4344,n4041,n4033);
or (n4345,n4346,n4347);
and (n4346,n4054,n4061);
and (n4347,n4055,n4058);
and (n4348,n4341,n4344);
and (n4349,n4336,n4337);
not (n4350,n4351);
or (n4351,n4352,n4365);
and (n4352,n4353,n4364);
xor (n4353,n4354,n4355);
xor (n4354,n3513,n3533);
or (n4355,n4356,n4363);
and (n4356,n4357,n4360);
xor (n4357,n4358,n4359);
xor (n4358,n3535,n3549);
xor (n4359,n3517,n3526);
or (n4360,n4361,n4362);
and (n4361,n4018,n4031);
and (n4362,n4019,n4025);
and (n4363,n4358,n4359);
xor (n4364,n4335,n4338);
and (n4365,n4354,n4355);
nand (n4366,n4367,n4379);
not (n4367,n4368);
nor (n4368,n4369,n4370);
xor (n4369,n4353,n4364);
or (n4370,n4371,n4378);
and (n4371,n4372,n4377);
xor (n4372,n4373,n4374);
xor (n4373,n4340,n4345);
or (n4374,n4375,n4376);
and (n4375,n4046,n4053);
and (n4376,n4047,n4050);
xor (n4377,n4357,n4360);
and (n4378,n4373,n4374);
or (n4379,n4380,n4383);
or (n4380,n4381,n4382);
and (n4381,n4016,n4064);
and (n4382,n4017,n4045);
xor (n4383,n4372,n4377);
nand (n4384,n4385,n4387);
not (n4385,n4386);
xor (n4386,n3504,n3558);
not (n4387,n4388);
or (n4388,n4389,n4390);
and (n4389,n4330,n4333);
and (n4390,n4331,n4332);
nand (n4391,n4392,n4384);
nand (n4392,n4393,n4399);
or (n4393,n4326,n4394);
not (n4394,n4395);
nand (n4395,n4396,n4398);
or (n4396,n4368,n4397);
nand (n4397,n4380,n4383);
nand (n4398,n4369,n4370);
nand (n4399,n4329,n4351);
nand (n4400,n4386,n4388);
and (n4401,n4402,n4568,n4599);
nand (n4402,n4403,n4536);
not (n4403,n4404);
xor (n4404,n4405,n4523);
xor (n4405,n4406,n4407);
xor (n4406,n2679,n2688);
or (n4407,n4408,n4522);
and (n4408,n4409,n4505);
xor (n4409,n4410,n4482);
or (n4410,n4411,n4481);
and (n4411,n4412,n4453);
xor (n4412,n4413,n4424);
or (n4413,n4414,n4423);
and (n4414,n4415,n4420);
xor (n4415,n4416,n4419);
nand (n4416,n4417,n4418);
or (n4417,n137,n3779);
or (n4418,n155,n2661);
and (n4419,n3783,n3788);
or (n4420,n4421,n4422);
and (n4421,n3847,n3862);
and (n4422,n3848,n3855);
and (n4423,n4416,n4419);
xor (n4424,n4425,n4452);
xor (n4425,n4426,n4441);
or (n4426,n4427,n4440);
and (n4427,n4428,n4437);
xor (n4428,n4429,n4434);
nand (n4429,n4430,n4432);
or (n4430,n4431,n625);
not (n4431,n3834);
nand (n4432,n4433,n616);
not (n4433,n2655);
nand (n4434,n4435,n4436);
or (n4435,n56,n3843);
or (n4436,n57,n2636);
nand (n4437,n4438,n4439);
or (n4438,n480,n3773);
or (n4439,n481,n2629);
and (n4440,n4429,n4434);
or (n4441,n4442,n4451);
and (n4442,n4443,n4448);
xor (n4443,n4444,n4445);
nor (n4444,n212,n1189);
nand (n4445,n4446,n4447);
or (n4446,n3790,n1331);
or (n4447,n1469,n2559);
nand (n4448,n4449,n4450);
or (n4449,n509,n3752);
or (n4450,n639,n2577);
and (n4451,n4444,n4445);
xor (n4452,n2646,n2659);
or (n4453,n4454,n4480);
and (n4454,n4455,n4469);
xor (n4455,n4456,n4468);
xor (n4456,n4457,n4465);
xor (n4457,n4458,n4462);
nand (n4458,n4459,n4460);
or (n4459,n3859,n296);
nand (n4460,n4461,n298);
not (n4461,n2606);
nand (n4462,n4463,n4464);
or (n4463,n28,n3865);
or (n4464,n37,n2613);
nand (n4465,n4466,n4467);
or (n4466,n1199,n3827);
or (n4467,n2623,n1192);
xor (n4468,n4443,n4448);
xor (n4469,n4470,n4477);
xor (n4470,n4471,n4474);
nand (n4471,n4472,n4473);
or (n4472,n80,n3759);
or (n4473,n81,n2584);
nand (n4474,n4475,n4476);
or (n4475,n236,n3765);
or (n4476,n254,n2590);
nand (n4477,n4478,n4479);
or (n4478,n111,n3850);
or (n4479,n112,n2600);
and (n4480,n4456,n4468);
and (n4481,n4413,n4424);
xor (n4482,n4483,n4498);
xor (n4483,n4484,n4495);
or (n4484,n4485,n4494);
and (n4485,n4486,n4491);
xor (n4486,n4487,n4488);
xor (n4487,n2552,n2557);
or (n4488,n4489,n4490);
and (n4489,n4470,n4477);
and (n4490,n4471,n4474);
or (n4491,n4492,n4493);
and (n4492,n4457,n4465);
and (n4493,n4458,n4462);
and (n4494,n4487,n4488);
or (n4495,n4496,n4497);
and (n4496,n4425,n4452);
and (n4497,n4426,n4441);
or (n4498,n4499,n4504);
and (n4499,n4500,n4503);
xor (n4500,n4501,n4502);
xor (n4501,n2574,n2588);
xor (n4502,n2597,n2611);
xor (n4503,n2620,n2633);
and (n4504,n4501,n4502);
or (n4505,n4506,n4521);
and (n4506,n4507,n4520);
xor (n4507,n4508,n4519);
or (n4508,n4509,n4518);
and (n4509,n4510,n4517);
xor (n4510,n4511,n4514);
or (n4511,n4512,n4513);
and (n4512,n3823,n3837);
and (n4513,n3824,n3830);
or (n4514,n4515,n4516);
and (n4515,n3746,n3762);
and (n4516,n3747,n3755);
xor (n4517,n4428,n4437);
and (n4518,n4511,n4514);
xor (n4519,n4486,n4491);
xor (n4520,n4500,n4503);
and (n4521,n4508,n4519);
and (n4522,n4410,n4482);
xor (n4523,n4524,n4535);
xor (n4524,n4525,n4528);
or (n4525,n4526,n4527);
and (n4526,n4483,n4498);
and (n4527,n4484,n4495);
or (n4528,n4529,n4534);
and (n4529,n4530,n4533);
xor (n4530,n4531,n4532);
xor (n4531,n2571,n2618);
xor (n4532,n2682,n2685);
xor (n4533,n2643,n2667);
and (n4534,n4531,n4532);
xor (n4535,n2568,n2669);
not (n4536,n4537);
or (n4537,n4538,n4567);
and (n4538,n4539,n4566);
xor (n4539,n4540,n4541);
xor (n4540,n4530,n4533);
or (n4541,n4542,n4565);
and (n4542,n4543,n4564);
xor (n4543,n4544,n4555);
or (n4544,n4545,n4554);
and (n4545,n4546,n4553);
xor (n4546,n4547,n4550);
or (n4547,n4548,n4549);
and (n4548,n3769,n3782);
and (n4549,n3770,n3776);
or (n4550,n4551,n4552);
and (n4551,n3804,n3811);
and (n4552,n3805,n3808);
xor (n4553,n4415,n4420);
and (n4554,n4547,n4550);
or (n4555,n4556,n4563);
and (n4556,n4557,n4562);
xor (n4557,n4558,n4559);
xor (n4558,n4510,n4517);
or (n4559,n4560,n4561);
and (n4560,n3818,n3846);
and (n4561,n3819,n3822);
xor (n4562,n4455,n4469);
and (n4563,n4558,n4559);
xor (n4564,n4412,n4453);
and (n4565,n4544,n4555);
xor (n4566,n4409,n4505);
and (n4567,n4540,n4541);
nor (n4568,n4569,n4588);
nor (n4569,n4570,n4585);
xor (n4570,n4571,n4582);
xor (n4571,n4572,n4573);
xor (n4572,n4557,n4562);
xor (n4573,n4574,n4579);
xor (n4574,n4575,n4578);
or (n4575,n4576,n4577);
and (n4576,n3744,n3795);
and (n4577,n3745,n3768);
xor (n4578,n4546,n4553);
or (n4579,n4580,n4581);
and (n4580,n3802,n3817);
and (n4581,n3803,n3814);
or (n4582,n4583,n4584);
and (n4583,n3742,n3801);
and (n4584,n3743,n3798);
or (n4585,n4586,n4587);
and (n4586,n3734,n3741);
and (n4587,n3735,n3738);
nor (n4588,n4589,n4592);
or (n4589,n4590,n4591);
and (n4590,n4571,n4582);
and (n4591,n4572,n4573);
xor (n4592,n4593,n4598);
xor (n4593,n4594,n4595);
xor (n4594,n4507,n4520);
or (n4595,n4596,n4597);
and (n4596,n4574,n4579);
and (n4597,n4575,n4578);
xor (n4598,n4543,n4564);
not (n4599,n4600);
nor (n4600,n4601,n4602);
xor (n4601,n4539,n4566);
or (n4602,n4603,n4604);
and (n4603,n4593,n4598);
and (n4604,n4594,n4595);
nor (n4605,n4606,n4617);
nor (n4606,n4607,n4608);
xor (n4607,n2527,n2691);
or (n4608,n4609,n4616);
and (n4609,n4610,n4615);
xor (n4610,n4611,n4612);
xor (n4611,n2530,n2566);
or (n4612,n4613,n4614);
and (n4613,n4524,n4535);
and (n4614,n4525,n4528);
xor (n4615,n2674,n2677);
and (n4616,n4611,n4612);
nor (n4617,n4618,n4619);
xor (n4618,n4610,n4615);
or (n4619,n4620,n4621);
and (n4620,n4405,n4523);
and (n4621,n4406,n4407);
nand (n4622,n4623,n2507,n4605);
nand (n4623,n4624,n4634);
or (n4624,n4625,n4626);
not (n4625,n4402);
not (n4626,n4627);
nand (n4627,n4628,n4633);
or (n4628,n4629,n4600);
nor (n4629,n4630,n4632);
nor (n4630,n4588,n4631);
nand (n4631,n4570,n4585);
and (n4632,n4589,n4592);
nand (n4633,n4601,n4602);
nand (n4634,n4404,n4537);
nor (n4635,n4636,n4641);
and (n4636,n2507,n4637);
nand (n4637,n4638,n4640);
or (n4638,n4606,n4639);
nand (n4639,n4618,n4619);
nand (n4640,n4607,n4608);
nand (n4641,n4642,n4644);
or (n4642,n2508,n4643);
nand (n4643,n2524,n2525);
nand (n4644,n2509,n2510);
nor (n4645,n4646,n4647);
not (n4646,n2421);
nand (n4647,n2285,n4648);
nor (n4648,n1118,n4649);
nor (n4649,n2147,n2282);
or (n4650,n4651,n9041);
and (n4651,n4652,n9040);
wire s0n4652,s1n4652,notn4652;
or (n4652,s0n4652,s1n4652);
not(notn4652,n10);
and (s0n4652,notn4652,n3);
and (s1n4652,n10,n4653);
xor (n4653,n4654,n8883);
xor (n4654,n4655,n9038);
xor (n4655,n4656,n8878);
xor (n4656,n4657,n9031);
xor (n4657,n4658,n8872);
xor (n4658,n4659,n9019);
xor (n4659,n4660,n8866);
xor (n4660,n4661,n9002);
xor (n4661,n4662,n8860);
xor (n4662,n4663,n8980);
xor (n4663,n4664,n8854);
xor (n4664,n4665,n8953);
xor (n4665,n4666,n8848);
xor (n4666,n4667,n8921);
xor (n4667,n4668,n8842);
xor (n4668,n4669,n8884);
xor (n4669,n4670,n8836);
xor (n4670,n4671,n8833);
xor (n4671,n4672,n8832);
xor (n4672,n4673,n8775);
xor (n4673,n4674,n8774);
xor (n4674,n4675,n8711);
xor (n4675,n4676,n8710);
xor (n4676,n4677,n8641);
xor (n4677,n4678,n8640);
xor (n4678,n4679,n8565);
xor (n4679,n4680,n8564);
xor (n4680,n4681,n8484);
xor (n4681,n4682,n8483);
xor (n4682,n4683,n8398);
xor (n4683,n4684,n8397);
xor (n4684,n4685,n8304);
xor (n4685,n4686,n8303);
xor (n4686,n4687,n8204);
xor (n4687,n4688,n8203);
xor (n4688,n4689,n8098);
xor (n4689,n4690,n8097);
xor (n4690,n4691,n7986);
xor (n4691,n4692,n7985);
xor (n4692,n4693,n7869);
xor (n4693,n4694,n7868);
xor (n4694,n4695,n7749);
xor (n4695,n4696,n7748);
xor (n4696,n4697,n7619);
xor (n4697,n4698,n7618);
xor (n4698,n4699,n7483);
xor (n4699,n4700,n7482);
xor (n4700,n4701,n7341);
xor (n4701,n4702,n7340);
xor (n4702,n4703,n7195);
xor (n4703,n4704,n7194);
xor (n4704,n4705,n7041);
xor (n4705,n4706,n7040);
xor (n4706,n4707,n6881);
xor (n4707,n4708,n6880);
xor (n4708,n4709,n6715);
xor (n4709,n4710,n6714);
xor (n4710,n4711,n6544);
xor (n4711,n4712,n6543);
xor (n4712,n4713,n6367);
xor (n4713,n4714,n6366);
xor (n4714,n4715,n4748);
xor (n4715,n4716,n4747);
xor (n4716,n4717,n4746);
xor (n4717,n4718,n4745);
xor (n4718,n4719,n4744);
xor (n4719,n4720,n4743);
xor (n4720,n4721,n4742);
xor (n4721,n4722,n4741);
xor (n4722,n4723,n4740);
xor (n4723,n4724,n4739);
xor (n4724,n4725,n4738);
xor (n4725,n4726,n4737);
xor (n4726,n4727,n4736);
xor (n4727,n4728,n916);
xor (n4728,n4729,n4735);
xor (n4729,n4730,n4734);
xor (n4730,n4731,n4733);
xor (n4731,n4732,n1196);
and (n4732,n132,n1193);
and (n4733,n4732,n1196);
and (n4734,n132,n906);
and (n4735,n4730,n4734);
and (n4736,n4728,n916);
and (n4737,n132,n619);
and (n4738,n4726,n4737);
and (n4739,n132,n515);
and (n4740,n4724,n4739);
and (n4741,n132,n513);
and (n4742,n4722,n4741);
and (n4743,n132,n115);
and (n4744,n4720,n4743);
and (n4745,n132,n117);
and (n4746,n4718,n4745);
and (n4747,n132,n121);
or (n4748,n4749,n6189);
and (n4749,n4750,n6188);
xor (n4750,n4717,n4751);
or (n4751,n4752,n6010);
and (n4752,n4753,n6009);
xor (n4753,n4719,n4754);
or (n4754,n4755,n5836);
and (n4755,n4756,n5835);
xor (n4756,n4721,n4757);
or (n4757,n4758,n5657);
and (n4758,n4759,n5656);
xor (n4759,n4723,n4760);
or (n4760,n4761,n5482);
and (n4761,n4762,n5481);
xor (n4762,n4725,n4763);
or (n4763,n4764,n5303);
and (n4764,n4765,n5302);
xor (n4765,n4727,n4766);
or (n4766,n4767,n5129);
and (n4767,n4768,n5128);
xor (n4768,n4729,n4769);
or (n4769,n4770,n4950);
and (n4770,n4771,n4949);
xor (n4771,n4731,n4772);
or (n4772,n4773,n4775);
and (n4773,n4732,n4774);
and (n4774,n126,n908);
and (n4775,n4776,n4777);
xor (n4776,n4732,n4774);
or (n4777,n4778,n4780);
and (n4778,n4779,n1323);
and (n4779,n126,n1193);
and (n4780,n4781,n4782);
xor (n4781,n4779,n1323);
or (n4782,n4783,n4786);
and (n4783,n4784,n4785);
and (n4784,n329,n1193);
and (n4785,n324,n908);
and (n4786,n4787,n4788);
xor (n4787,n4784,n4785);
or (n4788,n4789,n4792);
and (n4789,n4790,n4791);
and (n4790,n324,n1193);
and (n4791,n158,n908);
and (n4792,n4793,n4794);
xor (n4793,n4790,n4791);
or (n4794,n4795,n4798);
and (n4795,n4796,n4797);
and (n4796,n158,n1193);
and (n4797,n151,n908);
and (n4798,n4799,n4800);
xor (n4799,n4796,n4797);
or (n4800,n4801,n4804);
and (n4801,n4802,n4803);
and (n4802,n151,n1193);
and (n4803,n195,n908);
and (n4804,n4805,n4806);
xor (n4805,n4802,n4803);
or (n4806,n4807,n4810);
and (n4807,n4808,n4809);
and (n4808,n195,n1193);
and (n4809,n103,n908);
and (n4810,n4811,n4812);
xor (n4811,n4808,n4809);
or (n4812,n4813,n4816);
and (n4813,n4814,n4815);
and (n4814,n103,n1193);
and (n4815,n97,n908);
and (n4816,n4817,n4818);
xor (n4817,n4814,n4815);
or (n4818,n4819,n4822);
and (n4819,n4820,n4821);
and (n4820,n97,n1193);
and (n4821,n257,n908);
and (n4822,n4823,n4824);
xor (n4823,n4820,n4821);
or (n4824,n4825,n4828);
and (n4825,n4826,n4827);
and (n4826,n257,n1193);
and (n4827,n250,n908);
and (n4828,n4829,n4830);
xor (n4829,n4826,n4827);
or (n4830,n4831,n4834);
and (n4831,n4832,n4833);
and (n4832,n250,n1193);
and (n4833,n315,n908);
and (n4834,n4835,n4836);
xor (n4835,n4832,n4833);
or (n4836,n4837,n4840);
and (n4837,n4838,n4839);
and (n4838,n315,n1193);
and (n4839,n308,n908);
and (n4840,n4841,n4842);
xor (n4841,n4838,n4839);
or (n4842,n4843,n4846);
and (n4843,n4844,n4845);
and (n4844,n308,n1193);
and (n4845,n51,n908);
and (n4846,n4847,n4848);
xor (n4847,n4844,n4845);
or (n4848,n4849,n4852);
and (n4849,n4850,n4851);
and (n4850,n51,n1193);
and (n4851,n45,n908);
and (n4852,n4853,n4854);
xor (n4853,n4850,n4851);
or (n4854,n4855,n4858);
and (n4855,n4856,n4857);
and (n4856,n45,n1193);
and (n4857,n75,n908);
and (n4858,n4859,n4860);
xor (n4859,n4856,n4857);
or (n4860,n4861,n4864);
and (n4861,n4862,n4863);
and (n4862,n75,n1193);
and (n4863,n69,n908);
and (n4864,n4865,n4866);
xor (n4865,n4862,n4863);
or (n4866,n4867,n4870);
and (n4867,n4868,n4869);
and (n4868,n69,n1193);
and (n4869,n226,n908);
and (n4870,n4871,n4872);
xor (n4871,n4868,n4869);
or (n4872,n4873,n4876);
and (n4873,n4874,n4875);
and (n4874,n226,n1193);
and (n4875,n351,n908);
and (n4876,n4877,n4878);
xor (n4877,n4874,n4875);
or (n4878,n4879,n4882);
and (n4879,n4880,n4881);
and (n4880,n351,n1193);
and (n4881,n345,n908);
and (n4882,n4883,n4884);
xor (n4883,n4880,n4881);
or (n4884,n4885,n4887);
and (n4885,n4886,n3546);
and (n4886,n345,n1193);
and (n4887,n4888,n4889);
xor (n4888,n4886,n3546);
or (n4889,n4890,n4893);
and (n4890,n4891,n4892);
and (n4891,n372,n1193);
and (n4892,n281,n908);
and (n4893,n4894,n4895);
xor (n4894,n4891,n4892);
or (n4895,n4896,n4899);
and (n4896,n4897,n4898);
and (n4897,n281,n1193);
and (n4898,n185,n908);
and (n4899,n4900,n4901);
xor (n4900,n4897,n4898);
or (n4901,n4902,n4905);
and (n4902,n4903,n4904);
and (n4903,n185,n1193);
and (n4904,n179,n908);
and (n4905,n4906,n4907);
xor (n4906,n4903,n4904);
or (n4907,n4908,n4911);
and (n4908,n4909,n4910);
and (n4909,n179,n1193);
and (n4910,n289,n908);
and (n4911,n4912,n4913);
xor (n4912,n4909,n4910);
or (n4913,n4914,n4916);
and (n4914,n4915,n4103);
and (n4915,n289,n1193);
and (n4916,n4917,n4918);
xor (n4917,n4915,n4103);
or (n4918,n4919,n4921);
and (n4919,n4920,n4164);
and (n4920,n545,n1193);
and (n4921,n4922,n4923);
xor (n4922,n4920,n4164);
or (n4923,n4924,n4927);
and (n4924,n4925,n4926);
and (n4925,n719,n1193);
and (n4926,n837,n908);
and (n4927,n4928,n4929);
xor (n4928,n4925,n4926);
or (n4929,n4930,n4932);
and (n4930,n4931,n4261);
and (n4931,n837,n1193);
and (n4932,n4933,n4934);
xor (n4933,n4931,n4261);
or (n4934,n4935,n4938);
and (n4935,n4936,n4937);
and (n4936,n1175,n1193);
and (n4937,n1147,n908);
and (n4938,n4939,n4940);
xor (n4939,n4936,n4937);
or (n4940,n4941,n4944);
and (n4941,n4942,n4943);
and (n4942,n1147,n1193);
and (n4943,n1141,n908);
and (n4944,n4945,n4946);
xor (n4945,n4942,n4943);
and (n4946,n4947,n4948);
and (n4947,n1141,n1193);
and (n4948,n1187,n908);
and (n4949,n126,n906);
and (n4950,n4951,n4952);
xor (n4951,n4771,n4949);
or (n4952,n4953,n4956);
and (n4953,n4954,n4955);
xor (n4954,n4776,n4777);
and (n4955,n329,n906);
and (n4956,n4957,n4958);
xor (n4957,n4954,n4955);
or (n4958,n4959,n4962);
and (n4959,n4960,n4961);
xor (n4960,n4781,n4782);
and (n4961,n324,n906);
and (n4962,n4963,n4964);
xor (n4963,n4960,n4961);
or (n4964,n4965,n4968);
and (n4965,n4966,n4967);
xor (n4966,n4787,n4788);
and (n4967,n158,n906);
and (n4968,n4969,n4970);
xor (n4969,n4966,n4967);
or (n4970,n4971,n4974);
and (n4971,n4972,n4973);
xor (n4972,n4793,n4794);
and (n4973,n151,n906);
and (n4974,n4975,n4976);
xor (n4975,n4972,n4973);
or (n4976,n4977,n4980);
and (n4977,n4978,n4979);
xor (n4978,n4799,n4800);
and (n4979,n195,n906);
and (n4980,n4981,n4982);
xor (n4981,n4978,n4979);
or (n4982,n4983,n4986);
and (n4983,n4984,n4985);
xor (n4984,n4805,n4806);
and (n4985,n103,n906);
and (n4986,n4987,n4988);
xor (n4987,n4984,n4985);
or (n4988,n4989,n4992);
and (n4989,n4990,n4991);
xor (n4990,n4811,n4812);
and (n4991,n97,n906);
and (n4992,n4993,n4994);
xor (n4993,n4990,n4991);
or (n4994,n4995,n4998);
and (n4995,n4996,n4997);
xor (n4996,n4817,n4818);
and (n4997,n257,n906);
and (n4998,n4999,n5000);
xor (n4999,n4996,n4997);
or (n5000,n5001,n5004);
and (n5001,n5002,n5003);
xor (n5002,n4823,n4824);
and (n5003,n250,n906);
and (n5004,n5005,n5006);
xor (n5005,n5002,n5003);
or (n5006,n5007,n5010);
and (n5007,n5008,n5009);
xor (n5008,n4829,n4830);
and (n5009,n315,n906);
and (n5010,n5011,n5012);
xor (n5011,n5008,n5009);
or (n5012,n5013,n5016);
and (n5013,n5014,n5015);
xor (n5014,n4835,n4836);
and (n5015,n308,n906);
and (n5016,n5017,n5018);
xor (n5017,n5014,n5015);
or (n5018,n5019,n5022);
and (n5019,n5020,n5021);
xor (n5020,n4841,n4842);
and (n5021,n51,n906);
and (n5022,n5023,n5024);
xor (n5023,n5020,n5021);
or (n5024,n5025,n5028);
and (n5025,n5026,n5027);
xor (n5026,n4847,n4848);
and (n5027,n45,n906);
and (n5028,n5029,n5030);
xor (n5029,n5026,n5027);
or (n5030,n5031,n5034);
and (n5031,n5032,n5033);
xor (n5032,n4853,n4854);
and (n5033,n75,n906);
and (n5034,n5035,n5036);
xor (n5035,n5032,n5033);
or (n5036,n5037,n5040);
and (n5037,n5038,n5039);
xor (n5038,n4859,n4860);
and (n5039,n69,n906);
and (n5040,n5041,n5042);
xor (n5041,n5038,n5039);
or (n5042,n5043,n5046);
and (n5043,n5044,n5045);
xor (n5044,n4865,n4866);
and (n5045,n226,n906);
and (n5046,n5047,n5048);
xor (n5047,n5044,n5045);
or (n5048,n5049,n5052);
and (n5049,n5050,n5051);
xor (n5050,n4871,n4872);
and (n5051,n351,n906);
and (n5052,n5053,n5054);
xor (n5053,n5050,n5051);
or (n5054,n5055,n5058);
and (n5055,n5056,n5057);
xor (n5056,n4877,n4878);
and (n5057,n345,n906);
and (n5058,n5059,n5060);
xor (n5059,n5056,n5057);
or (n5060,n5061,n5064);
and (n5061,n5062,n5063);
xor (n5062,n4883,n4884);
and (n5063,n372,n906);
and (n5064,n5065,n5066);
xor (n5065,n5062,n5063);
or (n5066,n5067,n5070);
and (n5067,n5068,n5069);
xor (n5068,n4888,n4889);
and (n5069,n281,n906);
and (n5070,n5071,n5072);
xor (n5071,n5068,n5069);
or (n5072,n5073,n5076);
and (n5073,n5074,n5075);
xor (n5074,n4894,n4895);
and (n5075,n185,n906);
and (n5076,n5077,n5078);
xor (n5077,n5074,n5075);
or (n5078,n5079,n5082);
and (n5079,n5080,n5081);
xor (n5080,n4900,n4901);
and (n5081,n179,n906);
and (n5082,n5083,n5084);
xor (n5083,n5080,n5081);
or (n5084,n5085,n5088);
and (n5085,n5086,n5087);
xor (n5086,n4906,n4907);
and (n5087,n289,n906);
and (n5088,n5089,n5090);
xor (n5089,n5086,n5087);
or (n5090,n5091,n5094);
and (n5091,n5092,n5093);
xor (n5092,n4912,n4913);
and (n5093,n545,n906);
and (n5094,n5095,n5096);
xor (n5095,n5092,n5093);
or (n5096,n5097,n5100);
and (n5097,n5098,n5099);
xor (n5098,n4917,n4918);
and (n5099,n719,n906);
and (n5100,n5101,n5102);
xor (n5101,n5098,n5099);
or (n5102,n5103,n5106);
and (n5103,n5104,n5105);
xor (n5104,n4922,n4923);
and (n5105,n837,n906);
and (n5106,n5107,n5108);
xor (n5107,n5104,n5105);
or (n5108,n5109,n5112);
and (n5109,n5110,n5111);
xor (n5110,n4928,n4929);
and (n5111,n1175,n906);
and (n5112,n5113,n5114);
xor (n5113,n5110,n5111);
or (n5114,n5115,n5118);
and (n5115,n5116,n5117);
xor (n5116,n4933,n4934);
and (n5117,n1147,n906);
and (n5118,n5119,n5120);
xor (n5119,n5116,n5117);
or (n5120,n5121,n5124);
and (n5121,n5122,n5123);
xor (n5122,n4939,n4940);
and (n5123,n1141,n906);
and (n5124,n5125,n5126);
xor (n5125,n5122,n5123);
and (n5126,n5127,n4275);
xor (n5127,n4945,n4946);
and (n5128,n126,n621);
and (n5129,n5130,n5131);
xor (n5130,n4768,n5128);
or (n5131,n5132,n5135);
and (n5132,n5133,n5134);
xor (n5133,n4951,n4952);
and (n5134,n329,n621);
and (n5135,n5136,n5137);
xor (n5136,n5133,n5134);
or (n5137,n5138,n5140);
and (n5138,n5139,n1334);
xor (n5139,n4957,n4958);
and (n5140,n5141,n5142);
xor (n5141,n5139,n1334);
or (n5142,n5143,n5146);
and (n5143,n5144,n5145);
xor (n5144,n4963,n4964);
and (n5145,n158,n621);
and (n5146,n5147,n5148);
xor (n5147,n5144,n5145);
or (n5148,n5149,n5152);
and (n5149,n5150,n5151);
xor (n5150,n4969,n4970);
and (n5151,n151,n621);
and (n5152,n5153,n5154);
xor (n5153,n5150,n5151);
or (n5154,n5155,n5158);
and (n5155,n5156,n5157);
xor (n5156,n4975,n4976);
and (n5157,n195,n621);
and (n5158,n5159,n5160);
xor (n5159,n5156,n5157);
or (n5160,n5161,n5164);
and (n5161,n5162,n5163);
xor (n5162,n4981,n4982);
and (n5163,n103,n621);
and (n5164,n5165,n5166);
xor (n5165,n5162,n5163);
or (n5166,n5167,n5170);
and (n5167,n5168,n5169);
xor (n5168,n4987,n4988);
and (n5169,n97,n621);
and (n5170,n5171,n5172);
xor (n5171,n5168,n5169);
or (n5172,n5173,n5176);
and (n5173,n5174,n5175);
xor (n5174,n4993,n4994);
and (n5175,n257,n621);
and (n5176,n5177,n5178);
xor (n5177,n5174,n5175);
or (n5178,n5179,n5182);
and (n5179,n5180,n5181);
xor (n5180,n4999,n5000);
and (n5181,n250,n621);
and (n5182,n5183,n5184);
xor (n5183,n5180,n5181);
or (n5184,n5185,n5188);
and (n5185,n5186,n5187);
xor (n5186,n5005,n5006);
and (n5187,n315,n621);
and (n5188,n5189,n5190);
xor (n5189,n5186,n5187);
or (n5190,n5191,n5193);
and (n5191,n5192,n3045);
xor (n5192,n5011,n5012);
and (n5193,n5194,n5195);
xor (n5194,n5192,n3045);
or (n5195,n5196,n5199);
and (n5196,n5197,n5198);
xor (n5197,n5017,n5018);
and (n5198,n51,n621);
and (n5199,n5200,n5201);
xor (n5200,n5197,n5198);
or (n5201,n5202,n5205);
and (n5202,n5203,n5204);
xor (n5203,n5023,n5024);
and (n5204,n45,n621);
and (n5205,n5206,n5207);
xor (n5206,n5203,n5204);
or (n5207,n5208,n5211);
and (n5208,n5209,n5210);
xor (n5209,n5029,n5030);
and (n5210,n75,n621);
and (n5211,n5212,n5213);
xor (n5212,n5209,n5210);
or (n5213,n5214,n5217);
and (n5214,n5215,n5216);
xor (n5215,n5035,n5036);
and (n5216,n69,n621);
and (n5217,n5218,n5219);
xor (n5218,n5215,n5216);
or (n5219,n5220,n5223);
and (n5220,n5221,n5222);
xor (n5221,n5041,n5042);
and (n5222,n226,n621);
and (n5223,n5224,n5225);
xor (n5224,n5221,n5222);
or (n5225,n5226,n5229);
and (n5226,n5227,n5228);
xor (n5227,n5047,n5048);
and (n5228,n351,n621);
and (n5229,n5230,n5231);
xor (n5230,n5227,n5228);
or (n5231,n5232,n5235);
and (n5232,n5233,n5234);
xor (n5233,n5053,n5054);
and (n5234,n345,n621);
and (n5235,n5236,n5237);
xor (n5236,n5233,n5234);
or (n5237,n5238,n5241);
and (n5238,n5239,n5240);
xor (n5239,n5059,n5060);
and (n5240,n372,n621);
and (n5241,n5242,n5243);
xor (n5242,n5239,n5240);
or (n5243,n5244,n5247);
and (n5244,n5245,n5246);
xor (n5245,n5065,n5066);
and (n5246,n281,n621);
and (n5247,n5248,n5249);
xor (n5248,n5245,n5246);
or (n5249,n5250,n5253);
and (n5250,n5251,n5252);
xor (n5251,n5071,n5072);
and (n5252,n185,n621);
and (n5253,n5254,n5255);
xor (n5254,n5251,n5252);
or (n5255,n5256,n5259);
and (n5256,n5257,n5258);
xor (n5257,n5077,n5078);
and (n5258,n179,n621);
and (n5259,n5260,n5261);
xor (n5260,n5257,n5258);
or (n5261,n5262,n5265);
and (n5262,n5263,n5264);
xor (n5263,n5083,n5084);
and (n5264,n289,n621);
and (n5265,n5266,n5267);
xor (n5266,n5263,n5264);
or (n5267,n5268,n5271);
and (n5268,n5269,n5270);
xor (n5269,n5089,n5090);
and (n5270,n545,n621);
and (n5271,n5272,n5273);
xor (n5272,n5269,n5270);
or (n5273,n5274,n5277);
and (n5274,n5275,n5276);
xor (n5275,n5095,n5096);
and (n5276,n719,n621);
and (n5277,n5278,n5279);
xor (n5278,n5275,n5276);
or (n5279,n5280,n5282);
and (n5280,n5281,n4130);
xor (n5281,n5101,n5102);
and (n5282,n5283,n5284);
xor (n5283,n5281,n4130);
or (n5284,n5285,n5287);
and (n5285,n5286,n4172);
xor (n5286,n5107,n5108);
and (n5287,n5288,n5289);
xor (n5288,n5286,n4172);
or (n5289,n5290,n5292);
and (n5290,n5291,n4226);
xor (n5291,n5113,n5114);
and (n5292,n5293,n5294);
xor (n5293,n5291,n4226);
or (n5294,n5295,n5297);
and (n5295,n5296,n4253);
xor (n5296,n5119,n5120);
and (n5297,n5298,n5299);
xor (n5298,n5296,n4253);
and (n5299,n5300,n5301);
xor (n5300,n5125,n5126);
and (n5301,n1187,n621);
and (n5302,n126,n619);
and (n5303,n5304,n5305);
xor (n5304,n4765,n5302);
or (n5305,n5306,n5309);
and (n5306,n5307,n5308);
xor (n5307,n5130,n5131);
and (n5308,n329,n619);
and (n5309,n5310,n5311);
xor (n5310,n5307,n5308);
or (n5311,n5312,n5315);
and (n5312,n5313,n5314);
xor (n5313,n5136,n5137);
and (n5314,n324,n619);
and (n5315,n5316,n5317);
xor (n5316,n5313,n5314);
or (n5317,n5318,n5321);
and (n5318,n5319,n5320);
xor (n5319,n5141,n5142);
and (n5320,n158,n619);
and (n5321,n5322,n5323);
xor (n5322,n5319,n5320);
or (n5323,n5324,n5327);
and (n5324,n5325,n5326);
xor (n5325,n5147,n5148);
and (n5326,n151,n619);
and (n5327,n5328,n5329);
xor (n5328,n5325,n5326);
or (n5329,n5330,n5333);
and (n5330,n5331,n5332);
xor (n5331,n5153,n5154);
and (n5332,n195,n619);
and (n5333,n5334,n5335);
xor (n5334,n5331,n5332);
or (n5335,n5336,n5339);
and (n5336,n5337,n5338);
xor (n5337,n5159,n5160);
and (n5338,n103,n619);
and (n5339,n5340,n5341);
xor (n5340,n5337,n5338);
or (n5341,n5342,n5345);
and (n5342,n5343,n5344);
xor (n5343,n5165,n5166);
and (n5344,n97,n619);
and (n5345,n5346,n5347);
xor (n5346,n5343,n5344);
or (n5347,n5348,n5351);
and (n5348,n5349,n5350);
xor (n5349,n5171,n5172);
and (n5350,n257,n619);
and (n5351,n5352,n5353);
xor (n5352,n5349,n5350);
or (n5353,n5354,n5357);
and (n5354,n5355,n5356);
xor (n5355,n5177,n5178);
and (n5356,n250,n619);
and (n5357,n5358,n5359);
xor (n5358,n5355,n5356);
or (n5359,n5360,n5363);
and (n5360,n5361,n5362);
xor (n5361,n5183,n5184);
and (n5362,n315,n619);
and (n5363,n5364,n5365);
xor (n5364,n5361,n5362);
or (n5365,n5366,n5369);
and (n5366,n5367,n5368);
xor (n5367,n5189,n5190);
and (n5368,n308,n619);
and (n5369,n5370,n5371);
xor (n5370,n5367,n5368);
or (n5371,n5372,n5375);
and (n5372,n5373,n5374);
xor (n5373,n5194,n5195);
and (n5374,n51,n619);
and (n5375,n5376,n5377);
xor (n5376,n5373,n5374);
or (n5377,n5378,n5381);
and (n5378,n5379,n5380);
xor (n5379,n5200,n5201);
and (n5380,n45,n619);
and (n5381,n5382,n5383);
xor (n5382,n5379,n5380);
or (n5383,n5384,n5387);
and (n5384,n5385,n5386);
xor (n5385,n5206,n5207);
and (n5386,n75,n619);
and (n5387,n5388,n5389);
xor (n5388,n5385,n5386);
or (n5389,n5390,n5393);
and (n5390,n5391,n5392);
xor (n5391,n5212,n5213);
and (n5392,n69,n619);
and (n5393,n5394,n5395);
xor (n5394,n5391,n5392);
or (n5395,n5396,n5399);
and (n5396,n5397,n5398);
xor (n5397,n5218,n5219);
and (n5398,n226,n619);
and (n5399,n5400,n5401);
xor (n5400,n5397,n5398);
or (n5401,n5402,n5405);
and (n5402,n5403,n5404);
xor (n5403,n5224,n5225);
and (n5404,n351,n619);
and (n5405,n5406,n5407);
xor (n5406,n5403,n5404);
or (n5407,n5408,n5411);
and (n5408,n5409,n5410);
xor (n5409,n5230,n5231);
and (n5410,n345,n619);
and (n5411,n5412,n5413);
xor (n5412,n5409,n5410);
or (n5413,n5414,n5417);
and (n5414,n5415,n5416);
xor (n5415,n5236,n5237);
and (n5416,n372,n619);
and (n5417,n5418,n5419);
xor (n5418,n5415,n5416);
or (n5419,n5420,n5423);
and (n5420,n5421,n5422);
xor (n5421,n5242,n5243);
and (n5422,n281,n619);
and (n5423,n5424,n5425);
xor (n5424,n5421,n5422);
or (n5425,n5426,n5429);
and (n5426,n5427,n5428);
xor (n5427,n5248,n5249);
and (n5428,n185,n619);
and (n5429,n5430,n5431);
xor (n5430,n5427,n5428);
or (n5431,n5432,n5435);
and (n5432,n5433,n5434);
xor (n5433,n5254,n5255);
and (n5434,n179,n619);
and (n5435,n5436,n5437);
xor (n5436,n5433,n5434);
or (n5437,n5438,n5441);
and (n5438,n5439,n5440);
xor (n5439,n5260,n5261);
and (n5440,n289,n619);
and (n5441,n5442,n5443);
xor (n5442,n5439,n5440);
or (n5443,n5444,n5447);
and (n5444,n5445,n5446);
xor (n5445,n5266,n5267);
and (n5446,n545,n619);
and (n5447,n5448,n5449);
xor (n5448,n5445,n5446);
or (n5449,n5450,n5453);
and (n5450,n5451,n5452);
xor (n5451,n5272,n5273);
and (n5452,n719,n619);
and (n5453,n5454,n5455);
xor (n5454,n5451,n5452);
or (n5455,n5456,n5459);
and (n5456,n5457,n5458);
xor (n5457,n5278,n5279);
and (n5458,n837,n619);
and (n5459,n5460,n5461);
xor (n5460,n5457,n5458);
or (n5461,n5462,n5465);
and (n5462,n5463,n5464);
xor (n5463,n5283,n5284);
and (n5464,n1175,n619);
and (n5465,n5466,n5467);
xor (n5466,n5463,n5464);
or (n5467,n5468,n5471);
and (n5468,n5469,n5470);
xor (n5469,n5288,n5289);
and (n5470,n1147,n619);
and (n5471,n5472,n5473);
xor (n5472,n5469,n5470);
or (n5473,n5474,n5477);
and (n5474,n5475,n5476);
xor (n5475,n5293,n5294);
and (n5476,n1141,n619);
and (n5477,n5478,n5479);
xor (n5478,n5475,n5476);
and (n5479,n5480,n4199);
xor (n5480,n5298,n5299);
and (n5481,n126,n515);
and (n5482,n5483,n5484);
xor (n5483,n4762,n5481);
or (n5484,n5485,n5487);
and (n5485,n5486,n922);
xor (n5486,n5304,n5305);
and (n5487,n5488,n5489);
xor (n5488,n5486,n922);
or (n5489,n5490,n5493);
and (n5490,n5491,n5492);
xor (n5491,n5310,n5311);
and (n5492,n324,n515);
and (n5493,n5494,n5495);
xor (n5494,n5491,n5492);
or (n5495,n5496,n5499);
and (n5496,n5497,n5498);
xor (n5497,n5316,n5317);
and (n5498,n158,n515);
and (n5499,n5500,n5501);
xor (n5500,n5497,n5498);
or (n5501,n5502,n5505);
and (n5502,n5503,n5504);
xor (n5503,n5322,n5323);
and (n5504,n151,n515);
and (n5505,n5506,n5507);
xor (n5506,n5503,n5504);
or (n5507,n5508,n5511);
and (n5508,n5509,n5510);
xor (n5509,n5328,n5329);
and (n5510,n195,n515);
and (n5511,n5512,n5513);
xor (n5512,n5509,n5510);
or (n5513,n5514,n5517);
and (n5514,n5515,n5516);
xor (n5515,n5334,n5335);
and (n5516,n103,n515);
and (n5517,n5518,n5519);
xor (n5518,n5515,n5516);
or (n5519,n5520,n5523);
and (n5520,n5521,n5522);
xor (n5521,n5340,n5341);
and (n5522,n97,n515);
and (n5523,n5524,n5525);
xor (n5524,n5521,n5522);
or (n5525,n5526,n5529);
and (n5526,n5527,n5528);
xor (n5527,n5346,n5347);
and (n5528,n257,n515);
and (n5529,n5530,n5531);
xor (n5530,n5527,n5528);
or (n5531,n5532,n5535);
and (n5532,n5533,n5534);
xor (n5533,n5352,n5353);
and (n5534,n250,n515);
and (n5535,n5536,n5537);
xor (n5536,n5533,n5534);
or (n5537,n5538,n5541);
and (n5538,n5539,n5540);
xor (n5539,n5358,n5359);
and (n5540,n315,n515);
and (n5541,n5542,n5543);
xor (n5542,n5539,n5540);
or (n5543,n5544,n5547);
and (n5544,n5545,n5546);
xor (n5545,n5364,n5365);
and (n5546,n308,n515);
and (n5547,n5548,n5549);
xor (n5548,n5545,n5546);
or (n5549,n5550,n5552);
and (n5550,n5551,n3637);
xor (n5551,n5370,n5371);
and (n5552,n5553,n5554);
xor (n5553,n5551,n3637);
or (n5554,n5555,n5557);
and (n5555,n5556,n3070);
xor (n5556,n5376,n5377);
and (n5557,n5558,n5559);
xor (n5558,n5556,n3070);
or (n5559,n5560,n5563);
and (n5560,n5561,n5562);
xor (n5561,n5382,n5383);
and (n5562,n75,n515);
and (n5563,n5564,n5565);
xor (n5564,n5561,n5562);
or (n5565,n5566,n5569);
and (n5566,n5567,n5568);
xor (n5567,n5388,n5389);
and (n5568,n69,n515);
and (n5569,n5570,n5571);
xor (n5570,n5567,n5568);
or (n5571,n5572,n5575);
and (n5572,n5573,n5574);
xor (n5573,n5394,n5395);
and (n5574,n226,n515);
and (n5575,n5576,n5577);
xor (n5576,n5573,n5574);
or (n5577,n5578,n5581);
and (n5578,n5579,n5580);
xor (n5579,n5400,n5401);
and (n5580,n351,n515);
and (n5581,n5582,n5583);
xor (n5582,n5579,n5580);
or (n5583,n5584,n5587);
and (n5584,n5585,n5586);
xor (n5585,n5406,n5407);
and (n5586,n345,n515);
and (n5587,n5588,n5589);
xor (n5588,n5585,n5586);
or (n5589,n5590,n5593);
and (n5590,n5591,n5592);
xor (n5591,n5412,n5413);
and (n5592,n372,n515);
and (n5593,n5594,n5595);
xor (n5594,n5591,n5592);
or (n5595,n5596,n5599);
and (n5596,n5597,n5598);
xor (n5597,n5418,n5419);
and (n5598,n281,n515);
and (n5599,n5600,n5601);
xor (n5600,n5597,n5598);
or (n5601,n5602,n5605);
and (n5602,n5603,n5604);
xor (n5603,n5424,n5425);
and (n5604,n185,n515);
and (n5605,n5606,n5607);
xor (n5606,n5603,n5604);
or (n5607,n5608,n5611);
and (n5608,n5609,n5610);
xor (n5609,n5430,n5431);
and (n5610,n179,n515);
and (n5611,n5612,n5613);
xor (n5612,n5609,n5610);
or (n5613,n5614,n5617);
and (n5614,n5615,n5616);
xor (n5615,n5436,n5437);
and (n5616,n289,n515);
and (n5617,n5618,n5619);
xor (n5618,n5615,n5616);
or (n5619,n5620,n5623);
and (n5620,n5621,n5622);
xor (n5621,n5442,n5443);
and (n5622,n545,n515);
and (n5623,n5624,n5625);
xor (n5624,n5621,n5622);
or (n5625,n5626,n5629);
and (n5626,n5627,n5628);
xor (n5627,n5448,n5449);
and (n5628,n719,n515);
and (n5629,n5630,n5631);
xor (n5630,n5627,n5628);
or (n5631,n5632,n5635);
and (n5632,n5633,n5634);
xor (n5633,n5454,n5455);
and (n5634,n837,n515);
and (n5635,n5636,n5637);
xor (n5636,n5633,n5634);
or (n5637,n5638,n5641);
and (n5638,n5639,n5640);
xor (n5639,n5460,n5461);
and (n5640,n1175,n515);
and (n5641,n5642,n5643);
xor (n5642,n5639,n5640);
or (n5643,n5644,n5646);
and (n5644,n5645,n4137);
xor (n5645,n5466,n5467);
and (n5646,n5647,n5648);
xor (n5647,n5645,n4137);
or (n5648,n5649,n5651);
and (n5649,n5650,n4192);
xor (n5650,n5472,n5473);
and (n5651,n5652,n5653);
xor (n5652,n5650,n4192);
and (n5653,n5654,n5655);
xor (n5654,n5478,n5479);
and (n5655,n1187,n515);
and (n5656,n126,n513);
and (n5657,n5658,n5659);
xor (n5658,n4759,n5656);
or (n5659,n5660,n5663);
and (n5660,n5661,n5662);
xor (n5661,n5483,n5484);
and (n5662,n329,n513);
and (n5663,n5664,n5665);
xor (n5664,n5661,n5662);
or (n5665,n5666,n5669);
and (n5666,n5667,n5668);
xor (n5667,n5488,n5489);
and (n5668,n324,n513);
and (n5669,n5670,n5671);
xor (n5670,n5667,n5668);
or (n5671,n5672,n5675);
and (n5672,n5673,n5674);
xor (n5673,n5494,n5495);
and (n5674,n158,n513);
and (n5675,n5676,n5677);
xor (n5676,n5673,n5674);
or (n5677,n5678,n5681);
and (n5678,n5679,n5680);
xor (n5679,n5500,n5501);
and (n5680,n151,n513);
and (n5681,n5682,n5683);
xor (n5682,n5679,n5680);
or (n5683,n5684,n5687);
and (n5684,n5685,n5686);
xor (n5685,n5506,n5507);
and (n5686,n195,n513);
and (n5687,n5688,n5689);
xor (n5688,n5685,n5686);
or (n5689,n5690,n5693);
and (n5690,n5691,n5692);
xor (n5691,n5512,n5513);
and (n5692,n103,n513);
and (n5693,n5694,n5695);
xor (n5694,n5691,n5692);
or (n5695,n5696,n5699);
and (n5696,n5697,n5698);
xor (n5697,n5518,n5519);
and (n5698,n97,n513);
and (n5699,n5700,n5701);
xor (n5700,n5697,n5698);
or (n5701,n5702,n5705);
and (n5702,n5703,n5704);
xor (n5703,n5524,n5525);
and (n5704,n257,n513);
and (n5705,n5706,n5707);
xor (n5706,n5703,n5704);
or (n5707,n5708,n5711);
and (n5708,n5709,n5710);
xor (n5709,n5530,n5531);
and (n5710,n250,n513);
and (n5711,n5712,n5713);
xor (n5712,n5709,n5710);
or (n5713,n5714,n5717);
and (n5714,n5715,n5716);
xor (n5715,n5536,n5537);
and (n5716,n315,n513);
and (n5717,n5718,n5719);
xor (n5718,n5715,n5716);
or (n5719,n5720,n5723);
and (n5720,n5721,n5722);
xor (n5721,n5542,n5543);
and (n5722,n308,n513);
and (n5723,n5724,n5725);
xor (n5724,n5721,n5722);
or (n5725,n5726,n5729);
and (n5726,n5727,n5728);
xor (n5727,n5548,n5549);
and (n5728,n51,n513);
and (n5729,n5730,n5731);
xor (n5730,n5727,n5728);
or (n5731,n5732,n5735);
and (n5732,n5733,n5734);
xor (n5733,n5553,n5554);
and (n5734,n45,n513);
and (n5735,n5736,n5737);
xor (n5736,n5733,n5734);
or (n5737,n5738,n5741);
and (n5738,n5739,n5740);
xor (n5739,n5558,n5559);
and (n5740,n75,n513);
and (n5741,n5742,n5743);
xor (n5742,n5739,n5740);
or (n5743,n5744,n5747);
and (n5744,n5745,n5746);
xor (n5745,n5564,n5565);
and (n5746,n69,n513);
and (n5747,n5748,n5749);
xor (n5748,n5745,n5746);
or (n5749,n5750,n5753);
and (n5750,n5751,n5752);
xor (n5751,n5570,n5571);
and (n5752,n226,n513);
and (n5753,n5754,n5755);
xor (n5754,n5751,n5752);
or (n5755,n5756,n5759);
and (n5756,n5757,n5758);
xor (n5757,n5576,n5577);
and (n5758,n351,n513);
and (n5759,n5760,n5761);
xor (n5760,n5757,n5758);
or (n5761,n5762,n5765);
and (n5762,n5763,n5764);
xor (n5763,n5582,n5583);
and (n5764,n345,n513);
and (n5765,n5766,n5767);
xor (n5766,n5763,n5764);
or (n5767,n5768,n5771);
and (n5768,n5769,n5770);
xor (n5769,n5588,n5589);
and (n5770,n372,n513);
and (n5771,n5772,n5773);
xor (n5772,n5769,n5770);
or (n5773,n5774,n5777);
and (n5774,n5775,n5776);
xor (n5775,n5594,n5595);
and (n5776,n281,n513);
and (n5777,n5778,n5779);
xor (n5778,n5775,n5776);
or (n5779,n5780,n5783);
and (n5780,n5781,n5782);
xor (n5781,n5600,n5601);
and (n5782,n185,n513);
and (n5783,n5784,n5785);
xor (n5784,n5781,n5782);
or (n5785,n5786,n5789);
and (n5786,n5787,n5788);
xor (n5787,n5606,n5607);
and (n5788,n179,n513);
and (n5789,n5790,n5791);
xor (n5790,n5787,n5788);
or (n5791,n5792,n5795);
and (n5792,n5793,n5794);
xor (n5793,n5612,n5613);
and (n5794,n289,n513);
and (n5795,n5796,n5797);
xor (n5796,n5793,n5794);
or (n5797,n5798,n5801);
and (n5798,n5799,n5800);
xor (n5799,n5618,n5619);
and (n5800,n545,n513);
and (n5801,n5802,n5803);
xor (n5802,n5799,n5800);
or (n5803,n5804,n5807);
and (n5804,n5805,n5806);
xor (n5805,n5624,n5625);
and (n5806,n719,n513);
and (n5807,n5808,n5809);
xor (n5808,n5805,n5806);
or (n5809,n5810,n5813);
and (n5810,n5811,n5812);
xor (n5811,n5630,n5631);
and (n5812,n837,n513);
and (n5813,n5814,n5815);
xor (n5814,n5811,n5812);
or (n5815,n5816,n5819);
and (n5816,n5817,n5818);
xor (n5817,n5636,n5637);
and (n5818,n1175,n513);
and (n5819,n5820,n5821);
xor (n5820,n5817,n5818);
or (n5821,n5822,n5825);
and (n5822,n5823,n5824);
xor (n5823,n5642,n5643);
and (n5824,n1147,n513);
and (n5825,n5826,n5827);
xor (n5826,n5823,n5824);
or (n5827,n5828,n5831);
and (n5828,n5829,n5830);
xor (n5829,n5647,n5648);
and (n5830,n1141,n513);
and (n5831,n5832,n5833);
xor (n5832,n5829,n5830);
and (n5833,n5834,n4096);
xor (n5834,n5652,n5653);
and (n5835,n126,n115);
and (n5836,n5837,n5838);
xor (n5837,n4756,n5835);
or (n5838,n5839,n5842);
and (n5839,n5840,n5841);
xor (n5840,n5658,n5659);
and (n5841,n329,n115);
and (n5842,n5843,n5844);
xor (n5843,n5840,n5841);
or (n5844,n5845,n5848);
and (n5845,n5846,n5847);
xor (n5846,n5664,n5665);
and (n5847,n324,n115);
and (n5848,n5849,n5850);
xor (n5849,n5846,n5847);
or (n5850,n5851,n5854);
and (n5851,n5852,n5853);
xor (n5852,n5670,n5671);
and (n5853,n158,n115);
and (n5854,n5855,n5856);
xor (n5855,n5852,n5853);
or (n5856,n5857,n5860);
and (n5857,n5858,n5859);
xor (n5858,n5676,n5677);
and (n5859,n151,n115);
and (n5860,n5861,n5862);
xor (n5861,n5858,n5859);
or (n5862,n5863,n5866);
and (n5863,n5864,n5865);
xor (n5864,n5682,n5683);
and (n5865,n195,n115);
and (n5866,n5867,n5868);
xor (n5867,n5864,n5865);
or (n5868,n5869,n5872);
and (n5869,n5870,n5871);
xor (n5870,n5688,n5689);
and (n5871,n103,n115);
and (n5872,n5873,n5874);
xor (n5873,n5870,n5871);
or (n5874,n5875,n5878);
and (n5875,n5876,n5877);
xor (n5876,n5694,n5695);
and (n5877,n97,n115);
and (n5878,n5879,n5880);
xor (n5879,n5876,n5877);
or (n5880,n5881,n5884);
and (n5881,n5882,n5883);
xor (n5882,n5700,n5701);
and (n5883,n257,n115);
and (n5884,n5885,n5886);
xor (n5885,n5882,n5883);
or (n5886,n5887,n5890);
and (n5887,n5888,n5889);
xor (n5888,n5706,n5707);
and (n5889,n250,n115);
and (n5890,n5891,n5892);
xor (n5891,n5888,n5889);
or (n5892,n5893,n5896);
and (n5893,n5894,n5895);
xor (n5894,n5712,n5713);
and (n5895,n315,n115);
and (n5896,n5897,n5898);
xor (n5897,n5894,n5895);
or (n5898,n5899,n5902);
and (n5899,n5900,n5901);
xor (n5900,n5718,n5719);
and (n5901,n308,n115);
and (n5902,n5903,n5904);
xor (n5903,n5900,n5901);
or (n5904,n5905,n5908);
and (n5905,n5906,n5907);
xor (n5906,n5724,n5725);
and (n5907,n51,n115);
and (n5908,n5909,n5910);
xor (n5909,n5906,n5907);
or (n5910,n5911,n5914);
and (n5911,n5912,n5913);
xor (n5912,n5730,n5731);
and (n5913,n45,n115);
and (n5914,n5915,n5916);
xor (n5915,n5912,n5913);
or (n5916,n5917,n5920);
and (n5917,n5918,n5919);
xor (n5918,n5736,n5737);
and (n5919,n75,n115);
and (n5920,n5921,n5922);
xor (n5921,n5918,n5919);
or (n5922,n5923,n5925);
and (n5923,n5924,n2955);
xor (n5924,n5742,n5743);
and (n5925,n5926,n5927);
xor (n5926,n5924,n2955);
or (n5927,n5928,n5930);
and (n5928,n5929,n2891);
xor (n5929,n5748,n5749);
and (n5930,n5931,n5932);
xor (n5931,n5929,n2891);
or (n5932,n5933,n5935);
and (n5933,n5934,n2856);
xor (n5934,n5754,n5755);
and (n5935,n5936,n5937);
xor (n5936,n5934,n2856);
or (n5937,n5938,n5940);
and (n5938,n5939,n2760);
xor (n5939,n5760,n5761);
and (n5940,n5941,n5942);
xor (n5941,n5939,n2760);
or (n5942,n5943,n5946);
and (n5943,n5944,n5945);
xor (n5944,n5766,n5767);
and (n5945,n372,n115);
and (n5946,n5947,n5948);
xor (n5947,n5944,n5945);
or (n5948,n5949,n5952);
and (n5949,n5950,n5951);
xor (n5950,n5772,n5773);
and (n5951,n281,n115);
and (n5952,n5953,n5954);
xor (n5953,n5950,n5951);
or (n5954,n5955,n5958);
and (n5955,n5956,n5957);
xor (n5956,n5778,n5779);
and (n5957,n185,n115);
and (n5958,n5959,n5960);
xor (n5959,n5956,n5957);
or (n5960,n5961,n5964);
and (n5961,n5962,n5963);
xor (n5962,n5784,n5785);
and (n5963,n179,n115);
and (n5964,n5965,n5966);
xor (n5965,n5962,n5963);
or (n5966,n5967,n5969);
and (n5967,n5968,n3393);
xor (n5968,n5790,n5791);
and (n5969,n5970,n5971);
xor (n5970,n5968,n3393);
or (n5971,n5972,n5975);
and (n5972,n5973,n5974);
xor (n5973,n5796,n5797);
and (n5974,n545,n115);
and (n5975,n5976,n5977);
xor (n5976,n5973,n5974);
or (n5977,n5978,n5981);
and (n5978,n5979,n5980);
xor (n5979,n5802,n5803);
and (n5980,n719,n115);
and (n5981,n5982,n5983);
xor (n5982,n5979,n5980);
or (n5983,n5984,n5987);
and (n5984,n5985,n5986);
xor (n5985,n5808,n5809);
and (n5986,n837,n115);
and (n5987,n5988,n5989);
xor (n5988,n5985,n5986);
or (n5989,n5990,n5993);
and (n5990,n5991,n5992);
xor (n5991,n5814,n5815);
and (n5992,n1175,n115);
and (n5993,n5994,n5995);
xor (n5994,n5991,n5992);
or (n5995,n5996,n5999);
and (n5996,n5997,n5998);
xor (n5997,n5820,n5821);
and (n5998,n1147,n115);
and (n5999,n6000,n6001);
xor (n6000,n5997,n5998);
or (n6001,n6002,n6004);
and (n6002,n6003,n3966);
xor (n6003,n5826,n5827);
and (n6004,n6005,n6006);
xor (n6005,n6003,n3966);
and (n6006,n6007,n6008);
xor (n6007,n5832,n5833);
and (n6008,n1187,n115);
and (n6009,n126,n117);
and (n6010,n6011,n6012);
xor (n6011,n4753,n6009);
or (n6012,n6013,n6016);
and (n6013,n6014,n6015);
xor (n6014,n5837,n5838);
and (n6015,n329,n117);
and (n6016,n6017,n6018);
xor (n6017,n6014,n6015);
or (n6018,n6019,n6022);
and (n6019,n6020,n6021);
xor (n6020,n5843,n5844);
and (n6021,n324,n117);
and (n6022,n6023,n6024);
xor (n6023,n6020,n6021);
or (n6024,n6025,n6028);
and (n6025,n6026,n6027);
xor (n6026,n5849,n5850);
and (n6027,n158,n117);
and (n6028,n6029,n6030);
xor (n6029,n6026,n6027);
or (n6030,n6031,n6034);
and (n6031,n6032,n6033);
xor (n6032,n5855,n5856);
and (n6033,n151,n117);
and (n6034,n6035,n6036);
xor (n6035,n6032,n6033);
or (n6036,n6037,n6040);
and (n6037,n6038,n6039);
xor (n6038,n5861,n5862);
and (n6039,n195,n117);
and (n6040,n6041,n6042);
xor (n6041,n6038,n6039);
or (n6042,n6043,n6046);
and (n6043,n6044,n6045);
xor (n6044,n5867,n5868);
and (n6045,n103,n117);
and (n6046,n6047,n6048);
xor (n6047,n6044,n6045);
or (n6048,n6049,n6052);
and (n6049,n6050,n6051);
xor (n6050,n5873,n5874);
and (n6051,n97,n117);
and (n6052,n6053,n6054);
xor (n6053,n6050,n6051);
or (n6054,n6055,n6058);
and (n6055,n6056,n6057);
xor (n6056,n5879,n5880);
and (n6057,n257,n117);
and (n6058,n6059,n6060);
xor (n6059,n6056,n6057);
or (n6060,n6061,n6064);
and (n6061,n6062,n6063);
xor (n6062,n5885,n5886);
and (n6063,n250,n117);
and (n6064,n6065,n6066);
xor (n6065,n6062,n6063);
or (n6066,n6067,n6070);
and (n6067,n6068,n6069);
xor (n6068,n5891,n5892);
and (n6069,n315,n117);
and (n6070,n6071,n6072);
xor (n6071,n6068,n6069);
or (n6072,n6073,n6076);
and (n6073,n6074,n6075);
xor (n6074,n5897,n5898);
and (n6075,n308,n117);
and (n6076,n6077,n6078);
xor (n6077,n6074,n6075);
or (n6078,n6079,n6082);
and (n6079,n6080,n6081);
xor (n6080,n5903,n5904);
and (n6081,n51,n117);
and (n6082,n6083,n6084);
xor (n6083,n6080,n6081);
or (n6084,n6085,n6088);
and (n6085,n6086,n6087);
xor (n6086,n5909,n5910);
and (n6087,n45,n117);
and (n6088,n6089,n6090);
xor (n6089,n6086,n6087);
or (n6090,n6091,n6094);
and (n6091,n6092,n6093);
xor (n6092,n5915,n5916);
and (n6093,n75,n117);
and (n6094,n6095,n6096);
xor (n6095,n6092,n6093);
or (n6096,n6097,n6100);
and (n6097,n6098,n6099);
xor (n6098,n5921,n5922);
and (n6099,n69,n117);
and (n6100,n6101,n6102);
xor (n6101,n6098,n6099);
or (n6102,n6103,n6106);
and (n6103,n6104,n6105);
xor (n6104,n5926,n5927);
and (n6105,n226,n117);
and (n6106,n6107,n6108);
xor (n6107,n6104,n6105);
or (n6108,n6109,n6112);
and (n6109,n6110,n6111);
xor (n6110,n5931,n5932);
and (n6111,n351,n117);
and (n6112,n6113,n6114);
xor (n6113,n6110,n6111);
or (n6114,n6115,n6118);
and (n6115,n6116,n6117);
xor (n6116,n5936,n5937);
and (n6117,n345,n117);
and (n6118,n6119,n6120);
xor (n6119,n6116,n6117);
or (n6120,n6121,n6124);
and (n6121,n6122,n6123);
xor (n6122,n5941,n5942);
and (n6123,n372,n117);
and (n6124,n6125,n6126);
xor (n6125,n6122,n6123);
or (n6126,n6127,n6130);
and (n6127,n6128,n6129);
xor (n6128,n5947,n5948);
and (n6129,n281,n117);
and (n6130,n6131,n6132);
xor (n6131,n6128,n6129);
or (n6132,n6133,n6136);
and (n6133,n6134,n6135);
xor (n6134,n5953,n5954);
and (n6135,n185,n117);
and (n6136,n6137,n6138);
xor (n6137,n6134,n6135);
or (n6138,n6139,n6142);
and (n6139,n6140,n6141);
xor (n6140,n5959,n5960);
and (n6141,n179,n117);
and (n6142,n6143,n6144);
xor (n6143,n6140,n6141);
or (n6144,n6145,n6148);
and (n6145,n6146,n6147);
xor (n6146,n5965,n5966);
and (n6147,n289,n117);
and (n6148,n6149,n6150);
xor (n6149,n6146,n6147);
or (n6150,n6151,n6154);
and (n6151,n6152,n6153);
xor (n6152,n5970,n5971);
and (n6153,n545,n117);
and (n6154,n6155,n6156);
xor (n6155,n6152,n6153);
or (n6156,n6157,n6160);
and (n6157,n6158,n6159);
xor (n6158,n5976,n5977);
and (n6159,n719,n117);
and (n6160,n6161,n6162);
xor (n6161,n6158,n6159);
or (n6162,n6163,n6166);
and (n6163,n6164,n6165);
xor (n6164,n5982,n5983);
and (n6165,n837,n117);
and (n6166,n6167,n6168);
xor (n6167,n6164,n6165);
or (n6168,n6169,n6172);
and (n6169,n6170,n6171);
xor (n6170,n5988,n5989);
and (n6171,n1175,n117);
and (n6172,n6173,n6174);
xor (n6173,n6170,n6171);
or (n6174,n6175,n6178);
and (n6175,n6176,n6177);
xor (n6176,n5994,n5995);
and (n6177,n1147,n117);
and (n6178,n6179,n6180);
xor (n6179,n6176,n6177);
or (n6180,n6181,n6184);
and (n6181,n6182,n6183);
xor (n6182,n6000,n6001);
and (n6183,n1141,n117);
and (n6184,n6185,n6186);
xor (n6185,n6182,n6183);
and (n6186,n6187,n3939);
xor (n6187,n6005,n6006);
and (n6188,n126,n121);
and (n6189,n6190,n6191);
xor (n6190,n4750,n6188);
or (n6191,n6192,n6195);
and (n6192,n6193,n6194);
xor (n6193,n6011,n6012);
and (n6194,n329,n121);
and (n6195,n6196,n6197);
xor (n6196,n6193,n6194);
or (n6197,n6198,n6201);
and (n6198,n6199,n6200);
xor (n6199,n6017,n6018);
and (n6200,n324,n121);
and (n6201,n6202,n6203);
xor (n6202,n6199,n6200);
or (n6203,n6204,n6207);
and (n6204,n6205,n6206);
xor (n6205,n6023,n6024);
and (n6206,n158,n121);
and (n6207,n6208,n6209);
xor (n6208,n6205,n6206);
or (n6209,n6210,n6213);
and (n6210,n6211,n6212);
xor (n6211,n6029,n6030);
and (n6212,n151,n121);
and (n6213,n6214,n6215);
xor (n6214,n6211,n6212);
or (n6215,n6216,n6219);
and (n6216,n6217,n6218);
xor (n6217,n6035,n6036);
and (n6218,n195,n121);
and (n6219,n6220,n6221);
xor (n6220,n6217,n6218);
or (n6221,n6222,n6225);
and (n6222,n6223,n6224);
xor (n6223,n6041,n6042);
and (n6224,n103,n121);
and (n6225,n6226,n6227);
xor (n6226,n6223,n6224);
or (n6227,n6228,n6231);
and (n6228,n6229,n6230);
xor (n6229,n6047,n6048);
and (n6230,n97,n121);
and (n6231,n6232,n6233);
xor (n6232,n6229,n6230);
or (n6233,n6234,n6237);
and (n6234,n6235,n6236);
xor (n6235,n6053,n6054);
and (n6236,n257,n121);
and (n6237,n6238,n6239);
xor (n6238,n6235,n6236);
or (n6239,n6240,n6242);
and (n6240,n6241,n1214);
xor (n6241,n6059,n6060);
and (n6242,n6243,n6244);
xor (n6243,n6241,n1214);
or (n6244,n6245,n6248);
and (n6245,n6246,n6247);
xor (n6246,n6065,n6066);
and (n6247,n315,n121);
and (n6248,n6249,n6250);
xor (n6249,n6246,n6247);
or (n6250,n6251,n6254);
and (n6251,n6252,n6253);
xor (n6252,n6071,n6072);
and (n6253,n308,n121);
and (n6254,n6255,n6256);
xor (n6255,n6252,n6253);
or (n6256,n6257,n6260);
and (n6257,n6258,n6259);
xor (n6258,n6077,n6078);
and (n6259,n51,n121);
and (n6260,n6261,n6262);
xor (n6261,n6258,n6259);
or (n6262,n6263,n6266);
and (n6263,n6264,n6265);
xor (n6264,n6083,n6084);
and (n6265,n45,n121);
and (n6266,n6267,n6268);
xor (n6267,n6264,n6265);
or (n6268,n6269,n6272);
and (n6269,n6270,n6271);
xor (n6270,n6089,n6090);
and (n6271,n75,n121);
and (n6272,n6273,n6274);
xor (n6273,n6270,n6271);
or (n6274,n6275,n6278);
and (n6275,n6276,n6277);
xor (n6276,n6095,n6096);
and (n6277,n69,n121);
and (n6278,n6279,n6280);
xor (n6279,n6276,n6277);
or (n6280,n6281,n6284);
and (n6281,n6282,n6283);
xor (n6282,n6101,n6102);
and (n6283,n226,n121);
and (n6284,n6285,n6286);
xor (n6285,n6282,n6283);
or (n6286,n6287,n6290);
and (n6287,n6288,n6289);
xor (n6288,n6107,n6108);
and (n6289,n351,n121);
and (n6290,n6291,n6292);
xor (n6291,n6288,n6289);
or (n6292,n6293,n6296);
and (n6293,n6294,n6295);
xor (n6294,n6113,n6114);
and (n6295,n345,n121);
and (n6296,n6297,n6298);
xor (n6297,n6294,n6295);
or (n6298,n6299,n6302);
and (n6299,n6300,n6301);
xor (n6300,n6119,n6120);
and (n6301,n372,n121);
and (n6302,n6303,n6304);
xor (n6303,n6300,n6301);
or (n6304,n6305,n6307);
and (n6305,n6306,n2810);
xor (n6306,n6125,n6126);
and (n6307,n6308,n6309);
xor (n6308,n6306,n2810);
or (n6309,n6310,n6313);
and (n6310,n6311,n6312);
xor (n6311,n6131,n6132);
and (n6312,n185,n121);
and (n6313,n6314,n6315);
xor (n6314,n6311,n6312);
or (n6315,n6316,n6319);
and (n6316,n6317,n6318);
xor (n6317,n6137,n6138);
and (n6318,n179,n121);
and (n6319,n6320,n6321);
xor (n6320,n6317,n6318);
or (n6321,n6322,n6325);
and (n6322,n6323,n6324);
xor (n6323,n6143,n6144);
and (n6324,n289,n121);
and (n6325,n6326,n6327);
xor (n6326,n6323,n6324);
or (n6327,n6328,n6331);
and (n6328,n6329,n6330);
xor (n6329,n6149,n6150);
and (n6330,n545,n121);
and (n6331,n6332,n6333);
xor (n6332,n6329,n6330);
or (n6333,n6334,n6337);
and (n6334,n6335,n6336);
xor (n6335,n6155,n6156);
and (n6336,n719,n121);
and (n6337,n6338,n6339);
xor (n6338,n6335,n6336);
or (n6339,n6340,n6343);
and (n6340,n6341,n6342);
xor (n6341,n6161,n6162);
and (n6342,n837,n121);
and (n6343,n6344,n6345);
xor (n6344,n6341,n6342);
or (n6345,n6346,n6349);
and (n6346,n6347,n6348);
xor (n6347,n6167,n6168);
and (n6348,n1175,n121);
and (n6349,n6350,n6351);
xor (n6350,n6347,n6348);
or (n6351,n6352,n6355);
and (n6352,n6353,n6354);
xor (n6353,n6173,n6174);
and (n6354,n1147,n121);
and (n6355,n6356,n6357);
xor (n6356,n6353,n6354);
or (n6357,n6358,n6361);
and (n6358,n6359,n6360);
xor (n6359,n6179,n6180);
and (n6360,n1141,n121);
and (n6361,n6362,n6363);
xor (n6362,n6359,n6360);
and (n6363,n6364,n6365);
xor (n6364,n6185,n6186);
and (n6365,n1187,n121);
and (n6366,n126,n483);
or (n6367,n6368,n6371);
and (n6368,n6369,n6370);
xor (n6369,n6190,n6191);
and (n6370,n329,n483);
and (n6371,n6372,n6373);
xor (n6372,n6369,n6370);
or (n6373,n6374,n6377);
and (n6374,n6375,n6376);
xor (n6375,n6196,n6197);
and (n6376,n324,n483);
and (n6377,n6378,n6379);
xor (n6378,n6375,n6376);
or (n6379,n6380,n6383);
and (n6380,n6381,n6382);
xor (n6381,n6202,n6203);
and (n6382,n158,n483);
and (n6383,n6384,n6385);
xor (n6384,n6381,n6382);
or (n6385,n6386,n6389);
and (n6386,n6387,n6388);
xor (n6387,n6208,n6209);
and (n6388,n151,n483);
and (n6389,n6390,n6391);
xor (n6390,n6387,n6388);
or (n6391,n6392,n6395);
and (n6392,n6393,n6394);
xor (n6393,n6214,n6215);
and (n6394,n195,n483);
and (n6395,n6396,n6397);
xor (n6396,n6393,n6394);
or (n6397,n6398,n6401);
and (n6398,n6399,n6400);
xor (n6399,n6220,n6221);
and (n6400,n103,n483);
and (n6401,n6402,n6403);
xor (n6402,n6399,n6400);
or (n6403,n6404,n6407);
and (n6404,n6405,n6406);
xor (n6405,n6226,n6227);
and (n6406,n97,n483);
and (n6407,n6408,n6409);
xor (n6408,n6405,n6406);
or (n6409,n6410,n6413);
and (n6410,n6411,n6412);
xor (n6411,n6232,n6233);
and (n6412,n257,n483);
and (n6413,n6414,n6415);
xor (n6414,n6411,n6412);
or (n6415,n6416,n6419);
and (n6416,n6417,n6418);
xor (n6417,n6238,n6239);
and (n6418,n250,n483);
and (n6419,n6420,n6421);
xor (n6420,n6417,n6418);
or (n6421,n6422,n6425);
and (n6422,n6423,n6424);
xor (n6423,n6243,n6244);
and (n6424,n315,n483);
and (n6425,n6426,n6427);
xor (n6426,n6423,n6424);
or (n6427,n6428,n6431);
and (n6428,n6429,n6430);
xor (n6429,n6249,n6250);
and (n6430,n308,n483);
and (n6431,n6432,n6433);
xor (n6432,n6429,n6430);
or (n6433,n6434,n6437);
and (n6434,n6435,n6436);
xor (n6435,n6255,n6256);
and (n6436,n51,n483);
and (n6437,n6438,n6439);
xor (n6438,n6435,n6436);
or (n6439,n6440,n6443);
and (n6440,n6441,n6442);
xor (n6441,n6261,n6262);
and (n6442,n45,n483);
and (n6443,n6444,n6445);
xor (n6444,n6441,n6442);
or (n6445,n6446,n6449);
and (n6446,n6447,n6448);
xor (n6447,n6267,n6268);
and (n6448,n75,n483);
and (n6449,n6450,n6451);
xor (n6450,n6447,n6448);
or (n6451,n6452,n6455);
and (n6452,n6453,n6454);
xor (n6453,n6273,n6274);
and (n6454,n69,n483);
and (n6455,n6456,n6457);
xor (n6456,n6453,n6454);
or (n6457,n6458,n6461);
and (n6458,n6459,n6460);
xor (n6459,n6279,n6280);
and (n6460,n226,n483);
and (n6461,n6462,n6463);
xor (n6462,n6459,n6460);
or (n6463,n6464,n6467);
and (n6464,n6465,n6466);
xor (n6465,n6285,n6286);
and (n6466,n351,n483);
and (n6467,n6468,n6469);
xor (n6468,n6465,n6466);
or (n6469,n6470,n6473);
and (n6470,n6471,n6472);
xor (n6471,n6291,n6292);
and (n6472,n345,n483);
and (n6473,n6474,n6475);
xor (n6474,n6471,n6472);
or (n6475,n6476,n6479);
and (n6476,n6477,n6478);
xor (n6477,n6297,n6298);
and (n6478,n372,n483);
and (n6479,n6480,n6481);
xor (n6480,n6477,n6478);
or (n6481,n6482,n6485);
and (n6482,n6483,n6484);
xor (n6483,n6303,n6304);
and (n6484,n281,n483);
and (n6485,n6486,n6487);
xor (n6486,n6483,n6484);
or (n6487,n6488,n6491);
and (n6488,n6489,n6490);
xor (n6489,n6308,n6309);
and (n6490,n185,n483);
and (n6491,n6492,n6493);
xor (n6492,n6489,n6490);
or (n6493,n6494,n6497);
and (n6494,n6495,n6496);
xor (n6495,n6314,n6315);
and (n6496,n179,n483);
and (n6497,n6498,n6499);
xor (n6498,n6495,n6496);
or (n6499,n6500,n6503);
and (n6500,n6501,n6502);
xor (n6501,n6320,n6321);
and (n6502,n289,n483);
and (n6503,n6504,n6505);
xor (n6504,n6501,n6502);
or (n6505,n6506,n6509);
and (n6506,n6507,n6508);
xor (n6507,n6326,n6327);
and (n6508,n545,n483);
and (n6509,n6510,n6511);
xor (n6510,n6507,n6508);
or (n6511,n6512,n6515);
and (n6512,n6513,n6514);
xor (n6513,n6332,n6333);
and (n6514,n719,n483);
and (n6515,n6516,n6517);
xor (n6516,n6513,n6514);
or (n6517,n6518,n6521);
and (n6518,n6519,n6520);
xor (n6519,n6338,n6339);
and (n6520,n837,n483);
and (n6521,n6522,n6523);
xor (n6522,n6519,n6520);
or (n6523,n6524,n6527);
and (n6524,n6525,n6526);
xor (n6525,n6344,n6345);
and (n6526,n1175,n483);
and (n6527,n6528,n6529);
xor (n6528,n6525,n6526);
or (n6529,n6530,n6533);
and (n6530,n6531,n6532);
xor (n6531,n6350,n6351);
and (n6532,n1147,n483);
and (n6533,n6534,n6535);
xor (n6534,n6531,n6532);
or (n6535,n6536,n6539);
and (n6536,n6537,n6538);
xor (n6537,n6356,n6357);
and (n6538,n1141,n483);
and (n6539,n6540,n6541);
xor (n6540,n6537,n6538);
and (n6541,n6542,n4039);
xor (n6542,n6362,n6363);
and (n6543,n329,n143);
or (n6544,n6545,n6548);
and (n6545,n6546,n6547);
xor (n6546,n6372,n6373);
and (n6547,n324,n143);
and (n6548,n6549,n6550);
xor (n6549,n6546,n6547);
or (n6550,n6551,n6554);
and (n6551,n6552,n6553);
xor (n6552,n6378,n6379);
and (n6553,n158,n143);
and (n6554,n6555,n6556);
xor (n6555,n6552,n6553);
or (n6556,n6557,n6560);
and (n6557,n6558,n6559);
xor (n6558,n6384,n6385);
and (n6559,n151,n143);
and (n6560,n6561,n6562);
xor (n6561,n6558,n6559);
or (n6562,n6563,n6566);
and (n6563,n6564,n6565);
xor (n6564,n6390,n6391);
and (n6565,n195,n143);
and (n6566,n6567,n6568);
xor (n6567,n6564,n6565);
or (n6568,n6569,n6572);
and (n6569,n6570,n6571);
xor (n6570,n6396,n6397);
and (n6571,n103,n143);
and (n6572,n6573,n6574);
xor (n6573,n6570,n6571);
or (n6574,n6575,n6578);
and (n6575,n6576,n6577);
xor (n6576,n6402,n6403);
and (n6577,n97,n143);
and (n6578,n6579,n6580);
xor (n6579,n6576,n6577);
or (n6580,n6581,n6584);
and (n6581,n6582,n6583);
xor (n6582,n6408,n6409);
and (n6583,n257,n143);
and (n6584,n6585,n6586);
xor (n6585,n6582,n6583);
or (n6586,n6587,n6590);
and (n6587,n6588,n6589);
xor (n6588,n6414,n6415);
and (n6589,n250,n143);
and (n6590,n6591,n6592);
xor (n6591,n6588,n6589);
or (n6592,n6593,n6596);
and (n6593,n6594,n6595);
xor (n6594,n6420,n6421);
and (n6595,n315,n143);
and (n6596,n6597,n6598);
xor (n6597,n6594,n6595);
or (n6598,n6599,n6602);
and (n6599,n6600,n6601);
xor (n6600,n6426,n6427);
and (n6601,n308,n143);
and (n6602,n6603,n6604);
xor (n6603,n6600,n6601);
or (n6604,n6605,n6608);
and (n6605,n6606,n6607);
xor (n6606,n6432,n6433);
and (n6607,n51,n143);
and (n6608,n6609,n6610);
xor (n6609,n6606,n6607);
or (n6610,n6611,n6613);
and (n6611,n6612,n1958);
xor (n6612,n6438,n6439);
and (n6613,n6614,n6615);
xor (n6614,n6612,n1958);
or (n6615,n6616,n6619);
and (n6616,n6617,n6618);
xor (n6617,n6444,n6445);
and (n6618,n75,n143);
and (n6619,n6620,n6621);
xor (n6620,n6617,n6618);
or (n6621,n6622,n6625);
and (n6622,n6623,n6624);
xor (n6623,n6450,n6451);
and (n6624,n69,n143);
and (n6625,n6626,n6627);
xor (n6626,n6623,n6624);
or (n6627,n6628,n6631);
and (n6628,n6629,n6630);
xor (n6629,n6456,n6457);
and (n6630,n226,n143);
and (n6631,n6632,n6633);
xor (n6632,n6629,n6630);
or (n6633,n6634,n6637);
and (n6634,n6635,n6636);
xor (n6635,n6462,n6463);
and (n6636,n351,n143);
and (n6637,n6638,n6639);
xor (n6638,n6635,n6636);
or (n6639,n6640,n6643);
and (n6640,n6641,n6642);
xor (n6641,n6468,n6469);
and (n6642,n345,n143);
and (n6643,n6644,n6645);
xor (n6644,n6641,n6642);
or (n6645,n6646,n6649);
and (n6646,n6647,n6648);
xor (n6647,n6474,n6475);
and (n6648,n372,n143);
and (n6649,n6650,n6651);
xor (n6650,n6647,n6648);
or (n6651,n6652,n6655);
and (n6652,n6653,n6654);
xor (n6653,n6480,n6481);
and (n6654,n281,n143);
and (n6655,n6656,n6657);
xor (n6656,n6653,n6654);
or (n6657,n6658,n6661);
and (n6658,n6659,n6660);
xor (n6659,n6486,n6487);
and (n6660,n185,n143);
and (n6661,n6662,n6663);
xor (n6662,n6659,n6660);
or (n6663,n6664,n6667);
and (n6664,n6665,n6666);
xor (n6665,n6492,n6493);
and (n6666,n179,n143);
and (n6667,n6668,n6669);
xor (n6668,n6665,n6666);
or (n6669,n6670,n6673);
and (n6670,n6671,n6672);
xor (n6671,n6498,n6499);
and (n6672,n289,n143);
and (n6673,n6674,n6675);
xor (n6674,n6671,n6672);
or (n6675,n6676,n6679);
and (n6676,n6677,n6678);
xor (n6677,n6504,n6505);
and (n6678,n545,n143);
and (n6679,n6680,n6681);
xor (n6680,n6677,n6678);
or (n6681,n6682,n6685);
and (n6682,n6683,n6684);
xor (n6683,n6510,n6511);
and (n6684,n719,n143);
and (n6685,n6686,n6687);
xor (n6686,n6683,n6684);
or (n6687,n6688,n6691);
and (n6688,n6689,n6690);
xor (n6689,n6516,n6517);
and (n6690,n837,n143);
and (n6691,n6692,n6693);
xor (n6692,n6689,n6690);
or (n6693,n6694,n6697);
and (n6694,n6695,n6696);
xor (n6695,n6522,n6523);
and (n6696,n1175,n143);
and (n6697,n6698,n6699);
xor (n6698,n6695,n6696);
or (n6699,n6700,n6703);
and (n6700,n6701,n6702);
xor (n6701,n6528,n6529);
and (n6702,n1147,n143);
and (n6703,n6704,n6705);
xor (n6704,n6701,n6702);
or (n6705,n6706,n6709);
and (n6706,n6707,n6708);
xor (n6707,n6534,n6535);
and (n6708,n1141,n143);
and (n6709,n6710,n6711);
xor (n6710,n6707,n6708);
and (n6711,n6712,n6713);
xor (n6712,n6540,n6541);
and (n6713,n1187,n143);
and (n6714,n324,n141);
or (n6715,n6716,n6719);
and (n6716,n6717,n6718);
xor (n6717,n6549,n6550);
and (n6718,n158,n141);
and (n6719,n6720,n6721);
xor (n6720,n6717,n6718);
or (n6721,n6722,n6725);
and (n6722,n6723,n6724);
xor (n6723,n6555,n6556);
and (n6724,n151,n141);
and (n6725,n6726,n6727);
xor (n6726,n6723,n6724);
or (n6727,n6728,n6731);
and (n6728,n6729,n6730);
xor (n6729,n6561,n6562);
and (n6730,n195,n141);
and (n6731,n6732,n6733);
xor (n6732,n6729,n6730);
or (n6733,n6734,n6737);
and (n6734,n6735,n6736);
xor (n6735,n6567,n6568);
and (n6736,n103,n141);
and (n6737,n6738,n6739);
xor (n6738,n6735,n6736);
or (n6739,n6740,n6743);
and (n6740,n6741,n6742);
xor (n6741,n6573,n6574);
and (n6742,n97,n141);
and (n6743,n6744,n6745);
xor (n6744,n6741,n6742);
or (n6745,n6746,n6749);
and (n6746,n6747,n6748);
xor (n6747,n6579,n6580);
and (n6748,n257,n141);
and (n6749,n6750,n6751);
xor (n6750,n6747,n6748);
or (n6751,n6752,n6755);
and (n6752,n6753,n6754);
xor (n6753,n6585,n6586);
and (n6754,n250,n141);
and (n6755,n6756,n6757);
xor (n6756,n6753,n6754);
or (n6757,n6758,n6761);
and (n6758,n6759,n6760);
xor (n6759,n6591,n6592);
and (n6760,n315,n141);
and (n6761,n6762,n6763);
xor (n6762,n6759,n6760);
or (n6763,n6764,n6767);
and (n6764,n6765,n6766);
xor (n6765,n6597,n6598);
and (n6766,n308,n141);
and (n6767,n6768,n6769);
xor (n6768,n6765,n6766);
or (n6769,n6770,n6773);
and (n6770,n6771,n6772);
xor (n6771,n6603,n6604);
and (n6772,n51,n141);
and (n6773,n6774,n6775);
xor (n6774,n6771,n6772);
or (n6775,n6776,n6779);
and (n6776,n6777,n6778);
xor (n6777,n6609,n6610);
and (n6778,n45,n141);
and (n6779,n6780,n6781);
xor (n6780,n6777,n6778);
or (n6781,n6782,n6785);
and (n6782,n6783,n6784);
xor (n6783,n6614,n6615);
and (n6784,n75,n141);
and (n6785,n6786,n6787);
xor (n6786,n6783,n6784);
or (n6787,n6788,n6791);
and (n6788,n6789,n6790);
xor (n6789,n6620,n6621);
and (n6790,n69,n141);
and (n6791,n6792,n6793);
xor (n6792,n6789,n6790);
or (n6793,n6794,n6797);
and (n6794,n6795,n6796);
xor (n6795,n6626,n6627);
and (n6796,n226,n141);
and (n6797,n6798,n6799);
xor (n6798,n6795,n6796);
or (n6799,n6800,n6803);
and (n6800,n6801,n6802);
xor (n6801,n6632,n6633);
and (n6802,n351,n141);
and (n6803,n6804,n6805);
xor (n6804,n6801,n6802);
or (n6805,n6806,n6809);
and (n6806,n6807,n6808);
xor (n6807,n6638,n6639);
and (n6808,n345,n141);
and (n6809,n6810,n6811);
xor (n6810,n6807,n6808);
or (n6811,n6812,n6815);
and (n6812,n6813,n6814);
xor (n6813,n6644,n6645);
and (n6814,n372,n141);
and (n6815,n6816,n6817);
xor (n6816,n6813,n6814);
or (n6817,n6818,n6821);
and (n6818,n6819,n6820);
xor (n6819,n6650,n6651);
and (n6820,n281,n141);
and (n6821,n6822,n6823);
xor (n6822,n6819,n6820);
or (n6823,n6824,n6827);
and (n6824,n6825,n6826);
xor (n6825,n6656,n6657);
and (n6826,n185,n141);
and (n6827,n6828,n6829);
xor (n6828,n6825,n6826);
or (n6829,n6830,n6833);
and (n6830,n6831,n6832);
xor (n6831,n6662,n6663);
and (n6832,n179,n141);
and (n6833,n6834,n6835);
xor (n6834,n6831,n6832);
or (n6835,n6836,n6839);
and (n6836,n6837,n6838);
xor (n6837,n6668,n6669);
and (n6838,n289,n141);
and (n6839,n6840,n6841);
xor (n6840,n6837,n6838);
or (n6841,n6842,n6845);
and (n6842,n6843,n6844);
xor (n6843,n6674,n6675);
and (n6844,n545,n141);
and (n6845,n6846,n6847);
xor (n6846,n6843,n6844);
or (n6847,n6848,n6851);
and (n6848,n6849,n6850);
xor (n6849,n6680,n6681);
and (n6850,n719,n141);
and (n6851,n6852,n6853);
xor (n6852,n6849,n6850);
or (n6853,n6854,n6857);
and (n6854,n6855,n6856);
xor (n6855,n6686,n6687);
and (n6856,n837,n141);
and (n6857,n6858,n6859);
xor (n6858,n6855,n6856);
or (n6859,n6860,n6863);
and (n6860,n6861,n6862);
xor (n6861,n6692,n6693);
and (n6862,n1175,n141);
and (n6863,n6864,n6865);
xor (n6864,n6861,n6862);
or (n6865,n6866,n6869);
and (n6866,n6867,n6868);
xor (n6867,n6698,n6699);
and (n6868,n1147,n141);
and (n6869,n6870,n6871);
xor (n6870,n6867,n6868);
or (n6871,n6872,n6875);
and (n6872,n6873,n6874);
xor (n6873,n6704,n6705);
and (n6874,n1141,n141);
and (n6875,n6876,n6877);
xor (n6876,n6873,n6874);
and (n6877,n6878,n6879);
xor (n6878,n6710,n6711);
not (n6879,n3327);
and (n6880,n158,n85);
or (n6881,n6882,n6885);
and (n6882,n6883,n6884);
xor (n6883,n6720,n6721);
and (n6884,n151,n85);
and (n6885,n6886,n6887);
xor (n6886,n6883,n6884);
or (n6887,n6888,n6891);
and (n6888,n6889,n6890);
xor (n6889,n6726,n6727);
and (n6890,n195,n85);
and (n6891,n6892,n6893);
xor (n6892,n6889,n6890);
or (n6893,n6894,n6897);
and (n6894,n6895,n6896);
xor (n6895,n6732,n6733);
and (n6896,n103,n85);
and (n6897,n6898,n6899);
xor (n6898,n6895,n6896);
or (n6899,n6900,n6903);
and (n6900,n6901,n6902);
xor (n6901,n6738,n6739);
and (n6902,n97,n85);
and (n6903,n6904,n6905);
xor (n6904,n6901,n6902);
or (n6905,n6906,n6909);
and (n6906,n6907,n6908);
xor (n6907,n6744,n6745);
and (n6908,n257,n85);
and (n6909,n6910,n6911);
xor (n6910,n6907,n6908);
or (n6911,n6912,n6915);
and (n6912,n6913,n6914);
xor (n6913,n6750,n6751);
and (n6914,n250,n85);
and (n6915,n6916,n6917);
xor (n6916,n6913,n6914);
or (n6917,n6918,n6921);
and (n6918,n6919,n6920);
xor (n6919,n6756,n6757);
and (n6920,n315,n85);
and (n6921,n6922,n6923);
xor (n6922,n6919,n6920);
or (n6923,n6924,n6927);
and (n6924,n6925,n6926);
xor (n6925,n6762,n6763);
and (n6926,n308,n85);
and (n6927,n6928,n6929);
xor (n6928,n6925,n6926);
or (n6929,n6930,n6933);
and (n6930,n6931,n6932);
xor (n6931,n6768,n6769);
and (n6932,n51,n85);
and (n6933,n6934,n6935);
xor (n6934,n6931,n6932);
or (n6935,n6936,n6939);
and (n6936,n6937,n6938);
xor (n6937,n6774,n6775);
and (n6938,n45,n85);
and (n6939,n6940,n6941);
xor (n6940,n6937,n6938);
or (n6941,n6942,n6945);
and (n6942,n6943,n6944);
xor (n6943,n6780,n6781);
and (n6944,n75,n85);
and (n6945,n6946,n6947);
xor (n6946,n6943,n6944);
or (n6947,n6948,n6951);
and (n6948,n6949,n6950);
xor (n6949,n6786,n6787);
and (n6950,n69,n85);
and (n6951,n6952,n6953);
xor (n6952,n6949,n6950);
or (n6953,n6954,n6957);
and (n6954,n6955,n6956);
xor (n6955,n6792,n6793);
and (n6956,n226,n85);
and (n6957,n6958,n6959);
xor (n6958,n6955,n6956);
or (n6959,n6960,n6963);
and (n6960,n6961,n6962);
xor (n6961,n6798,n6799);
and (n6962,n351,n85);
and (n6963,n6964,n6965);
xor (n6964,n6961,n6962);
or (n6965,n6966,n6969);
and (n6966,n6967,n6968);
xor (n6967,n6804,n6805);
and (n6968,n345,n85);
and (n6969,n6970,n6971);
xor (n6970,n6967,n6968);
or (n6971,n6972,n6975);
and (n6972,n6973,n6974);
xor (n6973,n6810,n6811);
and (n6974,n372,n85);
and (n6975,n6976,n6977);
xor (n6976,n6973,n6974);
or (n6977,n6978,n6981);
and (n6978,n6979,n6980);
xor (n6979,n6816,n6817);
and (n6980,n281,n85);
and (n6981,n6982,n6983);
xor (n6982,n6979,n6980);
or (n6983,n6984,n6987);
and (n6984,n6985,n6986);
xor (n6985,n6822,n6823);
and (n6986,n185,n85);
and (n6987,n6988,n6989);
xor (n6988,n6985,n6986);
or (n6989,n6990,n6993);
and (n6990,n6991,n6992);
xor (n6991,n6828,n6829);
and (n6992,n179,n85);
and (n6993,n6994,n6995);
xor (n6994,n6991,n6992);
or (n6995,n6996,n6999);
and (n6996,n6997,n6998);
xor (n6997,n6834,n6835);
and (n6998,n289,n85);
and (n6999,n7000,n7001);
xor (n7000,n6997,n6998);
or (n7001,n7002,n7005);
and (n7002,n7003,n7004);
xor (n7003,n6840,n6841);
and (n7004,n545,n85);
and (n7005,n7006,n7007);
xor (n7006,n7003,n7004);
or (n7007,n7008,n7011);
and (n7008,n7009,n7010);
xor (n7009,n6846,n6847);
and (n7010,n719,n85);
and (n7011,n7012,n7013);
xor (n7012,n7009,n7010);
or (n7013,n7014,n7017);
and (n7014,n7015,n7016);
xor (n7015,n6852,n6853);
and (n7016,n837,n85);
and (n7017,n7018,n7019);
xor (n7018,n7015,n7016);
or (n7019,n7020,n7023);
and (n7020,n7021,n7022);
xor (n7021,n6858,n6859);
and (n7022,n1175,n85);
and (n7023,n7024,n7025);
xor (n7024,n7021,n7022);
or (n7025,n7026,n7029);
and (n7026,n7027,n7028);
xor (n7027,n6864,n6865);
and (n7028,n1147,n85);
and (n7029,n7030,n7031);
xor (n7030,n7027,n7028);
or (n7031,n7032,n7035);
and (n7032,n7033,n7034);
xor (n7033,n6870,n6871);
and (n7034,n1141,n85);
and (n7035,n7036,n7037);
xor (n7036,n7033,n7034);
and (n7037,n7038,n7039);
xor (n7038,n6876,n6877);
and (n7039,n1187,n85);
and (n7040,n151,n86);
or (n7041,n7042,n7045);
and (n7042,n7043,n7044);
xor (n7043,n6886,n6887);
and (n7044,n195,n86);
and (n7045,n7046,n7047);
xor (n7046,n7043,n7044);
or (n7047,n7048,n7051);
and (n7048,n7049,n7050);
xor (n7049,n6892,n6893);
and (n7050,n103,n86);
and (n7051,n7052,n7053);
xor (n7052,n7049,n7050);
or (n7053,n7054,n7057);
and (n7054,n7055,n7056);
xor (n7055,n6898,n6899);
and (n7056,n97,n86);
and (n7057,n7058,n7059);
xor (n7058,n7055,n7056);
or (n7059,n7060,n7063);
and (n7060,n7061,n7062);
xor (n7061,n6904,n6905);
and (n7062,n257,n86);
and (n7063,n7064,n7065);
xor (n7064,n7061,n7062);
or (n7065,n7066,n7069);
and (n7066,n7067,n7068);
xor (n7067,n6910,n6911);
and (n7068,n250,n86);
and (n7069,n7070,n7071);
xor (n7070,n7067,n7068);
or (n7071,n7072,n7075);
and (n7072,n7073,n7074);
xor (n7073,n6916,n6917);
and (n7074,n315,n86);
and (n7075,n7076,n7077);
xor (n7076,n7073,n7074);
or (n7077,n7078,n7081);
and (n7078,n7079,n7080);
xor (n7079,n6922,n6923);
and (n7080,n308,n86);
and (n7081,n7082,n7083);
xor (n7082,n7079,n7080);
or (n7083,n7084,n7087);
and (n7084,n7085,n7086);
xor (n7085,n6928,n6929);
and (n7086,n51,n86);
and (n7087,n7088,n7089);
xor (n7088,n7085,n7086);
or (n7089,n7090,n7093);
and (n7090,n7091,n7092);
xor (n7091,n6934,n6935);
and (n7092,n45,n86);
and (n7093,n7094,n7095);
xor (n7094,n7091,n7092);
or (n7095,n7096,n7099);
and (n7096,n7097,n7098);
xor (n7097,n6940,n6941);
and (n7098,n75,n86);
and (n7099,n7100,n7101);
xor (n7100,n7097,n7098);
or (n7101,n7102,n7105);
and (n7102,n7103,n7104);
xor (n7103,n6946,n6947);
and (n7104,n69,n86);
and (n7105,n7106,n7107);
xor (n7106,n7103,n7104);
or (n7107,n7108,n7111);
and (n7108,n7109,n7110);
xor (n7109,n6952,n6953);
and (n7110,n226,n86);
and (n7111,n7112,n7113);
xor (n7112,n7109,n7110);
or (n7113,n7114,n7117);
and (n7114,n7115,n7116);
xor (n7115,n6958,n6959);
and (n7116,n351,n86);
and (n7117,n7118,n7119);
xor (n7118,n7115,n7116);
or (n7119,n7120,n7123);
and (n7120,n7121,n7122);
xor (n7121,n6964,n6965);
and (n7122,n345,n86);
and (n7123,n7124,n7125);
xor (n7124,n7121,n7122);
or (n7125,n7126,n7129);
and (n7126,n7127,n7128);
xor (n7127,n6970,n6971);
and (n7128,n372,n86);
and (n7129,n7130,n7131);
xor (n7130,n7127,n7128);
or (n7131,n7132,n7135);
and (n7132,n7133,n7134);
xor (n7133,n6976,n6977);
and (n7134,n281,n86);
and (n7135,n7136,n7137);
xor (n7136,n7133,n7134);
or (n7137,n7138,n7141);
and (n7138,n7139,n7140);
xor (n7139,n6982,n6983);
and (n7140,n185,n86);
and (n7141,n7142,n7143);
xor (n7142,n7139,n7140);
or (n7143,n7144,n7147);
and (n7144,n7145,n7146);
xor (n7145,n6988,n6989);
and (n7146,n179,n86);
and (n7147,n7148,n7149);
xor (n7148,n7145,n7146);
or (n7149,n7150,n7153);
and (n7150,n7151,n7152);
xor (n7151,n6994,n6995);
and (n7152,n289,n86);
and (n7153,n7154,n7155);
xor (n7154,n7151,n7152);
or (n7155,n7156,n7159);
and (n7156,n7157,n7158);
xor (n7157,n7000,n7001);
and (n7158,n545,n86);
and (n7159,n7160,n7161);
xor (n7160,n7157,n7158);
or (n7161,n7162,n7165);
and (n7162,n7163,n7164);
xor (n7163,n7006,n7007);
and (n7164,n719,n86);
and (n7165,n7166,n7167);
xor (n7166,n7163,n7164);
or (n7167,n7168,n7171);
and (n7168,n7169,n7170);
xor (n7169,n7012,n7013);
and (n7170,n837,n86);
and (n7171,n7172,n7173);
xor (n7172,n7169,n7170);
or (n7173,n7174,n7177);
and (n7174,n7175,n7176);
xor (n7175,n7018,n7019);
and (n7176,n1175,n86);
and (n7177,n7178,n7179);
xor (n7178,n7175,n7176);
or (n7179,n7180,n7183);
and (n7180,n7181,n7182);
xor (n7181,n7024,n7025);
and (n7182,n1147,n86);
and (n7183,n7184,n7185);
xor (n7184,n7181,n7182);
or (n7185,n7186,n7189);
and (n7186,n7187,n7188);
xor (n7187,n7030,n7031);
and (n7188,n1141,n86);
and (n7189,n7190,n7191);
xor (n7190,n7187,n7188);
and (n7191,n7192,n7193);
xor (n7192,n7036,n7037);
not (n7193,n3348);
and (n7194,n195,n92);
or (n7195,n7196,n7199);
and (n7196,n7197,n7198);
xor (n7197,n7046,n7047);
and (n7198,n103,n92);
and (n7199,n7200,n7201);
xor (n7200,n7197,n7198);
or (n7201,n7202,n7205);
and (n7202,n7203,n7204);
xor (n7203,n7052,n7053);
and (n7204,n97,n92);
and (n7205,n7206,n7207);
xor (n7206,n7203,n7204);
or (n7207,n7208,n7211);
and (n7208,n7209,n7210);
xor (n7209,n7058,n7059);
and (n7210,n257,n92);
and (n7211,n7212,n7213);
xor (n7212,n7209,n7210);
or (n7213,n7214,n7217);
and (n7214,n7215,n7216);
xor (n7215,n7064,n7065);
and (n7216,n250,n92);
and (n7217,n7218,n7219);
xor (n7218,n7215,n7216);
or (n7219,n7220,n7223);
and (n7220,n7221,n7222);
xor (n7221,n7070,n7071);
and (n7222,n315,n92);
and (n7223,n7224,n7225);
xor (n7224,n7221,n7222);
or (n7225,n7226,n7229);
and (n7226,n7227,n7228);
xor (n7227,n7076,n7077);
and (n7228,n308,n92);
and (n7229,n7230,n7231);
xor (n7230,n7227,n7228);
or (n7231,n7232,n7235);
and (n7232,n7233,n7234);
xor (n7233,n7082,n7083);
and (n7234,n51,n92);
and (n7235,n7236,n7237);
xor (n7236,n7233,n7234);
or (n7237,n7238,n7241);
and (n7238,n7239,n7240);
xor (n7239,n7088,n7089);
and (n7240,n45,n92);
and (n7241,n7242,n7243);
xor (n7242,n7239,n7240);
or (n7243,n7244,n7247);
and (n7244,n7245,n7246);
xor (n7245,n7094,n7095);
and (n7246,n75,n92);
and (n7247,n7248,n7249);
xor (n7248,n7245,n7246);
or (n7249,n7250,n7253);
and (n7250,n7251,n7252);
xor (n7251,n7100,n7101);
and (n7252,n69,n92);
and (n7253,n7254,n7255);
xor (n7254,n7251,n7252);
or (n7255,n7256,n7259);
and (n7256,n7257,n7258);
xor (n7257,n7106,n7107);
and (n7258,n226,n92);
and (n7259,n7260,n7261);
xor (n7260,n7257,n7258);
or (n7261,n7262,n7265);
and (n7262,n7263,n7264);
xor (n7263,n7112,n7113);
and (n7264,n351,n92);
and (n7265,n7266,n7267);
xor (n7266,n7263,n7264);
or (n7267,n7268,n7271);
and (n7268,n7269,n7270);
xor (n7269,n7118,n7119);
and (n7270,n345,n92);
and (n7271,n7272,n7273);
xor (n7272,n7269,n7270);
or (n7273,n7274,n7277);
and (n7274,n7275,n7276);
xor (n7275,n7124,n7125);
and (n7276,n372,n92);
and (n7277,n7278,n7279);
xor (n7278,n7275,n7276);
or (n7279,n7280,n7283);
and (n7280,n7281,n7282);
xor (n7281,n7130,n7131);
and (n7282,n281,n92);
and (n7283,n7284,n7285);
xor (n7284,n7281,n7282);
or (n7285,n7286,n7289);
and (n7286,n7287,n7288);
xor (n7287,n7136,n7137);
and (n7288,n185,n92);
and (n7289,n7290,n7291);
xor (n7290,n7287,n7288);
or (n7291,n7292,n7294);
and (n7292,n7293,n3658);
xor (n7293,n7142,n7143);
and (n7294,n7295,n7296);
xor (n7295,n7293,n3658);
or (n7296,n7297,n7300);
and (n7297,n7298,n7299);
xor (n7298,n7148,n7149);
and (n7299,n289,n92);
and (n7300,n7301,n7302);
xor (n7301,n7298,n7299);
or (n7302,n7303,n7306);
and (n7303,n7304,n7305);
xor (n7304,n7154,n7155);
and (n7305,n545,n92);
and (n7306,n7307,n7308);
xor (n7307,n7304,n7305);
or (n7308,n7309,n7311);
and (n7309,n7310,n2862);
xor (n7310,n7160,n7161);
and (n7311,n7312,n7313);
xor (n7312,n7310,n2862);
or (n7313,n7314,n7317);
and (n7314,n7315,n7316);
xor (n7315,n7166,n7167);
and (n7316,n837,n92);
and (n7317,n7318,n7319);
xor (n7318,n7315,n7316);
or (n7319,n7320,n7323);
and (n7320,n7321,n7322);
xor (n7321,n7172,n7173);
and (n7322,n1175,n92);
and (n7323,n7324,n7325);
xor (n7324,n7321,n7322);
or (n7325,n7326,n7329);
and (n7326,n7327,n7328);
xor (n7327,n7178,n7179);
and (n7328,n1147,n92);
and (n7329,n7330,n7331);
xor (n7330,n7327,n7328);
or (n7331,n7332,n7335);
and (n7332,n7333,n7334);
xor (n7333,n7184,n7185);
and (n7334,n1141,n92);
and (n7335,n7336,n7337);
xor (n7336,n7333,n7334);
and (n7337,n7338,n7339);
xor (n7338,n7190,n7191);
and (n7339,n1187,n92);
and (n7340,n103,n242);
or (n7341,n7342,n7345);
and (n7342,n7343,n7344);
xor (n7343,n7200,n7201);
and (n7344,n97,n242);
and (n7345,n7346,n7347);
xor (n7346,n7343,n7344);
or (n7347,n7348,n7351);
and (n7348,n7349,n7350);
xor (n7349,n7206,n7207);
and (n7350,n257,n242);
and (n7351,n7352,n7353);
xor (n7352,n7349,n7350);
or (n7353,n7354,n7357);
and (n7354,n7355,n7356);
xor (n7355,n7212,n7213);
and (n7356,n250,n242);
and (n7357,n7358,n7359);
xor (n7358,n7355,n7356);
or (n7359,n7360,n7363);
and (n7360,n7361,n7362);
xor (n7361,n7218,n7219);
and (n7362,n315,n242);
and (n7363,n7364,n7365);
xor (n7364,n7361,n7362);
or (n7365,n7366,n7369);
and (n7366,n7367,n7368);
xor (n7367,n7224,n7225);
and (n7368,n308,n242);
and (n7369,n7370,n7371);
xor (n7370,n7367,n7368);
or (n7371,n7372,n7375);
and (n7372,n7373,n7374);
xor (n7373,n7230,n7231);
and (n7374,n51,n242);
and (n7375,n7376,n7377);
xor (n7376,n7373,n7374);
or (n7377,n7378,n7381);
and (n7378,n7379,n7380);
xor (n7379,n7236,n7237);
and (n7380,n45,n242);
and (n7381,n7382,n7383);
xor (n7382,n7379,n7380);
or (n7383,n7384,n7387);
and (n7384,n7385,n7386);
xor (n7385,n7242,n7243);
and (n7386,n75,n242);
and (n7387,n7388,n7389);
xor (n7388,n7385,n7386);
or (n7389,n7390,n7393);
and (n7390,n7391,n7392);
xor (n7391,n7248,n7249);
and (n7392,n69,n242);
and (n7393,n7394,n7395);
xor (n7394,n7391,n7392);
or (n7395,n7396,n7399);
and (n7396,n7397,n7398);
xor (n7397,n7254,n7255);
and (n7398,n226,n242);
and (n7399,n7400,n7401);
xor (n7400,n7397,n7398);
or (n7401,n7402,n7405);
and (n7402,n7403,n7404);
xor (n7403,n7260,n7261);
and (n7404,n351,n242);
and (n7405,n7406,n7407);
xor (n7406,n7403,n7404);
or (n7407,n7408,n7411);
and (n7408,n7409,n7410);
xor (n7409,n7266,n7267);
and (n7410,n345,n242);
and (n7411,n7412,n7413);
xor (n7412,n7409,n7410);
or (n7413,n7414,n7417);
and (n7414,n7415,n7416);
xor (n7415,n7272,n7273);
and (n7416,n372,n242);
and (n7417,n7418,n7419);
xor (n7418,n7415,n7416);
or (n7419,n7420,n7423);
and (n7420,n7421,n7422);
xor (n7421,n7278,n7279);
and (n7422,n281,n242);
and (n7423,n7424,n7425);
xor (n7424,n7421,n7422);
or (n7425,n7426,n7429);
and (n7426,n7427,n7428);
xor (n7427,n7284,n7285);
and (n7428,n185,n242);
and (n7429,n7430,n7431);
xor (n7430,n7427,n7428);
or (n7431,n7432,n7435);
and (n7432,n7433,n7434);
xor (n7433,n7290,n7291);
and (n7434,n179,n242);
and (n7435,n7436,n7437);
xor (n7436,n7433,n7434);
or (n7437,n7438,n7441);
and (n7438,n7439,n7440);
xor (n7439,n7295,n7296);
and (n7440,n289,n242);
and (n7441,n7442,n7443);
xor (n7442,n7439,n7440);
or (n7443,n7444,n7447);
and (n7444,n7445,n7446);
xor (n7445,n7301,n7302);
and (n7446,n545,n242);
and (n7447,n7448,n7449);
xor (n7448,n7445,n7446);
or (n7449,n7450,n7453);
and (n7450,n7451,n7452);
xor (n7451,n7307,n7308);
and (n7452,n719,n242);
and (n7453,n7454,n7455);
xor (n7454,n7451,n7452);
or (n7455,n7456,n7459);
and (n7456,n7457,n7458);
xor (n7457,n7312,n7313);
and (n7458,n837,n242);
and (n7459,n7460,n7461);
xor (n7460,n7457,n7458);
or (n7461,n7462,n7465);
and (n7462,n7463,n7464);
xor (n7463,n7318,n7319);
and (n7464,n1175,n242);
and (n7465,n7466,n7467);
xor (n7466,n7463,n7464);
or (n7467,n7468,n7471);
and (n7468,n7469,n7470);
xor (n7469,n7324,n7325);
and (n7470,n1147,n242);
and (n7471,n7472,n7473);
xor (n7472,n7469,n7470);
or (n7473,n7474,n7477);
and (n7474,n7475,n7476);
xor (n7475,n7330,n7331);
and (n7476,n1141,n242);
and (n7477,n7478,n7479);
xor (n7478,n7475,n7476);
and (n7479,n7480,n7481);
xor (n7480,n7336,n7337);
not (n7481,n3105);
and (n7482,n97,n241);
or (n7483,n7484,n7487);
and (n7484,n7485,n7486);
xor (n7485,n7346,n7347);
and (n7486,n257,n241);
and (n7487,n7488,n7489);
xor (n7488,n7485,n7486);
or (n7489,n7490,n7493);
and (n7490,n7491,n7492);
xor (n7491,n7352,n7353);
and (n7492,n250,n241);
and (n7493,n7494,n7495);
xor (n7494,n7491,n7492);
or (n7495,n7496,n7499);
and (n7496,n7497,n7498);
xor (n7497,n7358,n7359);
and (n7498,n315,n241);
and (n7499,n7500,n7501);
xor (n7500,n7497,n7498);
or (n7501,n7502,n7505);
and (n7502,n7503,n7504);
xor (n7503,n7364,n7365);
and (n7504,n308,n241);
and (n7505,n7506,n7507);
xor (n7506,n7503,n7504);
or (n7507,n7508,n7511);
and (n7508,n7509,n7510);
xor (n7509,n7370,n7371);
and (n7510,n51,n241);
and (n7511,n7512,n7513);
xor (n7512,n7509,n7510);
or (n7513,n7514,n7517);
and (n7514,n7515,n7516);
xor (n7515,n7376,n7377);
and (n7516,n45,n241);
and (n7517,n7518,n7519);
xor (n7518,n7515,n7516);
or (n7519,n7520,n7523);
and (n7520,n7521,n7522);
xor (n7521,n7382,n7383);
and (n7522,n75,n241);
and (n7523,n7524,n7525);
xor (n7524,n7521,n7522);
or (n7525,n7526,n7529);
and (n7526,n7527,n7528);
xor (n7527,n7388,n7389);
and (n7528,n69,n241);
and (n7529,n7530,n7531);
xor (n7530,n7527,n7528);
or (n7531,n7532,n7535);
and (n7532,n7533,n7534);
xor (n7533,n7394,n7395);
and (n7534,n226,n241);
and (n7535,n7536,n7537);
xor (n7536,n7533,n7534);
or (n7537,n7538,n7541);
and (n7538,n7539,n7540);
xor (n7539,n7400,n7401);
and (n7540,n351,n241);
and (n7541,n7542,n7543);
xor (n7542,n7539,n7540);
or (n7543,n7544,n7547);
and (n7544,n7545,n7546);
xor (n7545,n7406,n7407);
and (n7546,n345,n241);
and (n7547,n7548,n7549);
xor (n7548,n7545,n7546);
or (n7549,n7550,n7553);
and (n7550,n7551,n7552);
xor (n7551,n7412,n7413);
and (n7552,n372,n241);
and (n7553,n7554,n7555);
xor (n7554,n7551,n7552);
or (n7555,n7556,n7559);
and (n7556,n7557,n7558);
xor (n7557,n7418,n7419);
and (n7558,n281,n241);
and (n7559,n7560,n7561);
xor (n7560,n7557,n7558);
or (n7561,n7562,n7565);
and (n7562,n7563,n7564);
xor (n7563,n7424,n7425);
and (n7564,n185,n241);
and (n7565,n7566,n7567);
xor (n7566,n7563,n7564);
or (n7567,n7568,n7571);
and (n7568,n7569,n7570);
xor (n7569,n7430,n7431);
and (n7570,n179,n241);
and (n7571,n7572,n7573);
xor (n7572,n7569,n7570);
or (n7573,n7574,n7577);
and (n7574,n7575,n7576);
xor (n7575,n7436,n7437);
and (n7576,n289,n241);
and (n7577,n7578,n7579);
xor (n7578,n7575,n7576);
or (n7579,n7580,n7583);
and (n7580,n7581,n7582);
xor (n7581,n7442,n7443);
and (n7582,n545,n241);
and (n7583,n7584,n7585);
xor (n7584,n7581,n7582);
or (n7585,n7586,n7589);
and (n7586,n7587,n7588);
xor (n7587,n7448,n7449);
and (n7588,n719,n241);
and (n7589,n7590,n7591);
xor (n7590,n7587,n7588);
or (n7591,n7592,n7595);
and (n7592,n7593,n7594);
xor (n7593,n7454,n7455);
and (n7594,n837,n241);
and (n7595,n7596,n7597);
xor (n7596,n7593,n7594);
or (n7597,n7598,n7601);
and (n7598,n7599,n7600);
xor (n7599,n7460,n7461);
and (n7600,n1175,n241);
and (n7601,n7602,n7603);
xor (n7602,n7599,n7600);
or (n7603,n7604,n7607);
and (n7604,n7605,n7606);
xor (n7605,n7466,n7467);
and (n7606,n1147,n241);
and (n7607,n7608,n7609);
xor (n7608,n7605,n7606);
or (n7609,n7610,n7613);
and (n7610,n7611,n7612);
xor (n7611,n7472,n7473);
and (n7612,n1141,n241);
and (n7613,n7614,n7615);
xor (n7614,n7611,n7612);
and (n7615,n7616,n7617);
xor (n7616,n7478,n7479);
and (n7617,n1187,n241);
and (n7618,n257,n300);
or (n7619,n7620,n7623);
and (n7620,n7621,n7622);
xor (n7621,n7488,n7489);
and (n7622,n250,n300);
and (n7623,n7624,n7625);
xor (n7624,n7621,n7622);
or (n7625,n7626,n7629);
and (n7626,n7627,n7628);
xor (n7627,n7494,n7495);
and (n7628,n315,n300);
and (n7629,n7630,n7631);
xor (n7630,n7627,n7628);
or (n7631,n7632,n7635);
and (n7632,n7633,n7634);
xor (n7633,n7500,n7501);
and (n7634,n308,n300);
and (n7635,n7636,n7637);
xor (n7636,n7633,n7634);
or (n7637,n7638,n7641);
and (n7638,n7639,n7640);
xor (n7639,n7506,n7507);
and (n7640,n51,n300);
and (n7641,n7642,n7643);
xor (n7642,n7639,n7640);
or (n7643,n7644,n7647);
and (n7644,n7645,n7646);
xor (n7645,n7512,n7513);
and (n7646,n45,n300);
and (n7647,n7648,n7649);
xor (n7648,n7645,n7646);
or (n7649,n7650,n7653);
and (n7650,n7651,n7652);
xor (n7651,n7518,n7519);
and (n7652,n75,n300);
and (n7653,n7654,n7655);
xor (n7654,n7651,n7652);
or (n7655,n7656,n7659);
and (n7656,n7657,n7658);
xor (n7657,n7524,n7525);
and (n7658,n69,n300);
and (n7659,n7660,n7661);
xor (n7660,n7657,n7658);
or (n7661,n7662,n7665);
and (n7662,n7663,n7664);
xor (n7663,n7530,n7531);
and (n7664,n226,n300);
and (n7665,n7666,n7667);
xor (n7666,n7663,n7664);
or (n7667,n7668,n7671);
and (n7668,n7669,n7670);
xor (n7669,n7536,n7537);
and (n7670,n351,n300);
and (n7671,n7672,n7673);
xor (n7672,n7669,n7670);
or (n7673,n7674,n7677);
and (n7674,n7675,n7676);
xor (n7675,n7542,n7543);
and (n7676,n345,n300);
and (n7677,n7678,n7679);
xor (n7678,n7675,n7676);
or (n7679,n7680,n7683);
and (n7680,n7681,n7682);
xor (n7681,n7548,n7549);
and (n7682,n372,n300);
and (n7683,n7684,n7685);
xor (n7684,n7681,n7682);
or (n7685,n7686,n7689);
and (n7686,n7687,n7688);
xor (n7687,n7554,n7555);
and (n7688,n281,n300);
and (n7689,n7690,n7691);
xor (n7690,n7687,n7688);
or (n7691,n7692,n7695);
and (n7692,n7693,n7694);
xor (n7693,n7560,n7561);
and (n7694,n185,n300);
and (n7695,n7696,n7697);
xor (n7696,n7693,n7694);
or (n7697,n7698,n7701);
and (n7698,n7699,n7700);
xor (n7699,n7566,n7567);
and (n7700,n179,n300);
and (n7701,n7702,n7703);
xor (n7702,n7699,n7700);
or (n7703,n7704,n7707);
and (n7704,n7705,n7706);
xor (n7705,n7572,n7573);
and (n7706,n289,n300);
and (n7707,n7708,n7709);
xor (n7708,n7705,n7706);
or (n7709,n7710,n7713);
and (n7710,n7711,n7712);
xor (n7711,n7578,n7579);
and (n7712,n545,n300);
and (n7713,n7714,n7715);
xor (n7714,n7711,n7712);
or (n7715,n7716,n7719);
and (n7716,n7717,n7718);
xor (n7717,n7584,n7585);
and (n7718,n719,n300);
and (n7719,n7720,n7721);
xor (n7720,n7717,n7718);
or (n7721,n7722,n7725);
and (n7722,n7723,n7724);
xor (n7723,n7590,n7591);
and (n7724,n837,n300);
and (n7725,n7726,n7727);
xor (n7726,n7723,n7724);
or (n7727,n7728,n7731);
and (n7728,n7729,n7730);
xor (n7729,n7596,n7597);
and (n7730,n1175,n300);
and (n7731,n7732,n7733);
xor (n7732,n7729,n7730);
or (n7733,n7734,n7737);
and (n7734,n7735,n7736);
xor (n7735,n7602,n7603);
and (n7736,n1147,n300);
and (n7737,n7738,n7739);
xor (n7738,n7735,n7736);
or (n7739,n7740,n7743);
and (n7740,n7741,n7742);
xor (n7741,n7608,n7609);
and (n7742,n1141,n300);
and (n7743,n7744,n7745);
xor (n7744,n7741,n7742);
and (n7745,n7746,n7747);
xor (n7746,n7614,n7615);
not (n7747,n2727);
and (n7748,n250,n41);
or (n7749,n7750,n7753);
and (n7750,n7751,n7752);
xor (n7751,n7624,n7625);
and (n7752,n315,n41);
and (n7753,n7754,n7755);
xor (n7754,n7751,n7752);
or (n7755,n7756,n7759);
and (n7756,n7757,n7758);
xor (n7757,n7630,n7631);
and (n7758,n308,n41);
and (n7759,n7760,n7761);
xor (n7760,n7757,n7758);
or (n7761,n7762,n7765);
and (n7762,n7763,n7764);
xor (n7763,n7636,n7637);
and (n7764,n51,n41);
and (n7765,n7766,n7767);
xor (n7766,n7763,n7764);
or (n7767,n7768,n7771);
and (n7768,n7769,n7770);
xor (n7769,n7642,n7643);
and (n7770,n45,n41);
and (n7771,n7772,n7773);
xor (n7772,n7769,n7770);
or (n7773,n7774,n7777);
and (n7774,n7775,n7776);
xor (n7775,n7648,n7649);
and (n7776,n75,n41);
and (n7777,n7778,n7779);
xor (n7778,n7775,n7776);
or (n7779,n7780,n7783);
and (n7780,n7781,n7782);
xor (n7781,n7654,n7655);
and (n7782,n69,n41);
and (n7783,n7784,n7785);
xor (n7784,n7781,n7782);
or (n7785,n7786,n7789);
and (n7786,n7787,n7788);
xor (n7787,n7660,n7661);
and (n7788,n226,n41);
and (n7789,n7790,n7791);
xor (n7790,n7787,n7788);
or (n7791,n7792,n7795);
and (n7792,n7793,n7794);
xor (n7793,n7666,n7667);
and (n7794,n351,n41);
and (n7795,n7796,n7797);
xor (n7796,n7793,n7794);
or (n7797,n7798,n7801);
and (n7798,n7799,n7800);
xor (n7799,n7672,n7673);
and (n7800,n345,n41);
and (n7801,n7802,n7803);
xor (n7802,n7799,n7800);
or (n7803,n7804,n7807);
and (n7804,n7805,n7806);
xor (n7805,n7678,n7679);
and (n7806,n372,n41);
and (n7807,n7808,n7809);
xor (n7808,n7805,n7806);
or (n7809,n7810,n7812);
and (n7810,n7811,n1705);
xor (n7811,n7684,n7685);
and (n7812,n7813,n7814);
xor (n7813,n7811,n1705);
or (n7814,n7815,n7817);
and (n7815,n7816,n1877);
xor (n7816,n7690,n7691);
and (n7817,n7818,n7819);
xor (n7818,n7816,n1877);
or (n7819,n7820,n7823);
and (n7820,n7821,n7822);
xor (n7821,n7696,n7697);
and (n7822,n179,n41);
and (n7823,n7824,n7825);
xor (n7824,n7821,n7822);
or (n7825,n7826,n7829);
and (n7826,n7827,n7828);
xor (n7827,n7702,n7703);
and (n7828,n289,n41);
and (n7829,n7830,n7831);
xor (n7830,n7827,n7828);
or (n7831,n7832,n7835);
and (n7832,n7833,n7834);
xor (n7833,n7708,n7709);
and (n7834,n545,n41);
and (n7835,n7836,n7837);
xor (n7836,n7833,n7834);
or (n7837,n7838,n7841);
and (n7838,n7839,n7840);
xor (n7839,n7714,n7715);
and (n7840,n719,n41);
and (n7841,n7842,n7843);
xor (n7842,n7839,n7840);
or (n7843,n7844,n7846);
and (n7844,n7845,n3683);
xor (n7845,n7720,n7721);
and (n7846,n7847,n7848);
xor (n7847,n7845,n3683);
or (n7848,n7849,n7851);
and (n7849,n7850,n2983);
xor (n7850,n7726,n7727);
and (n7851,n7852,n7853);
xor (n7852,n7850,n2983);
or (n7853,n7854,n7857);
and (n7854,n7855,n7856);
xor (n7855,n7732,n7733);
and (n7856,n1147,n41);
and (n7857,n7858,n7859);
xor (n7858,n7855,n7856);
or (n7859,n7860,n7863);
and (n7860,n7861,n7862);
xor (n7861,n7738,n7739);
and (n7862,n1141,n41);
and (n7863,n7864,n7865);
xor (n7864,n7861,n7862);
and (n7865,n7866,n7867);
xor (n7866,n7744,n7745);
and (n7867,n1187,n41);
and (n7868,n315,n33);
or (n7869,n7870,n7873);
and (n7870,n7871,n7872);
xor (n7871,n7754,n7755);
and (n7872,n308,n33);
and (n7873,n7874,n7875);
xor (n7874,n7871,n7872);
or (n7875,n7876,n7879);
and (n7876,n7877,n7878);
xor (n7877,n7760,n7761);
and (n7878,n51,n33);
and (n7879,n7880,n7881);
xor (n7880,n7877,n7878);
or (n7881,n7882,n7885);
and (n7882,n7883,n7884);
xor (n7883,n7766,n7767);
and (n7884,n45,n33);
and (n7885,n7886,n7887);
xor (n7886,n7883,n7884);
or (n7887,n7888,n7891);
and (n7888,n7889,n7890);
xor (n7889,n7772,n7773);
and (n7890,n75,n33);
and (n7891,n7892,n7893);
xor (n7892,n7889,n7890);
or (n7893,n7894,n7897);
and (n7894,n7895,n7896);
xor (n7895,n7778,n7779);
and (n7896,n69,n33);
and (n7897,n7898,n7899);
xor (n7898,n7895,n7896);
or (n7899,n7900,n7903);
and (n7900,n7901,n7902);
xor (n7901,n7784,n7785);
and (n7902,n226,n33);
and (n7903,n7904,n7905);
xor (n7904,n7901,n7902);
or (n7905,n7906,n7909);
and (n7906,n7907,n7908);
xor (n7907,n7790,n7791);
and (n7908,n351,n33);
and (n7909,n7910,n7911);
xor (n7910,n7907,n7908);
or (n7911,n7912,n7915);
and (n7912,n7913,n7914);
xor (n7913,n7796,n7797);
and (n7914,n345,n33);
and (n7915,n7916,n7917);
xor (n7916,n7913,n7914);
or (n7917,n7918,n7921);
and (n7918,n7919,n7920);
xor (n7919,n7802,n7803);
and (n7920,n372,n33);
and (n7921,n7922,n7923);
xor (n7922,n7919,n7920);
or (n7923,n7924,n7927);
and (n7924,n7925,n7926);
xor (n7925,n7808,n7809);
and (n7926,n281,n33);
and (n7927,n7928,n7929);
xor (n7928,n7925,n7926);
or (n7929,n7930,n7933);
and (n7930,n7931,n7932);
xor (n7931,n7813,n7814);
and (n7932,n185,n33);
and (n7933,n7934,n7935);
xor (n7934,n7931,n7932);
or (n7935,n7936,n7939);
and (n7936,n7937,n7938);
xor (n7937,n7818,n7819);
and (n7938,n179,n33);
and (n7939,n7940,n7941);
xor (n7940,n7937,n7938);
or (n7941,n7942,n7945);
and (n7942,n7943,n7944);
xor (n7943,n7824,n7825);
and (n7944,n289,n33);
and (n7945,n7946,n7947);
xor (n7946,n7943,n7944);
or (n7947,n7948,n7951);
and (n7948,n7949,n7950);
xor (n7949,n7830,n7831);
and (n7950,n545,n33);
and (n7951,n7952,n7953);
xor (n7952,n7949,n7950);
or (n7953,n7954,n7957);
and (n7954,n7955,n7956);
xor (n7955,n7836,n7837);
and (n7956,n719,n33);
and (n7957,n7958,n7959);
xor (n7958,n7955,n7956);
or (n7959,n7960,n7963);
and (n7960,n7961,n7962);
xor (n7961,n7842,n7843);
and (n7962,n837,n33);
and (n7963,n7964,n7965);
xor (n7964,n7961,n7962);
or (n7965,n7966,n7969);
and (n7966,n7967,n7968);
xor (n7967,n7847,n7848);
and (n7968,n1175,n33);
and (n7969,n7970,n7971);
xor (n7970,n7967,n7968);
or (n7971,n7972,n7975);
and (n7972,n7973,n7974);
xor (n7973,n7852,n7853);
and (n7974,n1147,n33);
and (n7975,n7976,n7977);
xor (n7976,n7973,n7974);
or (n7977,n7978,n7981);
and (n7978,n7979,n7980);
xor (n7979,n7858,n7859);
and (n7980,n1141,n33);
and (n7981,n7982,n7983);
xor (n7982,n7979,n7980);
and (n7983,n7984,n3040);
xor (n7984,n7864,n7865);
and (n7985,n308,n34);
or (n7986,n7987,n7990);
and (n7987,n7988,n7989);
xor (n7988,n7874,n7875);
and (n7989,n51,n34);
and (n7990,n7991,n7992);
xor (n7991,n7988,n7989);
or (n7992,n7993,n7996);
and (n7993,n7994,n7995);
xor (n7994,n7880,n7881);
and (n7995,n45,n34);
and (n7996,n7997,n7998);
xor (n7997,n7994,n7995);
or (n7998,n7999,n8002);
and (n7999,n8000,n8001);
xor (n8000,n7886,n7887);
and (n8001,n75,n34);
and (n8002,n8003,n8004);
xor (n8003,n8000,n8001);
or (n8004,n8005,n8008);
and (n8005,n8006,n8007);
xor (n8006,n7892,n7893);
and (n8007,n69,n34);
and (n8008,n8009,n8010);
xor (n8009,n8006,n8007);
or (n8010,n8011,n8014);
and (n8011,n8012,n8013);
xor (n8012,n7898,n7899);
and (n8013,n226,n34);
and (n8014,n8015,n8016);
xor (n8015,n8012,n8013);
or (n8016,n8017,n8020);
and (n8017,n8018,n8019);
xor (n8018,n7904,n7905);
and (n8019,n351,n34);
and (n8020,n8021,n8022);
xor (n8021,n8018,n8019);
or (n8022,n8023,n8026);
and (n8023,n8024,n8025);
xor (n8024,n7910,n7911);
and (n8025,n345,n34);
and (n8026,n8027,n8028);
xor (n8027,n8024,n8025);
or (n8028,n8029,n8032);
and (n8029,n8030,n8031);
xor (n8030,n7916,n7917);
and (n8031,n372,n34);
and (n8032,n8033,n8034);
xor (n8033,n8030,n8031);
or (n8034,n8035,n8038);
and (n8035,n8036,n8037);
xor (n8036,n7922,n7923);
and (n8037,n281,n34);
and (n8038,n8039,n8040);
xor (n8039,n8036,n8037);
or (n8040,n8041,n8044);
and (n8041,n8042,n8043);
xor (n8042,n7928,n7929);
and (n8043,n185,n34);
and (n8044,n8045,n8046);
xor (n8045,n8042,n8043);
or (n8046,n8047,n8050);
and (n8047,n8048,n8049);
xor (n8048,n7934,n7935);
and (n8049,n179,n34);
and (n8050,n8051,n8052);
xor (n8051,n8048,n8049);
or (n8052,n8053,n8056);
and (n8053,n8054,n8055);
xor (n8054,n7940,n7941);
and (n8055,n289,n34);
and (n8056,n8057,n8058);
xor (n8057,n8054,n8055);
or (n8058,n8059,n8062);
and (n8059,n8060,n8061);
xor (n8060,n7946,n7947);
and (n8061,n545,n34);
and (n8062,n8063,n8064);
xor (n8063,n8060,n8061);
or (n8064,n8065,n8068);
and (n8065,n8066,n8067);
xor (n8066,n7952,n7953);
and (n8067,n719,n34);
and (n8068,n8069,n8070);
xor (n8069,n8066,n8067);
or (n8070,n8071,n8074);
and (n8071,n8072,n8073);
xor (n8072,n7958,n7959);
and (n8073,n837,n34);
and (n8074,n8075,n8076);
xor (n8075,n8072,n8073);
or (n8076,n8077,n8080);
and (n8077,n8078,n8079);
xor (n8078,n7964,n7965);
and (n8079,n1175,n34);
and (n8080,n8081,n8082);
xor (n8081,n8078,n8079);
or (n8082,n8083,n8086);
and (n8083,n8084,n8085);
xor (n8084,n7970,n7971);
and (n8085,n1147,n34);
and (n8086,n8087,n8088);
xor (n8087,n8084,n8085);
or (n8088,n8089,n8092);
and (n8089,n8090,n8091);
xor (n8090,n7976,n7977);
and (n8091,n1141,n34);
and (n8092,n8093,n8094);
xor (n8093,n8090,n8091);
and (n8094,n8095,n8096);
xor (n8095,n7982,n7983);
and (n8096,n1187,n34);
and (n8097,n51,n59);
or (n8098,n8099,n8102);
and (n8099,n8100,n8101);
xor (n8100,n7991,n7992);
and (n8101,n45,n59);
and (n8102,n8103,n8104);
xor (n8103,n8100,n8101);
or (n8104,n8105,n8108);
and (n8105,n8106,n8107);
xor (n8106,n7997,n7998);
and (n8107,n75,n59);
and (n8108,n8109,n8110);
xor (n8109,n8106,n8107);
or (n8110,n8111,n8114);
and (n8111,n8112,n8113);
xor (n8112,n8003,n8004);
and (n8113,n69,n59);
and (n8114,n8115,n8116);
xor (n8115,n8112,n8113);
or (n8116,n8117,n8120);
and (n8117,n8118,n8119);
xor (n8118,n8009,n8010);
and (n8119,n226,n59);
and (n8120,n8121,n8122);
xor (n8121,n8118,n8119);
or (n8122,n8123,n8126);
and (n8123,n8124,n8125);
xor (n8124,n8015,n8016);
and (n8125,n351,n59);
and (n8126,n8127,n8128);
xor (n8127,n8124,n8125);
or (n8128,n8129,n8132);
and (n8129,n8130,n8131);
xor (n8130,n8021,n8022);
and (n8131,n345,n59);
and (n8132,n8133,n8134);
xor (n8133,n8130,n8131);
or (n8134,n8135,n8138);
and (n8135,n8136,n8137);
xor (n8136,n8027,n8028);
and (n8137,n372,n59);
and (n8138,n8139,n8140);
xor (n8139,n8136,n8137);
or (n8140,n8141,n8144);
and (n8141,n8142,n8143);
xor (n8142,n8033,n8034);
and (n8143,n281,n59);
and (n8144,n8145,n8146);
xor (n8145,n8142,n8143);
or (n8146,n8147,n8150);
and (n8147,n8148,n8149);
xor (n8148,n8039,n8040);
and (n8149,n185,n59);
and (n8150,n8151,n8152);
xor (n8151,n8148,n8149);
or (n8152,n8153,n8156);
and (n8153,n8154,n8155);
xor (n8154,n8045,n8046);
and (n8155,n179,n59);
and (n8156,n8157,n8158);
xor (n8157,n8154,n8155);
or (n8158,n8159,n8162);
and (n8159,n8160,n8161);
xor (n8160,n8051,n8052);
and (n8161,n289,n59);
and (n8162,n8163,n8164);
xor (n8163,n8160,n8161);
or (n8164,n8165,n8168);
and (n8165,n8166,n8167);
xor (n8166,n8057,n8058);
and (n8167,n545,n59);
and (n8168,n8169,n8170);
xor (n8169,n8166,n8167);
or (n8170,n8171,n8174);
and (n8171,n8172,n8173);
xor (n8172,n8063,n8064);
and (n8173,n719,n59);
and (n8174,n8175,n8176);
xor (n8175,n8172,n8173);
or (n8176,n8177,n8180);
and (n8177,n8178,n8179);
xor (n8178,n8069,n8070);
and (n8179,n837,n59);
and (n8180,n8181,n8182);
xor (n8181,n8178,n8179);
or (n8182,n8183,n8186);
and (n8183,n8184,n8185);
xor (n8184,n8075,n8076);
and (n8185,n1175,n59);
and (n8186,n8187,n8188);
xor (n8187,n8184,n8185);
or (n8188,n8189,n8192);
and (n8189,n8190,n8191);
xor (n8190,n8081,n8082);
and (n8191,n1147,n59);
and (n8192,n8193,n8194);
xor (n8193,n8190,n8191);
or (n8194,n8195,n8198);
and (n8195,n8196,n8197);
xor (n8196,n8087,n8088);
and (n8197,n1141,n59);
and (n8198,n8199,n8200);
xor (n8199,n8196,n8197);
and (n8200,n8201,n8202);
xor (n8201,n8093,n8094);
not (n8202,n3786);
and (n8203,n45,n65);
or (n8204,n8205,n8208);
and (n8205,n8206,n8207);
xor (n8206,n8103,n8104);
and (n8207,n75,n65);
and (n8208,n8209,n8210);
xor (n8209,n8206,n8207);
or (n8210,n8211,n8214);
and (n8211,n8212,n8213);
xor (n8212,n8109,n8110);
and (n8213,n69,n65);
and (n8214,n8215,n8216);
xor (n8215,n8212,n8213);
or (n8216,n8217,n8220);
and (n8217,n8218,n8219);
xor (n8218,n8115,n8116);
and (n8219,n226,n65);
and (n8220,n8221,n8222);
xor (n8221,n8218,n8219);
or (n8222,n8223,n8226);
and (n8223,n8224,n8225);
xor (n8224,n8121,n8122);
and (n8225,n351,n65);
and (n8226,n8227,n8228);
xor (n8227,n8224,n8225);
or (n8228,n8229,n8232);
and (n8229,n8230,n8231);
xor (n8230,n8127,n8128);
and (n8231,n345,n65);
and (n8232,n8233,n8234);
xor (n8233,n8230,n8231);
or (n8234,n8235,n8238);
and (n8235,n8236,n8237);
xor (n8236,n8133,n8134);
and (n8237,n372,n65);
and (n8238,n8239,n8240);
xor (n8239,n8236,n8237);
or (n8240,n8241,n8244);
and (n8241,n8242,n8243);
xor (n8242,n8139,n8140);
and (n8243,n281,n65);
and (n8244,n8245,n8246);
xor (n8245,n8242,n8243);
or (n8246,n8247,n8250);
and (n8247,n8248,n8249);
xor (n8248,n8145,n8146);
and (n8249,n185,n65);
and (n8250,n8251,n8252);
xor (n8251,n8248,n8249);
or (n8252,n8253,n8256);
and (n8253,n8254,n8255);
xor (n8254,n8151,n8152);
and (n8255,n179,n65);
and (n8256,n8257,n8258);
xor (n8257,n8254,n8255);
or (n8258,n8259,n8262);
and (n8259,n8260,n8261);
xor (n8260,n8157,n8158);
and (n8261,n289,n65);
and (n8262,n8263,n8264);
xor (n8263,n8260,n8261);
or (n8264,n8265,n8268);
and (n8265,n8266,n8267);
xor (n8266,n8163,n8164);
and (n8267,n545,n65);
and (n8268,n8269,n8270);
xor (n8269,n8266,n8267);
or (n8270,n8271,n8274);
and (n8271,n8272,n8273);
xor (n8272,n8169,n8170);
and (n8273,n719,n65);
and (n8274,n8275,n8276);
xor (n8275,n8272,n8273);
or (n8276,n8277,n8280);
and (n8277,n8278,n8279);
xor (n8278,n8175,n8176);
and (n8279,n837,n65);
and (n8280,n8281,n8282);
xor (n8281,n8278,n8279);
or (n8282,n8283,n8286);
and (n8283,n8284,n8285);
xor (n8284,n8181,n8182);
and (n8285,n1175,n65);
and (n8286,n8287,n8288);
xor (n8287,n8284,n8285);
or (n8288,n8289,n8292);
and (n8289,n8290,n8291);
xor (n8290,n8187,n8188);
and (n8291,n1147,n65);
and (n8292,n8293,n8294);
xor (n8293,n8290,n8291);
or (n8294,n8295,n8298);
and (n8295,n8296,n8297);
xor (n8296,n8193,n8194);
and (n8297,n1141,n65);
and (n8298,n8299,n8300);
xor (n8299,n8296,n8297);
and (n8300,n8301,n8302);
xor (n8301,n8199,n8200);
and (n8302,n1187,n65);
and (n8303,n75,n215);
or (n8304,n8305,n8308);
and (n8305,n8306,n8307);
xor (n8306,n8209,n8210);
and (n8307,n69,n215);
and (n8308,n8309,n8310);
xor (n8309,n8306,n8307);
or (n8310,n8311,n8314);
and (n8311,n8312,n8313);
xor (n8312,n8215,n8216);
and (n8313,n226,n215);
and (n8314,n8315,n8316);
xor (n8315,n8312,n8313);
or (n8316,n8317,n8320);
and (n8317,n8318,n8319);
xor (n8318,n8221,n8222);
and (n8319,n351,n215);
and (n8320,n8321,n8322);
xor (n8321,n8318,n8319);
or (n8322,n8323,n8326);
and (n8323,n8324,n8325);
xor (n8324,n8227,n8228);
and (n8325,n345,n215);
and (n8326,n8327,n8328);
xor (n8327,n8324,n8325);
or (n8328,n8329,n8332);
and (n8329,n8330,n8331);
xor (n8330,n8233,n8234);
and (n8331,n372,n215);
and (n8332,n8333,n8334);
xor (n8333,n8330,n8331);
or (n8334,n8335,n8338);
and (n8335,n8336,n8337);
xor (n8336,n8239,n8240);
and (n8337,n281,n215);
and (n8338,n8339,n8340);
xor (n8339,n8336,n8337);
or (n8340,n8341,n8344);
and (n8341,n8342,n8343);
xor (n8342,n8245,n8246);
and (n8343,n185,n215);
and (n8344,n8345,n8346);
xor (n8345,n8342,n8343);
or (n8346,n8347,n8350);
and (n8347,n8348,n8349);
xor (n8348,n8251,n8252);
and (n8349,n179,n215);
and (n8350,n8351,n8352);
xor (n8351,n8348,n8349);
or (n8352,n8353,n8356);
and (n8353,n8354,n8355);
xor (n8354,n8257,n8258);
and (n8355,n289,n215);
and (n8356,n8357,n8358);
xor (n8357,n8354,n8355);
or (n8358,n8359,n8362);
and (n8359,n8360,n8361);
xor (n8360,n8263,n8264);
and (n8361,n545,n215);
and (n8362,n8363,n8364);
xor (n8363,n8360,n8361);
or (n8364,n8365,n8368);
and (n8365,n8366,n8367);
xor (n8366,n8269,n8270);
and (n8367,n719,n215);
and (n8368,n8369,n8370);
xor (n8369,n8366,n8367);
or (n8370,n8371,n8374);
and (n8371,n8372,n8373);
xor (n8372,n8275,n8276);
and (n8373,n837,n215);
and (n8374,n8375,n8376);
xor (n8375,n8372,n8373);
or (n8376,n8377,n8380);
and (n8377,n8378,n8379);
xor (n8378,n8281,n8282);
and (n8379,n1175,n215);
and (n8380,n8381,n8382);
xor (n8381,n8378,n8379);
or (n8382,n8383,n8386);
and (n8383,n8384,n8385);
xor (n8384,n8287,n8288);
and (n8385,n1147,n215);
and (n8386,n8387,n8388);
xor (n8387,n8384,n8385);
or (n8388,n8389,n8392);
and (n8389,n8390,n8391);
xor (n8390,n8293,n8294);
and (n8391,n1141,n215);
and (n8392,n8393,n8394);
xor (n8393,n8390,n8391);
and (n8394,n8395,n8396);
xor (n8395,n8299,n8300);
not (n8396,n2555);
and (n8397,n69,n209);
or (n8398,n8399,n8402);
and (n8399,n8400,n8401);
xor (n8400,n8309,n8310);
and (n8401,n226,n209);
and (n8402,n8403,n8404);
xor (n8403,n8400,n8401);
or (n8404,n8405,n8408);
and (n8405,n8406,n8407);
xor (n8406,n8315,n8316);
and (n8407,n351,n209);
and (n8408,n8409,n8410);
xor (n8409,n8406,n8407);
or (n8410,n8411,n8414);
and (n8411,n8412,n8413);
xor (n8412,n8321,n8322);
and (n8413,n345,n209);
and (n8414,n8415,n8416);
xor (n8415,n8412,n8413);
or (n8416,n8417,n8420);
and (n8417,n8418,n8419);
xor (n8418,n8327,n8328);
and (n8419,n372,n209);
and (n8420,n8421,n8422);
xor (n8421,n8418,n8419);
or (n8422,n8423,n8425);
and (n8423,n8424,n777);
xor (n8424,n8333,n8334);
and (n8425,n8426,n8427);
xor (n8426,n8424,n777);
or (n8427,n8428,n8430);
and (n8428,n8429,n885);
xor (n8429,n8339,n8340);
and (n8430,n8431,n8432);
xor (n8431,n8429,n885);
or (n8432,n8433,n8436);
and (n8433,n8434,n8435);
xor (n8434,n8345,n8346);
and (n8435,n179,n209);
and (n8436,n8437,n8438);
xor (n8437,n8434,n8435);
or (n8438,n8439,n8442);
and (n8439,n8440,n8441);
xor (n8440,n8351,n8352);
and (n8441,n289,n209);
and (n8442,n8443,n8444);
xor (n8443,n8440,n8441);
or (n8444,n8445,n8448);
and (n8445,n8446,n8447);
xor (n8446,n8357,n8358);
and (n8447,n545,n209);
and (n8448,n8449,n8450);
xor (n8449,n8446,n8447);
or (n8450,n8451,n8454);
and (n8451,n8452,n8453);
xor (n8452,n8363,n8364);
and (n8453,n719,n209);
and (n8454,n8455,n8456);
xor (n8455,n8452,n8453);
or (n8456,n8457,n8460);
and (n8457,n8458,n8459);
xor (n8458,n8369,n8370);
and (n8459,n837,n209);
and (n8460,n8461,n8462);
xor (n8461,n8458,n8459);
or (n8462,n8463,n8466);
and (n8463,n8464,n8465);
xor (n8464,n8375,n8376);
and (n8465,n1175,n209);
and (n8466,n8467,n8468);
xor (n8467,n8464,n8465);
or (n8468,n8469,n8472);
and (n8469,n8470,n8471);
xor (n8470,n8381,n8382);
and (n8471,n1147,n209);
and (n8472,n8473,n8474);
xor (n8473,n8470,n8471);
or (n8474,n8475,n8478);
and (n8475,n8476,n8477);
xor (n8476,n8387,n8388);
and (n8477,n1141,n209);
and (n8478,n8479,n8480);
xor (n8479,n8476,n8477);
and (n8480,n8481,n8482);
xor (n8481,n8393,n8394);
and (n8482,n1187,n209);
and (n8483,n226,n360);
or (n8484,n8485,n8488);
and (n8485,n8486,n8487);
xor (n8486,n8403,n8404);
and (n8487,n351,n360);
and (n8488,n8489,n8490);
xor (n8489,n8486,n8487);
or (n8490,n8491,n8494);
and (n8491,n8492,n8493);
xor (n8492,n8409,n8410);
and (n8493,n345,n360);
and (n8494,n8495,n8496);
xor (n8495,n8492,n8493);
or (n8496,n8497,n8500);
and (n8497,n8498,n8499);
xor (n8498,n8415,n8416);
and (n8499,n372,n360);
and (n8500,n8501,n8502);
xor (n8501,n8498,n8499);
or (n8502,n8503,n8506);
and (n8503,n8504,n8505);
xor (n8504,n8421,n8422);
and (n8505,n281,n360);
and (n8506,n8507,n8508);
xor (n8507,n8504,n8505);
or (n8508,n8509,n8512);
and (n8509,n8510,n8511);
xor (n8510,n8426,n8427);
and (n8511,n185,n360);
and (n8512,n8513,n8514);
xor (n8513,n8510,n8511);
or (n8514,n8515,n8518);
and (n8515,n8516,n8517);
xor (n8516,n8431,n8432);
and (n8517,n179,n360);
and (n8518,n8519,n8520);
xor (n8519,n8516,n8517);
or (n8520,n8521,n8524);
and (n8521,n8522,n8523);
xor (n8522,n8437,n8438);
and (n8523,n289,n360);
and (n8524,n8525,n8526);
xor (n8525,n8522,n8523);
or (n8526,n8527,n8530);
and (n8527,n8528,n8529);
xor (n8528,n8443,n8444);
and (n8529,n545,n360);
and (n8530,n8531,n8532);
xor (n8531,n8528,n8529);
or (n8532,n8533,n8536);
and (n8533,n8534,n8535);
xor (n8534,n8449,n8450);
and (n8535,n719,n360);
and (n8536,n8537,n8538);
xor (n8537,n8534,n8535);
or (n8538,n8539,n8542);
and (n8539,n8540,n8541);
xor (n8540,n8455,n8456);
and (n8541,n837,n360);
and (n8542,n8543,n8544);
xor (n8543,n8540,n8541);
or (n8544,n8545,n8548);
and (n8545,n8546,n8547);
xor (n8546,n8461,n8462);
and (n8547,n1175,n360);
and (n8548,n8549,n8550);
xor (n8549,n8546,n8547);
or (n8550,n8551,n8554);
and (n8551,n8552,n8553);
xor (n8552,n8467,n8468);
and (n8553,n1147,n360);
and (n8554,n8555,n8556);
xor (n8555,n8552,n8553);
or (n8556,n8557,n8560);
and (n8557,n8558,n8559);
xor (n8558,n8473,n8474);
and (n8559,n1141,n360);
and (n8560,n8561,n8562);
xor (n8561,n8558,n8559);
and (n8562,n8563,n2085);
xor (n8563,n8479,n8480);
and (n8564,n351,n272);
or (n8565,n8566,n8569);
and (n8566,n8567,n8568);
xor (n8567,n8489,n8490);
and (n8568,n345,n272);
and (n8569,n8570,n8571);
xor (n8570,n8567,n8568);
or (n8571,n8572,n8575);
and (n8572,n8573,n8574);
xor (n8573,n8495,n8496);
and (n8574,n372,n272);
and (n8575,n8576,n8577);
xor (n8576,n8573,n8574);
or (n8577,n8578,n8581);
and (n8578,n8579,n8580);
xor (n8579,n8501,n8502);
and (n8580,n281,n272);
and (n8581,n8582,n8583);
xor (n8582,n8579,n8580);
or (n8583,n8584,n8587);
and (n8584,n8585,n8586);
xor (n8585,n8507,n8508);
and (n8586,n185,n272);
and (n8587,n8588,n8589);
xor (n8588,n8585,n8586);
or (n8589,n8590,n8593);
and (n8590,n8591,n8592);
xor (n8591,n8513,n8514);
and (n8592,n179,n272);
and (n8593,n8594,n8595);
xor (n8594,n8591,n8592);
or (n8595,n8596,n8599);
and (n8596,n8597,n8598);
xor (n8597,n8519,n8520);
and (n8598,n289,n272);
and (n8599,n8600,n8601);
xor (n8600,n8597,n8598);
or (n8601,n8602,n8605);
and (n8602,n8603,n8604);
xor (n8603,n8525,n8526);
and (n8604,n545,n272);
and (n8605,n8606,n8607);
xor (n8606,n8603,n8604);
or (n8607,n8608,n8611);
and (n8608,n8609,n8610);
xor (n8609,n8531,n8532);
and (n8610,n719,n272);
and (n8611,n8612,n8613);
xor (n8612,n8609,n8610);
or (n8613,n8614,n8617);
and (n8614,n8615,n8616);
xor (n8615,n8537,n8538);
and (n8616,n837,n272);
and (n8617,n8618,n8619);
xor (n8618,n8615,n8616);
or (n8619,n8620,n8623);
and (n8620,n8621,n8622);
xor (n8621,n8543,n8544);
and (n8622,n1175,n272);
and (n8623,n8624,n8625);
xor (n8624,n8621,n8622);
or (n8625,n8626,n8629);
and (n8626,n8627,n8628);
xor (n8627,n8549,n8550);
and (n8628,n1147,n272);
and (n8629,n8630,n8631);
xor (n8630,n8627,n8628);
or (n8631,n8632,n8635);
and (n8632,n8633,n8634);
xor (n8633,n8555,n8556);
and (n8634,n1141,n272);
and (n8635,n8636,n8637);
xor (n8636,n8633,n8634);
and (n8637,n8638,n8639);
xor (n8638,n8561,n8562);
and (n8639,n1187,n272);
and (n8640,n345,n270);
or (n8641,n8642,n8645);
and (n8642,n8643,n8644);
xor (n8643,n8570,n8571);
and (n8644,n372,n270);
and (n8645,n8646,n8647);
xor (n8646,n8643,n8644);
or (n8647,n8648,n8651);
and (n8648,n8649,n8650);
xor (n8649,n8576,n8577);
and (n8650,n281,n270);
and (n8651,n8652,n8653);
xor (n8652,n8649,n8650);
or (n8653,n8654,n8657);
and (n8654,n8655,n8656);
xor (n8655,n8582,n8583);
and (n8656,n185,n270);
and (n8657,n8658,n8659);
xor (n8658,n8655,n8656);
or (n8659,n8660,n8663);
and (n8660,n8661,n8662);
xor (n8661,n8588,n8589);
and (n8662,n179,n270);
and (n8663,n8664,n8665);
xor (n8664,n8661,n8662);
or (n8665,n8666,n8669);
and (n8666,n8667,n8668);
xor (n8667,n8594,n8595);
and (n8668,n289,n270);
and (n8669,n8670,n8671);
xor (n8670,n8667,n8668);
or (n8671,n8672,n8675);
and (n8672,n8673,n8674);
xor (n8673,n8600,n8601);
and (n8674,n545,n270);
and (n8675,n8676,n8677);
xor (n8676,n8673,n8674);
or (n8677,n8678,n8681);
and (n8678,n8679,n8680);
xor (n8679,n8606,n8607);
and (n8680,n719,n270);
and (n8681,n8682,n8683);
xor (n8682,n8679,n8680);
or (n8683,n8684,n8687);
and (n8684,n8685,n8686);
xor (n8685,n8612,n8613);
and (n8686,n837,n270);
and (n8687,n8688,n8689);
xor (n8688,n8685,n8686);
or (n8689,n8690,n8693);
and (n8690,n8691,n8692);
xor (n8691,n8618,n8619);
and (n8692,n1175,n270);
and (n8693,n8694,n8695);
xor (n8694,n8691,n8692);
or (n8695,n8696,n8699);
and (n8696,n8697,n8698);
xor (n8697,n8624,n8625);
and (n8698,n1147,n270);
and (n8699,n8700,n8701);
xor (n8700,n8697,n8698);
or (n8701,n8702,n8705);
and (n8702,n8703,n8704);
xor (n8703,n8630,n8631);
and (n8704,n1141,n270);
and (n8705,n8706,n8707);
xor (n8706,n8703,n8704);
and (n8707,n8708,n8709);
xor (n8708,n8636,n8637);
not (n8709,n1779);
and (n8710,n372,n168);
or (n8711,n8712,n8715);
and (n8712,n8713,n8714);
xor (n8713,n8646,n8647);
and (n8714,n281,n168);
and (n8715,n8716,n8717);
xor (n8716,n8713,n8714);
or (n8717,n8718,n8721);
and (n8718,n8719,n8720);
xor (n8719,n8652,n8653);
and (n8720,n185,n168);
and (n8721,n8722,n8723);
xor (n8722,n8719,n8720);
or (n8723,n8724,n8727);
and (n8724,n8725,n8726);
xor (n8725,n8658,n8659);
and (n8726,n179,n168);
and (n8727,n8728,n8729);
xor (n8728,n8725,n8726);
or (n8729,n8730,n8733);
and (n8730,n8731,n8732);
xor (n8731,n8664,n8665);
and (n8732,n289,n168);
and (n8733,n8734,n8735);
xor (n8734,n8731,n8732);
or (n8735,n8736,n8739);
and (n8736,n8737,n8738);
xor (n8737,n8670,n8671);
and (n8738,n545,n168);
and (n8739,n8740,n8741);
xor (n8740,n8737,n8738);
or (n8741,n8742,n8745);
and (n8742,n8743,n8744);
xor (n8743,n8676,n8677);
and (n8744,n719,n168);
and (n8745,n8746,n8747);
xor (n8746,n8743,n8744);
or (n8747,n8748,n8751);
and (n8748,n8749,n8750);
xor (n8749,n8682,n8683);
and (n8750,n837,n168);
and (n8751,n8752,n8753);
xor (n8752,n8749,n8750);
or (n8753,n8754,n8757);
and (n8754,n8755,n8756);
xor (n8755,n8688,n8689);
and (n8756,n1175,n168);
and (n8757,n8758,n8759);
xor (n8758,n8755,n8756);
or (n8759,n8760,n8763);
and (n8760,n8761,n8762);
xor (n8761,n8694,n8695);
and (n8762,n1147,n168);
and (n8763,n8764,n8765);
xor (n8764,n8761,n8762);
or (n8765,n8766,n8769);
and (n8766,n8767,n8768);
xor (n8767,n8700,n8701);
and (n8768,n1141,n168);
and (n8769,n8770,n8771);
xor (n8770,n8767,n8768);
and (n8771,n8772,n8773);
xor (n8772,n8706,n8707);
and (n8773,n1187,n168);
and (n8774,n281,n169);
or (n8775,n8776,n8779);
and (n8776,n8777,n8778);
xor (n8777,n8716,n8717);
and (n8778,n185,n169);
and (n8779,n8780,n8781);
xor (n8780,n8777,n8778);
or (n8781,n8782,n8785);
and (n8782,n8783,n8784);
xor (n8783,n8722,n8723);
and (n8784,n179,n169);
and (n8785,n8786,n8787);
xor (n8786,n8783,n8784);
or (n8787,n8788,n8791);
and (n8788,n8789,n8790);
xor (n8789,n8728,n8729);
and (n8790,n289,n169);
and (n8791,n8792,n8793);
xor (n8792,n8789,n8790);
or (n8793,n8794,n8797);
and (n8794,n8795,n8796);
xor (n8795,n8734,n8735);
and (n8796,n545,n169);
and (n8797,n8798,n8799);
xor (n8798,n8795,n8796);
or (n8799,n8800,n8803);
and (n8800,n8801,n8802);
xor (n8801,n8740,n8741);
and (n8802,n719,n169);
and (n8803,n8804,n8805);
xor (n8804,n8801,n8802);
or (n8805,n8806,n8809);
and (n8806,n8807,n8808);
xor (n8807,n8746,n8747);
and (n8808,n837,n169);
and (n8809,n8810,n8811);
xor (n8810,n8807,n8808);
or (n8811,n8812,n8815);
and (n8812,n8813,n8814);
xor (n8813,n8752,n8753);
and (n8814,n1175,n169);
and (n8815,n8816,n8817);
xor (n8816,n8813,n8814);
or (n8817,n8818,n8821);
and (n8818,n8819,n8820);
xor (n8819,n8758,n8759);
and (n8820,n1147,n169);
and (n8821,n8822,n8823);
xor (n8822,n8819,n8820);
or (n8823,n8824,n8827);
and (n8824,n8825,n8826);
xor (n8825,n8764,n8765);
and (n8826,n1141,n169);
and (n8827,n8828,n8829);
xor (n8828,n8825,n8826);
and (n8829,n8830,n8831);
xor (n8830,n8770,n8771);
not (n8831,n1186);
and (n8832,n185,n175);
or (n8833,n8834,n8837);
and (n8834,n8835,n8836);
xor (n8835,n8780,n8781);
and (n8836,n179,n175);
and (n8837,n8838,n8839);
xor (n8838,n8835,n8836);
or (n8839,n8840,n8843);
and (n8840,n8841,n8842);
xor (n8841,n8786,n8787);
and (n8842,n289,n175);
and (n8843,n8844,n8845);
xor (n8844,n8841,n8842);
or (n8845,n8846,n8849);
and (n8846,n8847,n8848);
xor (n8847,n8792,n8793);
and (n8848,n545,n175);
and (n8849,n8850,n8851);
xor (n8850,n8847,n8848);
or (n8851,n8852,n8855);
and (n8852,n8853,n8854);
xor (n8853,n8798,n8799);
and (n8854,n719,n175);
and (n8855,n8856,n8857);
xor (n8856,n8853,n8854);
or (n8857,n8858,n8861);
and (n8858,n8859,n8860);
xor (n8859,n8804,n8805);
and (n8860,n837,n175);
and (n8861,n8862,n8863);
xor (n8862,n8859,n8860);
or (n8863,n8864,n8867);
and (n8864,n8865,n8866);
xor (n8865,n8810,n8811);
and (n8866,n1175,n175);
and (n8867,n8868,n8869);
xor (n8868,n8865,n8866);
or (n8869,n8870,n8873);
and (n8870,n8871,n8872);
xor (n8871,n8816,n8817);
and (n8872,n1147,n175);
and (n8873,n8874,n8875);
xor (n8874,n8871,n8872);
or (n8875,n8876,n8879);
and (n8876,n8877,n8878);
xor (n8877,n8822,n8823);
and (n8878,n1141,n175);
and (n8879,n8880,n8881);
xor (n8880,n8877,n8878);
and (n8881,n8882,n8883);
xor (n8882,n8828,n8829);
and (n8883,n1187,n175);
or (n8884,n8885,n8887);
and (n8885,n8886,n8842);
xor (n8886,n8838,n8839);
and (n8887,n8888,n8889);
xor (n8888,n8886,n8842);
or (n8889,n8890,n8892);
and (n8890,n8891,n8848);
xor (n8891,n8844,n8845);
and (n8892,n8893,n8894);
xor (n8893,n8891,n8848);
or (n8894,n8895,n8897);
and (n8895,n8896,n8854);
xor (n8896,n8850,n8851);
and (n8897,n8898,n8899);
xor (n8898,n8896,n8854);
or (n8899,n8900,n8902);
and (n8900,n8901,n8860);
xor (n8901,n8856,n8857);
and (n8902,n8903,n8904);
xor (n8903,n8901,n8860);
or (n8904,n8905,n8907);
and (n8905,n8906,n8866);
xor (n8906,n8862,n8863);
and (n8907,n8908,n8909);
xor (n8908,n8906,n8866);
or (n8909,n8910,n8912);
and (n8910,n8911,n8872);
xor (n8911,n8868,n8869);
and (n8912,n8913,n8914);
xor (n8913,n8911,n8872);
or (n8914,n8915,n8917);
and (n8915,n8916,n8878);
xor (n8916,n8874,n8875);
and (n8917,n8918,n8919);
xor (n8918,n8916,n8878);
and (n8919,n8920,n8883);
xor (n8920,n8880,n8881);
or (n8921,n8922,n8924);
and (n8922,n8923,n8848);
xor (n8923,n8888,n8889);
and (n8924,n8925,n8926);
xor (n8925,n8923,n8848);
or (n8926,n8927,n8929);
and (n8927,n8928,n8854);
xor (n8928,n8893,n8894);
and (n8929,n8930,n8931);
xor (n8930,n8928,n8854);
or (n8931,n8932,n8934);
and (n8932,n8933,n8860);
xor (n8933,n8898,n8899);
and (n8934,n8935,n8936);
xor (n8935,n8933,n8860);
or (n8936,n8937,n8939);
and (n8937,n8938,n8866);
xor (n8938,n8903,n8904);
and (n8939,n8940,n8941);
xor (n8940,n8938,n8866);
or (n8941,n8942,n8944);
and (n8942,n8943,n8872);
xor (n8943,n8908,n8909);
and (n8944,n8945,n8946);
xor (n8945,n8943,n8872);
or (n8946,n8947,n8949);
and (n8947,n8948,n8878);
xor (n8948,n8913,n8914);
and (n8949,n8950,n8951);
xor (n8950,n8948,n8878);
and (n8951,n8952,n8883);
xor (n8952,n8918,n8919);
or (n8953,n8954,n8956);
and (n8954,n8955,n8854);
xor (n8955,n8925,n8926);
and (n8956,n8957,n8958);
xor (n8957,n8955,n8854);
or (n8958,n8959,n8961);
and (n8959,n8960,n8860);
xor (n8960,n8930,n8931);
and (n8961,n8962,n8963);
xor (n8962,n8960,n8860);
or (n8963,n8964,n8966);
and (n8964,n8965,n8866);
xor (n8965,n8935,n8936);
and (n8966,n8967,n8968);
xor (n8967,n8965,n8866);
or (n8968,n8969,n8971);
and (n8969,n8970,n8872);
xor (n8970,n8940,n8941);
and (n8971,n8972,n8973);
xor (n8972,n8970,n8872);
or (n8973,n8974,n8976);
and (n8974,n8975,n8878);
xor (n8975,n8945,n8946);
and (n8976,n8977,n8978);
xor (n8977,n8975,n8878);
and (n8978,n8979,n8883);
xor (n8979,n8950,n8951);
or (n8980,n8981,n8983);
and (n8981,n8982,n8860);
xor (n8982,n8957,n8958);
and (n8983,n8984,n8985);
xor (n8984,n8982,n8860);
or (n8985,n8986,n8988);
and (n8986,n8987,n8866);
xor (n8987,n8962,n8963);
and (n8988,n8989,n8990);
xor (n8989,n8987,n8866);
or (n8990,n8991,n8993);
and (n8991,n8992,n8872);
xor (n8992,n8967,n8968);
and (n8993,n8994,n8995);
xor (n8994,n8992,n8872);
or (n8995,n8996,n8998);
and (n8996,n8997,n8878);
xor (n8997,n8972,n8973);
and (n8998,n8999,n9000);
xor (n8999,n8997,n8878);
and (n9000,n9001,n8883);
xor (n9001,n8977,n8978);
or (n9002,n9003,n9005);
and (n9003,n9004,n8866);
xor (n9004,n8984,n8985);
and (n9005,n9006,n9007);
xor (n9006,n9004,n8866);
or (n9007,n9008,n9010);
and (n9008,n9009,n8872);
xor (n9009,n8989,n8990);
and (n9010,n9011,n9012);
xor (n9011,n9009,n8872);
or (n9012,n9013,n9015);
and (n9013,n9014,n8878);
xor (n9014,n8994,n8995);
and (n9015,n9016,n9017);
xor (n9016,n9014,n8878);
and (n9017,n9018,n8883);
xor (n9018,n8999,n9000);
or (n9019,n9020,n9022);
and (n9020,n9021,n8872);
xor (n9021,n9006,n9007);
and (n9022,n9023,n9024);
xor (n9023,n9021,n8872);
or (n9024,n9025,n9027);
and (n9025,n9026,n8878);
xor (n9026,n9011,n9012);
and (n9027,n9028,n9029);
xor (n9028,n9026,n8878);
and (n9029,n9030,n8883);
xor (n9030,n9016,n9017);
or (n9031,n9032,n9034);
and (n9032,n9033,n8878);
xor (n9033,n9023,n9024);
and (n9034,n9035,n9036);
xor (n9035,n9033,n8878);
and (n9036,n9037,n8883);
xor (n9037,n9028,n9029);
and (n9038,n9039,n8883);
xor (n9039,n9035,n9036);
nor (n9040,n9,n7);
and (n9041,n3,n9042);
not (n9042,n9040);
endmodule
