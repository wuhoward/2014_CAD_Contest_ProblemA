module top (out,n23,n24,n28,n30,n37,n44,n51,n58,n65
        ,n72,n79,n86,n93,n99,n101,n168,n235,n302,n367
        ,n426,n479,n526,n567,n602,n652,n653,n657,n659,n666
        ,n673,n680,n687,n694,n701,n708,n715,n722,n728,n730
        ,n797,n864,n931,n996,n1055,n1108,n1155,n1196,n1231,n1259);
output out;
input n23;
input n24;
input n28;
input n30;
input n37;
input n44;
input n51;
input n58;
input n65;
input n72;
input n79;
input n86;
input n93;
input n99;
input n101;
input n168;
input n235;
input n302;
input n367;
input n426;
input n479;
input n526;
input n567;
input n602;
input n652;
input n653;
input n657;
input n659;
input n666;
input n673;
input n680;
input n687;
input n694;
input n701;
input n708;
input n715;
input n722;
input n728;
input n730;
input n797;
input n864;
input n931;
input n996;
input n1055;
input n1108;
input n1155;
input n1196;
input n1231;
input n1259;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n25;
wire n26;
wire n27;
wire n29;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n100;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n654;
wire n655;
wire n656;
wire n658;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n729;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
xor (out,n0,n1260);
wire s0n0,s1n0,notn0;
or (n0,s0n0,s1n0);
not(notn0,n1259);
and (s0n0,notn0,n1);
and (s1n0,n1259,n630);
xor (n1,n2,n603);
xor (n2,n3,n601);
xor (n3,n4,n568);
xor (n4,n5,n566);
xor (n5,n6,n527);
xor (n6,n7,n525);
xor (n7,n8,n480);
xor (n8,n9,n478);
xor (n9,n10,n427);
xor (n10,n11,n425);
xor (n11,n12,n368);
xor (n12,n13,n366);
xor (n13,n14,n303);
xor (n14,n15,n301);
or (n15,n16,n236);
and (n16,n17,n234);
or (n17,n18,n169);
and (n18,n19,n167);
or (n19,n20,n102);
and (n20,n21,n100);
and (n21,n22,n25);
and (n22,n23,n24);
or (n25,n26,n31);
and (n26,n27,n29);
and (n27,n23,n28);
and (n29,n30,n24);
and (n31,n32,n33);
xor (n32,n27,n29);
or (n33,n34,n38);
and (n34,n35,n36);
and (n35,n30,n28);
and (n36,n37,n24);
and (n38,n39,n40);
xor (n39,n35,n36);
or (n40,n41,n45);
and (n41,n42,n43);
and (n42,n37,n28);
and (n43,n44,n24);
and (n45,n46,n47);
xor (n46,n42,n43);
or (n47,n48,n52);
and (n48,n49,n50);
and (n49,n44,n28);
and (n50,n51,n24);
and (n52,n53,n54);
xor (n53,n49,n50);
or (n54,n55,n59);
and (n55,n56,n57);
and (n56,n51,n28);
and (n57,n58,n24);
and (n59,n60,n61);
xor (n60,n56,n57);
or (n61,n62,n66);
and (n62,n63,n64);
and (n63,n58,n28);
and (n64,n65,n24);
and (n66,n67,n68);
xor (n67,n63,n64);
or (n68,n69,n73);
and (n69,n70,n71);
and (n70,n65,n28);
and (n71,n72,n24);
and (n73,n74,n75);
xor (n74,n70,n71);
or (n75,n76,n80);
and (n76,n77,n78);
and (n77,n72,n28);
and (n78,n79,n24);
and (n80,n81,n82);
xor (n81,n77,n78);
or (n82,n83,n87);
and (n83,n84,n85);
and (n84,n79,n28);
and (n85,n86,n24);
and (n87,n88,n89);
xor (n88,n84,n85);
or (n89,n90,n94);
and (n90,n91,n92);
and (n91,n86,n28);
and (n92,n93,n24);
and (n94,n95,n96);
xor (n95,n91,n92);
and (n96,n97,n98);
and (n97,n93,n28);
and (n98,n99,n24);
and (n100,n23,n101);
and (n102,n103,n104);
xor (n103,n21,n100);
or (n104,n105,n108);
and (n105,n106,n107);
xor (n106,n22,n25);
and (n107,n30,n101);
and (n108,n109,n110);
xor (n109,n106,n107);
or (n110,n111,n114);
and (n111,n112,n113);
xor (n112,n32,n33);
and (n113,n37,n101);
and (n114,n115,n116);
xor (n115,n112,n113);
or (n116,n117,n120);
and (n117,n118,n119);
xor (n118,n39,n40);
and (n119,n44,n101);
and (n120,n121,n122);
xor (n121,n118,n119);
or (n122,n123,n126);
and (n123,n124,n125);
xor (n124,n46,n47);
and (n125,n51,n101);
and (n126,n127,n128);
xor (n127,n124,n125);
or (n128,n129,n132);
and (n129,n130,n131);
xor (n130,n53,n54);
and (n131,n58,n101);
and (n132,n133,n134);
xor (n133,n130,n131);
or (n134,n135,n138);
and (n135,n136,n137);
xor (n136,n60,n61);
and (n137,n65,n101);
and (n138,n139,n140);
xor (n139,n136,n137);
or (n140,n141,n144);
and (n141,n142,n143);
xor (n142,n67,n68);
and (n143,n72,n101);
and (n144,n145,n146);
xor (n145,n142,n143);
or (n146,n147,n150);
and (n147,n148,n149);
xor (n148,n74,n75);
and (n149,n79,n101);
and (n150,n151,n152);
xor (n151,n148,n149);
or (n152,n153,n156);
and (n153,n154,n155);
xor (n154,n81,n82);
and (n155,n86,n101);
and (n156,n157,n158);
xor (n157,n154,n155);
or (n158,n159,n162);
and (n159,n160,n161);
xor (n160,n88,n89);
and (n161,n93,n101);
and (n162,n163,n164);
xor (n163,n160,n161);
and (n164,n165,n166);
xor (n165,n95,n96);
and (n166,n99,n101);
and (n167,n23,n168);
and (n169,n170,n171);
xor (n170,n19,n167);
or (n171,n172,n175);
and (n172,n173,n174);
xor (n173,n103,n104);
and (n174,n30,n168);
and (n175,n176,n177);
xor (n176,n173,n174);
or (n177,n178,n181);
and (n178,n179,n180);
xor (n179,n109,n110);
and (n180,n37,n168);
and (n181,n182,n183);
xor (n182,n179,n180);
or (n183,n184,n187);
and (n184,n185,n186);
xor (n185,n115,n116);
and (n186,n44,n168);
and (n187,n188,n189);
xor (n188,n185,n186);
or (n189,n190,n193);
and (n190,n191,n192);
xor (n191,n121,n122);
and (n192,n51,n168);
and (n193,n194,n195);
xor (n194,n191,n192);
or (n195,n196,n199);
and (n196,n197,n198);
xor (n197,n127,n128);
and (n198,n58,n168);
and (n199,n200,n201);
xor (n200,n197,n198);
or (n201,n202,n205);
and (n202,n203,n204);
xor (n203,n133,n134);
and (n204,n65,n168);
and (n205,n206,n207);
xor (n206,n203,n204);
or (n207,n208,n211);
and (n208,n209,n210);
xor (n209,n139,n140);
and (n210,n72,n168);
and (n211,n212,n213);
xor (n212,n209,n210);
or (n213,n214,n217);
and (n214,n215,n216);
xor (n215,n145,n146);
and (n216,n79,n168);
and (n217,n218,n219);
xor (n218,n215,n216);
or (n219,n220,n223);
and (n220,n221,n222);
xor (n221,n151,n152);
and (n222,n86,n168);
and (n223,n224,n225);
xor (n224,n221,n222);
or (n225,n226,n229);
and (n226,n227,n228);
xor (n227,n157,n158);
and (n228,n93,n168);
and (n229,n230,n231);
xor (n230,n227,n228);
and (n231,n232,n233);
xor (n232,n163,n164);
and (n233,n99,n168);
and (n234,n23,n235);
and (n236,n237,n238);
xor (n237,n17,n234);
or (n238,n239,n242);
and (n239,n240,n241);
xor (n240,n170,n171);
and (n241,n30,n235);
and (n242,n243,n244);
xor (n243,n240,n241);
or (n244,n245,n248);
and (n245,n246,n247);
xor (n246,n176,n177);
and (n247,n37,n235);
and (n248,n249,n250);
xor (n249,n246,n247);
or (n250,n251,n254);
and (n251,n252,n253);
xor (n252,n182,n183);
and (n253,n44,n235);
and (n254,n255,n256);
xor (n255,n252,n253);
or (n256,n257,n260);
and (n257,n258,n259);
xor (n258,n188,n189);
and (n259,n51,n235);
and (n260,n261,n262);
xor (n261,n258,n259);
or (n262,n263,n266);
and (n263,n264,n265);
xor (n264,n194,n195);
and (n265,n58,n235);
and (n266,n267,n268);
xor (n267,n264,n265);
or (n268,n269,n272);
and (n269,n270,n271);
xor (n270,n200,n201);
and (n271,n65,n235);
and (n272,n273,n274);
xor (n273,n270,n271);
or (n274,n275,n278);
and (n275,n276,n277);
xor (n276,n206,n207);
and (n277,n72,n235);
and (n278,n279,n280);
xor (n279,n276,n277);
or (n280,n281,n284);
and (n281,n282,n283);
xor (n282,n212,n213);
and (n283,n79,n235);
and (n284,n285,n286);
xor (n285,n282,n283);
or (n286,n287,n290);
and (n287,n288,n289);
xor (n288,n218,n219);
and (n289,n86,n235);
and (n290,n291,n292);
xor (n291,n288,n289);
or (n292,n293,n296);
and (n293,n294,n295);
xor (n294,n224,n225);
and (n295,n93,n235);
and (n296,n297,n298);
xor (n297,n294,n295);
and (n298,n299,n300);
xor (n299,n230,n231);
and (n300,n99,n235);
and (n301,n23,n302);
or (n303,n304,n307);
and (n304,n305,n306);
xor (n305,n237,n238);
and (n306,n30,n302);
and (n307,n308,n309);
xor (n308,n305,n306);
or (n309,n310,n313);
and (n310,n311,n312);
xor (n311,n243,n244);
and (n312,n37,n302);
and (n313,n314,n315);
xor (n314,n311,n312);
or (n315,n316,n319);
and (n316,n317,n318);
xor (n317,n249,n250);
and (n318,n44,n302);
and (n319,n320,n321);
xor (n320,n317,n318);
or (n321,n322,n325);
and (n322,n323,n324);
xor (n323,n255,n256);
and (n324,n51,n302);
and (n325,n326,n327);
xor (n326,n323,n324);
or (n327,n328,n331);
and (n328,n329,n330);
xor (n329,n261,n262);
and (n330,n58,n302);
and (n331,n332,n333);
xor (n332,n329,n330);
or (n333,n334,n337);
and (n334,n335,n336);
xor (n335,n267,n268);
and (n336,n65,n302);
and (n337,n338,n339);
xor (n338,n335,n336);
or (n339,n340,n343);
and (n340,n341,n342);
xor (n341,n273,n274);
and (n342,n72,n302);
and (n343,n344,n345);
xor (n344,n341,n342);
or (n345,n346,n349);
and (n346,n347,n348);
xor (n347,n279,n280);
and (n348,n79,n302);
and (n349,n350,n351);
xor (n350,n347,n348);
or (n351,n352,n355);
and (n352,n353,n354);
xor (n353,n285,n286);
and (n354,n86,n302);
and (n355,n356,n357);
xor (n356,n353,n354);
or (n357,n358,n361);
and (n358,n359,n360);
xor (n359,n291,n292);
and (n360,n93,n302);
and (n361,n362,n363);
xor (n362,n359,n360);
and (n363,n364,n365);
xor (n364,n297,n298);
and (n365,n99,n302);
and (n366,n30,n367);
or (n368,n369,n372);
and (n369,n370,n371);
xor (n370,n308,n309);
and (n371,n37,n367);
and (n372,n373,n374);
xor (n373,n370,n371);
or (n374,n375,n378);
and (n375,n376,n377);
xor (n376,n314,n315);
and (n377,n44,n367);
and (n378,n379,n380);
xor (n379,n376,n377);
or (n380,n381,n384);
and (n381,n382,n383);
xor (n382,n320,n321);
and (n383,n51,n367);
and (n384,n385,n386);
xor (n385,n382,n383);
or (n386,n387,n390);
and (n387,n388,n389);
xor (n388,n326,n327);
and (n389,n58,n367);
and (n390,n391,n392);
xor (n391,n388,n389);
or (n392,n393,n396);
and (n393,n394,n395);
xor (n394,n332,n333);
and (n395,n65,n367);
and (n396,n397,n398);
xor (n397,n394,n395);
or (n398,n399,n402);
and (n399,n400,n401);
xor (n400,n338,n339);
and (n401,n72,n367);
and (n402,n403,n404);
xor (n403,n400,n401);
or (n404,n405,n408);
and (n405,n406,n407);
xor (n406,n344,n345);
and (n407,n79,n367);
and (n408,n409,n410);
xor (n409,n406,n407);
or (n410,n411,n414);
and (n411,n412,n413);
xor (n412,n350,n351);
and (n413,n86,n367);
and (n414,n415,n416);
xor (n415,n412,n413);
or (n416,n417,n420);
and (n417,n418,n419);
xor (n418,n356,n357);
and (n419,n93,n367);
and (n420,n421,n422);
xor (n421,n418,n419);
and (n422,n423,n424);
xor (n423,n362,n363);
and (n424,n99,n367);
and (n425,n37,n426);
or (n427,n428,n431);
and (n428,n429,n430);
xor (n429,n373,n374);
and (n430,n44,n426);
and (n431,n432,n433);
xor (n432,n429,n430);
or (n433,n434,n437);
and (n434,n435,n436);
xor (n435,n379,n380);
and (n436,n51,n426);
and (n437,n438,n439);
xor (n438,n435,n436);
or (n439,n440,n443);
and (n440,n441,n442);
xor (n441,n385,n386);
and (n442,n58,n426);
and (n443,n444,n445);
xor (n444,n441,n442);
or (n445,n446,n449);
and (n446,n447,n448);
xor (n447,n391,n392);
and (n448,n65,n426);
and (n449,n450,n451);
xor (n450,n447,n448);
or (n451,n452,n455);
and (n452,n453,n454);
xor (n453,n397,n398);
and (n454,n72,n426);
and (n455,n456,n457);
xor (n456,n453,n454);
or (n457,n458,n461);
and (n458,n459,n460);
xor (n459,n403,n404);
and (n460,n79,n426);
and (n461,n462,n463);
xor (n462,n459,n460);
or (n463,n464,n467);
and (n464,n465,n466);
xor (n465,n409,n410);
and (n466,n86,n426);
and (n467,n468,n469);
xor (n468,n465,n466);
or (n469,n470,n473);
and (n470,n471,n472);
xor (n471,n415,n416);
and (n472,n93,n426);
and (n473,n474,n475);
xor (n474,n471,n472);
and (n475,n476,n477);
xor (n476,n421,n422);
and (n477,n99,n426);
and (n478,n44,n479);
or (n480,n481,n484);
and (n481,n482,n483);
xor (n482,n432,n433);
and (n483,n51,n479);
and (n484,n485,n486);
xor (n485,n482,n483);
or (n486,n487,n490);
and (n487,n488,n489);
xor (n488,n438,n439);
and (n489,n58,n479);
and (n490,n491,n492);
xor (n491,n488,n489);
or (n492,n493,n496);
and (n493,n494,n495);
xor (n494,n444,n445);
and (n495,n65,n479);
and (n496,n497,n498);
xor (n497,n494,n495);
or (n498,n499,n502);
and (n499,n500,n501);
xor (n500,n450,n451);
and (n501,n72,n479);
and (n502,n503,n504);
xor (n503,n500,n501);
or (n504,n505,n508);
and (n505,n506,n507);
xor (n506,n456,n457);
and (n507,n79,n479);
and (n508,n509,n510);
xor (n509,n506,n507);
or (n510,n511,n514);
and (n511,n512,n513);
xor (n512,n462,n463);
and (n513,n86,n479);
and (n514,n515,n516);
xor (n515,n512,n513);
or (n516,n517,n520);
and (n517,n518,n519);
xor (n518,n468,n469);
and (n519,n93,n479);
and (n520,n521,n522);
xor (n521,n518,n519);
and (n522,n523,n524);
xor (n523,n474,n475);
and (n524,n99,n479);
and (n525,n51,n526);
or (n527,n528,n531);
and (n528,n529,n530);
xor (n529,n485,n486);
and (n530,n58,n526);
and (n531,n532,n533);
xor (n532,n529,n530);
or (n533,n534,n537);
and (n534,n535,n536);
xor (n535,n491,n492);
and (n536,n65,n526);
and (n537,n538,n539);
xor (n538,n535,n536);
or (n539,n540,n543);
and (n540,n541,n542);
xor (n541,n497,n498);
and (n542,n72,n526);
and (n543,n544,n545);
xor (n544,n541,n542);
or (n545,n546,n549);
and (n546,n547,n548);
xor (n547,n503,n504);
and (n548,n79,n526);
and (n549,n550,n551);
xor (n550,n547,n548);
or (n551,n552,n555);
and (n552,n553,n554);
xor (n553,n509,n510);
and (n554,n86,n526);
and (n555,n556,n557);
xor (n556,n553,n554);
or (n557,n558,n561);
and (n558,n559,n560);
xor (n559,n515,n516);
and (n560,n93,n526);
and (n561,n562,n563);
xor (n562,n559,n560);
and (n563,n564,n565);
xor (n564,n521,n522);
and (n565,n99,n526);
and (n566,n58,n567);
or (n568,n569,n572);
and (n569,n570,n571);
xor (n570,n532,n533);
and (n571,n65,n567);
and (n572,n573,n574);
xor (n573,n570,n571);
or (n574,n575,n578);
and (n575,n576,n577);
xor (n576,n538,n539);
and (n577,n72,n567);
and (n578,n579,n580);
xor (n579,n576,n577);
or (n580,n581,n584);
and (n581,n582,n583);
xor (n582,n544,n545);
and (n583,n79,n567);
and (n584,n585,n586);
xor (n585,n582,n583);
or (n586,n587,n590);
and (n587,n588,n589);
xor (n588,n550,n551);
and (n589,n86,n567);
and (n590,n591,n592);
xor (n591,n588,n589);
or (n592,n593,n596);
and (n593,n594,n595);
xor (n594,n556,n557);
and (n595,n93,n567);
and (n596,n597,n598);
xor (n597,n594,n595);
and (n598,n599,n600);
xor (n599,n562,n563);
and (n600,n99,n567);
and (n601,n65,n602);
or (n603,n604,n607);
and (n604,n605,n606);
xor (n605,n573,n574);
and (n606,n72,n602);
and (n607,n608,n609);
xor (n608,n605,n606);
or (n609,n610,n613);
and (n610,n611,n612);
xor (n611,n579,n580);
and (n612,n79,n602);
and (n613,n614,n615);
xor (n614,n611,n612);
or (n615,n616,n619);
and (n616,n617,n618);
xor (n617,n585,n586);
and (n618,n86,n602);
and (n619,n620,n621);
xor (n620,n617,n618);
or (n621,n622,n625);
and (n622,n623,n624);
xor (n623,n591,n592);
and (n624,n93,n602);
and (n625,n626,n627);
xor (n626,n623,n624);
and (n627,n628,n629);
xor (n628,n597,n598);
and (n629,n99,n602);
xor (n630,n631,n1232);
xor (n631,n632,n1230);
xor (n632,n633,n1197);
xor (n633,n634,n1195);
xor (n634,n635,n1156);
xor (n635,n636,n1154);
xor (n636,n637,n1109);
xor (n637,n638,n1107);
xor (n638,n639,n1056);
xor (n639,n640,n1054);
xor (n640,n641,n997);
xor (n641,n642,n995);
xor (n642,n643,n932);
xor (n643,n644,n930);
or (n644,n645,n865);
and (n645,n646,n863);
or (n646,n647,n798);
and (n647,n648,n796);
or (n648,n649,n731);
and (n649,n650,n729);
and (n650,n651,n654);
and (n651,n652,n653);
or (n654,n655,n660);
and (n655,n656,n658);
and (n656,n652,n657);
and (n658,n659,n653);
and (n660,n661,n662);
xor (n661,n656,n658);
or (n662,n663,n667);
and (n663,n664,n665);
and (n664,n659,n657);
and (n665,n666,n653);
and (n667,n668,n669);
xor (n668,n664,n665);
or (n669,n670,n674);
and (n670,n671,n672);
and (n671,n666,n657);
and (n672,n673,n653);
and (n674,n675,n676);
xor (n675,n671,n672);
or (n676,n677,n681);
and (n677,n678,n679);
and (n678,n673,n657);
and (n679,n680,n653);
and (n681,n682,n683);
xor (n682,n678,n679);
or (n683,n684,n688);
and (n684,n685,n686);
and (n685,n680,n657);
and (n686,n687,n653);
and (n688,n689,n690);
xor (n689,n685,n686);
or (n690,n691,n695);
and (n691,n692,n693);
and (n692,n687,n657);
and (n693,n694,n653);
and (n695,n696,n697);
xor (n696,n692,n693);
or (n697,n698,n702);
and (n698,n699,n700);
and (n699,n694,n657);
and (n700,n701,n653);
and (n702,n703,n704);
xor (n703,n699,n700);
or (n704,n705,n709);
and (n705,n706,n707);
and (n706,n701,n657);
and (n707,n708,n653);
and (n709,n710,n711);
xor (n710,n706,n707);
or (n711,n712,n716);
and (n712,n713,n714);
and (n713,n708,n657);
and (n714,n715,n653);
and (n716,n717,n718);
xor (n717,n713,n714);
or (n718,n719,n723);
and (n719,n720,n721);
and (n720,n715,n657);
and (n721,n722,n653);
and (n723,n724,n725);
xor (n724,n720,n721);
and (n725,n726,n727);
and (n726,n722,n657);
and (n727,n728,n653);
and (n729,n652,n730);
and (n731,n732,n733);
xor (n732,n650,n729);
or (n733,n734,n737);
and (n734,n735,n736);
xor (n735,n651,n654);
and (n736,n659,n730);
and (n737,n738,n739);
xor (n738,n735,n736);
or (n739,n740,n743);
and (n740,n741,n742);
xor (n741,n661,n662);
and (n742,n666,n730);
and (n743,n744,n745);
xor (n744,n741,n742);
or (n745,n746,n749);
and (n746,n747,n748);
xor (n747,n668,n669);
and (n748,n673,n730);
and (n749,n750,n751);
xor (n750,n747,n748);
or (n751,n752,n755);
and (n752,n753,n754);
xor (n753,n675,n676);
and (n754,n680,n730);
and (n755,n756,n757);
xor (n756,n753,n754);
or (n757,n758,n761);
and (n758,n759,n760);
xor (n759,n682,n683);
and (n760,n687,n730);
and (n761,n762,n763);
xor (n762,n759,n760);
or (n763,n764,n767);
and (n764,n765,n766);
xor (n765,n689,n690);
and (n766,n694,n730);
and (n767,n768,n769);
xor (n768,n765,n766);
or (n769,n770,n773);
and (n770,n771,n772);
xor (n771,n696,n697);
and (n772,n701,n730);
and (n773,n774,n775);
xor (n774,n771,n772);
or (n775,n776,n779);
and (n776,n777,n778);
xor (n777,n703,n704);
and (n778,n708,n730);
and (n779,n780,n781);
xor (n780,n777,n778);
or (n781,n782,n785);
and (n782,n783,n784);
xor (n783,n710,n711);
and (n784,n715,n730);
and (n785,n786,n787);
xor (n786,n783,n784);
or (n787,n788,n791);
and (n788,n789,n790);
xor (n789,n717,n718);
and (n790,n722,n730);
and (n791,n792,n793);
xor (n792,n789,n790);
and (n793,n794,n795);
xor (n794,n724,n725);
and (n795,n728,n730);
and (n796,n652,n797);
and (n798,n799,n800);
xor (n799,n648,n796);
or (n800,n801,n804);
and (n801,n802,n803);
xor (n802,n732,n733);
and (n803,n659,n797);
and (n804,n805,n806);
xor (n805,n802,n803);
or (n806,n807,n810);
and (n807,n808,n809);
xor (n808,n738,n739);
and (n809,n666,n797);
and (n810,n811,n812);
xor (n811,n808,n809);
or (n812,n813,n816);
and (n813,n814,n815);
xor (n814,n744,n745);
and (n815,n673,n797);
and (n816,n817,n818);
xor (n817,n814,n815);
or (n818,n819,n822);
and (n819,n820,n821);
xor (n820,n750,n751);
and (n821,n680,n797);
and (n822,n823,n824);
xor (n823,n820,n821);
or (n824,n825,n828);
and (n825,n826,n827);
xor (n826,n756,n757);
and (n827,n687,n797);
and (n828,n829,n830);
xor (n829,n826,n827);
or (n830,n831,n834);
and (n831,n832,n833);
xor (n832,n762,n763);
and (n833,n694,n797);
and (n834,n835,n836);
xor (n835,n832,n833);
or (n836,n837,n840);
and (n837,n838,n839);
xor (n838,n768,n769);
and (n839,n701,n797);
and (n840,n841,n842);
xor (n841,n838,n839);
or (n842,n843,n846);
and (n843,n844,n845);
xor (n844,n774,n775);
and (n845,n708,n797);
and (n846,n847,n848);
xor (n847,n844,n845);
or (n848,n849,n852);
and (n849,n850,n851);
xor (n850,n780,n781);
and (n851,n715,n797);
and (n852,n853,n854);
xor (n853,n850,n851);
or (n854,n855,n858);
and (n855,n856,n857);
xor (n856,n786,n787);
and (n857,n722,n797);
and (n858,n859,n860);
xor (n859,n856,n857);
and (n860,n861,n862);
xor (n861,n792,n793);
and (n862,n728,n797);
and (n863,n652,n864);
and (n865,n866,n867);
xor (n866,n646,n863);
or (n867,n868,n871);
and (n868,n869,n870);
xor (n869,n799,n800);
and (n870,n659,n864);
and (n871,n872,n873);
xor (n872,n869,n870);
or (n873,n874,n877);
and (n874,n875,n876);
xor (n875,n805,n806);
and (n876,n666,n864);
and (n877,n878,n879);
xor (n878,n875,n876);
or (n879,n880,n883);
and (n880,n881,n882);
xor (n881,n811,n812);
and (n882,n673,n864);
and (n883,n884,n885);
xor (n884,n881,n882);
or (n885,n886,n889);
and (n886,n887,n888);
xor (n887,n817,n818);
and (n888,n680,n864);
and (n889,n890,n891);
xor (n890,n887,n888);
or (n891,n892,n895);
and (n892,n893,n894);
xor (n893,n823,n824);
and (n894,n687,n864);
and (n895,n896,n897);
xor (n896,n893,n894);
or (n897,n898,n901);
and (n898,n899,n900);
xor (n899,n829,n830);
and (n900,n694,n864);
and (n901,n902,n903);
xor (n902,n899,n900);
or (n903,n904,n907);
and (n904,n905,n906);
xor (n905,n835,n836);
and (n906,n701,n864);
and (n907,n908,n909);
xor (n908,n905,n906);
or (n909,n910,n913);
and (n910,n911,n912);
xor (n911,n841,n842);
and (n912,n708,n864);
and (n913,n914,n915);
xor (n914,n911,n912);
or (n915,n916,n919);
and (n916,n917,n918);
xor (n917,n847,n848);
and (n918,n715,n864);
and (n919,n920,n921);
xor (n920,n917,n918);
or (n921,n922,n925);
and (n922,n923,n924);
xor (n923,n853,n854);
and (n924,n722,n864);
and (n925,n926,n927);
xor (n926,n923,n924);
and (n927,n928,n929);
xor (n928,n859,n860);
and (n929,n728,n864);
and (n930,n652,n931);
or (n932,n933,n936);
and (n933,n934,n935);
xor (n934,n866,n867);
and (n935,n659,n931);
and (n936,n937,n938);
xor (n937,n934,n935);
or (n938,n939,n942);
and (n939,n940,n941);
xor (n940,n872,n873);
and (n941,n666,n931);
and (n942,n943,n944);
xor (n943,n940,n941);
or (n944,n945,n948);
and (n945,n946,n947);
xor (n946,n878,n879);
and (n947,n673,n931);
and (n948,n949,n950);
xor (n949,n946,n947);
or (n950,n951,n954);
and (n951,n952,n953);
xor (n952,n884,n885);
and (n953,n680,n931);
and (n954,n955,n956);
xor (n955,n952,n953);
or (n956,n957,n960);
and (n957,n958,n959);
xor (n958,n890,n891);
and (n959,n687,n931);
and (n960,n961,n962);
xor (n961,n958,n959);
or (n962,n963,n966);
and (n963,n964,n965);
xor (n964,n896,n897);
and (n965,n694,n931);
and (n966,n967,n968);
xor (n967,n964,n965);
or (n968,n969,n972);
and (n969,n970,n971);
xor (n970,n902,n903);
and (n971,n701,n931);
and (n972,n973,n974);
xor (n973,n970,n971);
or (n974,n975,n978);
and (n975,n976,n977);
xor (n976,n908,n909);
and (n977,n708,n931);
and (n978,n979,n980);
xor (n979,n976,n977);
or (n980,n981,n984);
and (n981,n982,n983);
xor (n982,n914,n915);
and (n983,n715,n931);
and (n984,n985,n986);
xor (n985,n982,n983);
or (n986,n987,n990);
and (n987,n988,n989);
xor (n988,n920,n921);
and (n989,n722,n931);
and (n990,n991,n992);
xor (n991,n988,n989);
and (n992,n993,n994);
xor (n993,n926,n927);
and (n994,n728,n931);
and (n995,n659,n996);
or (n997,n998,n1001);
and (n998,n999,n1000);
xor (n999,n937,n938);
and (n1000,n666,n996);
and (n1001,n1002,n1003);
xor (n1002,n999,n1000);
or (n1003,n1004,n1007);
and (n1004,n1005,n1006);
xor (n1005,n943,n944);
and (n1006,n673,n996);
and (n1007,n1008,n1009);
xor (n1008,n1005,n1006);
or (n1009,n1010,n1013);
and (n1010,n1011,n1012);
xor (n1011,n949,n950);
and (n1012,n680,n996);
and (n1013,n1014,n1015);
xor (n1014,n1011,n1012);
or (n1015,n1016,n1019);
and (n1016,n1017,n1018);
xor (n1017,n955,n956);
and (n1018,n687,n996);
and (n1019,n1020,n1021);
xor (n1020,n1017,n1018);
or (n1021,n1022,n1025);
and (n1022,n1023,n1024);
xor (n1023,n961,n962);
and (n1024,n694,n996);
and (n1025,n1026,n1027);
xor (n1026,n1023,n1024);
or (n1027,n1028,n1031);
and (n1028,n1029,n1030);
xor (n1029,n967,n968);
and (n1030,n701,n996);
and (n1031,n1032,n1033);
xor (n1032,n1029,n1030);
or (n1033,n1034,n1037);
and (n1034,n1035,n1036);
xor (n1035,n973,n974);
and (n1036,n708,n996);
and (n1037,n1038,n1039);
xor (n1038,n1035,n1036);
or (n1039,n1040,n1043);
and (n1040,n1041,n1042);
xor (n1041,n979,n980);
and (n1042,n715,n996);
and (n1043,n1044,n1045);
xor (n1044,n1041,n1042);
or (n1045,n1046,n1049);
and (n1046,n1047,n1048);
xor (n1047,n985,n986);
and (n1048,n722,n996);
and (n1049,n1050,n1051);
xor (n1050,n1047,n1048);
and (n1051,n1052,n1053);
xor (n1052,n991,n992);
and (n1053,n728,n996);
and (n1054,n666,n1055);
or (n1056,n1057,n1060);
and (n1057,n1058,n1059);
xor (n1058,n1002,n1003);
and (n1059,n673,n1055);
and (n1060,n1061,n1062);
xor (n1061,n1058,n1059);
or (n1062,n1063,n1066);
and (n1063,n1064,n1065);
xor (n1064,n1008,n1009);
and (n1065,n680,n1055);
and (n1066,n1067,n1068);
xor (n1067,n1064,n1065);
or (n1068,n1069,n1072);
and (n1069,n1070,n1071);
xor (n1070,n1014,n1015);
and (n1071,n687,n1055);
and (n1072,n1073,n1074);
xor (n1073,n1070,n1071);
or (n1074,n1075,n1078);
and (n1075,n1076,n1077);
xor (n1076,n1020,n1021);
and (n1077,n694,n1055);
and (n1078,n1079,n1080);
xor (n1079,n1076,n1077);
or (n1080,n1081,n1084);
and (n1081,n1082,n1083);
xor (n1082,n1026,n1027);
and (n1083,n701,n1055);
and (n1084,n1085,n1086);
xor (n1085,n1082,n1083);
or (n1086,n1087,n1090);
and (n1087,n1088,n1089);
xor (n1088,n1032,n1033);
and (n1089,n708,n1055);
and (n1090,n1091,n1092);
xor (n1091,n1088,n1089);
or (n1092,n1093,n1096);
and (n1093,n1094,n1095);
xor (n1094,n1038,n1039);
and (n1095,n715,n1055);
and (n1096,n1097,n1098);
xor (n1097,n1094,n1095);
or (n1098,n1099,n1102);
and (n1099,n1100,n1101);
xor (n1100,n1044,n1045);
and (n1101,n722,n1055);
and (n1102,n1103,n1104);
xor (n1103,n1100,n1101);
and (n1104,n1105,n1106);
xor (n1105,n1050,n1051);
and (n1106,n728,n1055);
and (n1107,n673,n1108);
or (n1109,n1110,n1113);
and (n1110,n1111,n1112);
xor (n1111,n1061,n1062);
and (n1112,n680,n1108);
and (n1113,n1114,n1115);
xor (n1114,n1111,n1112);
or (n1115,n1116,n1119);
and (n1116,n1117,n1118);
xor (n1117,n1067,n1068);
and (n1118,n687,n1108);
and (n1119,n1120,n1121);
xor (n1120,n1117,n1118);
or (n1121,n1122,n1125);
and (n1122,n1123,n1124);
xor (n1123,n1073,n1074);
and (n1124,n694,n1108);
and (n1125,n1126,n1127);
xor (n1126,n1123,n1124);
or (n1127,n1128,n1131);
and (n1128,n1129,n1130);
xor (n1129,n1079,n1080);
and (n1130,n701,n1108);
and (n1131,n1132,n1133);
xor (n1132,n1129,n1130);
or (n1133,n1134,n1137);
and (n1134,n1135,n1136);
xor (n1135,n1085,n1086);
and (n1136,n708,n1108);
and (n1137,n1138,n1139);
xor (n1138,n1135,n1136);
or (n1139,n1140,n1143);
and (n1140,n1141,n1142);
xor (n1141,n1091,n1092);
and (n1142,n715,n1108);
and (n1143,n1144,n1145);
xor (n1144,n1141,n1142);
or (n1145,n1146,n1149);
and (n1146,n1147,n1148);
xor (n1147,n1097,n1098);
and (n1148,n722,n1108);
and (n1149,n1150,n1151);
xor (n1150,n1147,n1148);
and (n1151,n1152,n1153);
xor (n1152,n1103,n1104);
and (n1153,n728,n1108);
and (n1154,n680,n1155);
or (n1156,n1157,n1160);
and (n1157,n1158,n1159);
xor (n1158,n1114,n1115);
and (n1159,n687,n1155);
and (n1160,n1161,n1162);
xor (n1161,n1158,n1159);
or (n1162,n1163,n1166);
and (n1163,n1164,n1165);
xor (n1164,n1120,n1121);
and (n1165,n694,n1155);
and (n1166,n1167,n1168);
xor (n1167,n1164,n1165);
or (n1168,n1169,n1172);
and (n1169,n1170,n1171);
xor (n1170,n1126,n1127);
and (n1171,n701,n1155);
and (n1172,n1173,n1174);
xor (n1173,n1170,n1171);
or (n1174,n1175,n1178);
and (n1175,n1176,n1177);
xor (n1176,n1132,n1133);
and (n1177,n708,n1155);
and (n1178,n1179,n1180);
xor (n1179,n1176,n1177);
or (n1180,n1181,n1184);
and (n1181,n1182,n1183);
xor (n1182,n1138,n1139);
and (n1183,n715,n1155);
and (n1184,n1185,n1186);
xor (n1185,n1182,n1183);
or (n1186,n1187,n1190);
and (n1187,n1188,n1189);
xor (n1188,n1144,n1145);
and (n1189,n722,n1155);
and (n1190,n1191,n1192);
xor (n1191,n1188,n1189);
and (n1192,n1193,n1194);
xor (n1193,n1150,n1151);
and (n1194,n728,n1155);
and (n1195,n687,n1196);
or (n1197,n1198,n1201);
and (n1198,n1199,n1200);
xor (n1199,n1161,n1162);
and (n1200,n694,n1196);
and (n1201,n1202,n1203);
xor (n1202,n1199,n1200);
or (n1203,n1204,n1207);
and (n1204,n1205,n1206);
xor (n1205,n1167,n1168);
and (n1206,n701,n1196);
and (n1207,n1208,n1209);
xor (n1208,n1205,n1206);
or (n1209,n1210,n1213);
and (n1210,n1211,n1212);
xor (n1211,n1173,n1174);
and (n1212,n708,n1196);
and (n1213,n1214,n1215);
xor (n1214,n1211,n1212);
or (n1215,n1216,n1219);
and (n1216,n1217,n1218);
xor (n1217,n1179,n1180);
and (n1218,n715,n1196);
and (n1219,n1220,n1221);
xor (n1220,n1217,n1218);
or (n1221,n1222,n1225);
and (n1222,n1223,n1224);
xor (n1223,n1185,n1186);
and (n1224,n722,n1196);
and (n1225,n1226,n1227);
xor (n1226,n1223,n1224);
and (n1227,n1228,n1229);
xor (n1228,n1191,n1192);
and (n1229,n728,n1196);
and (n1230,n694,n1231);
or (n1232,n1233,n1236);
and (n1233,n1234,n1235);
xor (n1234,n1202,n1203);
and (n1235,n701,n1231);
and (n1236,n1237,n1238);
xor (n1237,n1234,n1235);
or (n1238,n1239,n1242);
and (n1239,n1240,n1241);
xor (n1240,n1208,n1209);
and (n1241,n708,n1231);
and (n1242,n1243,n1244);
xor (n1243,n1240,n1241);
or (n1244,n1245,n1248);
and (n1245,n1246,n1247);
xor (n1246,n1214,n1215);
and (n1247,n715,n1231);
and (n1248,n1249,n1250);
xor (n1249,n1246,n1247);
or (n1250,n1251,n1254);
and (n1251,n1252,n1253);
xor (n1252,n1220,n1221);
and (n1253,n722,n1231);
and (n1254,n1255,n1256);
xor (n1255,n1252,n1253);
and (n1256,n1257,n1258);
xor (n1257,n1226,n1227);
and (n1258,n728,n1231);
xor (n1260,n1261,n1862);
xor (n1261,n1262,n1860);
xor (n1262,n1263,n1827);
xor (n1263,n1264,n1825);
xor (n1264,n1265,n1786);
xor (n1265,n1266,n1784);
xor (n1266,n1267,n1739);
xor (n1267,n1268,n1737);
xor (n1268,n1269,n1686);
xor (n1269,n1270,n1684);
xor (n1270,n1271,n1627);
xor (n1271,n1272,n1625);
xor (n1272,n1273,n1562);
xor (n1273,n1274,n1560);
or (n1274,n1275,n1495);
and (n1275,n1276,n1493);
or (n1276,n1277,n1428);
and (n1277,n1278,n1426);
or (n1278,n1279,n1361);
and (n1279,n1280,n1359);
and (n1280,n1281,n1284);
and (n1281,n1282,n1283);
wire s0n1282,s1n1282,notn1282;
or (n1282,s0n1282,s1n1282);
not(notn1282,n1259);
and (s0n1282,notn1282,n23);
and (s1n1282,n1259,n652);
wire s0n1283,s1n1283,notn1283;
or (n1283,s0n1283,s1n1283);
not(notn1283,n1259);
and (s0n1283,notn1283,n24);
and (s1n1283,n1259,n653);
or (n1284,n1285,n1290);
and (n1285,n1286,n1288);
and (n1286,n1282,n1287);
wire s0n1287,s1n1287,notn1287;
or (n1287,s0n1287,s1n1287);
not(notn1287,n1259);
and (s0n1287,notn1287,n28);
and (s1n1287,n1259,n657);
and (n1288,n1289,n1283);
wire s0n1289,s1n1289,notn1289;
or (n1289,s0n1289,s1n1289);
not(notn1289,n1259);
and (s0n1289,notn1289,n30);
and (s1n1289,n1259,n659);
and (n1290,n1291,n1292);
xor (n1291,n1286,n1288);
or (n1292,n1293,n1297);
and (n1293,n1294,n1295);
and (n1294,n1289,n1287);
and (n1295,n1296,n1283);
wire s0n1296,s1n1296,notn1296;
or (n1296,s0n1296,s1n1296);
not(notn1296,n1259);
and (s0n1296,notn1296,n37);
and (s1n1296,n1259,n666);
and (n1297,n1298,n1299);
xor (n1298,n1294,n1295);
or (n1299,n1300,n1304);
and (n1300,n1301,n1302);
and (n1301,n1296,n1287);
and (n1302,n1303,n1283);
wire s0n1303,s1n1303,notn1303;
or (n1303,s0n1303,s1n1303);
not(notn1303,n1259);
and (s0n1303,notn1303,n44);
and (s1n1303,n1259,n673);
and (n1304,n1305,n1306);
xor (n1305,n1301,n1302);
or (n1306,n1307,n1311);
and (n1307,n1308,n1309);
and (n1308,n1303,n1287);
and (n1309,n1310,n1283);
wire s0n1310,s1n1310,notn1310;
or (n1310,s0n1310,s1n1310);
not(notn1310,n1259);
and (s0n1310,notn1310,n51);
and (s1n1310,n1259,n680);
and (n1311,n1312,n1313);
xor (n1312,n1308,n1309);
or (n1313,n1314,n1318);
and (n1314,n1315,n1316);
and (n1315,n1310,n1287);
and (n1316,n1317,n1283);
wire s0n1317,s1n1317,notn1317;
or (n1317,s0n1317,s1n1317);
not(notn1317,n1259);
and (s0n1317,notn1317,n58);
and (s1n1317,n1259,n687);
and (n1318,n1319,n1320);
xor (n1319,n1315,n1316);
or (n1320,n1321,n1325);
and (n1321,n1322,n1323);
and (n1322,n1317,n1287);
and (n1323,n1324,n1283);
wire s0n1324,s1n1324,notn1324;
or (n1324,s0n1324,s1n1324);
not(notn1324,n1259);
and (s0n1324,notn1324,n65);
and (s1n1324,n1259,n694);
and (n1325,n1326,n1327);
xor (n1326,n1322,n1323);
or (n1327,n1328,n1332);
and (n1328,n1329,n1330);
and (n1329,n1324,n1287);
and (n1330,n1331,n1283);
wire s0n1331,s1n1331,notn1331;
or (n1331,s0n1331,s1n1331);
not(notn1331,n1259);
and (s0n1331,notn1331,n72);
and (s1n1331,n1259,n701);
and (n1332,n1333,n1334);
xor (n1333,n1329,n1330);
or (n1334,n1335,n1339);
and (n1335,n1336,n1337);
and (n1336,n1331,n1287);
and (n1337,n1338,n1283);
wire s0n1338,s1n1338,notn1338;
or (n1338,s0n1338,s1n1338);
not(notn1338,n1259);
and (s0n1338,notn1338,n79);
and (s1n1338,n1259,n708);
and (n1339,n1340,n1341);
xor (n1340,n1336,n1337);
or (n1341,n1342,n1346);
and (n1342,n1343,n1344);
and (n1343,n1338,n1287);
and (n1344,n1345,n1283);
wire s0n1345,s1n1345,notn1345;
or (n1345,s0n1345,s1n1345);
not(notn1345,n1259);
and (s0n1345,notn1345,n86);
and (s1n1345,n1259,n715);
and (n1346,n1347,n1348);
xor (n1347,n1343,n1344);
or (n1348,n1349,n1353);
and (n1349,n1350,n1351);
and (n1350,n1345,n1287);
and (n1351,n1352,n1283);
wire s0n1352,s1n1352,notn1352;
or (n1352,s0n1352,s1n1352);
not(notn1352,n1259);
and (s0n1352,notn1352,n93);
and (s1n1352,n1259,n722);
and (n1353,n1354,n1355);
xor (n1354,n1350,n1351);
and (n1355,n1356,n1357);
and (n1356,n1352,n1287);
and (n1357,n1358,n1283);
wire s0n1358,s1n1358,notn1358;
or (n1358,s0n1358,s1n1358);
not(notn1358,n1259);
and (s0n1358,notn1358,n99);
and (s1n1358,n1259,n728);
and (n1359,n1282,n1360);
wire s0n1360,s1n1360,notn1360;
or (n1360,s0n1360,s1n1360);
not(notn1360,n1259);
and (s0n1360,notn1360,n101);
and (s1n1360,n1259,n730);
and (n1361,n1362,n1363);
xor (n1362,n1280,n1359);
or (n1363,n1364,n1367);
and (n1364,n1365,n1366);
xor (n1365,n1281,n1284);
and (n1366,n1289,n1360);
and (n1367,n1368,n1369);
xor (n1368,n1365,n1366);
or (n1369,n1370,n1373);
and (n1370,n1371,n1372);
xor (n1371,n1291,n1292);
and (n1372,n1296,n1360);
and (n1373,n1374,n1375);
xor (n1374,n1371,n1372);
or (n1375,n1376,n1379);
and (n1376,n1377,n1378);
xor (n1377,n1298,n1299);
and (n1378,n1303,n1360);
and (n1379,n1380,n1381);
xor (n1380,n1377,n1378);
or (n1381,n1382,n1385);
and (n1382,n1383,n1384);
xor (n1383,n1305,n1306);
and (n1384,n1310,n1360);
and (n1385,n1386,n1387);
xor (n1386,n1383,n1384);
or (n1387,n1388,n1391);
and (n1388,n1389,n1390);
xor (n1389,n1312,n1313);
and (n1390,n1317,n1360);
and (n1391,n1392,n1393);
xor (n1392,n1389,n1390);
or (n1393,n1394,n1397);
and (n1394,n1395,n1396);
xor (n1395,n1319,n1320);
and (n1396,n1324,n1360);
and (n1397,n1398,n1399);
xor (n1398,n1395,n1396);
or (n1399,n1400,n1403);
and (n1400,n1401,n1402);
xor (n1401,n1326,n1327);
and (n1402,n1331,n1360);
and (n1403,n1404,n1405);
xor (n1404,n1401,n1402);
or (n1405,n1406,n1409);
and (n1406,n1407,n1408);
xor (n1407,n1333,n1334);
and (n1408,n1338,n1360);
and (n1409,n1410,n1411);
xor (n1410,n1407,n1408);
or (n1411,n1412,n1415);
and (n1412,n1413,n1414);
xor (n1413,n1340,n1341);
and (n1414,n1345,n1360);
and (n1415,n1416,n1417);
xor (n1416,n1413,n1414);
or (n1417,n1418,n1421);
and (n1418,n1419,n1420);
xor (n1419,n1347,n1348);
and (n1420,n1352,n1360);
and (n1421,n1422,n1423);
xor (n1422,n1419,n1420);
and (n1423,n1424,n1425);
xor (n1424,n1354,n1355);
and (n1425,n1358,n1360);
and (n1426,n1282,n1427);
wire s0n1427,s1n1427,notn1427;
or (n1427,s0n1427,s1n1427);
not(notn1427,n1259);
and (s0n1427,notn1427,n168);
and (s1n1427,n1259,n797);
and (n1428,n1429,n1430);
xor (n1429,n1278,n1426);
or (n1430,n1431,n1434);
and (n1431,n1432,n1433);
xor (n1432,n1362,n1363);
and (n1433,n1289,n1427);
and (n1434,n1435,n1436);
xor (n1435,n1432,n1433);
or (n1436,n1437,n1440);
and (n1437,n1438,n1439);
xor (n1438,n1368,n1369);
and (n1439,n1296,n1427);
and (n1440,n1441,n1442);
xor (n1441,n1438,n1439);
or (n1442,n1443,n1446);
and (n1443,n1444,n1445);
xor (n1444,n1374,n1375);
and (n1445,n1303,n1427);
and (n1446,n1447,n1448);
xor (n1447,n1444,n1445);
or (n1448,n1449,n1452);
and (n1449,n1450,n1451);
xor (n1450,n1380,n1381);
and (n1451,n1310,n1427);
and (n1452,n1453,n1454);
xor (n1453,n1450,n1451);
or (n1454,n1455,n1458);
and (n1455,n1456,n1457);
xor (n1456,n1386,n1387);
and (n1457,n1317,n1427);
and (n1458,n1459,n1460);
xor (n1459,n1456,n1457);
or (n1460,n1461,n1464);
and (n1461,n1462,n1463);
xor (n1462,n1392,n1393);
and (n1463,n1324,n1427);
and (n1464,n1465,n1466);
xor (n1465,n1462,n1463);
or (n1466,n1467,n1470);
and (n1467,n1468,n1469);
xor (n1468,n1398,n1399);
and (n1469,n1331,n1427);
and (n1470,n1471,n1472);
xor (n1471,n1468,n1469);
or (n1472,n1473,n1476);
and (n1473,n1474,n1475);
xor (n1474,n1404,n1405);
and (n1475,n1338,n1427);
and (n1476,n1477,n1478);
xor (n1477,n1474,n1475);
or (n1478,n1479,n1482);
and (n1479,n1480,n1481);
xor (n1480,n1410,n1411);
and (n1481,n1345,n1427);
and (n1482,n1483,n1484);
xor (n1483,n1480,n1481);
or (n1484,n1485,n1488);
and (n1485,n1486,n1487);
xor (n1486,n1416,n1417);
and (n1487,n1352,n1427);
and (n1488,n1489,n1490);
xor (n1489,n1486,n1487);
and (n1490,n1491,n1492);
xor (n1491,n1422,n1423);
and (n1492,n1358,n1427);
and (n1493,n1282,n1494);
wire s0n1494,s1n1494,notn1494;
or (n1494,s0n1494,s1n1494);
not(notn1494,n1259);
and (s0n1494,notn1494,n235);
and (s1n1494,n1259,n864);
and (n1495,n1496,n1497);
xor (n1496,n1276,n1493);
or (n1497,n1498,n1501);
and (n1498,n1499,n1500);
xor (n1499,n1429,n1430);
and (n1500,n1289,n1494);
and (n1501,n1502,n1503);
xor (n1502,n1499,n1500);
or (n1503,n1504,n1507);
and (n1504,n1505,n1506);
xor (n1505,n1435,n1436);
and (n1506,n1296,n1494);
and (n1507,n1508,n1509);
xor (n1508,n1505,n1506);
or (n1509,n1510,n1513);
and (n1510,n1511,n1512);
xor (n1511,n1441,n1442);
and (n1512,n1303,n1494);
and (n1513,n1514,n1515);
xor (n1514,n1511,n1512);
or (n1515,n1516,n1519);
and (n1516,n1517,n1518);
xor (n1517,n1447,n1448);
and (n1518,n1310,n1494);
and (n1519,n1520,n1521);
xor (n1520,n1517,n1518);
or (n1521,n1522,n1525);
and (n1522,n1523,n1524);
xor (n1523,n1453,n1454);
and (n1524,n1317,n1494);
and (n1525,n1526,n1527);
xor (n1526,n1523,n1524);
or (n1527,n1528,n1531);
and (n1528,n1529,n1530);
xor (n1529,n1459,n1460);
and (n1530,n1324,n1494);
and (n1531,n1532,n1533);
xor (n1532,n1529,n1530);
or (n1533,n1534,n1537);
and (n1534,n1535,n1536);
xor (n1535,n1465,n1466);
and (n1536,n1331,n1494);
and (n1537,n1538,n1539);
xor (n1538,n1535,n1536);
or (n1539,n1540,n1543);
and (n1540,n1541,n1542);
xor (n1541,n1471,n1472);
and (n1542,n1338,n1494);
and (n1543,n1544,n1545);
xor (n1544,n1541,n1542);
or (n1545,n1546,n1549);
and (n1546,n1547,n1548);
xor (n1547,n1477,n1478);
and (n1548,n1345,n1494);
and (n1549,n1550,n1551);
xor (n1550,n1547,n1548);
or (n1551,n1552,n1555);
and (n1552,n1553,n1554);
xor (n1553,n1483,n1484);
and (n1554,n1352,n1494);
and (n1555,n1556,n1557);
xor (n1556,n1553,n1554);
and (n1557,n1558,n1559);
xor (n1558,n1489,n1490);
and (n1559,n1358,n1494);
and (n1560,n1282,n1561);
wire s0n1561,s1n1561,notn1561;
or (n1561,s0n1561,s1n1561);
not(notn1561,n1259);
and (s0n1561,notn1561,n302);
and (s1n1561,n1259,n931);
or (n1562,n1563,n1566);
and (n1563,n1564,n1565);
xor (n1564,n1496,n1497);
and (n1565,n1289,n1561);
and (n1566,n1567,n1568);
xor (n1567,n1564,n1565);
or (n1568,n1569,n1572);
and (n1569,n1570,n1571);
xor (n1570,n1502,n1503);
and (n1571,n1296,n1561);
and (n1572,n1573,n1574);
xor (n1573,n1570,n1571);
or (n1574,n1575,n1578);
and (n1575,n1576,n1577);
xor (n1576,n1508,n1509);
and (n1577,n1303,n1561);
and (n1578,n1579,n1580);
xor (n1579,n1576,n1577);
or (n1580,n1581,n1584);
and (n1581,n1582,n1583);
xor (n1582,n1514,n1515);
and (n1583,n1310,n1561);
and (n1584,n1585,n1586);
xor (n1585,n1582,n1583);
or (n1586,n1587,n1590);
and (n1587,n1588,n1589);
xor (n1588,n1520,n1521);
and (n1589,n1317,n1561);
and (n1590,n1591,n1592);
xor (n1591,n1588,n1589);
or (n1592,n1593,n1596);
and (n1593,n1594,n1595);
xor (n1594,n1526,n1527);
and (n1595,n1324,n1561);
and (n1596,n1597,n1598);
xor (n1597,n1594,n1595);
or (n1598,n1599,n1602);
and (n1599,n1600,n1601);
xor (n1600,n1532,n1533);
and (n1601,n1331,n1561);
and (n1602,n1603,n1604);
xor (n1603,n1600,n1601);
or (n1604,n1605,n1608);
and (n1605,n1606,n1607);
xor (n1606,n1538,n1539);
and (n1607,n1338,n1561);
and (n1608,n1609,n1610);
xor (n1609,n1606,n1607);
or (n1610,n1611,n1614);
and (n1611,n1612,n1613);
xor (n1612,n1544,n1545);
and (n1613,n1345,n1561);
and (n1614,n1615,n1616);
xor (n1615,n1612,n1613);
or (n1616,n1617,n1620);
and (n1617,n1618,n1619);
xor (n1618,n1550,n1551);
and (n1619,n1352,n1561);
and (n1620,n1621,n1622);
xor (n1621,n1618,n1619);
and (n1622,n1623,n1624);
xor (n1623,n1556,n1557);
and (n1624,n1358,n1561);
and (n1625,n1289,n1626);
wire s0n1626,s1n1626,notn1626;
or (n1626,s0n1626,s1n1626);
not(notn1626,n1259);
and (s0n1626,notn1626,n367);
and (s1n1626,n1259,n996);
or (n1627,n1628,n1631);
and (n1628,n1629,n1630);
xor (n1629,n1567,n1568);
and (n1630,n1296,n1626);
and (n1631,n1632,n1633);
xor (n1632,n1629,n1630);
or (n1633,n1634,n1637);
and (n1634,n1635,n1636);
xor (n1635,n1573,n1574);
and (n1636,n1303,n1626);
and (n1637,n1638,n1639);
xor (n1638,n1635,n1636);
or (n1639,n1640,n1643);
and (n1640,n1641,n1642);
xor (n1641,n1579,n1580);
and (n1642,n1310,n1626);
and (n1643,n1644,n1645);
xor (n1644,n1641,n1642);
or (n1645,n1646,n1649);
and (n1646,n1647,n1648);
xor (n1647,n1585,n1586);
and (n1648,n1317,n1626);
and (n1649,n1650,n1651);
xor (n1650,n1647,n1648);
or (n1651,n1652,n1655);
and (n1652,n1653,n1654);
xor (n1653,n1591,n1592);
and (n1654,n1324,n1626);
and (n1655,n1656,n1657);
xor (n1656,n1653,n1654);
or (n1657,n1658,n1661);
and (n1658,n1659,n1660);
xor (n1659,n1597,n1598);
and (n1660,n1331,n1626);
and (n1661,n1662,n1663);
xor (n1662,n1659,n1660);
or (n1663,n1664,n1667);
and (n1664,n1665,n1666);
xor (n1665,n1603,n1604);
and (n1666,n1338,n1626);
and (n1667,n1668,n1669);
xor (n1668,n1665,n1666);
or (n1669,n1670,n1673);
and (n1670,n1671,n1672);
xor (n1671,n1609,n1610);
and (n1672,n1345,n1626);
and (n1673,n1674,n1675);
xor (n1674,n1671,n1672);
or (n1675,n1676,n1679);
and (n1676,n1677,n1678);
xor (n1677,n1615,n1616);
and (n1678,n1352,n1626);
and (n1679,n1680,n1681);
xor (n1680,n1677,n1678);
and (n1681,n1682,n1683);
xor (n1682,n1621,n1622);
and (n1683,n1358,n1626);
and (n1684,n1296,n1685);
wire s0n1685,s1n1685,notn1685;
or (n1685,s0n1685,s1n1685);
not(notn1685,n1259);
and (s0n1685,notn1685,n426);
and (s1n1685,n1259,n1055);
or (n1686,n1687,n1690);
and (n1687,n1688,n1689);
xor (n1688,n1632,n1633);
and (n1689,n1303,n1685);
and (n1690,n1691,n1692);
xor (n1691,n1688,n1689);
or (n1692,n1693,n1696);
and (n1693,n1694,n1695);
xor (n1694,n1638,n1639);
and (n1695,n1310,n1685);
and (n1696,n1697,n1698);
xor (n1697,n1694,n1695);
or (n1698,n1699,n1702);
and (n1699,n1700,n1701);
xor (n1700,n1644,n1645);
and (n1701,n1317,n1685);
and (n1702,n1703,n1704);
xor (n1703,n1700,n1701);
or (n1704,n1705,n1708);
and (n1705,n1706,n1707);
xor (n1706,n1650,n1651);
and (n1707,n1324,n1685);
and (n1708,n1709,n1710);
xor (n1709,n1706,n1707);
or (n1710,n1711,n1714);
and (n1711,n1712,n1713);
xor (n1712,n1656,n1657);
and (n1713,n1331,n1685);
and (n1714,n1715,n1716);
xor (n1715,n1712,n1713);
or (n1716,n1717,n1720);
and (n1717,n1718,n1719);
xor (n1718,n1662,n1663);
and (n1719,n1338,n1685);
and (n1720,n1721,n1722);
xor (n1721,n1718,n1719);
or (n1722,n1723,n1726);
and (n1723,n1724,n1725);
xor (n1724,n1668,n1669);
and (n1725,n1345,n1685);
and (n1726,n1727,n1728);
xor (n1727,n1724,n1725);
or (n1728,n1729,n1732);
and (n1729,n1730,n1731);
xor (n1730,n1674,n1675);
and (n1731,n1352,n1685);
and (n1732,n1733,n1734);
xor (n1733,n1730,n1731);
and (n1734,n1735,n1736);
xor (n1735,n1680,n1681);
and (n1736,n1358,n1685);
and (n1737,n1303,n1738);
wire s0n1738,s1n1738,notn1738;
or (n1738,s0n1738,s1n1738);
not(notn1738,n1259);
and (s0n1738,notn1738,n479);
and (s1n1738,n1259,n1108);
or (n1739,n1740,n1743);
and (n1740,n1741,n1742);
xor (n1741,n1691,n1692);
and (n1742,n1310,n1738);
and (n1743,n1744,n1745);
xor (n1744,n1741,n1742);
or (n1745,n1746,n1749);
and (n1746,n1747,n1748);
xor (n1747,n1697,n1698);
and (n1748,n1317,n1738);
and (n1749,n1750,n1751);
xor (n1750,n1747,n1748);
or (n1751,n1752,n1755);
and (n1752,n1753,n1754);
xor (n1753,n1703,n1704);
and (n1754,n1324,n1738);
and (n1755,n1756,n1757);
xor (n1756,n1753,n1754);
or (n1757,n1758,n1761);
and (n1758,n1759,n1760);
xor (n1759,n1709,n1710);
and (n1760,n1331,n1738);
and (n1761,n1762,n1763);
xor (n1762,n1759,n1760);
or (n1763,n1764,n1767);
and (n1764,n1765,n1766);
xor (n1765,n1715,n1716);
and (n1766,n1338,n1738);
and (n1767,n1768,n1769);
xor (n1768,n1765,n1766);
or (n1769,n1770,n1773);
and (n1770,n1771,n1772);
xor (n1771,n1721,n1722);
and (n1772,n1345,n1738);
and (n1773,n1774,n1775);
xor (n1774,n1771,n1772);
or (n1775,n1776,n1779);
and (n1776,n1777,n1778);
xor (n1777,n1727,n1728);
and (n1778,n1352,n1738);
and (n1779,n1780,n1781);
xor (n1780,n1777,n1778);
and (n1781,n1782,n1783);
xor (n1782,n1733,n1734);
and (n1783,n1358,n1738);
and (n1784,n1310,n1785);
wire s0n1785,s1n1785,notn1785;
or (n1785,s0n1785,s1n1785);
not(notn1785,n1259);
and (s0n1785,notn1785,n526);
and (s1n1785,n1259,n1155);
or (n1786,n1787,n1790);
and (n1787,n1788,n1789);
xor (n1788,n1744,n1745);
and (n1789,n1317,n1785);
and (n1790,n1791,n1792);
xor (n1791,n1788,n1789);
or (n1792,n1793,n1796);
and (n1793,n1794,n1795);
xor (n1794,n1750,n1751);
and (n1795,n1324,n1785);
and (n1796,n1797,n1798);
xor (n1797,n1794,n1795);
or (n1798,n1799,n1802);
and (n1799,n1800,n1801);
xor (n1800,n1756,n1757);
and (n1801,n1331,n1785);
and (n1802,n1803,n1804);
xor (n1803,n1800,n1801);
or (n1804,n1805,n1808);
and (n1805,n1806,n1807);
xor (n1806,n1762,n1763);
and (n1807,n1338,n1785);
and (n1808,n1809,n1810);
xor (n1809,n1806,n1807);
or (n1810,n1811,n1814);
and (n1811,n1812,n1813);
xor (n1812,n1768,n1769);
and (n1813,n1345,n1785);
and (n1814,n1815,n1816);
xor (n1815,n1812,n1813);
or (n1816,n1817,n1820);
and (n1817,n1818,n1819);
xor (n1818,n1774,n1775);
and (n1819,n1352,n1785);
and (n1820,n1821,n1822);
xor (n1821,n1818,n1819);
and (n1822,n1823,n1824);
xor (n1823,n1780,n1781);
and (n1824,n1358,n1785);
and (n1825,n1317,n1826);
wire s0n1826,s1n1826,notn1826;
or (n1826,s0n1826,s1n1826);
not(notn1826,n1259);
and (s0n1826,notn1826,n567);
and (s1n1826,n1259,n1196);
or (n1827,n1828,n1831);
and (n1828,n1829,n1830);
xor (n1829,n1791,n1792);
and (n1830,n1324,n1826);
and (n1831,n1832,n1833);
xor (n1832,n1829,n1830);
or (n1833,n1834,n1837);
and (n1834,n1835,n1836);
xor (n1835,n1797,n1798);
and (n1836,n1331,n1826);
and (n1837,n1838,n1839);
xor (n1838,n1835,n1836);
or (n1839,n1840,n1843);
and (n1840,n1841,n1842);
xor (n1841,n1803,n1804);
and (n1842,n1338,n1826);
and (n1843,n1844,n1845);
xor (n1844,n1841,n1842);
or (n1845,n1846,n1849);
and (n1846,n1847,n1848);
xor (n1847,n1809,n1810);
and (n1848,n1345,n1826);
and (n1849,n1850,n1851);
xor (n1850,n1847,n1848);
or (n1851,n1852,n1855);
and (n1852,n1853,n1854);
xor (n1853,n1815,n1816);
and (n1854,n1352,n1826);
and (n1855,n1856,n1857);
xor (n1856,n1853,n1854);
and (n1857,n1858,n1859);
xor (n1858,n1821,n1822);
and (n1859,n1358,n1826);
and (n1860,n1324,n1861);
wire s0n1861,s1n1861,notn1861;
or (n1861,s0n1861,s1n1861);
not(notn1861,n1259);
and (s0n1861,notn1861,n602);
and (s1n1861,n1259,n1231);
or (n1862,n1863,n1866);
and (n1863,n1864,n1865);
xor (n1864,n1832,n1833);
and (n1865,n1331,n1861);
and (n1866,n1867,n1868);
xor (n1867,n1864,n1865);
or (n1868,n1869,n1872);
and (n1869,n1870,n1871);
xor (n1870,n1838,n1839);
and (n1871,n1338,n1861);
and (n1872,n1873,n1874);
xor (n1873,n1870,n1871);
or (n1874,n1875,n1878);
and (n1875,n1876,n1877);
xor (n1876,n1844,n1845);
and (n1877,n1345,n1861);
and (n1878,n1879,n1880);
xor (n1879,n1876,n1877);
or (n1880,n1881,n1884);
and (n1881,n1882,n1883);
xor (n1882,n1850,n1851);
and (n1883,n1352,n1861);
and (n1884,n1885,n1886);
xor (n1885,n1882,n1883);
and (n1886,n1887,n1888);
xor (n1887,n1856,n1857);
and (n1888,n1358,n1861);
endmodule
