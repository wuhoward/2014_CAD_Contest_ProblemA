module top (out,n13,n23,n25,n26,n28,n33,n36,n38,n43
        ,n47,n55,n59,n60,n61,n73,n77,n78,n79,n94
        ,n95,n96,n97,n98,n102,n103,n104,n109,n111,n113
        ,n150,n152,n153,n154,n165,n166,n167,n168,n180,n181
        ,n182,n183,n197,n203,n205,n206,n210,n211,n214,n216
        ,n217,n218,n291,n346,n349,n351,n439,n441,n442,n557
        ,n558,n559,n560,n567,n569,n573,n584,n587,n589,n590
        ,n592,n596,n602,n605,n607,n609,n613,n616,n618,n620
        ,n624,n627,n629,n631,n633,n639,n642,n644,n646,n650
        ,n653,n655,n657,n661,n664,n666,n668,n672,n675,n677
        ,n679,n686,n689,n691,n693,n697,n700,n702,n704,n708
        ,n711,n713,n715,n719,n722,n724,n726,n735,n739,n741
        ,n743,n765,n769,n771,n773,n783,n787,n789,n791,n801
        ,n805,n807,n809,n819,n823,n825,n827,n837,n841,n843
        ,n845,n856,n858,n860,n862,n935,n938,n940,n942,n946
        ,n949,n951,n953,n957,n960,n962,n964,n968,n971,n973
        ,n975,n982,n985,n987,n989,n993,n996,n998,n1000,n1004
        ,n1007,n1009,n1011,n1015,n1018,n1020,n1022,n1029,n1032,n1034
        ,n1036,n1040,n1043,n1045,n1047,n1051,n1054,n1056,n1058,n1062
        ,n1065,n1067,n1069,n1299,n1303,n1305,n1307,n1317,n1321,n1323
        ,n1325,n1337,n1339,n1341,n1343,n1355,n1357,n1359,n1361,n1371
        ,n1375,n1377,n1379,n1391,n1393,n1395,n1397,n1407,n1411,n1413
        ,n1415,n1424,n1428,n1430,n1432,n1762,n1766,n1768,n1770,n1779
        ,n1783,n1785,n1787,n1803,n1807,n1809,n1811,n1821,n1825,n1827
        ,n1829,n1839,n1843,n1845,n1847,n1859,n1861,n1863,n1865,n1877
        ,n1879,n1881,n1883,n1892,n1896,n1898,n1900,n2120,n2122,n2124
        ,n2126,n2138,n2140,n2142,n2144,n2156,n2158,n2160,n2162,n2174
        ,n2176,n2178,n2180,n2192,n2194,n2196,n2198,n2208,n2212,n2214
        ,n2216,n2228,n2230,n2232,n2234,n2245,n2247,n2249,n2251);
output out;
input n13;
input n23;
input n25;
input n26;
input n28;
input n33;
input n36;
input n38;
input n43;
input n47;
input n55;
input n59;
input n60;
input n61;
input n73;
input n77;
input n78;
input n79;
input n94;
input n95;
input n96;
input n97;
input n98;
input n102;
input n103;
input n104;
input n109;
input n111;
input n113;
input n150;
input n152;
input n153;
input n154;
input n165;
input n166;
input n167;
input n168;
input n180;
input n181;
input n182;
input n183;
input n197;
input n203;
input n205;
input n206;
input n210;
input n211;
input n214;
input n216;
input n217;
input n218;
input n291;
input n346;
input n349;
input n351;
input n439;
input n441;
input n442;
input n557;
input n558;
input n559;
input n560;
input n567;
input n569;
input n573;
input n584;
input n587;
input n589;
input n590;
input n592;
input n596;
input n602;
input n605;
input n607;
input n609;
input n613;
input n616;
input n618;
input n620;
input n624;
input n627;
input n629;
input n631;
input n633;
input n639;
input n642;
input n644;
input n646;
input n650;
input n653;
input n655;
input n657;
input n661;
input n664;
input n666;
input n668;
input n672;
input n675;
input n677;
input n679;
input n686;
input n689;
input n691;
input n693;
input n697;
input n700;
input n702;
input n704;
input n708;
input n711;
input n713;
input n715;
input n719;
input n722;
input n724;
input n726;
input n735;
input n739;
input n741;
input n743;
input n765;
input n769;
input n771;
input n773;
input n783;
input n787;
input n789;
input n791;
input n801;
input n805;
input n807;
input n809;
input n819;
input n823;
input n825;
input n827;
input n837;
input n841;
input n843;
input n845;
input n856;
input n858;
input n860;
input n862;
input n935;
input n938;
input n940;
input n942;
input n946;
input n949;
input n951;
input n953;
input n957;
input n960;
input n962;
input n964;
input n968;
input n971;
input n973;
input n975;
input n982;
input n985;
input n987;
input n989;
input n993;
input n996;
input n998;
input n1000;
input n1004;
input n1007;
input n1009;
input n1011;
input n1015;
input n1018;
input n1020;
input n1022;
input n1029;
input n1032;
input n1034;
input n1036;
input n1040;
input n1043;
input n1045;
input n1047;
input n1051;
input n1054;
input n1056;
input n1058;
input n1062;
input n1065;
input n1067;
input n1069;
input n1299;
input n1303;
input n1305;
input n1307;
input n1317;
input n1321;
input n1323;
input n1325;
input n1337;
input n1339;
input n1341;
input n1343;
input n1355;
input n1357;
input n1359;
input n1361;
input n1371;
input n1375;
input n1377;
input n1379;
input n1391;
input n1393;
input n1395;
input n1397;
input n1407;
input n1411;
input n1413;
input n1415;
input n1424;
input n1428;
input n1430;
input n1432;
input n1762;
input n1766;
input n1768;
input n1770;
input n1779;
input n1783;
input n1785;
input n1787;
input n1803;
input n1807;
input n1809;
input n1811;
input n1821;
input n1825;
input n1827;
input n1829;
input n1839;
input n1843;
input n1845;
input n1847;
input n1859;
input n1861;
input n1863;
input n1865;
input n1877;
input n1879;
input n1881;
input n1883;
input n1892;
input n1896;
input n1898;
input n1900;
input n2120;
input n2122;
input n2124;
input n2126;
input n2138;
input n2140;
input n2142;
input n2144;
input n2156;
input n2158;
input n2160;
input n2162;
input n2174;
input n2176;
input n2178;
input n2180;
input n2192;
input n2194;
input n2196;
input n2198;
input n2208;
input n2212;
input n2214;
input n2216;
input n2228;
input n2230;
input n2232;
input n2234;
input n2245;
input n2247;
input n2249;
input n2251;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n24;
wire n27;
wire n29;
wire n30;
wire n31;
wire n32;
wire n34;
wire n35;
wire n37;
wire n39;
wire n40;
wire n41;
wire n42;
wire n44;
wire n45;
wire n46;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n56;
wire n57;
wire n58;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n74;
wire n75;
wire n76;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n99;
wire n100;
wire n101;
wire n105;
wire n106;
wire n107;
wire n108;
wire n110;
wire n112;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n151;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n204;
wire n207;
wire n208;
wire n209;
wire n212;
wire n213;
wire n215;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n347;
wire n348;
wire n350;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n440;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n568;
wire n570;
wire n571;
wire n572;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n585;
wire n586;
wire n588;
wire n591;
wire n593;
wire n594;
wire n595;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n603;
wire n604;
wire n606;
wire n608;
wire n610;
wire n611;
wire n612;
wire n614;
wire n615;
wire n617;
wire n619;
wire n621;
wire n622;
wire n623;
wire n625;
wire n626;
wire n628;
wire n630;
wire n632;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n640;
wire n641;
wire n643;
wire n645;
wire n647;
wire n648;
wire n649;
wire n651;
wire n652;
wire n654;
wire n656;
wire n658;
wire n659;
wire n660;
wire n662;
wire n663;
wire n665;
wire n667;
wire n669;
wire n670;
wire n671;
wire n673;
wire n674;
wire n676;
wire n678;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n687;
wire n688;
wire n690;
wire n692;
wire n694;
wire n695;
wire n696;
wire n698;
wire n699;
wire n701;
wire n703;
wire n705;
wire n706;
wire n707;
wire n709;
wire n710;
wire n712;
wire n714;
wire n716;
wire n717;
wire n718;
wire n720;
wire n721;
wire n723;
wire n725;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n736;
wire n737;
wire n738;
wire n740;
wire n742;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n766;
wire n767;
wire n768;
wire n770;
wire n772;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n784;
wire n785;
wire n786;
wire n788;
wire n790;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n802;
wire n803;
wire n804;
wire n806;
wire n808;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n820;
wire n821;
wire n822;
wire n824;
wire n826;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n838;
wire n839;
wire n840;
wire n842;
wire n844;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n857;
wire n859;
wire n861;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n936;
wire n937;
wire n939;
wire n941;
wire n943;
wire n944;
wire n945;
wire n947;
wire n948;
wire n950;
wire n952;
wire n954;
wire n955;
wire n956;
wire n958;
wire n959;
wire n961;
wire n963;
wire n965;
wire n966;
wire n967;
wire n969;
wire n970;
wire n972;
wire n974;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n983;
wire n984;
wire n986;
wire n988;
wire n990;
wire n991;
wire n992;
wire n994;
wire n995;
wire n997;
wire n999;
wire n1001;
wire n1002;
wire n1003;
wire n1005;
wire n1006;
wire n1008;
wire n1010;
wire n1012;
wire n1013;
wire n1014;
wire n1016;
wire n1017;
wire n1019;
wire n1021;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1030;
wire n1031;
wire n1033;
wire n1035;
wire n1037;
wire n1038;
wire n1039;
wire n1041;
wire n1042;
wire n1044;
wire n1046;
wire n1048;
wire n1049;
wire n1050;
wire n1052;
wire n1053;
wire n1055;
wire n1057;
wire n1059;
wire n1060;
wire n1061;
wire n1063;
wire n1064;
wire n1066;
wire n1068;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1300;
wire n1301;
wire n1302;
wire n1304;
wire n1306;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1318;
wire n1319;
wire n1320;
wire n1322;
wire n1324;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1338;
wire n1340;
wire n1342;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1356;
wire n1358;
wire n1360;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1372;
wire n1373;
wire n1374;
wire n1376;
wire n1378;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1392;
wire n1394;
wire n1396;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1408;
wire n1409;
wire n1410;
wire n1412;
wire n1414;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1425;
wire n1426;
wire n1427;
wire n1429;
wire n1431;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1763;
wire n1764;
wire n1765;
wire n1767;
wire n1769;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1780;
wire n1781;
wire n1782;
wire n1784;
wire n1786;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1804;
wire n1805;
wire n1806;
wire n1808;
wire n1810;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1822;
wire n1823;
wire n1824;
wire n1826;
wire n1828;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1840;
wire n1841;
wire n1842;
wire n1844;
wire n1846;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1860;
wire n1862;
wire n1864;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1878;
wire n1880;
wire n1882;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1893;
wire n1894;
wire n1895;
wire n1897;
wire n1899;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2121;
wire n2123;
wire n2125;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2139;
wire n2141;
wire n2143;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2157;
wire n2159;
wire n2161;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2175;
wire n2177;
wire n2179;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2193;
wire n2195;
wire n2197;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2209;
wire n2210;
wire n2211;
wire n2213;
wire n2215;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2229;
wire n2231;
wire n2233;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2246;
wire n2248;
wire n2250;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2988;
wire n2989;
wire n2990;
wire n2991;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2996;
wire n2997;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3003;
wire n3004;
wire n3005;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3010;
wire n3011;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3038;
wire n3039;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
wire n3056;
wire n3057;
wire n3058;
wire n3059;
wire n3060;
wire n3061;
wire n3062;
wire n3063;
wire n3064;
wire n3065;
wire n3066;
wire n3067;
wire n3068;
wire n3069;
wire n3070;
wire n3071;
wire n3072;
wire n3073;
wire n3074;
wire n3075;
wire n3076;
wire n3077;
wire n3078;
wire n3079;
wire n3080;
wire n3081;
wire n3082;
wire n3083;
wire n3084;
wire n3085;
wire n3086;
wire n3087;
wire n3088;
wire n3089;
wire n3090;
wire n3091;
wire n3092;
wire n3093;
wire n3094;
wire n3095;
wire n3096;
wire n3097;
wire n3098;
wire n3099;
wire n3100;
wire n3101;
wire n3102;
wire n3103;
wire n3104;
wire n3105;
wire n3106;
wire n3107;
wire n3108;
wire n3109;
wire n3110;
wire n3111;
wire n3112;
wire n3113;
wire n3114;
wire n3115;
wire n3116;
wire n3117;
wire n3118;
wire n3119;
wire n3120;
wire n3121;
wire n3122;
wire n3123;
wire n3124;
wire n3125;
wire n3126;
wire n3127;
wire n3128;
wire n3129;
wire n3130;
wire n3131;
wire n3132;
wire n3133;
wire n3134;
wire n3135;
wire n3136;
wire n3137;
wire n3138;
wire n3139;
wire n3140;
wire n3141;
wire n3142;
wire n3143;
wire n3144;
wire n3145;
wire n3146;
wire n3147;
wire n3148;
wire n3149;
wire n3150;
wire n3151;
wire n3152;
wire n3153;
wire n3154;
wire n3155;
wire n3156;
wire n3157;
wire n3158;
wire n3159;
wire n3160;
wire n3161;
wire n3162;
wire n3163;
wire n3164;
wire n3165;
wire n3166;
wire n3167;
wire n3168;
wire n3169;
wire n3170;
wire n3171;
wire n3172;
wire n3173;
wire n3174;
wire n3175;
wire n3176;
wire n3177;
wire n3178;
wire n3179;
wire n3180;
wire n3181;
wire n3182;
wire n3183;
wire n3184;
wire n3185;
wire n3186;
wire n3187;
wire n3188;
wire n3189;
wire n3190;
wire n3191;
wire n3192;
wire n3193;
wire n3194;
wire n3195;
wire n3196;
wire n3197;
wire n3198;
wire n3199;
wire n3200;
wire n3201;
wire n3202;
wire n3203;
wire n3204;
wire n3205;
wire n3206;
wire n3207;
wire n3208;
wire n3209;
wire n3210;
wire n3211;
wire n3212;
wire n3213;
wire n3214;
wire n3215;
wire n3216;
wire n3217;
wire n3218;
wire n3219;
wire n3220;
wire n3221;
wire n3222;
wire n3223;
wire n3224;
wire n3225;
wire n3226;
wire n3227;
wire n3228;
wire n3229;
wire n3230;
wire n3231;
wire n3232;
wire n3233;
wire n3234;
wire n3235;
wire n3236;
wire n3237;
wire n3238;
wire n3239;
wire n3240;
wire n3241;
wire n3242;
wire n3243;
wire n3244;
wire n3245;
wire n3246;
wire n3247;
wire n3248;
wire n3249;
wire n3250;
wire n3251;
wire n3252;
wire n3253;
wire n3254;
wire n3255;
wire n3256;
wire n3257;
wire n3258;
wire n3259;
wire n3260;
wire n3261;
wire n3262;
wire n3263;
wire n3264;
wire n3265;
wire n3266;
wire n3267;
wire n3268;
wire n3269;
wire n3270;
wire n3271;
wire n3272;
wire n3273;
wire n3274;
wire n3275;
wire n3276;
wire n3277;
wire n3278;
wire n3279;
wire n3280;
wire n3281;
wire n3282;
wire n3283;
wire n3284;
wire n3285;
wire n3286;
wire n3287;
wire n3288;
wire n3289;
wire n3290;
wire n3291;
wire n3292;
wire n3293;
wire n3294;
wire n3295;
wire n3296;
wire n3297;
wire n3298;
wire n3299;
wire n3300;
wire n3301;
wire n3302;
wire n3303;
wire n3304;
wire n3305;
wire n3306;
wire n3307;
wire n3308;
wire n3309;
wire n3310;
wire n3311;
wire n3312;
wire n3313;
wire n3314;
wire n3315;
wire n3316;
wire n3317;
wire n3318;
wire n3319;
wire n3320;
wire n3321;
wire n3322;
wire n3323;
wire n3324;
wire n3325;
wire n3326;
wire n3327;
wire n3328;
wire n3329;
wire n3330;
wire n3331;
wire n3332;
wire n3333;
wire n3334;
wire n3335;
wire n3336;
wire n3337;
wire n3338;
wire n3339;
wire n3340;
wire n3341;
wire n3342;
wire n3343;
wire n3344;
wire n3345;
wire n3346;
wire n3347;
wire n3348;
wire n3349;
wire n3350;
wire n3351;
wire n3352;
wire n3353;
wire n3354;
wire n3355;
wire n3356;
wire n3357;
wire n3358;
wire n3359;
wire n3360;
wire n3361;
wire n3362;
wire n3363;
wire n3364;
wire n3365;
wire n3366;
wire n3367;
wire n3368;
wire n3369;
wire n3370;
wire n3371;
wire n3372;
wire n3373;
wire n3374;
wire n3375;
wire n3376;
wire n3377;
wire n3378;
wire n3379;
wire n3380;
wire n3381;
wire n3382;
wire n3383;
wire n3384;
wire n3385;
wire n3386;
wire n3387;
wire n3388;
wire n3389;
wire n3390;
wire n3391;
wire n3392;
wire n3393;
wire n3394;
wire n3395;
wire n3396;
wire n3397;
wire n3398;
wire n3399;
wire n3400;
wire n3401;
wire n3402;
wire n3403;
wire n3404;
wire n3405;
wire n3406;
wire n3407;
wire n3408;
wire n3409;
wire n3410;
wire n3411;
wire n3412;
wire n3413;
wire n3414;
wire n3415;
wire n3416;
wire n3417;
wire n3418;
wire n3419;
wire n3420;
wire n3421;
wire n3422;
wire n3423;
wire n3424;
wire n3425;
wire n3426;
wire n3427;
wire n3428;
wire n3429;
wire n3430;
wire n3431;
wire n3432;
wire n3433;
wire n3434;
wire n3435;
wire n3436;
wire n3437;
wire n3438;
wire n3439;
wire n3440;
wire n3441;
wire n3442;
wire n3443;
wire n3444;
wire n3445;
wire n3446;
wire n3447;
wire n3448;
wire n3449;
wire n3450;
wire n3451;
wire n3452;
wire n3453;
wire n3454;
wire n3455;
wire n3456;
wire n3457;
wire n3458;
wire n3459;
wire n3460;
wire n3461;
wire n3462;
wire n3463;
wire n3464;
wire n3465;
wire n3466;
wire n3467;
wire n3468;
wire n3469;
wire n3470;
wire n3471;
wire n3472;
wire n3473;
wire n3474;
wire n3475;
wire n3476;
wire n3477;
wire n3478;
wire n3479;
wire n3480;
wire n3481;
wire n3482;
wire n3483;
wire n3484;
wire n3485;
wire n3486;
wire n3487;
wire n3488;
wire n3489;
wire n3490;
wire n3491;
wire n3492;
wire n3493;
wire n3494;
wire n3495;
wire n3496;
wire n3497;
wire n3498;
wire n3499;
wire n3500;
wire n3501;
wire n3502;
wire n3503;
wire n3504;
wire n3505;
wire n3506;
wire n3507;
wire n3508;
wire n3509;
wire n3510;
wire n3511;
wire n3512;
wire n3513;
wire n3514;
wire n3515;
wire n3516;
wire n3517;
wire n3518;
wire n3519;
wire n3520;
wire n3521;
wire n3522;
wire n3523;
wire n3524;
wire n3525;
wire n3526;
wire n3527;
wire n3528;
wire n3529;
wire n3530;
wire n3531;
wire n3532;
wire n3533;
wire n3534;
wire n3535;
wire n3536;
wire n3537;
wire n3538;
wire n3539;
wire n3540;
wire n3541;
wire n3542;
wire n3543;
wire n3544;
wire n3545;
wire n3546;
wire n3547;
wire n3548;
wire n3549;
wire n3550;
wire n3551;
wire n3552;
xor (out,n0,n2670);
xor (n0,n1,n2647);
xor (n1,n2,n2548);
xor (n2,n3,n1752);
xor (n3,n4,n1657);
xor (n4,n5,n1291);
xor (n5,n6,n1071);
wire s0n6,s1n6,notn6;
or (n6,s0n6,s1n6);
not(notn6,n929);
and (s0n6,notn6,1'b0);
and (s1n6,n929,n8);
xor (n8,n9,n728);
wire s0n9,s1n9,notn9;
or (n9,s0n9,s1n9);
not(notn9,n578);
and (s0n9,notn9,1'b0);
and (s1n9,n578,n10);
nand (n10,n11,n563);
or (n11,n12,n14);
not (n12,n13);
not (n14,n15);
and (n15,n16,n561);
nor (n16,n17,n554);
not (n17,n18);
nor (n18,n19,n52);
nor (n19,n20,n39);
and (n20,n21,n38);
or (n21,n22,n27,n32,n35);
and (n22,n23,n24);
and (n24,n25,n26);
and (n27,n28,n29);
not (n29,n30);
nand (n30,n31,n26);
not (n31,n25);
and (n32,n33,n34);
nor (n34,n31,n26);
and (n35,n36,n37);
nor (n37,n25,n26);
nor (n39,n40,n48,n38);
and (n40,n41,n46);
nand (n41,n42,n44);
or (n42,n43,n36);
or (n44,n45,n28);
not (n45,n43);
not (n46,n47);
and (n48,n49,n47);
nand (n49,n50,n51);
or (n50,n43,n33);
or (n51,n45,n23);
nand (n52,n53,n62);
or (n53,n54,n56);
not (n54,n55);
not (n56,n57);
nand (n57,n58,n61);
nor (n58,n59,n60);
nand (n62,n63,n518);
nand (n63,n64,n510);
or (n64,n65,n434);
not (n65,n66);
or (n66,1'b0,n67,n354,n432);
and (n67,n68,n353);
wire s0n68,s1n68,notn68;
or (n68,s0n68,s1n68);
not(notn68,n344);
and (s0n68,notn68,n69);
and (s1n68,n344,1'b0);
wire s0n69,s1n69,notn69;
or (n69,s0n69,s1n69);
not(notn69,n280);
and (s0n69,notn69,1'b0);
and (s1n69,n280,n70);
or (n70,n71,n254,n260,n266,n271,1'b0,1'b0,1'b0);
and (n71,n72,n80);
xnor (n72,n73,n74);
not (n74,n75);
nor (n75,n76,n79);
or (n76,n77,n78);
and (n80,n81,n223,n242,n250);
wire s0n81,s1n81,notn81;
or (n81,s0n81,s1n81);
not(notn81,n114);
and (s0n81,notn81,n82);
and (s1n81,n114,1'b0);
wire s0n82,s1n82,notn82;
or (n82,s0n82,s1n82);
not(notn82,n112);
and (s0n82,notn82,n83);
and (s1n82,n112,n110);
wire s0n83,s1n83,notn83;
or (n83,s0n83,s1n83);
not(notn83,n105);
and (s0n83,notn83,n84);
and (s1n83,n105,n99);
wire s0n84,s1n84,notn84;
or (n84,s0n84,s1n84);
not(notn84,n98);
and (s0n84,notn84,n85);
and (s1n84,n98,1'b0);
wire s0n85,s1n85,notn85;
or (n85,s0n85,s1n85);
not(notn85,n97);
and (s0n85,notn85,n86);
and (s1n85,n97,1'b1);
wire s0n86,s1n86,notn86;
or (n86,s0n86,s1n86);
not(notn86,n96);
and (s0n86,notn86,n87);
and (s1n86,n96,1'b0);
wire s0n87,s1n87,notn87;
or (n87,s0n87,s1n87);
not(notn87,n95);
and (s0n87,notn87,n88);
and (s1n87,n95,1'b1);
wire s0n88,s1n88,notn88;
or (n88,s0n88,s1n88);
not(notn88,n94);
and (s0n88,notn88,n89);
and (s1n88,n94,1'b0);
wire s0n89,s1n89,notn89;
or (n89,s0n89,s1n89);
not(notn89,n73);
and (s0n89,notn89,n90);
and (s1n89,n73,1'b1);
wire s0n90,s1n90,notn90;
or (n90,s0n90,s1n90);
not(notn90,n79);
and (s0n90,notn90,n91);
and (s1n90,n79,1'b0);
wire s0n91,s1n91,notn91;
or (n91,s0n91,s1n91);
not(notn91,n77);
and (s0n91,notn91,n92);
and (s1n91,n77,1'b1);
not (n92,n78);
wire s0n99,s1n99,notn99;
or (n99,s0n99,s1n99);
not(notn99,n104);
and (s0n99,notn99,n100);
and (s1n99,n104,1'b0);
wire s0n100,s1n100,notn100;
or (n100,s0n100,s1n100);
not(notn100,n103);
and (s0n100,notn100,n101);
and (s1n100,n103,1'b1);
not (n101,n102);
or (n105,n106,n109);
or (n106,n104,n107);
not (n107,n108);
nor (n108,n103,n102);
not (n110,n111);
or (n112,n111,n113);
not (n114,n115);
or (n115,n116,n221);
or (n116,n117,n219);
or (n117,n118,n213);
or (n118,n119,n212);
or (n119,n120,n208);
or (n120,n121,n207);
or (n121,n122,n202);
or (n122,n123,n201);
or (n123,n124,n200);
or (n124,n125,n198);
or (n125,n126,n195);
or (n126,n127,n194);
or (n127,n128,n193);
or (n128,n129,n192);
or (n129,n130,n191);
or (n130,n131,n189);
or (n131,n132,n187);
or (n132,n133,n186);
or (n133,n134,n184);
or (n134,n135,n178);
or (n135,n136,n177);
or (n136,n137,n176);
or (n137,n138,n175);
or (n138,n139,n174);
or (n139,n140,n173);
or (n140,n141,n171);
or (n141,n142,n169);
or (n142,n143,n163);
or (n143,n144,n162);
or (n144,n145,n161);
or (n145,n146,n160);
or (n146,n147,n159);
or (n147,n148,n157);
or (n148,n149,n155);
nor (n149,n150,n151,n153,n154);
not (n151,n152);
nor (n155,n150,n151,n156,n154);
not (n156,n153);
and (n157,n150,n152,n153,n158);
not (n158,n154);
and (n159,n150,n151,n153,n158);
nor (n160,n150,n152,n156,n154);
and (n161,n150,n151,n153,n154);
and (n162,n150,n152,n153,n154);
nor (n163,n164,n166,n167,n168);
not (n164,n165);
nor (n169,n164,n170,n167,n168);
not (n170,n166);
and (n171,n164,n166,n167,n172);
not (n172,n168);
and (n173,n165,n166,n167,n172);
and (n174,n165,n170,n167,n172);
and (n175,n164,n170,n167,n168);
and (n176,n165,n170,n167,n168);
and (n177,n165,n166,n167,n168);
nor (n178,n179,n181,n182,n183);
not (n179,n180);
nor (n184,n179,n185,n182,n183);
not (n185,n181);
nor (n186,n180,n185,n182,n183);
nor (n187,n179,n185,n188,n183);
not (n188,n182);
nor (n189,n180,n181,n188,n190);
not (n190,n183);
and (n191,n179,n181,n182,n183);
and (n192,n179,n181,n188,n183);
and (n193,n180,n181,n188,n183);
and (n194,n180,n185,n188,n183);
nor (n195,n196,n61,n59,n60);
not (n196,n197);
nor (n198,n197,n199,n59,n60);
not (n199,n61);
and (n200,n196,n199,n59,n60);
and (n201,n197,n199,n59,n60);
nor (n202,n203,n204,n206);
not (n204,n205);
and (n207,n203,n205,n206);
nor (n208,n209,n211);
not (n209,n210);
and (n212,n209,n211);
nor (n213,n214,n215,n217,n218);
not (n215,n216);
and (n219,n214,n216,n217,n220);
not (n220,n218);
and (n221,n222,n215,n217,n220);
not (n222,n214);
not (n223,n224);
or (n224,n114,n225);
nand (n225,n226,n241);
or (n226,n227,n240);
nor (n227,n228,n238);
nor (n228,n229,n235);
and (n229,n230,n234);
nand (n230,n231,n232);
or (n231,n77,n79);
wire s0n232,s1n232,notn232;
or (n232,s0n232,s1n232);
not(notn232,n94);
and (s0n232,notn232,n233);
and (s1n232,n94,1'b0);
not (n233,n73);
nor (n234,n95,n96);
not (n235,n236);
wire s0n236,s1n236,notn236;
or (n236,s0n236,s1n236);
not(notn236,n98);
and (s0n236,notn236,n237);
and (s1n236,n98,1'b0);
not (n237,n97);
nand (n238,n239,n101);
not (n239,n109);
or (n240,n104,n103);
not (n241,n112);
wire s0n242,s1n242,notn242;
or (n242,s0n242,s1n242);
not(notn242,n114);
and (s0n242,notn242,n243);
and (s1n242,n114,1'b0);
wire s0n243,s1n243,notn243;
or (n243,s0n243,s1n243);
not(notn243,n112);
and (s0n243,notn243,n244);
and (s1n243,n112,1'b0);
wire s0n244,s1n244,notn244;
or (n244,s0n244,s1n244);
not(notn244,n105);
and (s0n244,notn244,n245);
and (s1n244,n105,n249);
wire s0n245,s1n245,notn245;
or (n245,s0n245,s1n245);
not(notn245,n98);
and (s0n245,notn245,n246);
and (s1n245,n98,1'b1);
wire s0n246,s1n246,notn246;
or (n246,s0n246,s1n246);
not(notn246,n97);
and (s0n246,notn246,n247);
and (s1n246,n97,1'b1);
wire s0n247,s1n247,notn247;
or (n247,s0n247,s1n247);
not(notn247,n96);
and (s0n247,notn247,n248);
and (s1n247,n96,1'b0);
wire s0n248,s1n248,notn248;
or (n248,s0n248,s1n248);
not(notn248,n95);
and (s0n248,notn248,n232);
and (s1n248,n95,1'b0);
not (n249,n240);
not (n250,n251);
wire s0n251,s1n251,notn251;
or (n251,s0n251,s1n251);
not(notn251,n114);
and (s0n251,notn251,n252);
and (s1n251,n114,1'b0);
wire s0n252,s1n252,notn252;
or (n252,s0n252,s1n252);
not(notn252,n112);
and (s0n252,notn252,n253);
and (s1n252,n112,1'b0);
wire s0n253,s1n253,notn253;
or (n253,s0n253,s1n253);
not(notn253,n105);
and (s0n253,notn253,n236);
and (s1n253,n105,1'b0);
and (n254,n255,n258);
xnor (n255,n95,n256);
or (n256,n94,n257);
or (n257,n73,n79);
and (n258,n259,n223,n242,n250);
not (n259,n81);
and (n260,n261,n265);
xnor (n261,n97,n262);
not (n262,n263);
nor (n263,n264,n96);
or (n264,n95,n94);
and (n265,n81,n224,n242,n250);
and (n266,n267,n270);
xnor (n267,n109,n268);
or (n268,n98,n269);
or (n269,n97,n96);
and (n270,n259,n224,n242,n250);
and (n271,n272,n275);
not (n272,n273);
nand (n273,n274,n250,n81,n223);
not (n274,n242);
not (n275,n276);
nand (n276,n277,n103);
or (n277,n102,n278);
not (n278,n279);
nor (n279,n98,n109);
or (n280,n281,n327);
or (n281,n282,n303,n311,n317);
nand (n282,n283,n294);
or (n283,n284,n203);
nand (n284,n285,n292,n205);
nor (n285,n286,n60);
not (n286,n287);
and (n287,n288,n289,n190);
nor (n288,n182,n181);
nor (n289,n290,n180);
not (n290,n291);
nor (n292,n293,n197);
nand (n293,n199,n59);
nor (n294,n295,n297);
and (n295,n285,n296,n210);
nor (n296,n196,n293);
nand (n297,n298,n302);
or (n298,n299,n301);
nor (n299,n300,n288);
and (n300,n181,n190);
nand (n301,n180,n291);
nand (n302,n188,n289,n181);
nor (n303,n304,n309,n168);
nand (n304,n285,n305);
and (n305,n306,n308,n199);
not (n306,n307);
or (n307,n150,n152,n153,n154);
nor (n308,n59,n197);
nor (n309,n310,n165);
and (n310,n167,n166);
nor (n311,n312,n313,n314,n306);
not (n312,n308);
not (n313,n285);
nor (n314,n315,n316);
and (n315,n153,n150);
nor (n316,n150,n154);
nor (n317,n318,n325);
nor (n318,n319,n292);
and (n319,n320,n324);
not (n320,n321);
nor (n321,n322,n323);
and (n322,n308,n61);
and (n323,n197,n199);
not (n324,n60);
nand (n325,n326,n287);
or (n326,n293,n60);
wire s0n327,s1n327,notn327;
or (n327,s0n327,s1n327);
not(notn327,n290);
and (s0n327,notn327,n328);
and (s1n327,n290,1'b0);
wire s0n328,s1n328,notn328;
or (n328,s0n328,s1n328);
not(notn328,n343);
and (s0n328,notn328,n329);
and (s1n328,n343,n342);
wire s0n329,s1n329,notn329;
or (n329,s0n329,s1n329);
not(notn329,n341);
and (s0n329,notn329,n330);
and (s1n329,n341,n333);
wire s0n330,s1n330,notn330;
or (n330,s0n330,s1n330);
not(notn330,n307);
and (s0n330,notn330,n331);
and (s1n330,n307,1'b0);
or (n331,n332,n177);
or (n332,n175,n176);
or (n333,1'b0,n201,n334,n339,1'b0);
and (n334,n335,n338);
or (n335,1'b0,n207,n336,1'b0);
and (n336,n337,n205,n206);
not (n337,n203);
and (n338,n196,n199,n59,n324);
and (n339,n211,n340);
and (n340,n197,n199,n59,n324);
or (n341,n197,n61,n59,n60);
or (n342,n191,n193);
or (n343,n180,n181,n182,n183);
nor (n344,n345,n347,n350);
not (n345,n346);
not (n347,n348);
xor (n348,n349,n346);
xor (n350,n351,n352);
and (n352,n349,n346);
and (n353,n281,n327);
and (n354,n355,n430);
wire s0n355,s1n355,notn355;
or (n355,s0n355,s1n355);
not(notn355,n415);
and (s0n355,notn355,n356);
and (s1n355,n415,n411);
xor (n356,n357,n373);
not (n357,n358);
wire s0n358,s1n358,notn358;
or (n358,s0n358,s1n358);
not(notn358,n280);
and (s0n358,notn358,1'b0);
and (s1n358,n280,n359);
or (n359,n360,n363,n366,n370,1'b0,1'b0,1'b0,1'b0);
and (n360,n361,n80);
xnor (n361,n94,n362);
or (n362,n76,n257);
and (n363,n364,n258);
xnor (n364,n96,n365);
or (n365,n95,n256);
and (n366,n367,n265);
xnor (n367,n98,n368);
not (n368,n369);
and (n369,n263,n237);
and (n370,n371,n270);
xnor (n371,n102,n372);
or (n372,n109,n268);
and (n373,n374,n375);
not (n374,n69);
and (n375,n376,n393);
not (n376,n377);
wire s0n377,s1n377,notn377;
or (n377,s0n377,s1n377);
not(notn377,n280);
and (s0n377,notn377,1'b0);
and (s1n377,n280,n378);
or (n378,n379,n381,n383,n385,n387,n390,1'b0,1'b0);
and (n379,n380,n80);
xnor (n380,n79,n76);
and (n381,n382,n258);
xnor (n382,n94,n257);
and (n383,n384,n265);
xnor (n384,n96,n264);
and (n385,n386,n270);
xnor (n386,n98,n269);
nor (n387,n388,n273);
not (n388,n389);
xnor (n389,n102,n278);
and (n390,n391,n392);
xnor (n391,n104,n107);
nor (n392,n81,n224,n242,n251);
not (n393,n394);
wire s0n394,s1n394,notn394;
or (n394,s0n394,s1n394);
not(notn394,n280);
and (s0n394,notn394,1'b0);
and (s1n394,n280,n395);
or (n395,n396,n398,n400,n402,n404,n406,n408,1'b0);
and (n396,n397,n80);
xnor (n397,n77,n78);
and (n398,n399,n258);
xnor (n399,n73,n79);
and (n400,n401,n265);
xnor (n401,n95,n94);
and (n402,n403,n270);
xnor (n403,n97,n96);
and (n404,n405,n272);
xnor (n405,n109,n98);
and (n406,n407,n392);
xnor (n407,n103,n102);
and (n408,n409,n410);
xnor (n409,n113,n104);
nor (n410,n259,n223,n242,n251);
xor (n411,n358,n412);
and (n412,n69,n413);
and (n413,n377,n414);
and (n414,n394,n415);
wire s0n415,s1n415,notn415;
or (n415,s0n415,s1n415);
not(notn415,n280);
and (s0n415,notn415,1'b0);
and (s1n415,n280,n416);
or (n416,n417,n418,n420,n422,n424,n427,n428,1'b0);
and (n417,n92,n80);
and (n418,n419,n258);
not (n419,n79);
and (n420,n421,n265);
not (n421,n94);
and (n422,n423,n270);
not (n423,n96);
not (n424,n425);
nand (n425,n272,n426);
not (n426,n98);
and (n427,n101,n392);
and (n428,n429,n410);
not (n429,n104);
nor (n430,n431,n281);
not (n431,n327);
and (n432,n69,n433);
and (n433,n281,n431);
not (n434,n435);
nand (n435,n436,n460);
or (n436,n437,n444);
or (n437,n438,n443);
nor (n438,n439,n440,n442);
not (n440,n441);
and (n443,n439,n441,n442);
not (n444,n445);
nand (n445,n446,n454);
or (n446,1'b0,n447,n449,n453);
and (n447,n448,n353);
wire s0n448,s1n448,notn448;
or (n448,s0n448,s1n448);
not(notn448,n344);
and (s0n448,notn448,n377);
and (s1n448,n344,1'b0);
and (n449,n450,n430);
wire s0n450,s1n450,notn450;
or (n450,s0n450,s1n450);
not(notn450,n415);
and (s0n450,notn450,n451);
and (s1n450,n415,n452);
xor (n451,n374,n375);
xor (n452,n69,n413);
and (n453,n377,n433);
or (n454,1'b0,n455,n457,n459);
and (n455,n456,n353);
wire s0n456,s1n456,notn456;
or (n456,s0n456,s1n456);
not(notn456,n344);
and (s0n456,notn456,n394);
and (s1n456,n344,1'b0);
and (n457,n458,n430);
xor (n458,n376,n393);
and (n459,n394,n433);
nor (n460,n461,n484);
not (n461,n462);
or (n462,1'b0,n463,n465,n483);
and (n463,n464,n353);
wire s0n464,s1n464,notn464;
or (n464,s0n464,s1n464);
not(notn464,n344);
and (s0n464,notn464,n358);
and (s1n464,n344,1'b0);
and (n465,n466,n430);
wire s0n466,s1n466,notn466;
or (n466,s0n466,s1n466);
not(notn466,n415);
and (s0n466,notn466,n467);
and (s1n466,n415,n481);
xor (n467,n468,n480);
not (n468,n469);
wire s0n469,s1n469,notn469;
or (n469,s0n469,s1n469);
not(notn469,n280);
and (s0n469,notn469,1'b0);
and (s1n469,n280,n470);
or (n470,n471,n474,n477,1'b0,1'b0,1'b0,1'b0,1'b0);
and (n471,n472,n80);
xnor (n472,n95,n473);
or (n473,n362,n94);
and (n474,n475,n258);
xnor (n475,n97,n476);
or (n476,n96,n365);
and (n477,n478,n265);
xnor (n478,n109,n479);
or (n479,n98,n368);
and (n480,n357,n373);
xor (n481,n469,n482);
and (n482,n358,n412);
and (n483,n358,n433);
nor (n484,n485,n488);
nand (n485,n486,n487);
not (n486,n446);
not (n487,n454);
or (n488,1'b0,n489,n507,n509);
and (n489,n490,n353);
wire s0n490,s1n490,notn490;
or (n490,s0n490,s1n490);
not(notn490,n344);
and (s0n490,notn490,n415);
and (s1n490,n344,n491);
not (n491,n492);
nor (n492,n415,n394,n377,n69,n358,n469,n493,n504);
wire s0n493,s1n493,notn493;
or (n493,s0n493,s1n493);
not(notn493,n280);
and (s0n493,notn493,1'b0);
and (s1n493,n280,n494);
or (n494,n495,n501,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0);
and (n495,n496,n80);
nand (n496,n497,n499);
or (n497,n498,n423);
nor (n498,n362,n264);
nand (n499,n500,n263);
not (n500,n362);
and (n501,n502,n258);
xnor (n502,n98,n503);
or (n503,n97,n476);
wire s0n504,s1n504,notn504;
or (n504,s0n504,s1n504);
not(notn504,n280);
and (s0n504,notn504,1'b0);
and (s1n504,n280,n505);
and (n505,n506,n80);
xnor (n506,n97,n499);
and (n507,n508,n430);
xor (n508,n394,n415);
and (n509,n415,n433);
nand (n510,n511,n65);
or (n511,n512,n514);
not (n512,n513);
nor (n513,n462,n437);
not (n514,n515);
nand (n515,n516,n446);
nand (n516,n517,n487);
not (n517,n488);
nor (n518,n519,n553);
nand (n519,n520,n535,n544);
not (n520,n521);
or (n521,1'b0,n522,n524,n534);
and (n522,n523,n353);
wire s0n523,s1n523,notn523;
or (n523,s0n523,s1n523);
not(notn523,n344);
and (s0n523,notn523,n493);
and (s1n523,n344,1'b0);
and (n524,n525,n430);
wire s0n525,s1n525,notn525;
or (n525,s0n525,s1n525);
not(notn525,n415);
and (s0n525,notn525,n526);
and (s1n525,n415,n531);
xor (n526,n527,n528);
not (n527,n504);
and (n528,n529,n530);
not (n529,n493);
and (n530,n468,n480);
xor (n531,n504,n532);
and (n532,n493,n533);
and (n533,n469,n482);
and (n534,n493,n433);
not (n535,n536);
or (n536,1'b0,n537,n539,n543);
and (n537,n538,n353);
wire s0n538,s1n538,notn538;
or (n538,s0n538,s1n538);
not(notn538,n344);
and (s0n538,notn538,n469);
and (s1n538,n344,1'b0);
and (n539,n540,n430);
wire s0n540,s1n540,notn540;
or (n540,s0n540,s1n540);
not(notn540,n415);
and (s0n540,notn540,n541);
and (s1n540,n415,n542);
xor (n541,n529,n530);
xor (n542,n493,n533);
and (n543,n469,n433);
not (n544,n545);
or (n545,1'b0,n546,n548,n552);
and (n546,n547,n353);
wire s0n547,s1n547,notn547;
or (n547,s0n547,s1n547);
not(notn547,n344);
and (s0n547,notn547,n504);
and (s1n547,n344,1'b0);
and (n548,n549,n430);
wire s0n549,s1n549,notn549;
or (n549,s0n549,s1n549);
not(notn549,n415);
and (s0n549,notn549,n550);
and (s1n549,n415,1'b0);
not (n550,n551);
and (n551,n527,n528);
and (n552,n504,n433);
not (n553,n198);
not (n554,n555);
nor (n555,n556,n558,n559,n560);
not (n556,n557);
and (n561,n562,n38);
not (n562,n52);
nand (n563,n564,n565);
and (n564,n17,n561);
or (n565,1'b0,n566,n568,n572,n575);
and (n566,n567,n555);
and (n568,n569,n570);
nor (n570,n557,n571,n559,n560);
not (n571,n558);
and (n572,n573,n574);
nor (n574,n556,n571,n559,n560);
and (n575,n13,n576);
nor (n576,n557,n558,n577,n560);
not (n577,n559);
nor (n578,n579,n634,n681);
wire s0n579,s1n579,notn579;
or (n579,s0n579,s1n579);
not(notn579,n561);
and (s0n579,notn579,1'b0);
and (s1n579,n561,n580);
wire s0n580,s1n580,notn580;
or (n580,s0n580,s1n580);
not(notn580,n633);
and (s0n580,notn580,n581);
and (s1n580,n633,n624);
or (n581,n582,n600,n611,n622);
and (n582,n583,n24);
wire s0n583,s1n583,notn583;
or (n583,s0n583,s1n583);
not(notn583,n18);
and (s0n583,notn583,n584);
and (s1n583,n18,n585);
or (n585,n586,n591,n595,n598);
and (n586,n587,n588);
nor (n588,n589,n590);
and (n591,n592,n593);
and (n593,n589,n594);
not (n594,n590);
and (n595,n596,n597);
nor (n597,n589,n594);
and (n598,n584,n599);
and (n599,n589,n590);
and (n600,n601,n29);
wire s0n601,s1n601,notn601;
or (n601,s0n601,s1n601);
not(notn601,n18);
and (s0n601,notn601,n602);
and (s1n601,n18,n603);
or (n603,n604,n606,n608,n610);
and (n604,n605,n588);
and (n606,n607,n593);
and (n608,n609,n597);
and (n610,n602,n599);
and (n611,n612,n34);
wire s0n612,s1n612,notn612;
or (n612,s0n612,s1n612);
not(notn612,n18);
and (s0n612,notn612,n613);
and (s1n612,n18,n614);
or (n614,n615,n617,n619,n621);
and (n615,n616,n588);
and (n617,n618,n593);
and (n619,n620,n597);
and (n621,n613,n599);
and (n622,n623,n37);
wire s0n623,s1n623,notn623;
or (n623,s0n623,s1n623);
not(notn623,n18);
and (s0n623,notn623,n624);
and (s1n623,n18,n625);
or (n625,n626,n628,n630,n632);
and (n626,n627,n588);
and (n628,n629,n593);
and (n630,n631,n597);
and (n632,n624,n599);
wire s0n634,s1n634,notn634;
or (n634,s0n634,s1n634);
not(notn634,n561);
and (s0n634,notn634,1'b0);
and (s1n634,n561,n635);
wire s0n635,s1n635,notn635;
or (n635,s0n635,s1n635);
not(notn635,n633);
and (s0n635,notn635,n636);
and (s1n635,n633,n672);
or (n636,n637,n648,n659,n670);
and (n637,n638,n24);
wire s0n638,s1n638,notn638;
or (n638,s0n638,s1n638);
not(notn638,n18);
and (s0n638,notn638,n639);
and (s1n638,n18,n640);
or (n640,n641,n643,n645,n647);
and (n641,n642,n588);
and (n643,n644,n593);
and (n645,n646,n597);
and (n647,n639,n599);
and (n648,n649,n29);
wire s0n649,s1n649,notn649;
or (n649,s0n649,s1n649);
not(notn649,n18);
and (s0n649,notn649,n650);
and (s1n649,n18,n651);
or (n651,n652,n654,n656,n658);
and (n652,n653,n588);
and (n654,n655,n593);
and (n656,n657,n597);
and (n658,n650,n599);
and (n659,n660,n34);
wire s0n660,s1n660,notn660;
or (n660,s0n660,s1n660);
not(notn660,n18);
and (s0n660,notn660,n661);
and (s1n660,n18,n662);
or (n662,n663,n665,n667,n669);
and (n663,n664,n588);
and (n665,n666,n593);
and (n667,n668,n597);
and (n669,n661,n599);
and (n670,n671,n37);
wire s0n671,s1n671,notn671;
or (n671,s0n671,s1n671);
not(notn671,n18);
and (s0n671,notn671,n672);
and (s1n671,n18,n673);
or (n673,n674,n676,n678,n680);
and (n674,n675,n588);
and (n676,n677,n593);
and (n678,n679,n597);
and (n680,n672,n599);
wire s0n681,s1n681,notn681;
or (n681,s0n681,s1n681);
not(notn681,n561);
and (s0n681,notn681,1'b0);
and (s1n681,n561,n682);
wire s0n682,s1n682,notn682;
or (n682,s0n682,s1n682);
not(notn682,n633);
and (s0n682,notn682,n683);
and (s1n682,n633,n719);
or (n683,n684,n695,n706,n717);
and (n684,n685,n24);
wire s0n685,s1n685,notn685;
or (n685,s0n685,s1n685);
not(notn685,n18);
and (s0n685,notn685,n686);
and (s1n685,n18,n687);
or (n687,n688,n690,n692,n694);
and (n688,n689,n588);
and (n690,n691,n593);
and (n692,n693,n597);
and (n694,n686,n599);
and (n695,n696,n29);
wire s0n696,s1n696,notn696;
or (n696,s0n696,s1n696);
not(notn696,n18);
and (s0n696,notn696,n697);
and (s1n696,n18,n698);
or (n698,n699,n701,n703,n705);
and (n699,n700,n588);
and (n701,n702,n593);
and (n703,n704,n597);
and (n705,n697,n599);
and (n706,n707,n34);
wire s0n707,s1n707,notn707;
or (n707,s0n707,s1n707);
not(notn707,n18);
and (s0n707,notn707,n708);
and (s1n707,n18,n709);
or (n709,n710,n712,n714,n716);
and (n710,n711,n588);
and (n712,n713,n593);
and (n714,n715,n597);
and (n716,n708,n599);
and (n717,n718,n37);
wire s0n718,s1n718,notn718;
or (n718,s0n718,s1n718);
not(notn718,n18);
and (s0n718,notn718,n719);
and (s1n718,n18,n720);
or (n720,n721,n723,n725,n727);
and (n721,n722,n588);
and (n723,n724,n593);
and (n725,n726,n597);
and (n727,n719,n599);
or (n728,n729,n870,n928);
and (n729,n730,n751);
xor (n730,n731,n745);
wire s0n731,s1n731,notn731;
or (n731,s0n731,s1n731);
not(notn731,n578);
and (s0n731,notn731,1'b0);
and (s1n731,n578,n732);
nand (n732,n733,n736);
or (n733,n734,n14);
not (n734,n735);
nand (n736,n564,n737);
or (n737,1'b0,n738,n740,n742,n744);
and (n738,n739,n555);
and (n740,n741,n570);
and (n742,n743,n574);
and (n744,n735,n576);
wire s0n745,s1n745,notn745;
or (n745,s0n745,s1n745);
not(notn745,n746);
and (s0n745,notn745,1'b0);
and (s1n745,n746,n10);
xor (n746,n747,n748);
not (n747,n681);
and (n748,n749,n750);
not (n749,n634);
not (n750,n579);
and (n751,n752,n754);
wire s0n752,s1n752,notn752;
or (n752,s0n752,s1n752);
not(notn752,n753);
and (s0n752,notn752,1'b0);
and (s1n752,n753,n10);
xor (n753,n749,n750);
or (n754,n755,n758,n869);
and (n755,n756,n757);
wire s0n756,s1n756,notn756;
or (n756,s0n756,s1n756);
not(notn756,n753);
and (s0n756,notn756,1'b0);
and (s1n756,n753,n732);
wire s0n757,s1n757,notn757;
or (n757,s0n757,s1n757);
not(notn757,n579);
and (s0n757,notn757,1'b0);
and (s1n757,n579,n10);
and (n758,n757,n759);
or (n759,n760,n776,n868);
and (n760,n761,n775);
wire s0n761,s1n761,notn761;
or (n761,s0n761,s1n761);
not(notn761,n753);
and (s0n761,notn761,1'b0);
and (s1n761,n753,n762);
nand (n762,n763,n766);
or (n763,n764,n14);
not (n764,n765);
nand (n766,n564,n767);
or (n767,1'b0,n768,n770,n772,n774);
and (n768,n769,n555);
and (n770,n771,n570);
and (n772,n773,n574);
and (n774,n765,n576);
wire s0n775,s1n775,notn775;
or (n775,s0n775,s1n775);
not(notn775,n579);
and (s0n775,notn775,1'b0);
and (s1n775,n579,n732);
and (n776,n775,n777);
or (n777,n778,n794,n867);
and (n778,n779,n793);
wire s0n779,s1n779,notn779;
or (n779,s0n779,s1n779);
not(notn779,n753);
and (s0n779,notn779,1'b0);
and (s1n779,n753,n780);
nand (n780,n781,n784);
or (n781,n782,n14);
not (n782,n783);
nand (n784,n564,n785);
or (n785,1'b0,n786,n788,n790,n792);
and (n786,n787,n555);
and (n788,n789,n570);
and (n790,n791,n574);
and (n792,n783,n576);
wire s0n793,s1n793,notn793;
or (n793,s0n793,s1n793);
not(notn793,n579);
and (s0n793,notn793,1'b0);
and (s1n793,n579,n762);
and (n794,n793,n795);
or (n795,n796,n812,n866);
and (n796,n797,n811);
wire s0n797,s1n797,notn797;
or (n797,s0n797,s1n797);
not(notn797,n753);
and (s0n797,notn797,1'b0);
and (s1n797,n753,n798);
nand (n798,n799,n802);
or (n799,n800,n14);
not (n800,n801);
nand (n802,n564,n803);
or (n803,1'b0,n804,n806,n808,n810);
and (n804,n805,n555);
and (n806,n807,n570);
and (n808,n809,n574);
and (n810,n801,n576);
wire s0n811,s1n811,notn811;
or (n811,s0n811,s1n811);
not(notn811,n579);
and (s0n811,notn811,1'b0);
and (s1n811,n579,n780);
and (n812,n811,n813);
or (n813,n814,n830,n832);
and (n814,n815,n829);
wire s0n815,s1n815,notn815;
or (n815,s0n815,s1n815);
not(notn815,n753);
and (s0n815,notn815,1'b0);
and (s1n815,n753,n816);
nand (n816,n817,n820);
or (n817,n818,n14);
not (n818,n819);
nand (n820,n564,n821);
or (n821,1'b0,n822,n824,n826,n828);
and (n822,n823,n555);
and (n824,n825,n570);
and (n826,n827,n574);
and (n828,n819,n576);
wire s0n829,s1n829,notn829;
or (n829,s0n829,s1n829);
not(notn829,n579);
and (s0n829,notn829,1'b0);
and (s1n829,n579,n798);
and (n830,n829,n831);
or (n831,n832,n848,n849);
and (n832,n833,n847);
wire s0n833,s1n833,notn833;
or (n833,s0n833,s1n833);
not(notn833,n753);
and (s0n833,notn833,1'b0);
and (s1n833,n753,n834);
nand (n834,n835,n838);
or (n835,n836,n14);
not (n836,n837);
nand (n838,n564,n839);
or (n839,1'b0,n840,n842,n844,n846);
and (n840,n841,n555);
and (n842,n843,n570);
and (n844,n845,n574);
and (n846,n837,n576);
wire s0n847,s1n847,notn847;
or (n847,s0n847,s1n847);
not(notn847,n579);
and (s0n847,notn847,1'b0);
and (s1n847,n579,n816);
and (n848,n847,n849);
and (n849,n850,n865);
wire s0n850,s1n850,notn850;
or (n850,s0n850,s1n850);
not(notn850,n753);
and (s0n850,notn850,1'b0);
and (s1n850,n753,n851);
nand (n851,n852,n864);
or (n852,n853,n863);
not (n853,n854);
or (n854,1'b0,n855,n857,n859,n861);
and (n855,n856,n555);
and (n857,n858,n570);
and (n859,n860,n574);
and (n861,n862,n576);
not (n863,n564);
nand (n864,n15,n862);
wire s0n865,s1n865,notn865;
or (n865,s0n865,s1n865);
not(notn865,n579);
and (s0n865,notn865,1'b0);
and (s1n865,n579,n834);
and (n866,n797,n813);
and (n867,n779,n795);
and (n868,n761,n777);
and (n869,n756,n759);
and (n870,n751,n871);
or (n871,n872,n877,n927);
and (n872,n873,n876);
xor (n873,n874,n875);
wire s0n874,s1n874,notn874;
or (n874,s0n874,s1n874);
not(notn874,n578);
and (s0n874,notn874,1'b0);
and (s1n874,n578,n762);
wire s0n875,s1n875,notn875;
or (n875,s0n875,s1n875);
not(notn875,n746);
and (s0n875,notn875,1'b0);
and (s1n875,n746,n732);
xor (n876,n752,n754);
and (n877,n876,n878);
or (n878,n879,n885,n926);
and (n879,n880,n883);
xor (n880,n881,n882);
wire s0n881,s1n881,notn881;
or (n881,s0n881,s1n881);
not(notn881,n578);
and (s0n881,notn881,1'b0);
and (s1n881,n578,n780);
wire s0n882,s1n882,notn882;
or (n882,s0n882,s1n882);
not(notn882,n746);
and (s0n882,notn882,1'b0);
and (s1n882,n746,n762);
xor (n883,n884,n759);
xor (n884,n756,n757);
and (n885,n883,n886);
or (n886,n887,n893,n925);
and (n887,n888,n891);
xor (n888,n889,n890);
wire s0n889,s1n889,notn889;
or (n889,s0n889,s1n889);
not(notn889,n578);
and (s0n889,notn889,1'b0);
and (s1n889,n578,n798);
wire s0n890,s1n890,notn890;
or (n890,s0n890,s1n890);
not(notn890,n746);
and (s0n890,notn890,1'b0);
and (s1n890,n746,n780);
xor (n891,n892,n777);
xor (n892,n761,n775);
and (n893,n891,n894);
or (n894,n895,n901,n924);
and (n895,n896,n899);
xor (n896,n897,n898);
wire s0n897,s1n897,notn897;
or (n897,s0n897,s1n897);
not(notn897,n578);
and (s0n897,notn897,1'b0);
and (s1n897,n578,n816);
wire s0n898,s1n898,notn898;
or (n898,s0n898,s1n898);
not(notn898,n746);
and (s0n898,notn898,1'b0);
and (s1n898,n746,n798);
xor (n899,n900,n795);
xor (n900,n779,n793);
and (n901,n899,n902);
or (n902,n903,n909,n923);
and (n903,n904,n907);
xor (n904,n905,n906);
wire s0n905,s1n905,notn905;
or (n905,s0n905,s1n905);
not(notn905,n578);
and (s0n905,notn905,1'b0);
and (s1n905,n578,n834);
wire s0n906,s1n906,notn906;
or (n906,s0n906,s1n906);
not(notn906,n746);
and (s0n906,notn906,1'b0);
and (s1n906,n746,n816);
xor (n907,n908,n813);
xor (n908,n797,n811);
and (n909,n907,n910);
or (n910,n911,n917,n922);
and (n911,n912,n915);
xor (n912,n913,n914);
wire s0n913,s1n913,notn913;
or (n913,s0n913,s1n913);
not(notn913,n578);
and (s0n913,notn913,1'b0);
and (s1n913,n578,n851);
wire s0n914,s1n914,notn914;
or (n914,s0n914,s1n914);
not(notn914,n746);
and (s0n914,notn914,1'b0);
and (s1n914,n746,n834);
xor (n915,n916,n831);
xor (n916,n815,n829);
and (n917,n915,n918);
and (n918,n919,n920);
wire s0n919,s1n919,notn919;
or (n919,s0n919,s1n919);
not(notn919,n746);
and (s0n919,notn919,1'b0);
and (s1n919,n746,n851);
xor (n920,n921,n849);
xor (n921,n833,n847);
and (n922,n912,n918);
and (n923,n904,n910);
and (n924,n896,n902);
and (n925,n888,n894);
and (n926,n880,n886);
and (n927,n873,n878);
and (n928,n730,n871);
nor (n929,n930,n977,n1024);
wire s0n930,s1n930,notn930;
or (n930,s0n930,s1n930);
not(notn930,n561);
and (s0n930,notn930,1'b0);
and (s1n930,n561,n931);
wire s0n931,s1n931,notn931;
or (n931,s0n931,s1n931);
not(notn931,n633);
and (s0n931,notn931,n932);
and (s1n931,n633,n968);
or (n932,n933,n944,n955,n966);
and (n933,n934,n24);
wire s0n934,s1n934,notn934;
or (n934,s0n934,s1n934);
not(notn934,n18);
and (s0n934,notn934,n935);
and (s1n934,n18,n936);
or (n936,n937,n939,n941,n943);
and (n937,n938,n588);
and (n939,n940,n593);
and (n941,n942,n597);
and (n943,n935,n599);
and (n944,n945,n29);
wire s0n945,s1n945,notn945;
or (n945,s0n945,s1n945);
not(notn945,n18);
and (s0n945,notn945,n946);
and (s1n945,n18,n947);
or (n947,n948,n950,n952,n954);
and (n948,n949,n588);
and (n950,n951,n593);
and (n952,n953,n597);
and (n954,n946,n599);
and (n955,n956,n34);
wire s0n956,s1n956,notn956;
or (n956,s0n956,s1n956);
not(notn956,n18);
and (s0n956,notn956,n957);
and (s1n956,n18,n958);
or (n958,n959,n961,n963,n965);
and (n959,n960,n588);
and (n961,n962,n593);
and (n963,n964,n597);
and (n965,n957,n599);
and (n966,n967,n37);
wire s0n967,s1n967,notn967;
or (n967,s0n967,s1n967);
not(notn967,n18);
and (s0n967,notn967,n968);
and (s1n967,n18,n969);
or (n969,n970,n972,n974,n976);
and (n970,n971,n588);
and (n972,n973,n593);
and (n974,n975,n597);
and (n976,n968,n599);
wire s0n977,s1n977,notn977;
or (n977,s0n977,s1n977);
not(notn977,n561);
and (s0n977,notn977,1'b0);
and (s1n977,n561,n978);
wire s0n978,s1n978,notn978;
or (n978,s0n978,s1n978);
not(notn978,n633);
and (s0n978,notn978,n979);
and (s1n978,n633,n1015);
or (n979,n980,n991,n1002,n1013);
and (n980,n981,n24);
wire s0n981,s1n981,notn981;
or (n981,s0n981,s1n981);
not(notn981,n18);
and (s0n981,notn981,n982);
and (s1n981,n18,n983);
or (n983,n984,n986,n988,n990);
and (n984,n985,n588);
and (n986,n987,n593);
and (n988,n989,n597);
and (n990,n982,n599);
and (n991,n992,n29);
wire s0n992,s1n992,notn992;
or (n992,s0n992,s1n992);
not(notn992,n18);
and (s0n992,notn992,n993);
and (s1n992,n18,n994);
or (n994,n995,n997,n999,n1001);
and (n995,n996,n588);
and (n997,n998,n593);
and (n999,n1000,n597);
and (n1001,n993,n599);
and (n1002,n1003,n34);
wire s0n1003,s1n1003,notn1003;
or (n1003,s0n1003,s1n1003);
not(notn1003,n18);
and (s0n1003,notn1003,n1004);
and (s1n1003,n18,n1005);
or (n1005,n1006,n1008,n1010,n1012);
and (n1006,n1007,n588);
and (n1008,n1009,n593);
and (n1010,n1011,n597);
and (n1012,n1004,n599);
and (n1013,n1014,n37);
wire s0n1014,s1n1014,notn1014;
or (n1014,s0n1014,s1n1014);
not(notn1014,n18);
and (s0n1014,notn1014,n1015);
and (s1n1014,n18,n1016);
or (n1016,n1017,n1019,n1021,n1023);
and (n1017,n1018,n588);
and (n1019,n1020,n593);
and (n1021,n1022,n597);
and (n1023,n1015,n599);
wire s0n1024,s1n1024,notn1024;
or (n1024,s0n1024,s1n1024);
not(notn1024,n561);
and (s0n1024,notn1024,1'b0);
and (s1n1024,n561,n1025);
wire s0n1025,s1n1025,notn1025;
or (n1025,s0n1025,s1n1025);
not(notn1025,n633);
and (s0n1025,notn1025,n1026);
and (s1n1025,n633,n1062);
or (n1026,n1027,n1038,n1049,n1060);
and (n1027,n1028,n24);
wire s0n1028,s1n1028,notn1028;
or (n1028,s0n1028,s1n1028);
not(notn1028,n18);
and (s0n1028,notn1028,n1029);
and (s1n1028,n18,n1030);
or (n1030,n1031,n1033,n1035,n1037);
and (n1031,n1032,n588);
and (n1033,n1034,n593);
and (n1035,n1036,n597);
and (n1037,n1029,n599);
and (n1038,n1039,n29);
wire s0n1039,s1n1039,notn1039;
or (n1039,s0n1039,s1n1039);
not(notn1039,n18);
and (s0n1039,notn1039,n1040);
and (s1n1039,n18,n1041);
or (n1041,n1042,n1044,n1046,n1048);
and (n1042,n1043,n588);
and (n1044,n1045,n593);
and (n1046,n1047,n597);
and (n1048,n1040,n599);
and (n1049,n1050,n34);
wire s0n1050,s1n1050,notn1050;
or (n1050,s0n1050,s1n1050);
not(notn1050,n18);
and (s0n1050,notn1050,n1051);
and (s1n1050,n18,n1052);
or (n1052,n1053,n1055,n1057,n1059);
and (n1053,n1054,n588);
and (n1055,n1056,n593);
and (n1057,n1058,n597);
and (n1059,n1051,n599);
and (n1060,n1061,n37);
wire s0n1061,s1n1061,notn1061;
or (n1061,s0n1061,s1n1061);
not(notn1061,n18);
and (s0n1061,notn1061,n1062);
and (s1n1061,n18,n1063);
or (n1063,n1064,n1066,n1068,n1070);
and (n1064,n1065,n588);
and (n1066,n1067,n593);
and (n1068,n1069,n597);
and (n1070,n1062,n599);
or (n1071,n1072,n1205,n1290);
and (n1072,n1073,n1083);
xor (n1073,n1074,n1077);
wire s0n1074,s1n1074,notn1074;
or (n1074,s0n1074,s1n1074);
not(notn1074,n929);
and (s0n1074,notn1074,1'b0);
and (s1n1074,n929,n1075);
xor (n1075,n1076,n871);
xor (n1076,n730,n751);
wire s0n1077,s1n1077,notn1077;
or (n1077,s0n1077,s1n1077);
not(notn1077,n1078);
and (s0n1077,notn1077,1'b0);
and (s1n1077,n1078,n8);
xor (n1078,n1079,n1080);
not (n1079,n1024);
and (n1080,n1081,n1082);
not (n1081,n977);
not (n1082,n930);
and (n1083,n1084,n1086);
wire s0n1084,s1n1084,notn1084;
or (n1084,s0n1084,s1n1084);
not(notn1084,n1085);
and (s0n1084,notn1084,1'b0);
and (s1n1084,n1085,n8);
xor (n1085,n1081,n1082);
or (n1086,n1087,n1090,n1204);
and (n1087,n1088,n1089);
wire s0n1088,s1n1088,notn1088;
or (n1088,s0n1088,s1n1088);
not(notn1088,n1085);
and (s0n1088,notn1088,1'b0);
and (s1n1088,n1085,n1075);
wire s0n1089,s1n1089,notn1089;
or (n1089,s0n1089,s1n1089);
not(notn1089,n930);
and (s0n1089,notn1089,1'b0);
and (s1n1089,n930,n8);
and (n1090,n1089,n1091);
or (n1091,n1092,n1097,n1203);
and (n1092,n1093,n1096);
wire s0n1093,s1n1093,notn1093;
or (n1093,s0n1093,s1n1093);
not(notn1093,n1085);
and (s0n1093,notn1093,1'b0);
and (s1n1093,n1085,n1094);
xor (n1094,n1095,n878);
xor (n1095,n873,n876);
wire s0n1096,s1n1096,notn1096;
or (n1096,s0n1096,s1n1096);
not(notn1096,n930);
and (s0n1096,notn1096,1'b0);
and (s1n1096,n930,n1075);
and (n1097,n1096,n1098);
or (n1098,n1099,n1153,n1202);
and (n1099,n1100,n1152);
and (n1100,n1101,n1085);
xor (n1101,n1102,n1114);
nor (n1102,n1103,n1113);
not (n1103,n1104);
or (n1104,n1105,n1108);
xor (n1105,n1106,n760);
xor (n1106,n882,n1107);
xor (n1107,n884,n881);
or (n1108,n1109,n1112);
and (n1109,n1110,n778);
xor (n1110,n890,n1111);
xor (n1111,n892,n889);
and (n1112,n890,n1111);
and (n1113,n1105,n1108);
nand (n1114,n1115,n1151);
or (n1115,n1116,n1124);
not (n1116,n1117);
or (n1117,n1118,n1119);
xor (n1118,n1110,n778);
or (n1119,n1120,n1123);
and (n1120,n1121,n796);
xor (n1121,n898,n1122);
xor (n1122,n900,n897);
and (n1123,n898,n1122);
not (n1124,n1125);
nand (n1125,n1126,n1147,n1150);
nand (n1126,n1127,n1134,n1144);
or (n1127,n1128,n1129);
xor (n1128,n1121,n796);
or (n1129,n1130,n1133);
and (n1130,n1131,n1132);
xor (n1131,n906,n814);
xor (n1132,n908,n905);
and (n1133,n906,n814);
or (n1134,n1135,n1143);
and (n1135,n1136,n1141);
xor (n1136,n832,n1137);
or (n1137,n1138,n1140);
and (n1138,n1139,n921);
xor (n1139,n849,n919);
and (n1140,n849,n919);
xor (n1141,n1142,n914);
xor (n1142,n913,n916);
and (n1143,n832,n1137);
or (n1144,n1145,n1146);
xor (n1145,n1131,n1132);
and (n1146,n1142,n914);
nand (n1147,n1148,n1127);
not (n1148,n1149);
nand (n1149,n1145,n1146);
nand (n1150,n1128,n1129);
nand (n1151,n1118,n1119);
wire s0n1152,s1n1152,notn1152;
or (n1152,s0n1152,s1n1152);
not(notn1152,n930);
and (s0n1152,notn1152,1'b0);
and (s1n1152,n930,n1094);
and (n1153,n1152,n1154);
or (n1154,n1155,n1160,n1201);
and (n1155,n1156,n1159);
and (n1156,n1157,n1085);
xnor (n1157,n1125,n1158);
nand (n1158,n1117,n1151);
and (n1159,n1101,n930);
and (n1160,n1159,n1161);
or (n1161,n1162,n1167,n1200);
and (n1162,n1163,n1166);
wire s0n1163,s1n1163,notn1163;
or (n1163,s0n1163,s1n1163);
not(notn1163,n1085);
and (s0n1163,notn1163,1'b0);
and (s1n1163,n1085,n1164);
xor (n1164,n1165,n902);
xor (n1165,n896,n899);
and (n1166,n1157,n930);
and (n1167,n1166,n1168);
or (n1168,n1169,n1174,n1199);
and (n1169,n1170,n1173);
wire s0n1170,s1n1170,notn1170;
or (n1170,s0n1170,s1n1170);
not(notn1170,n1085);
and (s0n1170,notn1170,1'b0);
and (s1n1170,n1085,n1171);
xor (n1171,n1172,n910);
xor (n1172,n904,n907);
wire s0n1173,s1n1173,notn1173;
or (n1173,s0n1173,s1n1173);
not(notn1173,n930);
and (s0n1173,notn1173,1'b0);
and (s1n1173,n930,n1164);
and (n1174,n1173,n1175);
or (n1175,n1176,n1181,n1198);
and (n1176,n1177,n1180);
wire s0n1177,s1n1177,notn1177;
or (n1177,s0n1177,s1n1177);
not(notn1177,n1085);
and (s0n1177,notn1177,1'b0);
and (s1n1177,n1085,n1178);
xor (n1178,n1179,n918);
xor (n1179,n912,n915);
wire s0n1180,s1n1180,notn1180;
or (n1180,s0n1180,s1n1180);
not(notn1180,n930);
and (s0n1180,notn1180,1'b0);
and (s1n1180,n930,n1171);
and (n1181,n1180,n1182);
or (n1182,n1183,n1187,n1189);
and (n1183,n1184,n1186);
wire s0n1184,s1n1184,notn1184;
or (n1184,s0n1184,s1n1184);
not(notn1184,n1085);
and (s0n1184,notn1184,1'b0);
and (s1n1184,n1085,n1185);
xor (n1185,n919,n920);
wire s0n1186,s1n1186,notn1186;
or (n1186,s0n1186,s1n1186);
not(notn1186,n930);
and (s0n1186,notn1186,1'b0);
and (s1n1186,n930,n1178);
and (n1187,n1186,n1188);
or (n1188,n1189,n1193,n1194);
and (n1189,n1190,n1192);
wire s0n1190,s1n1190,notn1190;
or (n1190,s0n1190,s1n1190);
not(notn1190,n1085);
and (s0n1190,notn1190,1'b0);
and (s1n1190,n1085,n1191);
xor (n1191,n850,n865);
wire s0n1192,s1n1192,notn1192;
or (n1192,s0n1192,s1n1192);
not(notn1192,n930);
and (s0n1192,notn1192,1'b0);
and (s1n1192,n930,n1185);
and (n1193,n1192,n1194);
and (n1194,n1195,n1197);
wire s0n1195,s1n1195,notn1195;
or (n1195,s0n1195,s1n1195);
not(notn1195,n1085);
and (s0n1195,notn1195,1'b0);
and (s1n1195,n1085,n1196);
wire s0n1196,s1n1196,notn1196;
or (n1196,s0n1196,s1n1196);
not(notn1196,n579);
and (s0n1196,notn1196,1'b0);
and (s1n1196,n579,n851);
wire s0n1197,s1n1197,notn1197;
or (n1197,s0n1197,s1n1197);
not(notn1197,n930);
and (s0n1197,notn1197,1'b0);
and (s1n1197,n930,n1191);
and (n1198,n1177,n1182);
and (n1199,n1170,n1175);
and (n1200,n1163,n1168);
and (n1201,n1156,n1161);
and (n1202,n1100,n1154);
and (n1203,n1093,n1098);
and (n1204,n1088,n1091);
and (n1205,n1083,n1206);
or (n1206,n1207,n1212,n1289);
and (n1207,n1208,n1211);
xor (n1208,n1209,n1210);
wire s0n1209,s1n1209,notn1209;
or (n1209,s0n1209,s1n1209);
not(notn1209,n929);
and (s0n1209,notn1209,1'b0);
and (s1n1209,n929,n1094);
wire s0n1210,s1n1210,notn1210;
or (n1210,s0n1210,s1n1210);
not(notn1210,n1078);
and (s0n1210,notn1210,1'b0);
and (s1n1210,n1078,n1075);
xor (n1211,n1084,n1086);
and (n1212,n1211,n1213);
or (n1213,n1214,n1220,n1288);
and (n1214,n1215,n1218);
xor (n1215,n1216,n1217);
and (n1216,n1101,n929);
wire s0n1217,s1n1217,notn1217;
or (n1217,s0n1217,s1n1217);
not(notn1217,n1078);
and (s0n1217,notn1217,1'b0);
and (s1n1217,n1078,n1094);
xor (n1218,n1219,n1091);
xor (n1219,n1088,n1089);
and (n1220,n1218,n1221);
or (n1221,n1222,n1228,n1287);
and (n1222,n1223,n1226);
xor (n1223,n1224,n1225);
and (n1224,n1157,n929);
and (n1225,n1101,n1078);
xor (n1226,n1227,n1098);
xor (n1227,n1093,n1096);
and (n1228,n1226,n1229);
or (n1229,n1230,n1236,n1286);
and (n1230,n1231,n1234);
xor (n1231,n1232,n1233);
wire s0n1232,s1n1232,notn1232;
or (n1232,s0n1232,s1n1232);
not(notn1232,n929);
and (s0n1232,notn1232,1'b0);
and (s1n1232,n929,n1164);
and (n1233,n1157,n1078);
xor (n1234,n1235,n1154);
xor (n1235,n1100,n1152);
and (n1236,n1234,n1237);
or (n1237,n1238,n1244,n1285);
and (n1238,n1239,n1242);
xor (n1239,n1240,n1241);
wire s0n1240,s1n1240,notn1240;
or (n1240,s0n1240,s1n1240);
not(notn1240,n929);
and (s0n1240,notn1240,1'b0);
and (s1n1240,n929,n1171);
wire s0n1241,s1n1241,notn1241;
or (n1241,s0n1241,s1n1241);
not(notn1241,n1078);
and (s0n1241,notn1241,1'b0);
and (s1n1241,n1078,n1164);
xor (n1242,n1243,n1161);
xor (n1243,n1156,n1159);
and (n1244,n1242,n1245);
or (n1245,n1246,n1252,n1284);
and (n1246,n1247,n1250);
xor (n1247,n1248,n1249);
wire s0n1248,s1n1248,notn1248;
or (n1248,s0n1248,s1n1248);
not(notn1248,n929);
and (s0n1248,notn1248,1'b0);
and (s1n1248,n929,n1178);
wire s0n1249,s1n1249,notn1249;
or (n1249,s0n1249,s1n1249);
not(notn1249,n1078);
and (s0n1249,notn1249,1'b0);
and (s1n1249,n1078,n1171);
xor (n1250,n1251,n1168);
xor (n1251,n1163,n1166);
and (n1252,n1250,n1253);
or (n1253,n1254,n1260,n1283);
and (n1254,n1255,n1258);
xor (n1255,n1256,n1257);
wire s0n1256,s1n1256,notn1256;
or (n1256,s0n1256,s1n1256);
not(notn1256,n929);
and (s0n1256,notn1256,1'b0);
and (s1n1256,n929,n1185);
wire s0n1257,s1n1257,notn1257;
or (n1257,s0n1257,s1n1257);
not(notn1257,n1078);
and (s0n1257,notn1257,1'b0);
and (s1n1257,n1078,n1178);
xor (n1258,n1259,n1175);
xor (n1259,n1170,n1173);
and (n1260,n1258,n1261);
or (n1261,n1262,n1268,n1282);
and (n1262,n1263,n1266);
xor (n1263,n1264,n1265);
wire s0n1264,s1n1264,notn1264;
or (n1264,s0n1264,s1n1264);
not(notn1264,n929);
and (s0n1264,notn1264,1'b0);
and (s1n1264,n929,n1191);
wire s0n1265,s1n1265,notn1265;
or (n1265,s0n1265,s1n1265);
not(notn1265,n1078);
and (s0n1265,notn1265,1'b0);
and (s1n1265,n1078,n1185);
xor (n1266,n1267,n1182);
xor (n1267,n1177,n1180);
and (n1268,n1266,n1269);
or (n1269,n1270,n1276,n1281);
and (n1270,n1271,n1274);
xor (n1271,n1272,n1273);
wire s0n1272,s1n1272,notn1272;
or (n1272,s0n1272,s1n1272);
not(notn1272,n929);
and (s0n1272,notn1272,1'b0);
and (s1n1272,n929,n1196);
wire s0n1273,s1n1273,notn1273;
or (n1273,s0n1273,s1n1273);
not(notn1273,n1078);
and (s0n1273,notn1273,1'b0);
and (s1n1273,n1078,n1191);
xor (n1274,n1275,n1188);
xor (n1275,n1184,n1186);
and (n1276,n1274,n1277);
and (n1277,n1278,n1279);
wire s0n1278,s1n1278,notn1278;
or (n1278,s0n1278,s1n1278);
not(notn1278,n1078);
and (s0n1278,notn1278,1'b0);
and (s1n1278,n1078,n1196);
xor (n1279,n1280,n1194);
xor (n1280,n1190,n1192);
and (n1281,n1271,n1277);
and (n1282,n1263,n1269);
and (n1283,n1255,n1261);
and (n1284,n1247,n1253);
and (n1285,n1239,n1245);
and (n1286,n1231,n1237);
and (n1287,n1223,n1229);
and (n1288,n1215,n1221);
and (n1289,n1208,n1213);
and (n1290,n1073,n1206);
xor (n1291,n1292,n1492);
wire s0n1292,s1n1292,notn1292;
or (n1292,s0n1292,s1n1292);
not(notn1292,n929);
and (s0n1292,notn1292,1'b0);
and (s1n1292,n929,n1293);
or (n1293,n1294,n1439,n1491);
and (n1294,n1295,n1309);
and (n1295,n681,n1296);
nand (n1296,n1297,n1300);
or (n1297,n1298,n14);
not (n1298,n1299);
nand (n1300,n564,n1301);
or (n1301,1'b0,n1302,n1304,n1306,n1308);
and (n1302,n1303,n555);
and (n1304,n1305,n570);
and (n1306,n1307,n574);
and (n1308,n1299,n576);
and (n1309,n1310,n1311);
wire s0n1310,s1n1310,notn1310;
or (n1310,s0n1310,s1n1310);
not(notn1310,n634);
and (s0n1310,notn1310,1'b0);
and (s1n1310,n634,n1296);
or (n1311,n1312,n1328,n1438);
and (n1312,n1313,n1327);
wire s0n1313,s1n1313,notn1313;
or (n1313,s0n1313,s1n1313);
not(notn1313,n634);
and (s0n1313,notn1313,1'b0);
and (s1n1313,n634,n1314);
nand (n1314,n1315,n1318);
or (n1315,n1316,n14);
not (n1316,n1317);
nand (n1318,n564,n1319);
or (n1319,1'b0,n1320,n1322,n1324,n1326);
and (n1320,n1321,n555);
and (n1322,n1323,n570);
and (n1324,n1325,n574);
and (n1326,n1317,n576);
wire s0n1327,s1n1327,notn1327;
or (n1327,s0n1327,s1n1327);
not(notn1327,n579);
and (s0n1327,notn1327,1'b0);
and (s1n1327,n579,n1296);
and (n1328,n1327,n1329);
or (n1329,n1330,n1346,n1437);
and (n1330,n1331,n1345);
wire s0n1331,s1n1331,notn1331;
or (n1331,s0n1331,s1n1331);
not(notn1331,n634);
and (s0n1331,notn1331,1'b0);
and (s1n1331,n634,n1332);
nand (n1332,n1333,n1344);
or (n1333,n1334,n863);
not (n1334,n1335);
or (n1335,1'b0,n1336,n1338,n1340,n1342);
and (n1336,n1337,n555);
and (n1338,n1339,n570);
and (n1340,n1341,n574);
and (n1342,n1343,n576);
nand (n1344,n15,n1343);
wire s0n1345,s1n1345,notn1345;
or (n1345,s0n1345,s1n1345);
not(notn1345,n579);
and (s0n1345,notn1345,1'b0);
and (s1n1345,n579,n1314);
and (n1346,n1345,n1347);
or (n1347,n1348,n1364,n1436);
and (n1348,n1349,n1363);
wire s0n1349,s1n1349,notn1349;
or (n1349,s0n1349,s1n1349);
not(notn1349,n634);
and (s0n1349,notn1349,1'b0);
and (s1n1349,n634,n1350);
nand (n1350,n1351,n1362);
or (n1351,n1352,n863);
not (n1352,n1353);
or (n1353,1'b0,n1354,n1356,n1358,n1360);
and (n1354,n1355,n555);
and (n1356,n1357,n570);
and (n1358,n1359,n574);
and (n1360,n1361,n576);
nand (n1362,n15,n1361);
wire s0n1363,s1n1363,notn1363;
or (n1363,s0n1363,s1n1363);
not(notn1363,n579);
and (s0n1363,notn1363,1'b0);
and (s1n1363,n579,n1332);
and (n1364,n1363,n1365);
or (n1365,n1366,n1382,n1435);
and (n1366,n1367,n1381);
wire s0n1367,s1n1367,notn1367;
or (n1367,s0n1367,s1n1367);
not(notn1367,n634);
and (s0n1367,notn1367,1'b0);
and (s1n1367,n634,n1368);
nand (n1368,n1369,n1372);
or (n1369,n1370,n14);
not (n1370,n1371);
nand (n1372,n564,n1373);
or (n1373,1'b0,n1374,n1376,n1378,n1380);
and (n1374,n1375,n555);
and (n1376,n1377,n570);
and (n1378,n1379,n574);
and (n1380,n1371,n576);
wire s0n1381,s1n1381,notn1381;
or (n1381,s0n1381,s1n1381);
not(notn1381,n579);
and (s0n1381,notn1381,1'b0);
and (s1n1381,n579,n1350);
and (n1382,n1381,n1383);
or (n1383,n1384,n1400,n1402);
and (n1384,n1385,n1399);
wire s0n1385,s1n1385,notn1385;
or (n1385,s0n1385,s1n1385);
not(notn1385,n634);
and (s0n1385,notn1385,1'b0);
and (s1n1385,n634,n1386);
nand (n1386,n1387,n1398);
or (n1387,n1388,n863);
not (n1388,n1389);
or (n1389,1'b0,n1390,n1392,n1394,n1396);
and (n1390,n1391,n555);
and (n1392,n1393,n570);
and (n1394,n1395,n574);
and (n1396,n1397,n576);
nand (n1398,n15,n1397);
wire s0n1399,s1n1399,notn1399;
or (n1399,s0n1399,s1n1399);
not(notn1399,n579);
and (s0n1399,notn1399,1'b0);
and (s1n1399,n579,n1368);
and (n1400,n1399,n1401);
or (n1401,n1402,n1418,n1419);
and (n1402,n1403,n1417);
wire s0n1403,s1n1403,notn1403;
or (n1403,s0n1403,s1n1403);
not(notn1403,n634);
and (s0n1403,notn1403,1'b0);
and (s1n1403,n634,n1404);
nand (n1404,n1405,n1408);
or (n1405,n1406,n14);
not (n1406,n1407);
nand (n1408,n564,n1409);
or (n1409,1'b0,n1410,n1412,n1414,n1416);
and (n1410,n1411,n555);
and (n1412,n1413,n570);
and (n1414,n1415,n574);
and (n1416,n1407,n576);
wire s0n1417,s1n1417,notn1417;
or (n1417,s0n1417,s1n1417);
not(notn1417,n579);
and (s0n1417,notn1417,1'b0);
and (s1n1417,n579,n1386);
and (n1418,n1417,n1419);
and (n1419,n1420,n1434);
wire s0n1420,s1n1420,notn1420;
or (n1420,s0n1420,s1n1420);
not(notn1420,n634);
and (s0n1420,notn1420,1'b0);
and (s1n1420,n634,n1421);
nand (n1421,n1422,n1425);
or (n1422,n1423,n14);
not (n1423,n1424);
nand (n1425,n564,n1426);
or (n1426,1'b0,n1427,n1429,n1431,n1433);
and (n1427,n1428,n555);
and (n1429,n1430,n570);
and (n1431,n1432,n574);
and (n1433,n1424,n576);
wire s0n1434,s1n1434,notn1434;
or (n1434,s0n1434,s1n1434);
not(notn1434,n579);
and (s0n1434,notn1434,1'b0);
and (s1n1434,n579,n1404);
and (n1435,n1367,n1383);
and (n1436,n1349,n1365);
and (n1437,n1331,n1347);
and (n1438,n1313,n1329);
and (n1439,n1309,n1440);
or (n1440,n1441,n1445,n1490);
and (n1441,n1442,n1444);
not (n1442,n1443);
nand (n1443,n681,n1314);
xor (n1444,n1310,n1311);
and (n1445,n1444,n1446);
or (n1446,n1447,n1452,n1489);
and (n1447,n1448,n1450);
not (n1448,n1449);
nand (n1449,n681,n1332);
xor (n1450,n1451,n1329);
xor (n1451,n1313,n1327);
and (n1452,n1450,n1453);
or (n1453,n1454,n1459,n1488);
and (n1454,n1455,n1457);
not (n1455,n1456);
nand (n1456,n681,n1350);
xor (n1457,n1458,n1347);
xor (n1458,n1331,n1345);
and (n1459,n1457,n1460);
or (n1460,n1461,n1466,n1487);
and (n1461,n1462,n1464);
not (n1462,n1463);
nand (n1463,n681,n1368);
xor (n1464,n1465,n1365);
xor (n1465,n1349,n1363);
and (n1466,n1464,n1467);
or (n1467,n1468,n1473,n1486);
and (n1468,n1469,n1471);
not (n1469,n1470);
nand (n1470,n681,n1386);
xor (n1471,n1472,n1383);
xor (n1472,n1367,n1381);
and (n1473,n1471,n1474);
or (n1474,n1475,n1480,n1485);
and (n1475,n1476,n1478);
not (n1476,n1477);
nand (n1477,n681,n1404);
xor (n1478,n1479,n1401);
xor (n1479,n1385,n1399);
and (n1480,n1478,n1481);
and (n1481,n1482,n1483);
and (n1482,n681,n1421);
xor (n1483,n1484,n1419);
xor (n1484,n1403,n1417);
and (n1485,n1476,n1481);
and (n1486,n1469,n1474);
and (n1487,n1462,n1467);
and (n1488,n1455,n1460);
and (n1489,n1448,n1453);
and (n1490,n1442,n1446);
and (n1491,n1295,n1440);
or (n1492,n1493,n1571,n1656);
and (n1493,n1494,n1499);
xor (n1494,n1495,n1498);
wire s0n1495,s1n1495,notn1495;
or (n1495,s0n1495,s1n1495);
not(notn1495,n929);
and (s0n1495,notn1495,1'b0);
and (s1n1495,n929,n1496);
xor (n1496,n1497,n1440);
xor (n1497,n1295,n1309);
wire s0n1498,s1n1498,notn1498;
or (n1498,s0n1498,s1n1498);
not(notn1498,n1078);
and (s0n1498,notn1498,1'b0);
and (s1n1498,n1078,n1293);
and (n1499,n1500,n1501);
wire s0n1500,s1n1500,notn1500;
or (n1500,s0n1500,s1n1500);
not(notn1500,n1085);
and (s0n1500,notn1500,1'b0);
and (s1n1500,n1085,n1293);
or (n1501,n1502,n1505,n1570);
and (n1502,n1503,n1504);
wire s0n1503,s1n1503,notn1503;
or (n1503,s0n1503,s1n1503);
not(notn1503,n1085);
and (s0n1503,notn1503,1'b0);
and (s1n1503,n1085,n1496);
wire s0n1504,s1n1504,notn1504;
or (n1504,s0n1504,s1n1504);
not(notn1504,n930);
and (s0n1504,notn1504,1'b0);
and (s1n1504,n930,n1293);
and (n1505,n1504,n1506);
or (n1506,n1507,n1512,n1569);
and (n1507,n1508,n1511);
wire s0n1508,s1n1508,notn1508;
or (n1508,s0n1508,s1n1508);
not(notn1508,n1085);
and (s0n1508,notn1508,1'b0);
and (s1n1508,n1085,n1509);
xor (n1509,n1510,n1446);
xor (n1510,n1442,n1444);
wire s0n1511,s1n1511,notn1511;
or (n1511,s0n1511,s1n1511);
not(notn1511,n930);
and (s0n1511,notn1511,1'b0);
and (s1n1511,n930,n1496);
and (n1512,n1511,n1513);
or (n1513,n1514,n1519,n1568);
and (n1514,n1515,n1518);
wire s0n1515,s1n1515,notn1515;
or (n1515,s0n1515,s1n1515);
not(notn1515,n1085);
and (s0n1515,notn1515,1'b0);
and (s1n1515,n1085,n1516);
xor (n1516,n1517,n1453);
xor (n1517,n1448,n1450);
wire s0n1518,s1n1518,notn1518;
or (n1518,s0n1518,s1n1518);
not(notn1518,n930);
and (s0n1518,notn1518,1'b0);
and (s1n1518,n930,n1509);
and (n1519,n1518,n1520);
or (n1520,n1521,n1526,n1567);
and (n1521,n1522,n1525);
wire s0n1522,s1n1522,notn1522;
or (n1522,s0n1522,s1n1522);
not(notn1522,n1085);
and (s0n1522,notn1522,1'b0);
and (s1n1522,n1085,n1523);
xor (n1523,n1524,n1460);
xor (n1524,n1455,n1457);
wire s0n1525,s1n1525,notn1525;
or (n1525,s0n1525,s1n1525);
not(notn1525,n930);
and (s0n1525,notn1525,1'b0);
and (s1n1525,n930,n1516);
and (n1526,n1525,n1527);
or (n1527,n1528,n1533,n1566);
and (n1528,n1529,n1532);
wire s0n1529,s1n1529,notn1529;
or (n1529,s0n1529,s1n1529);
not(notn1529,n1085);
and (s0n1529,notn1529,1'b0);
and (s1n1529,n1085,n1530);
xor (n1530,n1531,n1467);
xor (n1531,n1462,n1464);
wire s0n1532,s1n1532,notn1532;
or (n1532,s0n1532,s1n1532);
not(notn1532,n930);
and (s0n1532,notn1532,1'b0);
and (s1n1532,n930,n1523);
and (n1533,n1532,n1534);
or (n1534,n1535,n1540,n1565);
and (n1535,n1536,n1539);
wire s0n1536,s1n1536,notn1536;
or (n1536,s0n1536,s1n1536);
not(notn1536,n1085);
and (s0n1536,notn1536,1'b0);
and (s1n1536,n1085,n1537);
xor (n1537,n1538,n1474);
xor (n1538,n1469,n1471);
wire s0n1539,s1n1539,notn1539;
or (n1539,s0n1539,s1n1539);
not(notn1539,n930);
and (s0n1539,notn1539,1'b0);
and (s1n1539,n930,n1530);
and (n1540,n1539,n1541);
or (n1541,n1542,n1547,n1564);
and (n1542,n1543,n1546);
wire s0n1543,s1n1543,notn1543;
or (n1543,s0n1543,s1n1543);
not(notn1543,n1085);
and (s0n1543,notn1543,1'b0);
and (s1n1543,n1085,n1544);
xor (n1544,n1545,n1481);
xor (n1545,n1476,n1478);
wire s0n1546,s1n1546,notn1546;
or (n1546,s0n1546,s1n1546);
not(notn1546,n930);
and (s0n1546,notn1546,1'b0);
and (s1n1546,n930,n1537);
and (n1547,n1546,n1548);
or (n1548,n1549,n1553,n1555);
and (n1549,n1550,n1552);
wire s0n1550,s1n1550,notn1550;
or (n1550,s0n1550,s1n1550);
not(notn1550,n1085);
and (s0n1550,notn1550,1'b0);
and (s1n1550,n1085,n1551);
xor (n1551,n1482,n1483);
wire s0n1552,s1n1552,notn1552;
or (n1552,s0n1552,s1n1552);
not(notn1552,n930);
and (s0n1552,notn1552,1'b0);
and (s1n1552,n930,n1544);
and (n1553,n1552,n1554);
or (n1554,n1555,n1559,n1560);
and (n1555,n1556,n1558);
wire s0n1556,s1n1556,notn1556;
or (n1556,s0n1556,s1n1556);
not(notn1556,n1085);
and (s0n1556,notn1556,1'b0);
and (s1n1556,n1085,n1557);
xor (n1557,n1420,n1434);
wire s0n1558,s1n1558,notn1558;
or (n1558,s0n1558,s1n1558);
not(notn1558,n930);
and (s0n1558,notn1558,1'b0);
and (s1n1558,n930,n1551);
and (n1559,n1558,n1560);
and (n1560,n1561,n1563);
wire s0n1561,s1n1561,notn1561;
or (n1561,s0n1561,s1n1561);
not(notn1561,n1085);
and (s0n1561,notn1561,1'b0);
and (s1n1561,n1085,n1562);
wire s0n1562,s1n1562,notn1562;
or (n1562,s0n1562,s1n1562);
not(notn1562,n579);
and (s0n1562,notn1562,1'b0);
and (s1n1562,n579,n1421);
wire s0n1563,s1n1563,notn1563;
or (n1563,s0n1563,s1n1563);
not(notn1563,n930);
and (s0n1563,notn1563,1'b0);
and (s1n1563,n930,n1557);
and (n1564,n1543,n1548);
and (n1565,n1536,n1541);
and (n1566,n1529,n1534);
and (n1567,n1522,n1527);
and (n1568,n1515,n1520);
and (n1569,n1508,n1513);
and (n1570,n1503,n1506);
and (n1571,n1499,n1572);
or (n1572,n1573,n1578,n1655);
and (n1573,n1574,n1577);
xor (n1574,n1575,n1576);
wire s0n1575,s1n1575,notn1575;
or (n1575,s0n1575,s1n1575);
not(notn1575,n929);
and (s0n1575,notn1575,1'b0);
and (s1n1575,n929,n1509);
wire s0n1576,s1n1576,notn1576;
or (n1576,s0n1576,s1n1576);
not(notn1576,n1078);
and (s0n1576,notn1576,1'b0);
and (s1n1576,n1078,n1496);
xor (n1577,n1500,n1501);
and (n1578,n1577,n1579);
or (n1579,n1580,n1586,n1654);
and (n1580,n1581,n1584);
xor (n1581,n1582,n1583);
wire s0n1582,s1n1582,notn1582;
or (n1582,s0n1582,s1n1582);
not(notn1582,n929);
and (s0n1582,notn1582,1'b0);
and (s1n1582,n929,n1516);
wire s0n1583,s1n1583,notn1583;
or (n1583,s0n1583,s1n1583);
not(notn1583,n1078);
and (s0n1583,notn1583,1'b0);
and (s1n1583,n1078,n1509);
xor (n1584,n1585,n1506);
xor (n1585,n1503,n1504);
and (n1586,n1584,n1587);
or (n1587,n1588,n1594,n1653);
and (n1588,n1589,n1592);
xor (n1589,n1590,n1591);
wire s0n1590,s1n1590,notn1590;
or (n1590,s0n1590,s1n1590);
not(notn1590,n929);
and (s0n1590,notn1590,1'b0);
and (s1n1590,n929,n1523);
wire s0n1591,s1n1591,notn1591;
or (n1591,s0n1591,s1n1591);
not(notn1591,n1078);
and (s0n1591,notn1591,1'b0);
and (s1n1591,n1078,n1516);
xor (n1592,n1593,n1513);
xor (n1593,n1508,n1511);
and (n1594,n1592,n1595);
or (n1595,n1596,n1602,n1652);
and (n1596,n1597,n1600);
xor (n1597,n1598,n1599);
wire s0n1598,s1n1598,notn1598;
or (n1598,s0n1598,s1n1598);
not(notn1598,n929);
and (s0n1598,notn1598,1'b0);
and (s1n1598,n929,n1530);
wire s0n1599,s1n1599,notn1599;
or (n1599,s0n1599,s1n1599);
not(notn1599,n1078);
and (s0n1599,notn1599,1'b0);
and (s1n1599,n1078,n1523);
xor (n1600,n1601,n1520);
xor (n1601,n1515,n1518);
and (n1602,n1600,n1603);
or (n1603,n1604,n1610,n1651);
and (n1604,n1605,n1608);
xor (n1605,n1606,n1607);
wire s0n1606,s1n1606,notn1606;
or (n1606,s0n1606,s1n1606);
not(notn1606,n929);
and (s0n1606,notn1606,1'b0);
and (s1n1606,n929,n1537);
wire s0n1607,s1n1607,notn1607;
or (n1607,s0n1607,s1n1607);
not(notn1607,n1078);
and (s0n1607,notn1607,1'b0);
and (s1n1607,n1078,n1530);
xor (n1608,n1609,n1527);
xor (n1609,n1522,n1525);
and (n1610,n1608,n1611);
or (n1611,n1612,n1618,n1650);
and (n1612,n1613,n1616);
xor (n1613,n1614,n1615);
wire s0n1614,s1n1614,notn1614;
or (n1614,s0n1614,s1n1614);
not(notn1614,n929);
and (s0n1614,notn1614,1'b0);
and (s1n1614,n929,n1544);
wire s0n1615,s1n1615,notn1615;
or (n1615,s0n1615,s1n1615);
not(notn1615,n1078);
and (s0n1615,notn1615,1'b0);
and (s1n1615,n1078,n1537);
xor (n1616,n1617,n1534);
xor (n1617,n1529,n1532);
and (n1618,n1616,n1619);
or (n1619,n1620,n1626,n1649);
and (n1620,n1621,n1624);
xor (n1621,n1622,n1623);
wire s0n1622,s1n1622,notn1622;
or (n1622,s0n1622,s1n1622);
not(notn1622,n929);
and (s0n1622,notn1622,1'b0);
and (s1n1622,n929,n1551);
wire s0n1623,s1n1623,notn1623;
or (n1623,s0n1623,s1n1623);
not(notn1623,n1078);
and (s0n1623,notn1623,1'b0);
and (s1n1623,n1078,n1544);
xor (n1624,n1625,n1541);
xor (n1625,n1536,n1539);
and (n1626,n1624,n1627);
or (n1627,n1628,n1634,n1648);
and (n1628,n1629,n1632);
xor (n1629,n1630,n1631);
wire s0n1630,s1n1630,notn1630;
or (n1630,s0n1630,s1n1630);
not(notn1630,n929);
and (s0n1630,notn1630,1'b0);
and (s1n1630,n929,n1557);
wire s0n1631,s1n1631,notn1631;
or (n1631,s0n1631,s1n1631);
not(notn1631,n1078);
and (s0n1631,notn1631,1'b0);
and (s1n1631,n1078,n1551);
xor (n1632,n1633,n1548);
xor (n1633,n1543,n1546);
and (n1634,n1632,n1635);
or (n1635,n1636,n1642,n1647);
and (n1636,n1637,n1640);
xor (n1637,n1638,n1639);
wire s0n1638,s1n1638,notn1638;
or (n1638,s0n1638,s1n1638);
not(notn1638,n929);
and (s0n1638,notn1638,1'b0);
and (s1n1638,n929,n1562);
wire s0n1639,s1n1639,notn1639;
or (n1639,s0n1639,s1n1639);
not(notn1639,n1078);
and (s0n1639,notn1639,1'b0);
and (s1n1639,n1078,n1557);
xor (n1640,n1641,n1554);
xor (n1641,n1550,n1552);
and (n1642,n1640,n1643);
and (n1643,n1644,n1645);
wire s0n1644,s1n1644,notn1644;
or (n1644,s0n1644,s1n1644);
not(notn1644,n1078);
and (s0n1644,notn1644,1'b0);
and (s1n1644,n1078,n1562);
xor (n1645,n1646,n1560);
xor (n1646,n1556,n1558);
and (n1647,n1637,n1643);
and (n1648,n1629,n1635);
and (n1649,n1621,n1627);
and (n1650,n1613,n1619);
and (n1651,n1605,n1611);
and (n1652,n1597,n1603);
and (n1653,n1589,n1595);
and (n1654,n1581,n1587);
and (n1655,n1574,n1579);
and (n1656,n1494,n1572);
or (n1657,n1658,n1663,n1751);
and (n1658,n1659,n1661);
xor (n1659,n1660,n1206);
xor (n1660,n1073,n1083);
xor (n1661,n1662,n1572);
xor (n1662,n1494,n1499);
and (n1663,n1661,n1664);
or (n1664,n1665,n1670,n1750);
and (n1665,n1666,n1668);
xor (n1666,n1667,n1213);
xor (n1667,n1208,n1211);
xor (n1668,n1669,n1579);
xor (n1669,n1574,n1577);
and (n1670,n1668,n1671);
or (n1671,n1672,n1677,n1749);
and (n1672,n1673,n1675);
xor (n1673,n1674,n1221);
xor (n1674,n1215,n1218);
xor (n1675,n1676,n1587);
xor (n1676,n1581,n1584);
and (n1677,n1675,n1678);
or (n1678,n1679,n1684,n1748);
and (n1679,n1680,n1682);
xor (n1680,n1681,n1229);
xor (n1681,n1223,n1226);
xor (n1682,n1683,n1595);
xor (n1683,n1589,n1592);
and (n1684,n1682,n1685);
or (n1685,n1686,n1691,n1747);
and (n1686,n1687,n1689);
xor (n1687,n1688,n1237);
xor (n1688,n1231,n1234);
xor (n1689,n1690,n1603);
xor (n1690,n1597,n1600);
and (n1691,n1689,n1692);
or (n1692,n1693,n1698,n1746);
and (n1693,n1694,n1696);
xor (n1694,n1695,n1245);
xor (n1695,n1239,n1242);
xor (n1696,n1697,n1611);
xor (n1697,n1605,n1608);
and (n1698,n1696,n1699);
or (n1699,n1700,n1705,n1745);
and (n1700,n1701,n1703);
xor (n1701,n1702,n1253);
xor (n1702,n1247,n1250);
xor (n1703,n1704,n1619);
xor (n1704,n1613,n1616);
and (n1705,n1703,n1706);
or (n1706,n1707,n1712,n1744);
and (n1707,n1708,n1710);
xor (n1708,n1709,n1261);
xor (n1709,n1255,n1258);
xor (n1710,n1711,n1627);
xor (n1711,n1621,n1624);
and (n1712,n1710,n1713);
or (n1713,n1714,n1719,n1743);
and (n1714,n1715,n1717);
xor (n1715,n1716,n1269);
xor (n1716,n1263,n1266);
xor (n1717,n1718,n1635);
xor (n1718,n1629,n1632);
and (n1719,n1717,n1720);
or (n1720,n1721,n1726,n1742);
and (n1721,n1722,n1724);
xor (n1722,n1723,n1277);
xor (n1723,n1271,n1274);
xor (n1724,n1725,n1643);
xor (n1725,n1637,n1640);
and (n1726,n1724,n1727);
or (n1727,n1728,n1731,n1741);
and (n1728,n1729,n1730);
xor (n1729,n1278,n1279);
xor (n1730,n1644,n1645);
and (n1731,n1730,n1732);
or (n1732,n1733,n1736,n1740);
and (n1733,n1734,n1735);
xor (n1734,n1195,n1197);
xor (n1735,n1561,n1563);
and (n1736,n1735,n1737);
and (n1737,n1738,n1739);
wire s0n1738,s1n1738,notn1738;
or (n1738,s0n1738,s1n1738);
not(notn1738,n930);
and (s0n1738,notn1738,1'b0);
and (s1n1738,n930,n1196);
wire s0n1739,s1n1739,notn1739;
or (n1739,s0n1739,s1n1739);
not(notn1739,n930);
and (s0n1739,notn1739,1'b0);
and (s1n1739,n930,n1562);
and (n1740,n1734,n1737);
and (n1741,n1729,n1732);
and (n1742,n1722,n1727);
and (n1743,n1715,n1720);
and (n1744,n1708,n1713);
and (n1745,n1701,n1706);
and (n1746,n1694,n1699);
and (n1747,n1687,n1692);
and (n1748,n1680,n1685);
and (n1749,n1673,n1678);
and (n1750,n1666,n1671);
and (n1751,n1659,n1664);
xor (n1752,n1753,n2453);
xor (n1753,n1754,n2108);
or (n1754,n1755,n2040,n2107);
and (n1755,n1756,n1966);
wire s0n1756,s1n1756,notn1756;
or (n1756,s0n1756,s1n1756);
not(notn1756,n1024);
and (s0n1756,notn1756,1'b0);
and (s1n1756,n1024,n1757);
xor (n1757,n1758,n1772);
wire s0n1758,s1n1758,notn1758;
or (n1758,s0n1758,s1n1758);
not(notn1758,n578);
and (s0n1758,notn1758,1'b0);
and (s1n1758,n578,n1759);
nand (n1759,n1760,n1763);
or (n1760,n1761,n14);
not (n1761,n1762);
nand (n1763,n564,n1764);
or (n1764,1'b0,n1765,n1767,n1769,n1771);
and (n1765,n1766,n555);
and (n1767,n1768,n570);
and (n1769,n1770,n574);
and (n1771,n1762,n576);
or (n1772,n1773,n1907,n1965);
and (n1773,n1774,n1790);
xor (n1774,n1775,n1789);
wire s0n1775,s1n1775,notn1775;
or (n1775,s0n1775,s1n1775);
not(notn1775,n578);
and (s0n1775,notn1775,1'b0);
and (s1n1775,n578,n1776);
nand (n1776,n1777,n1780);
or (n1777,n1778,n14);
not (n1778,n1779);
nand (n1780,n564,n1781);
or (n1781,1'b0,n1782,n1784,n1786,n1788);
and (n1782,n1783,n555);
and (n1784,n1785,n570);
and (n1786,n1787,n574);
and (n1788,n1779,n576);
wire s0n1789,s1n1789,notn1789;
or (n1789,s0n1789,s1n1789);
not(notn1789,n746);
and (s0n1789,notn1789,1'b0);
and (s1n1789,n746,n1759);
and (n1790,n1791,n1792);
wire s0n1791,s1n1791,notn1791;
or (n1791,s0n1791,s1n1791);
not(notn1791,n753);
and (s0n1791,notn1791,1'b0);
and (s1n1791,n753,n1759);
or (n1792,n1793,n1796,n1906);
and (n1793,n1794,n1795);
wire s0n1794,s1n1794,notn1794;
or (n1794,s0n1794,s1n1794);
not(notn1794,n753);
and (s0n1794,notn1794,1'b0);
and (s1n1794,n753,n1776);
wire s0n1795,s1n1795,notn1795;
or (n1795,s0n1795,s1n1795);
not(notn1795,n579);
and (s0n1795,notn1795,1'b0);
and (s1n1795,n579,n1759);
and (n1796,n1795,n1797);
or (n1797,n1798,n1814,n1905);
and (n1798,n1799,n1813);
wire s0n1799,s1n1799,notn1799;
or (n1799,s0n1799,s1n1799);
not(notn1799,n753);
and (s0n1799,notn1799,1'b0);
and (s1n1799,n753,n1800);
nand (n1800,n1801,n1804);
or (n1801,n1802,n14);
not (n1802,n1803);
nand (n1804,n564,n1805);
or (n1805,1'b0,n1806,n1808,n1810,n1812);
and (n1806,n1807,n555);
and (n1808,n1809,n570);
and (n1810,n1811,n574);
and (n1812,n1803,n576);
wire s0n1813,s1n1813,notn1813;
or (n1813,s0n1813,s1n1813);
not(notn1813,n579);
and (s0n1813,notn1813,1'b0);
and (s1n1813,n579,n1776);
and (n1814,n1813,n1815);
or (n1815,n1816,n1832,n1904);
and (n1816,n1817,n1831);
wire s0n1817,s1n1817,notn1817;
or (n1817,s0n1817,s1n1817);
not(notn1817,n753);
and (s0n1817,notn1817,1'b0);
and (s1n1817,n753,n1818);
nand (n1818,n1819,n1822);
or (n1819,n1820,n14);
not (n1820,n1821);
nand (n1822,n564,n1823);
or (n1823,1'b0,n1824,n1826,n1828,n1830);
and (n1824,n1825,n555);
and (n1826,n1827,n570);
and (n1828,n1829,n574);
and (n1830,n1821,n576);
wire s0n1831,s1n1831,notn1831;
or (n1831,s0n1831,s1n1831);
not(notn1831,n579);
and (s0n1831,notn1831,1'b0);
and (s1n1831,n579,n1800);
and (n1832,n1831,n1833);
or (n1833,n1834,n1850,n1903);
and (n1834,n1835,n1849);
wire s0n1835,s1n1835,notn1835;
or (n1835,s0n1835,s1n1835);
not(notn1835,n753);
and (s0n1835,notn1835,1'b0);
and (s1n1835,n753,n1836);
nand (n1836,n1837,n1840);
or (n1837,n1838,n14);
not (n1838,n1839);
nand (n1840,n564,n1841);
or (n1841,1'b0,n1842,n1844,n1846,n1848);
and (n1842,n1843,n555);
and (n1844,n1845,n570);
and (n1846,n1847,n574);
and (n1848,n1839,n576);
wire s0n1849,s1n1849,notn1849;
or (n1849,s0n1849,s1n1849);
not(notn1849,n579);
and (s0n1849,notn1849,1'b0);
and (s1n1849,n579,n1818);
and (n1850,n1849,n1851);
or (n1851,n1852,n1868,n1870);
and (n1852,n1853,n1867);
wire s0n1853,s1n1853,notn1853;
or (n1853,s0n1853,s1n1853);
not(notn1853,n753);
and (s0n1853,notn1853,1'b0);
and (s1n1853,n753,n1854);
nand (n1854,n1855,n1866);
or (n1855,n1856,n863);
not (n1856,n1857);
or (n1857,1'b0,n1858,n1860,n1862,n1864);
and (n1858,n1859,n555);
and (n1860,n1861,n570);
and (n1862,n1863,n574);
and (n1864,n1865,n576);
nand (n1866,n15,n1865);
wire s0n1867,s1n1867,notn1867;
or (n1867,s0n1867,s1n1867);
not(notn1867,n579);
and (s0n1867,notn1867,1'b0);
and (s1n1867,n579,n1836);
and (n1868,n1867,n1869);
or (n1869,n1870,n1886,n1887);
and (n1870,n1871,n1885);
wire s0n1871,s1n1871,notn1871;
or (n1871,s0n1871,s1n1871);
not(notn1871,n753);
and (s0n1871,notn1871,1'b0);
and (s1n1871,n753,n1872);
nand (n1872,n1873,n1884);
or (n1873,n1874,n863);
not (n1874,n1875);
or (n1875,1'b0,n1876,n1878,n1880,n1882);
and (n1876,n1877,n555);
and (n1878,n1879,n570);
and (n1880,n1881,n574);
and (n1882,n1883,n576);
nand (n1884,n15,n1883);
wire s0n1885,s1n1885,notn1885;
or (n1885,s0n1885,s1n1885);
not(notn1885,n579);
and (s0n1885,notn1885,1'b0);
and (s1n1885,n579,n1854);
and (n1886,n1885,n1887);
and (n1887,n1888,n1902);
wire s0n1888,s1n1888,notn1888;
or (n1888,s0n1888,s1n1888);
not(notn1888,n753);
and (s0n1888,notn1888,1'b0);
and (s1n1888,n753,n1889);
nand (n1889,n1890,n1893);
or (n1890,n1891,n14);
not (n1891,n1892);
nand (n1893,n564,n1894);
or (n1894,1'b0,n1895,n1897,n1899,n1901);
and (n1895,n1896,n555);
and (n1897,n1898,n570);
and (n1899,n1900,n574);
and (n1901,n1892,n576);
wire s0n1902,s1n1902,notn1902;
or (n1902,s0n1902,s1n1902);
not(notn1902,n579);
and (s0n1902,notn1902,1'b0);
and (s1n1902,n579,n1872);
and (n1903,n1835,n1851);
and (n1904,n1817,n1833);
and (n1905,n1799,n1815);
and (n1906,n1794,n1797);
and (n1907,n1790,n1908);
or (n1908,n1909,n1914,n1964);
and (n1909,n1910,n1913);
xor (n1910,n1911,n1912);
wire s0n1911,s1n1911,notn1911;
or (n1911,s0n1911,s1n1911);
not(notn1911,n578);
and (s0n1911,notn1911,1'b0);
and (s1n1911,n578,n1800);
wire s0n1912,s1n1912,notn1912;
or (n1912,s0n1912,s1n1912);
not(notn1912,n746);
and (s0n1912,notn1912,1'b0);
and (s1n1912,n746,n1776);
xor (n1913,n1791,n1792);
and (n1914,n1913,n1915);
or (n1915,n1916,n1922,n1963);
and (n1916,n1917,n1920);
xor (n1917,n1918,n1919);
wire s0n1918,s1n1918,notn1918;
or (n1918,s0n1918,s1n1918);
not(notn1918,n578);
and (s0n1918,notn1918,1'b0);
and (s1n1918,n578,n1818);
wire s0n1919,s1n1919,notn1919;
or (n1919,s0n1919,s1n1919);
not(notn1919,n746);
and (s0n1919,notn1919,1'b0);
and (s1n1919,n746,n1800);
xor (n1920,n1921,n1797);
xor (n1921,n1794,n1795);
and (n1922,n1920,n1923);
or (n1923,n1924,n1930,n1962);
and (n1924,n1925,n1928);
xor (n1925,n1926,n1927);
wire s0n1926,s1n1926,notn1926;
or (n1926,s0n1926,s1n1926);
not(notn1926,n578);
and (s0n1926,notn1926,1'b0);
and (s1n1926,n578,n1836);
wire s0n1927,s1n1927,notn1927;
or (n1927,s0n1927,s1n1927);
not(notn1927,n746);
and (s0n1927,notn1927,1'b0);
and (s1n1927,n746,n1818);
xor (n1928,n1929,n1815);
xor (n1929,n1799,n1813);
and (n1930,n1928,n1931);
or (n1931,n1932,n1938,n1961);
and (n1932,n1933,n1936);
xor (n1933,n1934,n1935);
wire s0n1934,s1n1934,notn1934;
or (n1934,s0n1934,s1n1934);
not(notn1934,n578);
and (s0n1934,notn1934,1'b0);
and (s1n1934,n578,n1854);
wire s0n1935,s1n1935,notn1935;
or (n1935,s0n1935,s1n1935);
not(notn1935,n746);
and (s0n1935,notn1935,1'b0);
and (s1n1935,n746,n1836);
xor (n1936,n1937,n1833);
xor (n1937,n1817,n1831);
and (n1938,n1936,n1939);
or (n1939,n1940,n1946,n1960);
and (n1940,n1941,n1944);
xor (n1941,n1942,n1943);
wire s0n1942,s1n1942,notn1942;
or (n1942,s0n1942,s1n1942);
not(notn1942,n578);
and (s0n1942,notn1942,1'b0);
and (s1n1942,n578,n1872);
wire s0n1943,s1n1943,notn1943;
or (n1943,s0n1943,s1n1943);
not(notn1943,n746);
and (s0n1943,notn1943,1'b0);
and (s1n1943,n746,n1854);
xor (n1944,n1945,n1851);
xor (n1945,n1835,n1849);
and (n1946,n1944,n1947);
or (n1947,n1948,n1954,n1959);
and (n1948,n1949,n1952);
xor (n1949,n1950,n1951);
wire s0n1950,s1n1950,notn1950;
or (n1950,s0n1950,s1n1950);
not(notn1950,n578);
and (s0n1950,notn1950,1'b0);
and (s1n1950,n578,n1889);
wire s0n1951,s1n1951,notn1951;
or (n1951,s0n1951,s1n1951);
not(notn1951,n746);
and (s0n1951,notn1951,1'b0);
and (s1n1951,n746,n1872);
xor (n1952,n1953,n1869);
xor (n1953,n1853,n1867);
and (n1954,n1952,n1955);
and (n1955,n1956,n1957);
wire s0n1956,s1n1956,notn1956;
or (n1956,s0n1956,s1n1956);
not(notn1956,n746);
and (s0n1956,notn1956,1'b0);
and (s1n1956,n746,n1889);
xor (n1957,n1958,n1887);
xor (n1958,n1871,n1885);
and (n1959,n1949,n1955);
and (n1960,n1941,n1947);
and (n1961,n1933,n1939);
and (n1962,n1925,n1931);
and (n1963,n1917,n1923);
and (n1964,n1910,n1915);
and (n1965,n1774,n1908);
and (n1966,n1967,n1968);
wire s0n1967,s1n1967,notn1967;
or (n1967,s0n1967,s1n1967);
not(notn1967,n977);
and (s0n1967,notn1967,1'b0);
and (s1n1967,n977,n1757);
or (n1968,n1969,n1974,n2039);
and (n1969,n1970,n1973);
wire s0n1970,s1n1970,notn1970;
or (n1970,s0n1970,s1n1970);
not(notn1970,n977);
and (s0n1970,notn1970,1'b0);
and (s1n1970,n977,n1971);
xor (n1971,n1972,n1908);
xor (n1972,n1774,n1790);
wire s0n1973,s1n1973,notn1973;
or (n1973,s0n1973,s1n1973);
not(notn1973,n930);
and (s0n1973,notn1973,1'b0);
and (s1n1973,n930,n1757);
and (n1974,n1973,n1975);
or (n1975,n1976,n1981,n2038);
and (n1976,n1977,n1980);
wire s0n1977,s1n1977,notn1977;
or (n1977,s0n1977,s1n1977);
not(notn1977,n977);
and (s0n1977,notn1977,1'b0);
and (s1n1977,n977,n1978);
xor (n1978,n1979,n1915);
xor (n1979,n1910,n1913);
wire s0n1980,s1n1980,notn1980;
or (n1980,s0n1980,s1n1980);
not(notn1980,n930);
and (s0n1980,notn1980,1'b0);
and (s1n1980,n930,n1971);
and (n1981,n1980,n1982);
or (n1982,n1983,n1988,n2037);
and (n1983,n1984,n1987);
wire s0n1984,s1n1984,notn1984;
or (n1984,s0n1984,s1n1984);
not(notn1984,n977);
and (s0n1984,notn1984,1'b0);
and (s1n1984,n977,n1985);
xor (n1985,n1986,n1923);
xor (n1986,n1917,n1920);
wire s0n1987,s1n1987,notn1987;
or (n1987,s0n1987,s1n1987);
not(notn1987,n930);
and (s0n1987,notn1987,1'b0);
and (s1n1987,n930,n1978);
and (n1988,n1987,n1989);
or (n1989,n1990,n1995,n2036);
and (n1990,n1991,n1994);
wire s0n1991,s1n1991,notn1991;
or (n1991,s0n1991,s1n1991);
not(notn1991,n977);
and (s0n1991,notn1991,1'b0);
and (s1n1991,n977,n1992);
xor (n1992,n1993,n1931);
xor (n1993,n1925,n1928);
wire s0n1994,s1n1994,notn1994;
or (n1994,s0n1994,s1n1994);
not(notn1994,n930);
and (s0n1994,notn1994,1'b0);
and (s1n1994,n930,n1985);
and (n1995,n1994,n1996);
or (n1996,n1997,n2002,n2035);
and (n1997,n1998,n2001);
wire s0n1998,s1n1998,notn1998;
or (n1998,s0n1998,s1n1998);
not(notn1998,n977);
and (s0n1998,notn1998,1'b0);
and (s1n1998,n977,n1999);
xor (n1999,n2000,n1939);
xor (n2000,n1933,n1936);
wire s0n2001,s1n2001,notn2001;
or (n2001,s0n2001,s1n2001);
not(notn2001,n930);
and (s0n2001,notn2001,1'b0);
and (s1n2001,n930,n1992);
and (n2002,n2001,n2003);
or (n2003,n2004,n2009,n2034);
and (n2004,n2005,n2008);
wire s0n2005,s1n2005,notn2005;
or (n2005,s0n2005,s1n2005);
not(notn2005,n977);
and (s0n2005,notn2005,1'b0);
and (s1n2005,n977,n2006);
xor (n2006,n2007,n1947);
xor (n2007,n1941,n1944);
wire s0n2008,s1n2008,notn2008;
or (n2008,s0n2008,s1n2008);
not(notn2008,n930);
and (s0n2008,notn2008,1'b0);
and (s1n2008,n930,n1999);
and (n2009,n2008,n2010);
or (n2010,n2011,n2016,n2033);
and (n2011,n2012,n2015);
wire s0n2012,s1n2012,notn2012;
or (n2012,s0n2012,s1n2012);
not(notn2012,n977);
and (s0n2012,notn2012,1'b0);
and (s1n2012,n977,n2013);
xor (n2013,n2014,n1955);
xor (n2014,n1949,n1952);
wire s0n2015,s1n2015,notn2015;
or (n2015,s0n2015,s1n2015);
not(notn2015,n930);
and (s0n2015,notn2015,1'b0);
and (s1n2015,n930,n2006);
and (n2016,n2015,n2017);
or (n2017,n2018,n2022,n2024);
and (n2018,n2019,n2021);
wire s0n2019,s1n2019,notn2019;
or (n2019,s0n2019,s1n2019);
not(notn2019,n977);
and (s0n2019,notn2019,1'b0);
and (s1n2019,n977,n2020);
xor (n2020,n1956,n1957);
wire s0n2021,s1n2021,notn2021;
or (n2021,s0n2021,s1n2021);
not(notn2021,n930);
and (s0n2021,notn2021,1'b0);
and (s1n2021,n930,n2013);
and (n2022,n2021,n2023);
or (n2023,n2024,n2028,n2029);
and (n2024,n2025,n2027);
wire s0n2025,s1n2025,notn2025;
or (n2025,s0n2025,s1n2025);
not(notn2025,n977);
and (s0n2025,notn2025,1'b0);
and (s1n2025,n977,n2026);
xor (n2026,n1888,n1902);
wire s0n2027,s1n2027,notn2027;
or (n2027,s0n2027,s1n2027);
not(notn2027,n930);
and (s0n2027,notn2027,1'b0);
and (s1n2027,n930,n2020);
and (n2028,n2027,n2029);
and (n2029,n2030,n2032);
wire s0n2030,s1n2030,notn2030;
or (n2030,s0n2030,s1n2030);
not(notn2030,n977);
and (s0n2030,notn2030,1'b0);
and (s1n2030,n977,n2031);
wire s0n2031,s1n2031,notn2031;
or (n2031,s0n2031,s1n2031);
not(notn2031,n579);
and (s0n2031,notn2031,1'b0);
and (s1n2031,n579,n1889);
wire s0n2032,s1n2032,notn2032;
or (n2032,s0n2032,s1n2032);
not(notn2032,n930);
and (s0n2032,notn2032,1'b0);
and (s1n2032,n930,n2026);
and (n2033,n2012,n2017);
and (n2034,n2005,n2010);
and (n2035,n1998,n2003);
and (n2036,n1991,n1996);
and (n2037,n1984,n1989);
and (n2038,n1977,n1982);
and (n2039,n1970,n1975);
and (n2040,n1966,n2041);
or (n2041,n2042,n2045,n2106);
and (n2042,n2043,n2044);
wire s0n2043,s1n2043,notn2043;
or (n2043,s0n2043,s1n2043);
not(notn2043,n1024);
and (s0n2043,notn2043,1'b0);
and (s1n2043,n1024,n1971);
xor (n2044,n1967,n1968);
and (n2045,n2044,n2046);
or (n2046,n2047,n2051,n2105);
and (n2047,n2048,n2049);
wire s0n2048,s1n2048,notn2048;
or (n2048,s0n2048,s1n2048);
not(notn2048,n1024);
and (s0n2048,notn2048,1'b0);
and (s1n2048,n1024,n1978);
xor (n2049,n2050,n1975);
xor (n2050,n1970,n1973);
and (n2051,n2049,n2052);
or (n2052,n2053,n2057,n2104);
and (n2053,n2054,n2055);
wire s0n2054,s1n2054,notn2054;
or (n2054,s0n2054,s1n2054);
not(notn2054,n1024);
and (s0n2054,notn2054,1'b0);
and (s1n2054,n1024,n1985);
xor (n2055,n2056,n1982);
xor (n2056,n1977,n1980);
and (n2057,n2055,n2058);
or (n2058,n2059,n2063,n2103);
and (n2059,n2060,n2061);
wire s0n2060,s1n2060,notn2060;
or (n2060,s0n2060,s1n2060);
not(notn2060,n1024);
and (s0n2060,notn2060,1'b0);
and (s1n2060,n1024,n1992);
xor (n2061,n2062,n1989);
xor (n2062,n1984,n1987);
and (n2063,n2061,n2064);
or (n2064,n2065,n2069,n2102);
and (n2065,n2066,n2067);
wire s0n2066,s1n2066,notn2066;
or (n2066,s0n2066,s1n2066);
not(notn2066,n1024);
and (s0n2066,notn2066,1'b0);
and (s1n2066,n1024,n1999);
xor (n2067,n2068,n1996);
xor (n2068,n1991,n1994);
and (n2069,n2067,n2070);
or (n2070,n2071,n2075,n2101);
and (n2071,n2072,n2073);
wire s0n2072,s1n2072,notn2072;
or (n2072,s0n2072,s1n2072);
not(notn2072,n1024);
and (s0n2072,notn2072,1'b0);
and (s1n2072,n1024,n2006);
xor (n2073,n2074,n2003);
xor (n2074,n1998,n2001);
and (n2075,n2073,n2076);
or (n2076,n2077,n2081,n2100);
and (n2077,n2078,n2079);
wire s0n2078,s1n2078,notn2078;
or (n2078,s0n2078,s1n2078);
not(notn2078,n1024);
and (s0n2078,notn2078,1'b0);
and (s1n2078,n1024,n2013);
xor (n2079,n2080,n2010);
xor (n2080,n2005,n2008);
and (n2081,n2079,n2082);
or (n2082,n2083,n2087,n2099);
and (n2083,n2084,n2085);
wire s0n2084,s1n2084,notn2084;
or (n2084,s0n2084,s1n2084);
not(notn2084,n1024);
and (s0n2084,notn2084,1'b0);
and (s1n2084,n1024,n2020);
xor (n2085,n2086,n2017);
xor (n2086,n2012,n2015);
and (n2087,n2085,n2088);
or (n2088,n2089,n2093,n2098);
and (n2089,n2090,n2091);
wire s0n2090,s1n2090,notn2090;
or (n2090,s0n2090,s1n2090);
not(notn2090,n1024);
and (s0n2090,notn2090,1'b0);
and (s1n2090,n1024,n2026);
xor (n2091,n2092,n2023);
xor (n2092,n2019,n2021);
and (n2093,n2091,n2094);
and (n2094,n2095,n2096);
wire s0n2095,s1n2095,notn2095;
or (n2095,s0n2095,s1n2095);
not(notn2095,n1024);
and (s0n2095,notn2095,1'b0);
and (s1n2095,n1024,n2031);
xor (n2096,n2097,n2029);
xor (n2097,n2025,n2027);
and (n2098,n2090,n2094);
and (n2099,n2084,n2088);
and (n2100,n2078,n2082);
and (n2101,n2072,n2076);
and (n2102,n2066,n2070);
and (n2103,n2060,n2064);
and (n2104,n2054,n2058);
and (n2105,n2048,n2052);
and (n2106,n2043,n2046);
and (n2107,n1756,n2041);
or (n2108,n2109,n2385,n2452);
and (n2109,n2110,n2311);
wire s0n2110,s1n2110,notn2110;
or (n2110,s0n2110,s1n2110);
not(notn2110,n1024);
and (s0n2110,notn2110,1'b0);
and (s1n2110,n1024,n2111);
or (n2111,n2112,n2258,n2310);
and (n2112,n2113,n2128);
not (n2113,n2114);
nand (n2114,n681,n2115);
nand (n2115,n2116,n2127);
or (n2116,n2117,n863);
not (n2117,n2118);
or (n2118,1'b0,n2119,n2121,n2123,n2125);
and (n2119,n2120,n555);
and (n2121,n2122,n570);
and (n2123,n2124,n574);
and (n2125,n2126,n576);
nand (n2127,n15,n2126);
and (n2128,n2129,n2130);
wire s0n2129,s1n2129,notn2129;
or (n2129,s0n2129,s1n2129);
not(notn2129,n634);
and (s0n2129,notn2129,1'b0);
and (s1n2129,n634,n2115);
or (n2130,n2131,n2147,n2257);
and (n2131,n2132,n2146);
wire s0n2132,s1n2132,notn2132;
or (n2132,s0n2132,s1n2132);
not(notn2132,n634);
and (s0n2132,notn2132,1'b0);
and (s1n2132,n634,n2133);
nand (n2133,n2134,n2145);
or (n2134,n2135,n863);
not (n2135,n2136);
or (n2136,1'b0,n2137,n2139,n2141,n2143);
and (n2137,n2138,n555);
and (n2139,n2140,n570);
and (n2141,n2142,n574);
and (n2143,n2144,n576);
nand (n2145,n15,n2144);
wire s0n2146,s1n2146,notn2146;
or (n2146,s0n2146,s1n2146);
not(notn2146,n579);
and (s0n2146,notn2146,1'b0);
and (s1n2146,n579,n2115);
and (n2147,n2146,n2148);
or (n2148,n2149,n2165,n2256);
and (n2149,n2150,n2164);
wire s0n2150,s1n2150,notn2150;
or (n2150,s0n2150,s1n2150);
not(notn2150,n634);
and (s0n2150,notn2150,1'b0);
and (s1n2150,n634,n2151);
nand (n2151,n2152,n2163);
or (n2152,n2153,n863);
not (n2153,n2154);
or (n2154,1'b0,n2155,n2157,n2159,n2161);
and (n2155,n2156,n555);
and (n2157,n2158,n570);
and (n2159,n2160,n574);
and (n2161,n2162,n576);
nand (n2163,n15,n2162);
wire s0n2164,s1n2164,notn2164;
or (n2164,s0n2164,s1n2164);
not(notn2164,n579);
and (s0n2164,notn2164,1'b0);
and (s1n2164,n579,n2133);
and (n2165,n2164,n2166);
or (n2166,n2167,n2183,n2255);
and (n2167,n2168,n2182);
wire s0n2168,s1n2168,notn2168;
or (n2168,s0n2168,s1n2168);
not(notn2168,n634);
and (s0n2168,notn2168,1'b0);
and (s1n2168,n634,n2169);
nand (n2169,n2170,n2181);
or (n2170,n2171,n863);
not (n2171,n2172);
or (n2172,1'b0,n2173,n2175,n2177,n2179);
and (n2173,n2174,n555);
and (n2175,n2176,n570);
and (n2177,n2178,n574);
and (n2179,n2180,n576);
nand (n2181,n15,n2180);
wire s0n2182,s1n2182,notn2182;
or (n2182,s0n2182,s1n2182);
not(notn2182,n579);
and (s0n2182,notn2182,1'b0);
and (s1n2182,n579,n2151);
and (n2183,n2182,n2184);
or (n2184,n2185,n2201,n2254);
and (n2185,n2186,n2200);
wire s0n2186,s1n2186,notn2186;
or (n2186,s0n2186,s1n2186);
not(notn2186,n634);
and (s0n2186,notn2186,1'b0);
and (s1n2186,n634,n2187);
nand (n2187,n2188,n2199);
or (n2188,n2189,n863);
not (n2189,n2190);
or (n2190,1'b0,n2191,n2193,n2195,n2197);
and (n2191,n2192,n555);
and (n2193,n2194,n570);
and (n2195,n2196,n574);
and (n2197,n2198,n576);
nand (n2199,n15,n2198);
wire s0n2200,s1n2200,notn2200;
or (n2200,s0n2200,s1n2200);
not(notn2200,n579);
and (s0n2200,notn2200,1'b0);
and (s1n2200,n579,n2169);
and (n2201,n2200,n2202);
or (n2202,n2203,n2219,n2221);
and (n2203,n2204,n2218);
wire s0n2204,s1n2204,notn2204;
or (n2204,s0n2204,s1n2204);
not(notn2204,n634);
and (s0n2204,notn2204,1'b0);
and (s1n2204,n634,n2205);
nand (n2205,n2206,n2209);
or (n2206,n2207,n14);
not (n2207,n2208);
nand (n2209,n564,n2210);
or (n2210,1'b0,n2211,n2213,n2215,n2217);
and (n2211,n2212,n555);
and (n2213,n2214,n570);
and (n2215,n2216,n574);
and (n2217,n2208,n576);
wire s0n2218,s1n2218,notn2218;
or (n2218,s0n2218,s1n2218);
not(notn2218,n579);
and (s0n2218,notn2218,1'b0);
and (s1n2218,n579,n2187);
and (n2219,n2218,n2220);
or (n2220,n2221,n2237,n2238);
and (n2221,n2222,n2236);
wire s0n2222,s1n2222,notn2222;
or (n2222,s0n2222,s1n2222);
not(notn2222,n634);
and (s0n2222,notn2222,1'b0);
and (s1n2222,n634,n2223);
nand (n2223,n2224,n2235);
or (n2224,n2225,n863);
not (n2225,n2226);
or (n2226,1'b0,n2227,n2229,n2231,n2233);
and (n2227,n2228,n555);
and (n2229,n2230,n570);
and (n2231,n2232,n574);
and (n2233,n2234,n576);
nand (n2235,n15,n2234);
wire s0n2236,s1n2236,notn2236;
or (n2236,s0n2236,s1n2236);
not(notn2236,n579);
and (s0n2236,notn2236,1'b0);
and (s1n2236,n579,n2205);
and (n2237,n2236,n2238);
and (n2238,n2239,n2253);
wire s0n2239,s1n2239,notn2239;
or (n2239,s0n2239,s1n2239);
not(notn2239,n634);
and (s0n2239,notn2239,1'b0);
and (s1n2239,n634,n2240);
nand (n2240,n2241,n2252);
or (n2241,n2242,n863);
not (n2242,n2243);
or (n2243,1'b0,n2244,n2246,n2248,n2250);
and (n2244,n2245,n555);
and (n2246,n2247,n570);
and (n2248,n2249,n574);
and (n2250,n2251,n576);
nand (n2252,n15,n2251);
wire s0n2253,s1n2253,notn2253;
or (n2253,s0n2253,s1n2253);
not(notn2253,n579);
and (s0n2253,notn2253,1'b0);
and (s1n2253,n579,n2223);
and (n2254,n2186,n2202);
and (n2255,n2168,n2184);
and (n2256,n2150,n2166);
and (n2257,n2132,n2148);
and (n2258,n2128,n2259);
or (n2259,n2260,n2264,n2309);
and (n2260,n2261,n2263);
not (n2261,n2262);
nand (n2262,n681,n2133);
xor (n2263,n2129,n2130);
and (n2264,n2263,n2265);
or (n2265,n2266,n2271,n2308);
and (n2266,n2267,n2269);
not (n2267,n2268);
nand (n2268,n681,n2151);
xor (n2269,n2270,n2148);
xor (n2270,n2132,n2146);
and (n2271,n2269,n2272);
or (n2272,n2273,n2278,n2307);
and (n2273,n2274,n2276);
not (n2274,n2275);
nand (n2275,n681,n2169);
xor (n2276,n2277,n2166);
xor (n2277,n2150,n2164);
and (n2278,n2276,n2279);
or (n2279,n2280,n2284,n2306);
and (n2280,n2281,n2282);
and (n2281,n681,n2187);
xor (n2282,n2283,n2184);
xor (n2283,n2168,n2182);
and (n2284,n2282,n2285);
or (n2285,n2286,n2291,n2305);
and (n2286,n2287,n2289);
not (n2287,n2288);
nand (n2288,n681,n2205);
xor (n2289,n2290,n2202);
xor (n2290,n2186,n2200);
and (n2291,n2289,n2292);
or (n2292,n2293,n2298,n2304);
and (n2293,n2294,n2296);
not (n2294,n2295);
nand (n2295,n681,n2223);
xor (n2296,n2297,n2220);
xor (n2297,n2204,n2218);
and (n2298,n2296,n2299);
and (n2299,n2300,n2302);
not (n2300,n2301);
nand (n2301,n681,n2240);
xor (n2302,n2303,n2238);
xor (n2303,n2222,n2236);
and (n2304,n2294,n2299);
and (n2305,n2287,n2292);
and (n2306,n2281,n2285);
and (n2307,n2274,n2279);
and (n2308,n2267,n2272);
and (n2309,n2261,n2265);
and (n2310,n2113,n2259);
and (n2311,n2312,n2313);
wire s0n2312,s1n2312,notn2312;
or (n2312,s0n2312,s1n2312);
not(notn2312,n977);
and (s0n2312,notn2312,1'b0);
and (s1n2312,n977,n2111);
or (n2313,n2314,n2319,n2384);
and (n2314,n2315,n2318);
wire s0n2315,s1n2315,notn2315;
or (n2315,s0n2315,s1n2315);
not(notn2315,n977);
and (s0n2315,notn2315,1'b0);
and (s1n2315,n977,n2316);
xor (n2316,n2317,n2259);
xor (n2317,n2113,n2128);
wire s0n2318,s1n2318,notn2318;
or (n2318,s0n2318,s1n2318);
not(notn2318,n930);
and (s0n2318,notn2318,1'b0);
and (s1n2318,n930,n2111);
and (n2319,n2318,n2320);
or (n2320,n2321,n2326,n2383);
and (n2321,n2322,n2325);
wire s0n2322,s1n2322,notn2322;
or (n2322,s0n2322,s1n2322);
not(notn2322,n977);
and (s0n2322,notn2322,1'b0);
and (s1n2322,n977,n2323);
xor (n2323,n2324,n2265);
xor (n2324,n2261,n2263);
wire s0n2325,s1n2325,notn2325;
or (n2325,s0n2325,s1n2325);
not(notn2325,n930);
and (s0n2325,notn2325,1'b0);
and (s1n2325,n930,n2316);
and (n2326,n2325,n2327);
or (n2327,n2328,n2333,n2382);
and (n2328,n2329,n2332);
wire s0n2329,s1n2329,notn2329;
or (n2329,s0n2329,s1n2329);
not(notn2329,n977);
and (s0n2329,notn2329,1'b0);
and (s1n2329,n977,n2330);
xor (n2330,n2331,n2272);
xor (n2331,n2267,n2269);
wire s0n2332,s1n2332,notn2332;
or (n2332,s0n2332,s1n2332);
not(notn2332,n930);
and (s0n2332,notn2332,1'b0);
and (s1n2332,n930,n2323);
and (n2333,n2332,n2334);
or (n2334,n2335,n2340,n2381);
and (n2335,n2336,n2339);
wire s0n2336,s1n2336,notn2336;
or (n2336,s0n2336,s1n2336);
not(notn2336,n977);
and (s0n2336,notn2336,1'b0);
and (s1n2336,n977,n2337);
xor (n2337,n2338,n2279);
xor (n2338,n2274,n2276);
wire s0n2339,s1n2339,notn2339;
or (n2339,s0n2339,s1n2339);
not(notn2339,n930);
and (s0n2339,notn2339,1'b0);
and (s1n2339,n930,n2330);
and (n2340,n2339,n2341);
or (n2341,n2342,n2347,n2380);
and (n2342,n2343,n2346);
wire s0n2343,s1n2343,notn2343;
or (n2343,s0n2343,s1n2343);
not(notn2343,n977);
and (s0n2343,notn2343,1'b0);
and (s1n2343,n977,n2344);
xor (n2344,n2345,n2285);
xor (n2345,n2281,n2282);
wire s0n2346,s1n2346,notn2346;
or (n2346,s0n2346,s1n2346);
not(notn2346,n930);
and (s0n2346,notn2346,1'b0);
and (s1n2346,n930,n2337);
and (n2347,n2346,n2348);
or (n2348,n2349,n2354,n2379);
and (n2349,n2350,n2353);
wire s0n2350,s1n2350,notn2350;
or (n2350,s0n2350,s1n2350);
not(notn2350,n977);
and (s0n2350,notn2350,1'b0);
and (s1n2350,n977,n2351);
xor (n2351,n2352,n2292);
xor (n2352,n2287,n2289);
wire s0n2353,s1n2353,notn2353;
or (n2353,s0n2353,s1n2353);
not(notn2353,n930);
and (s0n2353,notn2353,1'b0);
and (s1n2353,n930,n2344);
and (n2354,n2353,n2355);
or (n2355,n2356,n2361,n2378);
and (n2356,n2357,n2360);
wire s0n2357,s1n2357,notn2357;
or (n2357,s0n2357,s1n2357);
not(notn2357,n977);
and (s0n2357,notn2357,1'b0);
and (s1n2357,n977,n2358);
xor (n2358,n2359,n2299);
xor (n2359,n2294,n2296);
wire s0n2360,s1n2360,notn2360;
or (n2360,s0n2360,s1n2360);
not(notn2360,n930);
and (s0n2360,notn2360,1'b0);
and (s1n2360,n930,n2351);
and (n2361,n2360,n2362);
or (n2362,n2363,n2367,n2369);
and (n2363,n2364,n2366);
wire s0n2364,s1n2364,notn2364;
or (n2364,s0n2364,s1n2364);
not(notn2364,n977);
and (s0n2364,notn2364,1'b0);
and (s1n2364,n977,n2365);
xor (n2365,n2300,n2302);
wire s0n2366,s1n2366,notn2366;
or (n2366,s0n2366,s1n2366);
not(notn2366,n930);
and (s0n2366,notn2366,1'b0);
and (s1n2366,n930,n2358);
and (n2367,n2366,n2368);
or (n2368,n2369,n2373,n2374);
and (n2369,n2370,n2372);
wire s0n2370,s1n2370,notn2370;
or (n2370,s0n2370,s1n2370);
not(notn2370,n977);
and (s0n2370,notn2370,1'b0);
and (s1n2370,n977,n2371);
xor (n2371,n2239,n2253);
wire s0n2372,s1n2372,notn2372;
or (n2372,s0n2372,s1n2372);
not(notn2372,n930);
and (s0n2372,notn2372,1'b0);
and (s1n2372,n930,n2365);
and (n2373,n2372,n2374);
and (n2374,n2375,n2377);
wire s0n2375,s1n2375,notn2375;
or (n2375,s0n2375,s1n2375);
not(notn2375,n977);
and (s0n2375,notn2375,1'b0);
and (s1n2375,n977,n2376);
wire s0n2376,s1n2376,notn2376;
or (n2376,s0n2376,s1n2376);
not(notn2376,n579);
and (s0n2376,notn2376,1'b0);
and (s1n2376,n579,n2240);
wire s0n2377,s1n2377,notn2377;
or (n2377,s0n2377,s1n2377);
not(notn2377,n930);
and (s0n2377,notn2377,1'b0);
and (s1n2377,n930,n2371);
and (n2378,n2357,n2362);
and (n2379,n2350,n2355);
and (n2380,n2343,n2348);
and (n2381,n2336,n2341);
and (n2382,n2329,n2334);
and (n2383,n2322,n2327);
and (n2384,n2315,n2320);
and (n2385,n2311,n2386);
or (n2386,n2387,n2390,n2451);
and (n2387,n2388,n2389);
wire s0n2388,s1n2388,notn2388;
or (n2388,s0n2388,s1n2388);
not(notn2388,n1024);
and (s0n2388,notn2388,1'b0);
and (s1n2388,n1024,n2316);
xor (n2389,n2312,n2313);
and (n2390,n2389,n2391);
or (n2391,n2392,n2396,n2450);
and (n2392,n2393,n2394);
wire s0n2393,s1n2393,notn2393;
or (n2393,s0n2393,s1n2393);
not(notn2393,n1024);
and (s0n2393,notn2393,1'b0);
and (s1n2393,n1024,n2323);
xor (n2394,n2395,n2320);
xor (n2395,n2315,n2318);
and (n2396,n2394,n2397);
or (n2397,n2398,n2402,n2449);
and (n2398,n2399,n2400);
wire s0n2399,s1n2399,notn2399;
or (n2399,s0n2399,s1n2399);
not(notn2399,n1024);
and (s0n2399,notn2399,1'b0);
and (s1n2399,n1024,n2330);
xor (n2400,n2401,n2327);
xor (n2401,n2322,n2325);
and (n2402,n2400,n2403);
or (n2403,n2404,n2408,n2448);
and (n2404,n2405,n2406);
wire s0n2405,s1n2405,notn2405;
or (n2405,s0n2405,s1n2405);
not(notn2405,n1024);
and (s0n2405,notn2405,1'b0);
and (s1n2405,n1024,n2337);
xor (n2406,n2407,n2334);
xor (n2407,n2329,n2332);
and (n2408,n2406,n2409);
or (n2409,n2410,n2414,n2447);
and (n2410,n2411,n2412);
wire s0n2411,s1n2411,notn2411;
or (n2411,s0n2411,s1n2411);
not(notn2411,n1024);
and (s0n2411,notn2411,1'b0);
and (s1n2411,n1024,n2344);
xor (n2412,n2413,n2341);
xor (n2413,n2336,n2339);
and (n2414,n2412,n2415);
or (n2415,n2416,n2420,n2446);
and (n2416,n2417,n2418);
wire s0n2417,s1n2417,notn2417;
or (n2417,s0n2417,s1n2417);
not(notn2417,n1024);
and (s0n2417,notn2417,1'b0);
and (s1n2417,n1024,n2351);
xor (n2418,n2419,n2348);
xor (n2419,n2343,n2346);
and (n2420,n2418,n2421);
or (n2421,n2422,n2426,n2445);
and (n2422,n2423,n2424);
wire s0n2423,s1n2423,notn2423;
or (n2423,s0n2423,s1n2423);
not(notn2423,n1024);
and (s0n2423,notn2423,1'b0);
and (s1n2423,n1024,n2358);
xor (n2424,n2425,n2355);
xor (n2425,n2350,n2353);
and (n2426,n2424,n2427);
or (n2427,n2428,n2432,n2444);
and (n2428,n2429,n2430);
wire s0n2429,s1n2429,notn2429;
or (n2429,s0n2429,s1n2429);
not(notn2429,n1024);
and (s0n2429,notn2429,1'b0);
and (s1n2429,n1024,n2365);
xor (n2430,n2431,n2362);
xor (n2431,n2357,n2360);
and (n2432,n2430,n2433);
or (n2433,n2434,n2438,n2443);
and (n2434,n2435,n2436);
wire s0n2435,s1n2435,notn2435;
or (n2435,s0n2435,s1n2435);
not(notn2435,n1024);
and (s0n2435,notn2435,1'b0);
and (s1n2435,n1024,n2371);
xor (n2436,n2437,n2368);
xor (n2437,n2364,n2366);
and (n2438,n2436,n2439);
and (n2439,n2440,n2441);
wire s0n2440,s1n2440,notn2440;
or (n2440,s0n2440,s1n2440);
not(notn2440,n1024);
and (s0n2440,notn2440,1'b0);
and (s1n2440,n1024,n2376);
xor (n2441,n2442,n2374);
xor (n2442,n2370,n2372);
and (n2443,n2435,n2439);
and (n2444,n2429,n2433);
and (n2445,n2423,n2427);
and (n2446,n2417,n2421);
and (n2447,n2411,n2415);
and (n2448,n2405,n2409);
and (n2449,n2399,n2403);
and (n2450,n2393,n2397);
and (n2451,n2388,n2391);
and (n2452,n2110,n2386);
or (n2453,n2454,n2459,n2547);
and (n2454,n2455,n2457);
xor (n2455,n2456,n2041);
xor (n2456,n1756,n1966);
xor (n2457,n2458,n2386);
xor (n2458,n2110,n2311);
and (n2459,n2457,n2460);
or (n2460,n2461,n2466,n2546);
and (n2461,n2462,n2464);
xor (n2462,n2463,n2046);
xor (n2463,n2043,n2044);
xor (n2464,n2465,n2391);
xor (n2465,n2388,n2389);
and (n2466,n2464,n2467);
or (n2467,n2468,n2473,n2545);
and (n2468,n2469,n2471);
xor (n2469,n2470,n2052);
xor (n2470,n2048,n2049);
xor (n2471,n2472,n2397);
xor (n2472,n2393,n2394);
and (n2473,n2471,n2474);
or (n2474,n2475,n2480,n2544);
and (n2475,n2476,n2478);
xor (n2476,n2477,n2058);
xor (n2477,n2054,n2055);
xor (n2478,n2479,n2403);
xor (n2479,n2399,n2400);
and (n2480,n2478,n2481);
or (n2481,n2482,n2487,n2543);
and (n2482,n2483,n2485);
xor (n2483,n2484,n2064);
xor (n2484,n2060,n2061);
xor (n2485,n2486,n2409);
xor (n2486,n2405,n2406);
and (n2487,n2485,n2488);
or (n2488,n2489,n2494,n2542);
and (n2489,n2490,n2492);
xor (n2490,n2491,n2070);
xor (n2491,n2066,n2067);
xor (n2492,n2493,n2415);
xor (n2493,n2411,n2412);
and (n2494,n2492,n2495);
or (n2495,n2496,n2501,n2541);
and (n2496,n2497,n2499);
xor (n2497,n2498,n2076);
xor (n2498,n2072,n2073);
xor (n2499,n2500,n2421);
xor (n2500,n2417,n2418);
and (n2501,n2499,n2502);
or (n2502,n2503,n2508,n2540);
and (n2503,n2504,n2506);
xor (n2504,n2505,n2082);
xor (n2505,n2078,n2079);
xor (n2506,n2507,n2427);
xor (n2507,n2423,n2424);
and (n2508,n2506,n2509);
or (n2509,n2510,n2515,n2539);
and (n2510,n2511,n2513);
xor (n2511,n2512,n2088);
xor (n2512,n2084,n2085);
xor (n2513,n2514,n2433);
xor (n2514,n2429,n2430);
and (n2515,n2513,n2516);
or (n2516,n2517,n2522,n2538);
and (n2517,n2518,n2520);
xor (n2518,n2519,n2094);
xor (n2519,n2090,n2091);
xor (n2520,n2521,n2439);
xor (n2521,n2435,n2436);
and (n2522,n2520,n2523);
or (n2523,n2524,n2527,n2537);
and (n2524,n2525,n2526);
xor (n2525,n2095,n2096);
xor (n2526,n2440,n2441);
and (n2527,n2526,n2528);
or (n2528,n2529,n2532,n2536);
and (n2529,n2530,n2531);
xor (n2530,n2030,n2032);
xor (n2531,n2375,n2377);
and (n2532,n2531,n2533);
and (n2533,n2534,n2535);
wire s0n2534,s1n2534,notn2534;
or (n2534,s0n2534,s1n2534);
not(notn2534,n930);
and (s0n2534,notn2534,1'b0);
and (s1n2534,n930,n2031);
wire s0n2535,s1n2535,notn2535;
or (n2535,s0n2535,s1n2535);
not(notn2535,n930);
and (s0n2535,notn2535,1'b0);
and (s1n2535,n930,n2376);
and (n2536,n2530,n2533);
and (n2537,n2525,n2528);
and (n2538,n2518,n2523);
and (n2539,n2511,n2516);
and (n2540,n2504,n2509);
and (n2541,n2497,n2502);
and (n2542,n2490,n2495);
and (n2543,n2483,n2488);
and (n2544,n2476,n2481);
and (n2545,n2469,n2474);
and (n2546,n2462,n2467);
and (n2547,n2455,n2460);
or (n2548,n2549,n2554,n2646);
and (n2549,n2550,n2552);
xor (n2550,n2551,n1664);
xor (n2551,n1659,n1661);
xor (n2552,n2553,n2460);
xor (n2553,n2455,n2457);
and (n2554,n2552,n2555);
or (n2555,n2556,n2561,n2645);
and (n2556,n2557,n2559);
xor (n2557,n2558,n1671);
xor (n2558,n1666,n1668);
xor (n2559,n2560,n2467);
xor (n2560,n2462,n2464);
and (n2561,n2559,n2562);
or (n2562,n2563,n2568,n2644);
and (n2563,n2564,n2566);
xor (n2564,n2565,n1678);
xor (n2565,n1673,n1675);
xor (n2566,n2567,n2474);
xor (n2567,n2469,n2471);
and (n2568,n2566,n2569);
or (n2569,n2570,n2575,n2643);
and (n2570,n2571,n2573);
xor (n2571,n2572,n1685);
xor (n2572,n1680,n1682);
xor (n2573,n2574,n2481);
xor (n2574,n2476,n2478);
and (n2575,n2573,n2576);
or (n2576,n2577,n2582,n2642);
and (n2577,n2578,n2580);
xor (n2578,n2579,n1692);
xor (n2579,n1687,n1689);
xor (n2580,n2581,n2488);
xor (n2581,n2483,n2485);
and (n2582,n2580,n2583);
or (n2583,n2584,n2589,n2641);
and (n2584,n2585,n2587);
xor (n2585,n2586,n1699);
xor (n2586,n1694,n1696);
xor (n2587,n2588,n2495);
xor (n2588,n2490,n2492);
and (n2589,n2587,n2590);
or (n2590,n2591,n2596,n2640);
and (n2591,n2592,n2594);
xor (n2592,n2593,n1706);
xor (n2593,n1701,n1703);
xor (n2594,n2595,n2502);
xor (n2595,n2497,n2499);
and (n2596,n2594,n2597);
or (n2597,n2598,n2603,n2639);
and (n2598,n2599,n2601);
xor (n2599,n2600,n1713);
xor (n2600,n1708,n1710);
xor (n2601,n2602,n2509);
xor (n2602,n2504,n2506);
and (n2603,n2601,n2604);
or (n2604,n2605,n2610,n2638);
and (n2605,n2606,n2608);
xor (n2606,n2607,n1720);
xor (n2607,n1715,n1717);
xor (n2608,n2609,n2516);
xor (n2609,n2511,n2513);
and (n2610,n2608,n2611);
or (n2611,n2612,n2617,n2637);
and (n2612,n2613,n2615);
xor (n2613,n2614,n1727);
xor (n2614,n1722,n1724);
xor (n2615,n2616,n2523);
xor (n2616,n2518,n2520);
and (n2617,n2615,n2618);
or (n2618,n2619,n2624,n2636);
and (n2619,n2620,n2622);
xor (n2620,n2621,n1732);
xor (n2621,n1729,n1730);
xor (n2622,n2623,n2528);
xor (n2623,n2525,n2526);
and (n2624,n2622,n2625);
or (n2625,n2626,n2631,n2635);
and (n2626,n2627,n2629);
xor (n2627,n2628,n1737);
xor (n2628,n1734,n1735);
xor (n2629,n2630,n2533);
xor (n2630,n2530,n2531);
and (n2631,n2629,n2632);
and (n2632,n2633,n2634);
xor (n2633,n1738,n1739);
xor (n2634,n2534,n2535);
and (n2635,n2627,n2632);
and (n2636,n2620,n2625);
and (n2637,n2613,n2618);
and (n2638,n2606,n2611);
and (n2639,n2599,n2604);
and (n2640,n2592,n2597);
and (n2641,n2585,n2590);
and (n2642,n2578,n2583);
and (n2643,n2571,n2576);
and (n2644,n2564,n2569);
and (n2645,n2557,n2562);
and (n2646,n2550,n2555);
and (n2647,n2648,n2650);
xor (n2648,n2649,n2555);
xor (n2649,n2550,n2552);
and (n2650,n2651,n2653);
xor (n2651,n2652,n2562);
xor (n2652,n2557,n2559);
and (n2653,n2654,n2656);
xor (n2654,n2655,n2569);
xor (n2655,n2564,n2566);
and (n2656,n2657,n2659);
xor (n2657,n2658,n2576);
xor (n2658,n2571,n2573);
and (n2659,n2660,n2662);
xor (n2660,n2661,n2583);
xor (n2661,n2578,n2580);
and (n2662,n2663,n2665);
xor (n2663,n2664,n2590);
xor (n2664,n2585,n2587);
and (n2665,n2666,n2668);
xor (n2666,n2667,n2597);
xor (n2667,n2592,n2594);
xor (n2668,n2669,n2604);
xor (n2669,n2599,n2601);
nand (n2670,n2671,n3552);
or (n2671,n2672,n3073);
not (n2672,n2673);
nor (n2673,n2674,n2676);
and (n2674,n2675,n3048);
not (n2675,n2676);
or (n2676,n2677,n3047);
and (n2677,n2678,n2996);
xor (n2678,n2679,n2971);
or (n2679,n2680,n2970);
and (n2680,n2681,n2822);
xor (n2681,n2682,n2797);
xor (n2682,n2683,n2724);
xor (n2683,n2684,n2686);
xor (n2684,n2685,n1210);
xor (n2685,n1084,n2043);
xor (n2686,n2687,n2312);
xor (n2687,n2688,n2722);
or (n2688,n2689,n2721);
and (n2689,n2690,n2393);
xor (n2690,n2691,n1583);
and (n2691,n2692,n1591);
xor (n2692,n1590,n2693);
xor (n2693,n2694,n2701);
xor (n2694,n2695,n2700);
xor (n2695,n2696,n2699);
xor (n2696,n2697,n2698);
nor (n2697,n2114,n1082);
and (n2698,n1295,n930);
and (n2699,n2698,n1313);
and (n2700,n2697,n2132);
or (n2701,n2702,n2720);
and (n2702,n2703,n2712);
xor (n2703,n2704,n2707);
nor (n2704,n2705,n1082);
xnor (n2705,n2262,n2706);
not (n2706,n2129);
and (n2707,n2708,n930);
nand (n2708,n2709,n2711);
or (n2709,n2710,n1442);
not (n2710,n1310);
or (n2711,n1443,n1310);
and (n2712,n2713,n930);
or (n2713,n2714,n2718);
nor (n2714,n2715,n2717);
and (n2715,n2268,n2716);
not (n2716,n2146);
not (n2717,n2132);
nor (n2718,n2719,n2114);
not (n2719,n2182);
and (n2720,n2704,n2707);
and (n2721,n2691,n1583);
xor (n2722,n2723,n1576);
xor (n2723,n1500,n1575);
or (n2724,n2725,n2796);
and (n2725,n2726,n2732);
xor (n2726,n2727,n2731);
or (n2727,n2728,n2730);
and (n2728,n2729,n1225);
xor (n2729,n1977,n2054);
and (n2730,n1977,n2054);
xor (n2731,n2690,n2393);
and (n2732,n2733,n1093);
xor (n2733,n1224,n2734);
or (n2734,n2735,n2795);
and (n2735,n2736,n2769);
xor (n2736,n2405,n2737);
and (n2737,n2738,n2763);
or (n2738,n2739,n2762);
and (n2739,n2740,n2754);
xor (n2740,n2741,n2748);
and (n2741,n2742,n930);
nand (n2742,n2743,n2745,n2747);
or (n2743,n2744,n2268);
not (n2744,n2218);
or (n2745,n2275,n2746);
not (n2746,n2186);
not (n2747,n2167);
nor (n2748,n1082,n2749);
nor (n2749,n1348,n2750);
nor (n2750,n2751,n1463);
and (n2751,n2752,n2753);
not (n2752,n1363);
not (n2753,n1349);
nor (n2754,n2755,n1082);
nor (n2755,n2756,n2760);
and (n2756,n2757,n1331);
not (n2757,n2758);
xor (n2758,n1456,n2759);
not (n2759,n1345);
and (n2760,n2758,n2761);
not (n2761,n1331);
and (n2762,n2741,n2748);
and (n2763,n2764,n930);
nor (n2764,n2765,n2767);
and (n2765,n2766,n2132);
xor (n2766,n2268,n2716);
and (n2767,n2768,n2717);
not (n2768,n2766);
or (n2769,n2770,n2794);
and (n2770,n2771,n2411);
xor (n2771,n1607,n2772);
xor (n2772,n2773,n2786);
xor (n2773,n2774,n2779);
and (n2774,n2775,n930);
nand (n2775,n2776,n2777,n2778);
or (n2776,n1449,n2753);
not (n2777,n1330);
or (n2778,n1456,n2759);
and (n2779,n2780,n930);
nand (n2780,n2781,n2785);
or (n2781,n2782,n2275);
and (n2782,n2783,n2784);
not (n2783,n2150);
not (n2784,n2164);
not (n2785,n2149);
and (n2786,n2787,n930);
nor (n2787,n2788,n2791);
and (n2788,n2789,n1313);
xor (n2789,n2790,n1449);
not (n2790,n1327);
and (n2791,n2792,n2793);
not (n2792,n2789);
not (n2793,n1313);
and (n2794,n1607,n2772);
and (n2795,n2405,n2737);
and (n2796,n2727,n2731);
xor (n2797,n2798,n2818);
xor (n2798,n2799,n2808);
xor (n2799,n2800,n2388);
xor (n2800,n1209,n2801);
and (n2801,n2802,n2805);
or (n2802,n2803,n2804);
and (n2803,n2694,n2701);
and (n2804,n2695,n2700);
or (n2805,n2806,n2807);
and (n2806,n2696,n2699);
and (n2807,n2697,n2698);
or (n2808,n2809,n2817);
and (n2809,n2810,n1217);
xor (n2810,n2811,n2048);
or (n2811,n2812,n2816);
and (n2812,n2813,n2322);
xor (n2813,n2814,n2815);
xor (n2814,n2692,n1591);
and (n2815,n1597,n1515);
and (n2816,n2814,n2815);
and (n2817,n2811,n2048);
or (n2818,n2819,n2821);
and (n2819,n2820,n1088);
xor (n2820,n1089,n1973);
and (n2821,n1089,n1973);
or (n2822,n2823,n2969);
and (n2823,n2824,n2849);
xor (n2824,n2825,n2826);
xor (n2825,n2726,n2732);
or (n2826,n2827,n2848);
and (n2827,n2828,n2835);
xor (n2828,n2829,n2830);
xor (n2829,n2733,n1093);
or (n2830,n2831,n2834);
and (n2831,n2832,n1987);
xor (n2832,n1233,n2833);
xor (n2833,n2736,n2769);
and (n2834,n1233,n2833);
or (n2835,n2836,n2847);
and (n2836,n2837,n1100);
xor (n2837,n1984,n2838);
or (n2838,n2839,n2846);
and (n2839,n2840,n1240);
xor (n2840,n2841,n2843);
xor (n2841,n2842,n1606);
xor (n2842,n2738,n2763);
and (n2843,n2844,n2417);
xor (n2844,n2845,n1614);
xor (n2845,n2740,n2754);
and (n2846,n2841,n2843);
and (n2847,n1984,n2838);
and (n2848,n2829,n2830);
or (n2849,n2850,n2968);
and (n2850,n2851,n2950);
xor (n2851,n2852,n2949);
or (n2852,n2853,n2948);
and (n2853,n2854,n1152);
xor (n2854,n2855,n2882);
or (n2855,n2856,n2881);
and (n2856,n2857,n2066);
xor (n2857,n2858,n2859);
xor (n2858,n2771,n2411);
or (n2859,n2860,n2880);
and (n2860,n2861,n2343);
xor (n2861,n1529,n2862);
or (n2862,n2863,n2879);
and (n2863,n2864,n1623);
xor (n2864,n2865,n2875);
and (n2865,n2866,n930);
nand (n2866,n2867,n2873);
or (n2867,n2168,n2868);
not (n2868,n2869);
nand (n2869,n2870,n2872);
or (n2870,n2182,n2871);
not (n2871,n2281);
or (n2872,n2281,n2719);
or (n2873,n2869,n2874);
not (n2874,n2168);
and (n2875,n2876,n930);
nand (n2876,n2877,n2878);
or (n2877,n1463,n1465);
nand (n2878,n1465,n1463);
and (n2879,n2865,n2875);
and (n2880,n1529,n2862);
and (n2881,n2858,n2859);
or (n2882,n2883,n2947);
and (n2883,n2884,n1241);
xor (n2884,n2885,n2906);
xor (n2885,n2886,n2336);
xor (n2886,n1522,n2887);
or (n2887,n2888,n2905);
and (n2888,n2889,n1615);
xor (n2889,n2890,n2903);
or (n2890,n2891,n2898);
and (n2891,n2892,n930);
nand (n2892,n2893,n2895,n2897);
or (n2893,n1456,n2894);
not (n2894,n1417);
or (n2895,n1463,n2896);
not (n2896,n1385);
not (n2897,n1366);
and (n2898,n2899,n930);
or (n2899,n2900,n2185);
nor (n2900,n2901,n2288);
and (n2901,n2902,n2746);
not (n2902,n2200);
nor (n2903,n2904,n1082);
xor (n2904,n2277,n2275);
and (n2905,n2890,n2903);
and (n2906,n2907,n2946);
xor (n2907,n2908,n2944);
or (n2908,n2909,n2943);
and (n2909,n2910,n2423);
xor (n2910,n2911,n2921);
and (n2911,n2912,n2919);
xor (n2912,n2913,n1630);
and (n2913,n2914,n2916);
nor (n2914,n2915,n2288);
not (n2915,n2535);
and (n2916,n2917,n930);
nor (n2917,n2918,n2894);
not (n2918,n1482);
and (n2919,n2920,n930);
xnor (n2920,n2288,n2290);
or (n2921,n2922,n2942);
and (n2922,n2923,n2937);
xor (n2923,n2924,n2930);
and (n2924,n2925,n930);
nand (n2925,n2926,n2927,n2929);
or (n2926,n1477,n2896);
or (n2927,n1463,n2928);
not (n2928,n1434);
not (n2929,n1384);
and (n2930,n2931,n930);
not (n2931,n2932);
nor (n2932,n2933,n2934);
and (n2933,n2287,n2222);
nor (n2934,n2935,n2744);
and (n2935,n2295,n2936);
not (n2936,n2204);
and (n2937,n2938,n930);
xor (n2938,n2939,n2940);
not (n2939,n1367);
xnor (n2940,n1470,n2941);
not (n2941,n1381);
and (n2942,n2924,n2930);
and (n2943,n2911,n2921);
and (n2944,n2945,n1536);
xor (n2945,n2350,n1622);
xor (n2946,n2844,n2417);
and (n2947,n2885,n2906);
and (n2948,n2855,n2882);
xor (n2949,n2729,n1225);
xor (n2950,n2951,n1096);
xor (n2951,n1980,n2952);
xor (n2952,n2953,n2399);
xor (n2953,n1508,n2954);
or (n2954,n2955,n2967);
and (n2955,n2956,n2964);
xor (n2956,n2957,n2958);
xor (n2957,n2703,n2712);
and (n2958,n2959,n930);
nand (n2959,n2960,n2962);
or (n2960,n2961,n2793);
and (n2961,n2790,n1449);
or (n2962,n2752,n2963);
not (n2963,n1295);
or (n2964,n2965,n2966);
and (n2965,n2773,n2786);
and (n2966,n2774,n2779);
and (n2967,n2957,n2958);
and (n2968,n2852,n2949);
and (n2969,n2825,n2826);
and (n2970,n2682,n2797);
xor (n2971,n2972,n2989);
xor (n2972,n2973,n2976);
or (n2973,n2974,n2975);
and (n2974,n2798,n2818);
and (n2975,n2799,n2808);
and (n2976,n2977,n2984);
xor (n2977,n2978,n1967);
or (n2978,n2979,n2983);
and (n2979,n2980,n1970);
xor (n2980,n1503,n2981);
xor (n2981,n2982,n1582);
xor (n2982,n2802,n2805);
and (n2983,n1503,n2981);
and (n2984,n2985,n2315);
xor (n2985,n1216,n2986);
or (n2986,n2987,n2988);
and (n2987,n2953,n2399);
and (n2988,n1508,n2954);
xor (n2989,n2990,n2993);
xor (n2990,n2991,n2992);
and (n2991,n2800,n2388);
and (n2992,n2723,n1576);
or (n2993,n2994,n2995);
and (n2994,n2685,n1210);
and (n2995,n1084,n2043);
xor (n2996,n2997,n3009);
xor (n2997,n2998,n3001);
or (n2998,n2999,n3000);
and (n2999,n2683,n2724);
and (n3000,n2684,n2686);
xor (n3001,n3002,n3007);
xor (n3002,n3003,n3006);
or (n3003,n3004,n3005);
and (n3004,n2687,n2312);
and (n3005,n2688,n2722);
xor (n3006,n1494,n1074);
xor (n3007,n3008,n1077);
xor (n3008,n1756,n2110);
or (n3009,n3010,n3046);
and (n3010,n3011,n3022);
xor (n3011,n3012,n3021);
or (n3012,n3013,n3020);
and (n3013,n3014,n3017);
xor (n3014,n3015,n3016);
xor (n3015,n2810,n1217);
xor (n3016,n2980,n1970);
or (n3017,n3018,n3019);
and (n3018,n2951,n1096);
and (n3019,n1980,n2952);
and (n3020,n3015,n3016);
xor (n3021,n2977,n2984);
or (n3022,n3023,n3045);
and (n3023,n3024,n3044);
xor (n3024,n3025,n3026);
xor (n3025,n2985,n2315);
or (n3026,n3027,n3043);
and (n3027,n3028,n3038);
xor (n3028,n3029,n3030);
xor (n3029,n2813,n2322);
or (n3030,n3031,n3037);
and (n3031,n3032,n2329);
xor (n3032,n3033,n3036);
or (n3033,n3034,n3035);
and (n3034,n2886,n2336);
and (n3035,n1522,n2887);
xor (n3036,n2956,n2964);
and (n3037,n3033,n3036);
or (n3038,n3039,n3042);
and (n3039,n3040,n2060);
xor (n3040,n1232,n3041);
xor (n3041,n1597,n1515);
and (n3042,n1232,n3041);
and (n3043,n3029,n3030);
xor (n3044,n2820,n1088);
and (n3045,n3025,n3026);
and (n3046,n3012,n3021);
and (n3047,n2679,n2971);
not (n3048,n3049);
nor (n3049,n3050,n3052);
and (n3050,n3051,n3055);
not (n3051,n3052);
or (n3052,n3053,n3054);
and (n3053,n2997,n3009);
and (n3054,n2998,n3001);
not (n3055,n3056);
nor (n3056,n3057,n3070);
not (n3057,n3058);
nor (n3058,n3059,n3067);
not (n3059,n3060);
nor (n3060,n3061,n3062);
and (n3061,n3008,n1077);
not (n3062,n3063);
nor (n3063,n3064,n3065);
and (n3064,n1494,n1074);
not (n3065,n3066);
xnor (n3066,n6,n1292);
or (n3067,n3068,n3069);
and (n3068,n3002,n3007);
and (n3069,n3003,n3006);
or (n3070,n3071,n3072);
and (n3071,n2972,n2989);
and (n3072,n2973,n2976);
not (n3073,n3074);
or (n3074,n3075,n3551);
and (n3075,n3076,n3136);
xor (n3076,n3077,n3078);
xor (n3077,n2678,n2996);
or (n3078,n3079,n3135);
and (n3079,n3080,n3134);
xor (n3080,n3081,n3082);
xor (n3081,n3011,n3022);
or (n3082,n3083,n3133);
and (n3083,n3084,n3087);
xor (n3084,n3085,n3086);
xor (n3085,n3024,n3044);
xor (n3086,n3014,n3017);
or (n3087,n3088,n3132);
and (n3088,n3089,n3122);
xor (n3089,n3090,n3121);
or (n3090,n3091,n3120);
and (n3091,n3092,n3095);
xor (n3092,n3093,n3094);
xor (n3093,n3040,n2060);
xor (n3094,n3032,n2329);
or (n3095,n3096,n3119);
and (n3096,n3097,n1994);
xor (n3097,n3098,n3116);
or (n3098,n3099,n3115);
and (n3099,n3100,n1249);
xor (n3100,n3101,n3102);
xor (n3101,n2861,n2343);
or (n3102,n3103,n3114);
and (n3103,n3104,n3110);
xor (n3104,n3105,n3106);
xor (n3105,n2864,n1623);
nand (n3106,n3107,n2890);
or (n3107,n3108,n3109);
not (n3108,n2898);
not (n3109,n2891);
or (n3110,n3111,n3113);
and (n3111,n3112,n1543);
xor (n3112,n1631,n2429);
and (n3113,n1631,n2429);
and (n3114,n3105,n3106);
and (n3115,n3101,n3102);
and (n3116,n3117,n2072);
xor (n3117,n1248,n3118);
xor (n3118,n2889,n1615);
and (n3119,n3098,n3116);
and (n3120,n3093,n3094);
xor (n3121,n3028,n3038);
or (n3122,n3123,n3131);
and (n3123,n3124,n3130);
xor (n3124,n3125,n3126);
xor (n3125,n2832,n1987);
or (n3126,n3127,n3129);
and (n3127,n3128,n1159);
xor (n3128,n1156,n1991);
and (n3129,n1156,n1991);
xor (n3130,n2837,n1100);
and (n3131,n3125,n3126);
and (n3132,n3090,n3121);
and (n3133,n3085,n3086);
xor (n3134,n2681,n2822);
and (n3135,n3081,n3082);
or (n3136,n3137,n3550);
and (n3137,n3138,n3202);
xor (n3138,n3139,n3140);
xor (n3139,n3080,n3134);
or (n3140,n3141,n3201);
and (n3141,n3142,n3200);
xor (n3142,n3143,n3144);
xor (n3143,n2824,n2849);
or (n3144,n3145,n3199);
and (n3145,n3146,n3149);
xor (n3146,n3147,n3148);
xor (n3147,n2828,n2835);
xor (n3148,n2851,n2950);
or (n3149,n3150,n3198);
and (n3150,n3151,n3182);
xor (n3151,n3152,n3153);
xor (n3152,n2854,n1152);
or (n3153,n3154,n3181);
and (n3154,n3155,n3158);
xor (n3155,n3156,n3157);
xor (n3156,n2857,n2066);
xor (n3157,n2840,n1240);
or (n3158,n3159,n3180);
and (n3159,n3160,n1998);
xor (n3160,n3161,n1163);
and (n3161,n3162,n3163);
xor (n3162,n2910,n2423);
or (n3163,n3164,n3179);
and (n3164,n3165,n2357);
xor (n3165,n3166,n3178);
or (n3166,n3167,n3177);
and (n3167,n3168,n3170);
xor (n3168,n2435,n3169);
and (n3169,n2440,n2095);
and (n3170,n3171,n930);
nand (n3171,n3172,n3176);
or (n3172,n2936,n3173);
nand (n3173,n3174,n3175);
or (n3174,n2218,n2295);
nand (n3175,n2218,n2295);
nand (n3176,n3173,n2936);
and (n3177,n2435,n3169);
xor (n3178,n2923,n2937);
and (n3179,n3166,n3178);
and (n3180,n3161,n1163);
and (n3181,n3156,n3157);
or (n3182,n3183,n3197);
and (n3183,n3184,n3196);
xor (n3184,n3185,n3186);
xor (n3185,n2884,n1241);
or (n3186,n3187,n3195);
and (n3187,n3188,n1166);
xor (n3188,n3189,n3194);
or (n3189,n3190,n3193);
and (n3190,n3191,n1257);
xor (n3191,n3192,n2078);
xor (n3192,n2945,n1536);
and (n3193,n3192,n2078);
xor (n3194,n2907,n2946);
and (n3195,n3189,n3194);
xor (n3196,n3128,n1159);
and (n3197,n3185,n3186);
and (n3198,n3152,n3153);
and (n3199,n3147,n3148);
xor (n3200,n3084,n3087);
and (n3201,n3143,n3144);
or (n3202,n3203,n3549);
and (n3203,n3204,n3313);
xor (n3204,n3205,n3206);
xor (n3205,n3142,n3200);
or (n3206,n3207,n3312);
and (n3207,n3208,n3311);
xor (n3208,n3209,n3210);
xor (n3209,n3089,n3122);
or (n3210,n3211,n3310);
and (n3211,n3212,n3309);
xor (n3212,n3213,n3214);
xor (n3213,n3092,n3095);
or (n3214,n3215,n3308);
and (n3215,n3216,n3247);
xor (n3216,n3217,n3246);
or (n3217,n3218,n3245);
and (n3218,n3219,n3221);
xor (n3219,n3220,n2001);
xor (n3220,n3117,n2072);
or (n3221,n3222,n3244);
and (n3222,n3223,n1170);
xor (n3223,n3224,n3231);
or (n3224,n3225,n3230);
and (n3225,n3226,n1265);
xor (n3226,n2084,n3227);
and (n3227,n3228,n2364);
xor (n3228,n3229,n1638);
xor (n3229,n2914,n2916);
and (n3230,n2084,n3227);
or (n3231,n3232,n3243);
and (n3232,n3233,n1264);
xor (n3233,n3234,n3235);
xor (n3234,n2912,n2919);
and (n3235,n3236,n1639);
xor (n3236,n3237,n1272);
and (n3237,n3238,n930);
xnor (n3238,n3239,n2896);
nand (n3239,n3240,n3242);
or (n3240,n1476,n3241);
not (n3241,n1399);
nand (n3242,n1476,n3241);
and (n3243,n3234,n3235);
and (n3244,n3224,n3231);
and (n3245,n3220,n2001);
xor (n3246,n3097,n1994);
or (n3247,n3248,n3307);
and (n3248,n3249,n3306);
xor (n3249,n3250,n3305);
or (n3250,n3251,n3304);
and (n3251,n3252,n2005);
xor (n3252,n3253,n3254);
xor (n3253,n3104,n3110);
or (n3254,n3255,n3303);
and (n3255,n3256,n3282);
xor (n3256,n3257,n3258);
xor (n3257,n3112,n1543);
or (n3258,n3259,n3281);
and (n3259,n3260,n1550);
xor (n3260,n3261,n3270);
or (n3261,n3262,n3269);
and (n3262,n3263,n3265);
xor (n3263,n2370,n3264);
xor (n3264,n2440,n2095);
and (n3265,n3266,n930);
nand (n3266,n3267,n3268);
or (n3267,n1417,n2918);
or (n3268,n1482,n2894);
and (n3269,n2370,n3264);
or (n3270,n3271,n3280);
and (n3271,n3272,n3275);
xor (n3272,n3273,n3274);
and (n3273,n1403,n930);
and (n3274,n2222,n930);
and (n3275,n3276,n930);
nand (n3276,n3277,n3279);
or (n3277,n2300,n3278);
not (n3278,n2236);
nand (n3279,n2300,n3278);
and (n3280,n3273,n3274);
and (n3281,n3261,n3270);
or (n3282,n3283,n3302);
and (n3283,n3284,n2090);
xor (n3284,n3285,n3286);
xor (n3285,n3168,n3170);
or (n3286,n3287,n3301);
and (n3287,n3288,n1278);
xor (n3288,n3289,n3296);
or (n3289,n3290,n3295);
and (n3290,n3291,n3293);
xor (n3291,n3292,n2375);
nor (n3292,n2928,n1082);
nor (n3293,n3294,n1082);
not (n3294,n2253);
and (n3295,n3292,n2375);
and (n3296,n3297,n3299);
nor (n3297,n3298,n1082);
not (n3298,n1420);
nor (n3299,n3300,n1082);
not (n3300,n2239);
and (n3301,n3289,n3296);
and (n3302,n3285,n3286);
and (n3303,n3257,n3258);
and (n3304,n3253,n3254);
xor (n3305,n3100,n1249);
xor (n3306,n3160,n1998);
and (n3307,n3250,n3305);
and (n3308,n3217,n3246);
xor (n3309,n3124,n3130);
and (n3310,n3213,n3214);
xor (n3311,n3146,n3149);
and (n3312,n3209,n3210);
or (n3313,n3314,n3548);
and (n3314,n3315,n3365);
xor (n3315,n3316,n3317);
xor (n3316,n3208,n3311);
or (n3317,n3318,n3364);
and (n3318,n3319,n3363);
xor (n3319,n3320,n3321);
xor (n3320,n3151,n3182);
or (n3321,n3322,n3362);
and (n3322,n3323,n3361);
xor (n3323,n3324,n3325);
xor (n3324,n3155,n3158);
or (n3325,n3326,n3360);
and (n3326,n3327,n3359);
xor (n3327,n3328,n3334);
or (n3328,n3329,n3333);
and (n3329,n3330,n2008);
xor (n3330,n3331,n1173);
xor (n3331,n3332,n1256);
xor (n3332,n3162,n3163);
and (n3333,n3331,n1173);
or (n3334,n3335,n3358);
and (n3335,n3336,n3353);
xor (n3336,n3337,n3352);
or (n3337,n3338,n3351);
and (n3338,n3339,n1177);
xor (n3339,n3340,n3341);
xor (n3340,n3233,n1264);
or (n3341,n3342,n3350);
and (n3342,n3343,n3349);
xor (n3343,n1273,n3344);
or (n3344,n3345,n3348);
and (n3345,n3346,n1644);
xor (n3346,n3347,n1556);
xor (n3347,n3272,n3275);
and (n3348,n3347,n1556);
xor (n3349,n3228,n2364);
and (n3350,n1273,n3344);
and (n3351,n3340,n3341);
xor (n3352,n3191,n1257);
or (n3353,n3354,n3357);
and (n3354,n3355,n1180);
xor (n3355,n2012,n3356);
xor (n3356,n3165,n2357);
and (n3357,n2012,n3356);
and (n3358,n3337,n3352);
xor (n3359,n3188,n1166);
and (n3360,n3328,n3334);
xor (n3361,n3184,n3196);
and (n3362,n3324,n3325);
xor (n3363,n3212,n3309);
and (n3364,n3320,n3321);
or (n3365,n3366,n3547);
and (n3366,n3367,n3397);
xor (n3367,n3368,n3396);
or (n3368,n3369,n3395);
and (n3369,n3370,n3394);
xor (n3370,n3371,n3393);
or (n3371,n3372,n3392);
and (n3372,n3373,n3391);
xor (n3373,n3374,n3390);
or (n3374,n3375,n3389);
and (n3375,n3376,n3379);
xor (n3376,n3377,n3378);
xor (n3377,n3223,n1170);
xor (n3378,n3252,n2005);
or (n3379,n3380,n3388);
and (n3380,n3381,n2015);
xor (n3381,n3382,n3383);
xor (n3382,n3226,n1265);
or (n3383,n3384,n3387);
and (n3384,n3385,n1184);
xor (n3385,n3386,n2019);
xor (n3386,n3236,n1639);
and (n3387,n3386,n2019);
and (n3388,n3382,n3383);
and (n3389,n3377,n3378);
xor (n3390,n3219,n3221);
xor (n3391,n3249,n3306);
and (n3392,n3374,n3390);
xor (n3393,n3216,n3247);
xor (n3394,n3323,n3361);
and (n3395,n3371,n3393);
xor (n3396,n3319,n3363);
or (n3397,n3398,n3546);
and (n3398,n3399,n3455);
xor (n3399,n3400,n3454);
or (n3400,n3401,n3453);
and (n3401,n3402,n3452);
xor (n3402,n3403,n3451);
or (n3403,n3404,n3450);
and (n3404,n3405,n3443);
xor (n3405,n3406,n3442);
or (n3406,n3407,n3441);
and (n3407,n3408,n3427);
xor (n3408,n3409,n3426);
or (n3409,n3410,n3425);
and (n3410,n3411,n3424);
xor (n3411,n3412,n3423);
or (n3412,n3413,n3422);
and (n3413,n3414,n1190);
xor (n3414,n3415,n3416);
xor (n3415,n3263,n3265);
or (n3416,n3417,n3421);
and (n3417,n3418,n3420);
xor (n3418,n3419,n2030);
and (n3419,n1739,n2534);
xor (n3420,n3297,n3299);
and (n3421,n3419,n2030);
and (n3422,n3415,n3416);
xor (n3423,n3260,n1550);
xor (n3424,n3284,n2090);
and (n3425,n3412,n3423);
xor (n3426,n3256,n3282);
or (n3427,n3428,n3440);
and (n3428,n3429,n1186);
xor (n3429,n3430,n2021);
or (n3430,n3431,n3439);
and (n3431,n3432,n3438);
xor (n3432,n2025,n3433);
or (n3433,n3434,n3437);
and (n3434,n3435,n1561);
xor (n3435,n1195,n3436);
xor (n3436,n3291,n3293);
and (n3437,n1195,n3436);
xor (n3438,n3346,n1644);
and (n3439,n2025,n3433);
and (n3440,n3430,n2021);
and (n3441,n3409,n3426);
xor (n3442,n3330,n2008);
or (n3443,n3444,n3449);
and (n3444,n3445,n3448);
xor (n3445,n3446,n3447);
xor (n3446,n3339,n1177);
xor (n3447,n3355,n1180);
xor (n3448,n3381,n2015);
and (n3449,n3446,n3447);
and (n3450,n3406,n3442);
xor (n3451,n3327,n3359);
xor (n3452,n3373,n3391);
and (n3453,n3403,n3451);
xor (n3454,n3370,n3394);
or (n3455,n3456,n3545);
and (n3456,n3457,n3544);
xor (n3457,n3458,n3497);
or (n3458,n3459,n3496);
and (n3459,n3460,n3495);
xor (n3460,n3461,n3494);
or (n3461,n3462,n3493);
and (n3462,n3463,n3476);
xor (n3463,n3464,n3475);
or (n3464,n3465,n3474);
and (n3465,n3466,n3473);
xor (n3466,n3467,n3472);
or (n3467,n3468,n3471);
and (n3468,n3469,n1192);
xor (n3469,n2027,n3470);
xor (n3470,n3288,n1278);
and (n3471,n2027,n3470);
xor (n3472,n3343,n3349);
xor (n3473,n3385,n1184);
and (n3474,n3467,n3472);
xor (n3475,n3408,n3427);
or (n3476,n3477,n3492);
and (n3477,n3478,n3491);
xor (n3478,n3479,n3480);
xor (n3479,n3411,n3424);
or (n3480,n3481,n3490);
and (n3481,n3482,n3489);
xor (n3482,n3483,n3488);
or (n3483,n3484,n3487);
and (n3484,n3485,n2032);
xor (n3485,n1197,n3486);
xor (n3486,n3418,n3420);
and (n3487,n1197,n3486);
xor (n3488,n3414,n1190);
xor (n3489,n3432,n3438);
and (n3490,n3483,n3488);
xor (n3491,n3429,n1186);
and (n3492,n3479,n3480);
and (n3493,n3464,n3475);
xor (n3494,n3336,n3353);
xor (n3495,n3376,n3379);
and (n3496,n3461,n3494);
nand (n3497,n3498,n3540);
or (n3498,n3499,n3538);
not (n3499,n3500);
nand (n3500,n3501,n3503,n3537);
not (n3501,n3502);
xor (n3502,n3405,n3443);
nand (n3503,n3504,n3536);
or (n3504,n3505,n3506);
xor (n3505,n3463,n3476);
nand (n3506,n3507,n3533);
or (n3507,n3508,n3531);
not (n3508,n3509);
nand (n3509,n3510,n3528);
or (n3510,n3511,n3526);
not (n3511,n3512);
nand (n3512,n3513,n3523);
or (n3513,n3514,n3521);
not (n3514,n3515);
nand (n3515,n3516,n3518);
or (n3516,n2915,n3517);
not (n3517,n1738);
nand (n3518,n3519,n3520);
or (n3519,n1738,n2535);
xor (n3520,n1739,n2534);
not (n3521,n3522);
xor (n3522,n3435,n1561);
nand (n3523,n3524,n3525);
or (n3524,n3522,n3515);
xor (n3525,n3485,n2032);
not (n3526,n3527);
xor (n3527,n3469,n1192);
nand (n3528,n3529,n3530);
or (n3529,n3527,n3512);
xor (n3530,n3482,n3489);
not (n3531,n3532);
xor (n3532,n3466,n3473);
nand (n3533,n3534,n3535);
or (n3534,n3532,n3509);
xor (n3535,n3478,n3491);
xor (n3536,n3445,n3448);
nand (n3537,n3505,n3506);
not (n3538,n3539);
xor (n3539,n3460,n3495);
nand (n3540,n3541,n3502);
or (n3541,n3542,n3543);
not (n3542,n3537);
not (n3543,n3503);
xor (n3544,n3402,n3452);
and (n3545,n3458,n3497);
and (n3546,n3400,n3454);
and (n3547,n3368,n3396);
and (n3548,n3316,n3317);
and (n3549,n3205,n3206);
and (n3550,n3139,n3140);
and (n3551,n3077,n3078);
or (n3552,n3074,n2673);
endmodule
