module top (out,n20,n21,n25,n27,n29,n30,n33,n35,n37
        ,n39,n40,n41,n42,n43,n44,n45,n46,n47,n48
        ,n49,n50,n51,n52,n53,n54,n55,n56,n57,n58
        ,n59,n60,n61,n62,n63,n64,n65,n66,n67,n70
        ,n71,n75,n77,n79,n80,n81,n85,n86,n87,n94
        ,n95,n96,n105,n106,n107,n111,n112,n113,n119,n120
        ,n121,n129,n130,n131,n139,n140,n141,n164,n165,n166
        ,n169,n170,n171,n182,n183,n184,n194,n195,n196,n210
        ,n211,n212,n221,n222,n223,n229,n230,n231,n237,n238
        ,n239,n250,n251,n252,n260,n261,n262,n269,n270,n271
        ,n284,n285,n286,n289,n290,n291,n298,n299,n300,n307
        ,n308,n309,n334,n335,n336,n348,n349,n350,n360,n361
        ,n362,n435,n436,n437,n939,n940,n941,n959,n960,n961
        ,n1023,n1024,n1028,n1030,n1032,n1035,n1036,n1040,n1042,n1044
        ,n1045,n1048,n1050,n1052,n1054,n1055,n1056,n1057,n1058,n1059
        ,n1060,n1061,n1062,n1063,n1064,n1065,n1066,n1067,n1068,n1069
        ,n1070,n1071,n1072,n1073,n1074,n1075,n1076,n1077,n1078,n1079
        ,n1080,n1081,n1082);
output out;
input n20;
input n21;
input n25;
input n27;
input n29;
input n30;
input n33;
input n35;
input n37;
input n39;
input n40;
input n41;
input n42;
input n43;
input n44;
input n45;
input n46;
input n47;
input n48;
input n49;
input n50;
input n51;
input n52;
input n53;
input n54;
input n55;
input n56;
input n57;
input n58;
input n59;
input n60;
input n61;
input n62;
input n63;
input n64;
input n65;
input n66;
input n67;
input n70;
input n71;
input n75;
input n77;
input n79;
input n80;
input n81;
input n85;
input n86;
input n87;
input n94;
input n95;
input n96;
input n105;
input n106;
input n107;
input n111;
input n112;
input n113;
input n119;
input n120;
input n121;
input n129;
input n130;
input n131;
input n139;
input n140;
input n141;
input n164;
input n165;
input n166;
input n169;
input n170;
input n171;
input n182;
input n183;
input n184;
input n194;
input n195;
input n196;
input n210;
input n211;
input n212;
input n221;
input n222;
input n223;
input n229;
input n230;
input n231;
input n237;
input n238;
input n239;
input n250;
input n251;
input n252;
input n260;
input n261;
input n262;
input n269;
input n270;
input n271;
input n284;
input n285;
input n286;
input n289;
input n290;
input n291;
input n298;
input n299;
input n300;
input n307;
input n308;
input n309;
input n334;
input n335;
input n336;
input n348;
input n349;
input n350;
input n360;
input n361;
input n362;
input n435;
input n436;
input n437;
input n939;
input n940;
input n941;
input n959;
input n960;
input n961;
input n1023;
input n1024;
input n1028;
input n1030;
input n1032;
input n1035;
input n1036;
input n1040;
input n1042;
input n1044;
input n1045;
input n1048;
input n1050;
input n1052;
input n1054;
input n1055;
input n1056;
input n1057;
input n1058;
input n1059;
input n1060;
input n1061;
input n1062;
input n1063;
input n1064;
input n1065;
input n1066;
input n1067;
input n1068;
input n1069;
input n1070;
input n1071;
input n1072;
input n1073;
input n1074;
input n1075;
input n1076;
input n1077;
input n1078;
input n1079;
input n1080;
input n1081;
input n1082;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n22;
wire n23;
wire n24;
wire n26;
wire n28;
wire n31;
wire n32;
wire n34;
wire n36;
wire n38;
wire n68;
wire n69;
wire n72;
wire n73;
wire n74;
wire n76;
wire n78;
wire n82;
wire n83;
wire n84;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n108;
wire n109;
wire n110;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n167;
wire n168;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n287;
wire n288;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1025;
wire n1026;
wire n1027;
wire n1029;
wire n1031;
wire n1033;
wire n1034;
wire n1037;
wire n1038;
wire n1039;
wire n1041;
wire n1043;
wire n1046;
wire n1047;
wire n1049;
wire n1051;
wire n1053;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
xor (out,n0,n1084);
and (n0,n1,n1020);
nor (n1,n2,n1018);
and (n2,n3,n916);
nand (n3,n4,n911);
or (n4,n5,n597);
nand (n5,n6,n545);
not (n6,n7);
nor (n7,n8,n488);
xor (n8,n9,n388);
xor (n9,n10,n312);
xor (n10,n11,n200);
xor (n11,n12,n143);
xor (n12,n13,n97);
nor (n13,n14,n91);
and (n14,n15,n88);
nand (n15,n16,n82);
not (n16,n17);
and (n17,n18,n68);
wire s0n18,s1n18,notn18;
or (n18,s0n18,s1n18);
not(notn18,n31);
and (s0n18,notn18,n19);
and (s1n18,n31,n30);
wire s0n19,s1n19,notn19;
or (n19,s0n19,s1n19);
not(notn19,n22);
and (s0n19,notn19,n20);
and (s1n19,n22,n21);
and (n22,n23,n28);
and (n23,n24,n26);
not (n24,n25);
not (n26,n27);
not (n28,n29);
and (n31,n32,n34);
not (n32,n33);
or (n34,n35,n36);
and (n36,n37,n38);
or (n38,n39,n40,n41,n42,n43,n44,n45,n46,n47,n48,n49,n50,n51,n52,n53,n54,n55,n56,n57,n58,n59,n60,n61,n62,n63,n64,n65,n66,n67);
wire s0n68,s1n68,notn68;
or (n68,s0n68,s1n68);
not(notn68,n81);
and (s0n68,notn68,n69);
and (s1n68,n81,n80);
wire s0n69,s1n69,notn69;
or (n69,s0n69,s1n69);
not(notn69,n72);
and (s0n69,notn69,n70);
and (s1n69,n72,n71);
and (n72,n73,n78);
and (n73,n74,n76);
not (n74,n75);
not (n76,n77);
not (n78,n79);
not (n82,n83);
wire s0n83,s1n83,notn83;
or (n83,s0n83,s1n83);
not(notn83,n81);
and (s0n83,notn83,n84);
and (s1n83,n81,n87);
wire s0n84,s1n84,notn84;
or (n84,s0n84,s1n84);
not(notn84,n72);
and (s0n84,notn84,n85);
and (s1n84,n72,n86);
nand (n88,n89,n90);
not (n89,n18);
not (n90,n68);
not (n91,n92);
wire s0n92,s1n92,notn92;
or (n92,s0n92,s1n92);
not(notn92,n81);
and (s0n92,notn92,n93);
and (s1n92,n81,n96);
wire s0n93,s1n93,notn93;
or (n93,s0n93,s1n93);
not(notn93,n72);
and (s0n93,notn93,n94);
and (s1n93,n72,n95);
nand (n97,n98,n133);
or (n98,n99,n123);
nand (n99,n100,n115);
not (n100,n101);
nand (n101,n102,n114);
or (n102,n103,n108);
wire s0n103,s1n103,notn103;
or (n103,s0n103,s1n103);
not(notn103,n81);
and (s0n103,notn103,n104);
and (s1n103,n81,n107);
wire s0n104,s1n104,notn104;
or (n104,s0n104,s1n104);
not(notn104,n72);
and (s0n104,notn104,n105);
and (s1n104,n72,n106);
not (n108,n109);
wire s0n109,s1n109,notn109;
or (n109,s0n109,s1n109);
not(notn109,n81);
and (s0n109,notn109,n110);
and (s1n109,n81,n113);
wire s0n110,s1n110,notn110;
or (n110,s0n110,s1n110);
not(notn110,n72);
and (s0n110,notn110,n111);
and (s1n110,n72,n112);
nand (n114,n108,n103);
nand (n115,n116,n122);
or (n116,n108,n117);
wire s0n117,s1n117,notn117;
or (n117,s0n117,s1n117);
not(notn117,n81);
and (s0n117,notn117,n118);
and (s1n117,n81,n121);
wire s0n118,s1n118,notn118;
or (n118,s0n118,s1n118);
not(notn118,n72);
and (s0n118,notn118,n119);
and (s1n118,n72,n120);
nand (n122,n117,n108);
not (n123,n124);
nand (n124,n125,n132);
or (n125,n126,n127);
not (n126,n117);
wire s0n127,s1n127,notn127;
or (n127,s0n127,s1n127);
not(notn127,n31);
and (s0n127,notn127,n128);
and (s1n127,n31,n131);
wire s0n128,s1n128,notn128;
or (n128,s0n128,s1n128);
not(notn128,n22);
and (s0n128,notn128,n129);
and (s1n128,n22,n130);
nand (n132,n127,n126);
nand (n133,n134,n101);
nand (n134,n135,n142);
or (n135,n117,n136);
not (n136,n137);
wire s0n137,s1n137,notn137;
or (n137,s0n137,s1n137);
not(notn137,n31);
and (s0n137,notn137,n138);
and (s1n137,n31,n141);
wire s0n138,s1n138,notn138;
or (n138,s0n138,s1n138);
not(notn138,n22);
and (s0n138,notn138,n139);
and (s1n138,n22,n140);
nand (n142,n136,n117);
or (n143,n144,n199);
and (n144,n145,n186);
xor (n145,n146,n150);
nor (n146,n89,n147);
nor (n147,n148,n149);
and (n148,n82,n68);
and (n149,n83,n90);
nand (n150,n151,n176);
or (n151,n152,n157);
not (n152,n153);
nand (n153,n154,n156);
or (n154,n155,n137);
not (n155,n103);
nand (n156,n137,n155);
nand (n157,n158,n173);
not (n158,n159);
nand (n159,n160,n172);
or (n160,n161,n167);
not (n161,n162);
wire s0n162,s1n162,notn162;
or (n162,s0n162,s1n162);
not(notn162,n81);
and (s0n162,notn162,n163);
and (s1n162,n81,n166);
wire s0n163,s1n163,notn163;
or (n163,s0n163,s1n163);
not(notn163,n72);
and (s0n163,notn163,n164);
and (s1n163,n72,n165);
wire s0n167,s1n167,notn167;
or (n167,s0n167,s1n167);
not(notn167,n81);
and (s0n167,notn167,n168);
and (s1n167,n81,n171);
wire s0n168,s1n168,notn168;
or (n168,s0n168,s1n168);
not(notn168,n72);
and (s0n168,notn168,n169);
and (s1n168,n72,n170);
nand (n172,n167,n161);
nand (n173,n174,n175);
or (n174,n155,n162);
nand (n175,n155,n162);
nand (n176,n177,n159);
nand (n177,n178,n185);
or (n178,n103,n179);
not (n179,n180);
wire s0n180,s1n180,notn180;
or (n180,s0n180,s1n180);
not(notn180,n31);
and (s0n180,notn180,n181);
and (s1n180,n31,n184);
wire s0n181,s1n181,notn181;
or (n181,s0n181,s1n181);
not(notn181,n22);
and (s0n181,notn181,n182);
and (s1n181,n22,n183);
nand (n185,n179,n103);
nand (n186,n187,n198);
or (n187,n188,n99);
not (n188,n189);
nand (n189,n190,n197);
or (n190,n117,n191);
not (n191,n192);
wire s0n192,s1n192,notn192;
or (n192,s0n192,s1n192);
not(notn192,n31);
and (s0n192,notn192,n193);
and (s1n192,n31,n196);
wire s0n193,s1n193,notn193;
or (n193,s0n193,s1n193);
not(notn193,n22);
and (s0n193,notn193,n194);
and (s1n193,n22,n195);
nand (n197,n191,n117);
nand (n198,n124,n101);
and (n199,n146,n150);
or (n200,n201,n311);
and (n201,n202,n277);
xor (n202,n203,n242);
nand (n203,n204,n232);
or (n204,n205,n214);
not (n205,n206);
nand (n206,n207,n213);
or (n207,n82,n208);
wire s0n208,s1n208,notn208;
or (n208,s0n208,s1n208);
not(notn208,n31);
and (s0n208,notn208,n209);
and (s1n208,n31,n212);
wire s0n209,s1n209,notn209;
or (n209,s0n209,s1n209);
not(notn209,n22);
and (s0n209,notn209,n210);
and (s1n209,n22,n211);
nand (n213,n82,n208);
nand (n214,n215,n226);
or (n215,n216,n224);
not (n216,n217);
nand (n217,n83,n218);
not (n218,n219);
wire s0n219,s1n219,notn219;
or (n219,s0n219,s1n219);
not(notn219,n81);
and (s0n219,notn219,n220);
and (s1n219,n81,n223);
wire s0n220,s1n220,notn220;
or (n220,s0n220,s1n220);
not(notn220,n72);
and (s0n220,notn220,n221);
and (s1n220,n72,n222);
not (n224,n225);
nand (n225,n82,n219);
xnor (n226,n227,n219);
wire s0n227,s1n227,notn227;
or (n227,s0n227,s1n227);
not(notn227,n81);
and (s0n227,notn227,n228);
and (s1n227,n81,n231);
wire s0n228,s1n228,notn228;
or (n228,s0n228,s1n228);
not(notn228,n72);
and (s0n228,notn228,n229);
and (s1n228,n72,n230);
nand (n232,n233,n241);
nand (n233,n234,n240);
or (n234,n82,n235);
wire s0n235,s1n235,notn235;
or (n235,s0n235,s1n235);
not(notn235,n31);
and (s0n235,notn235,n236);
and (s1n235,n31,n239);
wire s0n236,s1n236,notn236;
or (n236,s0n236,s1n236);
not(notn236,n22);
and (s0n236,notn236,n237);
and (s1n236,n22,n238);
nand (n240,n235,n82);
not (n241,n226);
nand (n242,n243,n264);
or (n243,n244,n254);
not (n244,n245);
nand (n245,n246,n253);
or (n246,n247,n117);
not (n247,n248);
wire s0n248,s1n248,notn248;
or (n248,s0n248,s1n248);
not(notn248,n81);
and (s0n248,notn248,n249);
and (s1n248,n81,n252);
wire s0n249,s1n249,notn249;
or (n249,s0n249,s1n249);
not(notn249,n72);
and (s0n249,notn249,n250);
and (s1n249,n72,n251);
nand (n253,n117,n247);
not (n254,n255);
nand (n255,n256,n263);
or (n256,n257,n258);
not (n257,n227);
wire s0n258,s1n258,notn258;
or (n258,s0n258,s1n258);
not(notn258,n31);
and (s0n258,notn258,n259);
and (s1n258,n31,n262);
wire s0n259,s1n259,notn259;
or (n259,s0n259,s1n259);
not(notn259,n22);
and (s0n259,notn259,n260);
and (s1n259,n22,n261);
nand (n263,n258,n257);
nand (n264,n265,n273);
nand (n265,n266,n272);
or (n266,n257,n267);
wire s0n267,s1n267,notn267;
or (n267,s0n267,s1n267);
not(notn267,n31);
and (s0n267,notn267,n268);
and (s1n267,n31,n271);
wire s0n268,s1n268,notn268;
or (n268,s0n268,s1n268);
not(notn268,n22);
and (s0n268,notn268,n269);
and (s1n268,n22,n270);
nand (n272,n267,n257);
nor (n273,n274,n245);
nor (n274,n275,n276);
and (n275,n257,n248);
and (n276,n227,n247);
nand (n277,n278,n302);
or (n278,n279,n292);
not (n279,n280);
nor (n280,n281,n287);
not (n281,n282);
wire s0n282,s1n282,notn282;
or (n282,s0n282,s1n282);
not(notn282,n81);
and (s0n282,notn282,n283);
and (s1n282,n81,n286);
wire s0n283,s1n283,notn283;
or (n283,s0n283,s1n283);
not(notn283,n72);
and (s0n283,notn283,n284);
and (s1n283,n72,n285);
wire s0n287,s1n287,notn287;
or (n287,s0n287,s1n287);
not(notn287,n81);
and (s0n287,notn287,n288);
and (s1n287,n81,n291);
wire s0n288,s1n288,notn288;
or (n288,s0n288,s1n288);
not(notn288,n72);
and (s0n288,notn288,n289);
and (s1n288,n72,n290);
not (n292,n293);
nand (n293,n294,n301);
or (n294,n282,n295);
not (n295,n296);
wire s0n296,s1n296,notn296;
or (n296,s0n296,s1n296);
not(notn296,n31);
and (s0n296,notn296,n297);
and (s1n296,n31,n300);
wire s0n297,s1n297,notn297;
or (n297,s0n297,s1n297);
not(notn297,n22);
and (s0n297,notn297,n298);
and (s1n297,n22,n299);
nand (n301,n295,n282);
nand (n302,n303,n287);
nand (n303,n304,n310);
or (n304,n281,n305);
wire s0n305,s1n305,notn305;
or (n305,s0n305,s1n305);
not(notn305,n31);
and (s0n305,notn305,n306);
and (s1n305,n31,n309);
wire s0n306,s1n306,notn306;
or (n306,s0n306,s1n306);
not(notn306,n22);
and (s0n306,notn306,n307);
and (s1n306,n22,n308);
nand (n310,n305,n281);
and (n311,n203,n242);
or (n312,n313,n387);
and (n313,n314,n317);
xor (n314,n315,n316);
xor (n315,n202,n277);
xor (n316,n145,n186);
or (n317,n318,n386);
and (n318,n319,n365);
xor (n319,n320,n352);
nand (n320,n321,n343);
or (n321,n322,n327);
not (n322,n323);
nand (n323,n324,n326);
or (n324,n325,n180);
not (n325,n167);
nand (n326,n180,n325);
nand (n327,n328,n339);
or (n328,n329,n337);
not (n329,n330);
nand (n330,n167,n331);
not (n331,n332);
wire s0n332,s1n332,notn332;
or (n332,s0n332,s1n332);
not(notn332,n81);
and (s0n332,notn332,n333);
and (s1n332,n81,n336);
wire s0n333,s1n333,notn333;
or (n333,s0n333,s1n333);
not(notn333,n72);
and (s0n333,notn333,n334);
and (s1n333,n72,n335);
not (n337,n338);
nand (n338,n325,n332);
not (n339,n340);
nand (n340,n341,n342);
or (n341,n282,n331);
nand (n342,n331,n282);
nand (n343,n340,n344);
nand (n344,n345,n351);
or (n345,n325,n346);
wire s0n346,s1n346,notn346;
or (n346,s0n346,s1n346);
not(notn346,n31);
and (s0n346,notn346,n347);
and (s1n346,n31,n350);
wire s0n347,s1n347,notn347;
or (n347,s0n347,s1n347);
not(notn347,n22);
and (s0n347,notn347,n348);
and (s1n347,n22,n349);
nand (n351,n346,n325);
nand (n352,n353,n364);
or (n353,n354,n279);
not (n354,n355);
nand (n355,n356,n363);
or (n356,n282,n357);
not (n357,n358);
wire s0n358,s1n358,notn358;
or (n358,s0n358,s1n358);
not(notn358,n31);
and (s0n358,notn358,n359);
and (s1n358,n31,n362);
wire s0n359,s1n359,notn359;
or (n359,s0n359,s1n359);
not(notn359,n22);
and (s0n359,notn359,n360);
and (s1n359,n22,n361);
nand (n363,n357,n282);
nand (n364,n293,n287);
nand (n365,n366,n385);
or (n366,n367,n376);
not (n367,n368);
nand (n368,n369,n83);
or (n369,n370,n372);
not (n370,n371);
nand (n371,n89,n218);
not (n372,n373);
nand (n373,n374,n257);
not (n374,n375);
and (n375,n18,n219);
not (n376,n377);
nand (n377,n378,n384);
or (n378,n379,n157);
not (n379,n380);
nand (n380,n381,n383);
or (n381,n103,n382);
not (n382,n127);
nand (n383,n382,n103);
nand (n384,n153,n159);
or (n385,n368,n377);
and (n386,n320,n352);
and (n387,n315,n316);
xor (n388,n389,n454);
xor (n389,n390,n425);
xor (n390,n391,n415);
xor (n391,n392,n399);
nand (n392,n393,n395);
or (n393,n394,n214);
not (n394,n233);
nand (n395,n241,n396);
nand (n396,n397,n398);
or (n397,n82,n267);
nand (n398,n267,n82);
nand (n399,n400,n410);
or (n400,n401,n404);
nor (n401,n402,n403);
and (n402,n92,n89);
and (n403,n91,n18);
nand (n404,n405,n147);
or (n405,n406,n408);
not (n406,n407);
nand (n407,n92,n90);
not (n408,n409);
nand (n409,n91,n68);
nand (n410,n411,n414);
nand (n411,n412,n413);
or (n412,n91,n208);
nand (n413,n208,n91);
not (n414,n147);
nand (n415,n416,n421);
or (n416,n417,n327);
not (n417,n418);
nand (n418,n419,n420);
or (n419,n325,n358);
nand (n420,n358,n325);
nand (n421,n422,n340);
nand (n422,n423,n424);
or (n423,n325,n296);
nand (n424,n296,n325);
xor (n425,n426,n447);
xor (n426,n427,n439);
nand (n427,n428,n430);
or (n428,n429,n279);
not (n429,n303);
nand (n430,n431,n287);
nand (n431,n432,n438);
or (n432,n281,n433);
wire s0n433,s1n433,notn433;
or (n433,s0n433,s1n433);
not(notn433,n31);
and (s0n433,notn433,n434);
and (s1n433,n31,n437);
wire s0n434,s1n434,notn434;
or (n434,s0n434,s1n434);
not(notn434,n22);
and (s0n434,notn434,n435);
and (s1n434,n22,n436);
nand (n438,n433,n281);
nand (n439,n440,n442);
nand (n440,n441,n177);
not (n441,n157);
nand (n442,n159,n443);
nand (n443,n444,n446);
or (n444,n103,n445);
not (n445,n346);
nand (n446,n445,n103);
nand (n447,n448,n450);
or (n448,n449,n254);
not (n449,n273);
nand (n450,n451,n245);
nand (n451,n452,n453);
or (n452,n257,n192);
nand (n453,n192,n257);
or (n454,n455,n487);
and (n455,n456,n462);
xor (n456,n457,n461);
nand (n457,n458,n460);
or (n458,n459,n327);
not (n459,n344);
nand (n460,n418,n340);
nor (n461,n376,n368);
or (n462,n463,n486);
and (n463,n464,n479);
xor (n464,n465,n472);
nand (n465,n466,n467);
or (n466,n100,n188);
nand (n467,n468,n471);
nand (n468,n469,n470);
or (n469,n126,n258);
nand (n470,n258,n126);
not (n471,n99);
nand (n472,n473,n478);
or (n473,n474,n214);
not (n474,n475);
nor (n475,n476,n477);
and (n476,n82,n89);
and (n477,n18,n83);
nand (n478,n206,n241);
nand (n479,n480,n482);
or (n480,n244,n481);
not (n481,n265);
nand (n482,n483,n273);
nand (n483,n484,n485);
or (n484,n257,n235);
nand (n485,n235,n257);
and (n486,n465,n472);
and (n487,n457,n461);
or (n488,n489,n544);
and (n489,n490,n543);
xor (n490,n491,n492);
xor (n491,n456,n462);
or (n492,n493,n542);
and (n493,n494,n541);
xor (n494,n495,n522);
or (n495,n496,n521);
and (n496,n497,n514);
xor (n497,n498,n506);
nand (n498,n499,n505);
or (n499,n500,n449);
not (n500,n501);
nand (n501,n502,n504);
or (n502,n227,n503);
not (n503,n208);
nand (n504,n503,n227);
nand (n505,n483,n245);
nand (n506,n507,n509);
or (n507,n100,n508);
not (n508,n468);
nand (n509,n471,n510);
nand (n510,n511,n513);
or (n511,n117,n512);
not (n512,n267);
nand (n513,n512,n117);
nand (n514,n515,n520);
or (n515,n516,n327);
not (n516,n517);
nor (n517,n518,n519);
and (n518,n137,n167);
and (n519,n325,n136);
nand (n520,n323,n340);
and (n521,n498,n506);
or (n522,n523,n540);
and (n523,n524,n533);
xor (n524,n525,n526);
nor (n525,n89,n226);
nand (n526,n527,n532);
or (n527,n157,n528);
not (n528,n529);
nand (n529,n530,n531);
or (n530,n103,n191);
nand (n531,n191,n103);
nand (n532,n380,n159);
nand (n533,n534,n539);
or (n534,n535,n279);
not (n535,n536);
nand (n536,n537,n538);
or (n537,n282,n445);
nand (n538,n445,n282);
nand (n539,n355,n287);
and (n540,n525,n526);
xor (n541,n464,n479);
and (n542,n495,n522);
xor (n543,n314,n317);
and (n544,n491,n492);
or (n545,n546,n547);
xor (n546,n490,n543);
or (n547,n548,n596);
and (n548,n549,n552);
xor (n549,n550,n551);
xor (n550,n319,n365);
xor (n551,n494,n541);
or (n552,n553,n595);
and (n553,n554,n594);
xor (n554,n555,n569);
and (n555,n556,n562);
nor (n556,n557,n257);
and (n557,n558,n561);
nand (n558,n559,n126);
not (n559,n560);
and (n560,n18,n248);
nand (n561,n89,n247);
nand (n562,n563,n568);
or (n563,n157,n564);
not (n564,n565);
nand (n565,n566,n567);
or (n566,n155,n258);
nand (n567,n258,n155);
nand (n568,n529,n159);
or (n569,n570,n593);
and (n570,n571,n586);
xor (n571,n572,n579);
nand (n572,n573,n578);
or (n573,n279,n574);
not (n574,n575);
nand (n575,n576,n577);
or (n576,n282,n179);
nand (n577,n179,n282);
nand (n578,n536,n287);
nand (n579,n580,n585);
or (n580,n581,n327);
not (n581,n582);
nand (n582,n583,n584);
or (n583,n325,n127);
nand (n584,n127,n325);
nand (n585,n517,n340);
nand (n586,n587,n592);
or (n587,n588,n99);
not (n588,n589);
nand (n589,n590,n591);
or (n590,n126,n235);
nand (n591,n235,n126);
nand (n592,n510,n101);
and (n593,n572,n579);
xor (n594,n524,n533);
and (n595,n555,n569);
and (n596,n550,n551);
not (n597,n598);
nand (n598,n599,n895,n901);
nand (n599,n600,n641,n748);
nand (n600,n601,n603);
not (n601,n602);
xor (n602,n549,n552);
not (n603,n604);
or (n604,n605,n640);
and (n605,n606,n639);
xor (n606,n607,n608);
xor (n607,n497,n514);
or (n608,n609,n638);
and (n609,n610,n619);
xor (n610,n611,n618);
nand (n611,n612,n617);
or (n612,n449,n613);
not (n613,n614);
nor (n614,n615,n616);
and (n615,n18,n227);
and (n616,n257,n89);
nand (n617,n245,n501);
xor (n618,n556,n562);
or (n619,n620,n637);
and (n620,n621,n630);
xor (n621,n622,n623);
and (n622,n245,n18);
nand (n623,n624,n629);
or (n624,n327,n625);
not (n625,n626);
nand (n626,n627,n628);
or (n627,n167,n191);
nand (n628,n191,n167);
nand (n629,n582,n340);
nand (n630,n631,n636);
or (n631,n279,n632);
not (n632,n633);
nor (n633,n634,n635);
and (n634,n137,n282);
and (n635,n281,n136);
nand (n636,n575,n287);
and (n637,n622,n623);
and (n638,n611,n618);
xor (n639,n554,n594);
and (n640,n607,n608);
not (n641,n642);
nand (n642,n643,n741);
nor (n643,n644,n711);
nor (n644,n645,n681);
xor (n645,n646,n680);
xor (n646,n647,n648);
xor (n647,n571,n586);
or (n648,n649,n679);
and (n649,n650,n665);
xor (n650,n651,n658);
nand (n651,n652,n657);
or (n652,n653,n99);
not (n653,n654);
nand (n654,n655,n656);
or (n655,n126,n208);
nand (n656,n208,n126);
nand (n657,n589,n101);
nand (n658,n659,n664);
or (n659,n660,n157);
not (n660,n661);
nand (n661,n662,n663);
or (n662,n155,n267);
nand (n663,n267,n155);
nand (n664,n565,n159);
and (n665,n666,n673);
nand (n666,n667,n672);
or (n667,n668,n327);
not (n668,n669);
nand (n669,n670,n671);
or (n670,n325,n258);
nand (n671,n258,n325);
nand (n672,n626,n340);
nor (n673,n674,n126);
and (n674,n675,n678);
nand (n675,n676,n155);
not (n676,n677);
and (n677,n18,n109);
nand (n678,n89,n108);
and (n679,n651,n658);
xor (n680,n610,n619);
or (n681,n682,n710);
and (n682,n683,n709);
xor (n683,n684,n708);
or (n684,n685,n707);
and (n685,n686,n700);
xor (n686,n687,n693);
nand (n687,n688,n692);
nand (n688,n689,n280);
nand (n689,n690,n691);
or (n690,n281,n127);
nand (n691,n127,n281);
nand (n692,n633,n287);
nand (n693,n694,n699);
or (n694,n695,n99);
not (n695,n696);
nand (n696,n697,n698);
or (n697,n117,n89);
or (n698,n18,n126);
nand (n699,n654,n101);
nand (n700,n701,n706);
or (n701,n702,n157);
not (n702,n703);
nand (n703,n704,n705);
or (n704,n155,n235);
nand (n705,n235,n155);
nand (n706,n661,n159);
and (n707,n687,n693);
xor (n708,n621,n630);
xor (n709,n650,n665);
and (n710,n684,n708);
nor (n711,n712,n713);
xor (n712,n683,n709);
or (n713,n714,n740);
and (n714,n715,n739);
xor (n715,n716,n720);
nand (n716,n717,n719);
or (n717,n673,n718);
not (n718,n666);
nand (n719,n718,n673);
or (n720,n721,n738);
and (n721,n722,n731);
xor (n722,n723,n724);
nor (n723,n89,n100);
nand (n724,n725,n730);
or (n725,n726,n327);
not (n726,n727);
nand (n727,n728,n729);
or (n728,n167,n512);
nand (n729,n512,n167);
nand (n730,n669,n340);
nand (n731,n732,n737);
or (n732,n733,n157);
not (n733,n734);
nand (n734,n735,n736);
or (n735,n155,n208);
nand (n736,n208,n155);
nand (n737,n703,n159);
and (n738,n723,n724);
xor (n739,n686,n700);
and (n740,n716,n720);
nand (n741,n742,n744);
not (n742,n743);
xor (n743,n606,n639);
not (n744,n745);
or (n745,n746,n747);
and (n746,n646,n680);
and (n747,n647,n648);
nand (n748,n749,n894);
or (n749,n750,n781);
not (n750,n751);
nand (n751,n752,n754);
not (n752,n753);
xor (n753,n715,n739);
not (n754,n755);
or (n755,n756,n780);
and (n756,n757,n779);
xor (n757,n758,n765);
nand (n758,n759,n764);
or (n759,n279,n760);
not (n760,n761);
nand (n761,n762,n763);
or (n762,n282,n191);
nand (n763,n282,n191);
nand (n764,n689,n287);
and (n765,n766,n773);
nand (n766,n767,n768);
or (n767,n339,n726);
nand (n768,n769,n770);
not (n769,n327);
nand (n770,n771,n772);
or (n771,n325,n235);
nand (n772,n235,n325);
nor (n773,n774,n155);
and (n774,n775,n778);
nand (n775,n776,n325);
not (n776,n777);
and (n777,n18,n162);
nand (n778,n89,n161);
xor (n779,n722,n731);
and (n780,n758,n765);
not (n781,n782);
nand (n782,n783,n893);
or (n783,n784,n812);
not (n784,n785);
nand (n785,n786,n788);
not (n786,n787);
xor (n787,n757,n779);
not (n788,n789);
or (n789,n790,n811);
and (n790,n791,n807);
xor (n791,n792,n799);
nand (n792,n793,n798);
or (n793,n794,n157);
not (n794,n795);
nor (n795,n796,n797);
and (n796,n155,n89);
and (n797,n18,n103);
nand (n798,n159,n734);
nand (n799,n800,n802);
or (n800,n801,n760);
not (n801,n287);
nand (n802,n803,n280);
nand (n803,n804,n806);
or (n804,n282,n805);
not (n805,n258);
nand (n806,n282,n805);
nand (n807,n808,n810);
or (n808,n773,n809);
not (n809,n766);
nand (n810,n809,n773);
and (n811,n792,n799);
not (n812,n813);
nand (n813,n814,n892);
or (n814,n815,n887);
nor (n815,n816,n886);
and (n816,n817,n853);
nand (n817,n818,n836);
not (n818,n819);
xor (n819,n820,n829);
xor (n820,n821,n822);
and (n821,n159,n18);
nand (n822,n823,n825);
or (n823,n801,n824);
not (n824,n803);
nand (n825,n826,n280);
nand (n826,n827,n828);
or (n827,n282,n512);
nand (n828,n512,n282);
nand (n829,n830,n835);
or (n830,n831,n327);
not (n831,n832);
nand (n832,n833,n834);
or (n833,n325,n208);
nand (n834,n208,n325);
nand (n835,n770,n340);
nand (n836,n837,n846);
not (n837,n838);
nand (n838,n839,n167);
or (n839,n840,n842);
not (n840,n841);
nand (n841,n331,n89);
not (n842,n843);
nand (n843,n844,n281);
not (n844,n845);
and (n845,n18,n332);
nand (n846,n847,n849);
or (n847,n801,n848);
not (n848,n826);
nand (n849,n850,n280);
nand (n850,n851,n852);
or (n851,n281,n235);
nand (n852,n235,n281);
nand (n853,n854,n885);
nand (n854,n855,n866);
or (n855,n856,n859);
nand (n856,n857,n858);
or (n857,n838,n846);
nand (n858,n846,n838);
nand (n859,n860,n865);
or (n860,n861,n327);
not (n861,n862);
nor (n862,n863,n864);
and (n863,n325,n89);
and (n864,n18,n167);
nand (n865,n340,n832);
or (n866,n867,n884);
and (n867,n868,n877);
xor (n868,n869,n870);
and (n869,n18,n340);
nand (n870,n871,n873);
or (n871,n801,n872);
not (n872,n850);
nand (n873,n874,n280);
nand (n874,n875,n876);
or (n875,n281,n208);
nand (n876,n208,n281);
nor (n877,n878,n881);
nor (n878,n879,n880);
and (n879,n280,n89);
and (n880,n874,n287);
nand (n881,n882,n282);
not (n882,n883);
and (n883,n18,n287);
and (n884,n869,n870);
nand (n885,n856,n859);
nor (n886,n818,n836);
nor (n887,n888,n889);
xor (n888,n791,n807);
or (n889,n890,n891);
and (n890,n820,n829);
and (n891,n821,n822);
nand (n892,n888,n889);
nand (n893,n787,n789);
nand (n894,n753,n755);
nand (n895,n896,n600);
or (n896,n897,n899);
not (n897,n898);
nand (n898,n743,n745);
not (n899,n900);
nand (n900,n602,n604);
nand (n901,n600,n902);
nor (n902,n903,n910);
nand (n903,n904,n909);
or (n904,n905,n907);
not (n905,n906);
nand (n906,n712,n713);
not (n907,n908);
nand (n908,n645,n681);
not (n909,n644);
not (n910,n741);
not (n911,n912);
nand (n912,n913,n915);
or (n913,n7,n914);
nand (n914,n546,n547);
nand (n915,n8,n488);
not (n916,n917);
nand (n917,n918,n1016);
not (n918,n919);
nor (n919,n920,n1012);
not (n920,n921);
xor (n921,n922,n1009);
xor (n922,n923,n963);
xor (n923,n924,n931);
xor (n924,n925,n928);
or (n925,n926,n927);
and (n926,n391,n415);
and (n927,n392,n399);
or (n928,n929,n930);
and (n929,n426,n447);
and (n930,n427,n439);
xor (n931,n932,n950);
xor (n932,n933,n943);
and (n933,n934,n18);
nand (n934,n935,n942);
or (n935,n936,n92);
not (n936,n937);
wire s0n937,s1n937,notn937;
or (n937,s0n937,s1n937);
not(notn937,n81);
and (s0n937,notn937,n938);
and (s1n937,n81,n941);
wire s0n938,s1n938,notn938;
or (n938,s0n938,s1n938);
not(notn938,n72);
and (s0n938,notn938,n939);
and (s1n938,n72,n940);
nand (n942,n92,n936);
nand (n943,n944,n946);
or (n944,n945,n99);
not (n945,n134);
nand (n946,n947,n101);
nand (n947,n948,n949);
or (n948,n126,n180);
nand (n949,n180,n126);
nand (n950,n951,n953);
or (n951,n952,n279);
not (n952,n431);
nand (n953,n954,n287);
nor (n954,n955,n962);
and (n955,n281,n956);
not (n956,n957);
wire s0n957,s1n957,notn957;
or (n957,s0n957,s1n957);
not(notn957,n31);
and (s0n957,notn957,n958);
and (s1n957,n31,n961);
wire s0n958,s1n958,notn958;
or (n958,s0n958,s1n958);
not(notn958,n22);
and (s0n958,notn958,n959);
and (s1n958,n22,n960);
and (n962,n957,n282);
xor (n963,n964,n1006);
xor (n964,n965,n988);
xor (n965,n966,n981);
xor (n966,n967,n974);
nand (n967,n968,n970);
or (n968,n969,n157);
not (n969,n443);
nand (n970,n971,n159);
nand (n971,n972,n973);
or (n972,n103,n357);
nand (n973,n357,n103);
nand (n974,n975,n977);
or (n975,n449,n976);
not (n976,n451);
nand (n977,n978,n245);
nand (n978,n979,n980);
or (n979,n257,n127);
nand (n980,n127,n257);
nand (n981,n982,n984);
or (n982,n214,n983);
not (n983,n396);
nand (n984,n985,n241);
nand (n985,n986,n987);
or (n986,n82,n258);
nand (n987,n258,n82);
xor (n988,n989,n1005);
xor (n989,n990,n997);
nand (n990,n991,n993);
or (n991,n992,n404);
not (n992,n411);
nand (n993,n994,n414);
nand (n994,n995,n996);
or (n995,n91,n235);
nand (n996,n235,n91);
nand (n997,n998,n1000);
or (n998,n999,n327);
not (n999,n422);
nand (n1000,n1001,n340);
nand (n1001,n1002,n1004);
or (n1002,n167,n1003);
not (n1003,n305);
nand (n1004,n1003,n167);
and (n1005,n13,n97);
or (n1006,n1007,n1008);
and (n1007,n11,n200);
and (n1008,n12,n143);
or (n1009,n1010,n1011);
and (n1010,n389,n454);
and (n1011,n390,n425);
not (n1012,n1013);
or (n1013,n1014,n1015);
and (n1014,n9,n388);
and (n1015,n10,n312);
not (n1016,n1017);
nor (n1017,n921,n1013);
and (n1018,n1019,n917);
not (n1019,n3);
xor (n1020,n1021,n1083);
and (n1021,n1022,n1033);
wire s0n1022,s1n1022,notn1022;
or (n1022,s0n1022,s1n1022);
not(notn1022,n1025);
and (s0n1022,notn1022,n1023);
and (s1n1022,n1025,n1024);
and (n1025,n1026,n1031);
and (n1026,n1027,n1029);
not (n1027,n1028);
not (n1029,n1030);
not (n1031,n1032);
wire s0n1033,s1n1033,notn1033;
or (n1033,s0n1033,s1n1033);
not(notn1033,n1046);
and (s0n1033,notn1033,n1034);
and (s1n1033,n1046,n1045);
wire s0n1034,s1n1034,notn1034;
or (n1034,s0n1034,s1n1034);
not(notn1034,n1037);
and (s0n1034,notn1034,n1035);
and (s1n1034,n1037,n1036);
and (n1037,n1038,n1043);
and (n1038,n1039,n1041);
not (n1039,n1040);
not (n1041,n1042);
not (n1043,n1044);
and (n1046,n1047,n1049);
not (n1047,n1048);
or (n1049,n1050,n1051);
and (n1051,n1052,n1053);
or (n1053,n1054,n1055,n1056,n1057,n1058,n1059,n1060,n1061,n1062,n1063,n1064,n1065,n1066,n1067,n1068,n1069,n1070,n1071,n1072,n1073,n1074,n1075,n1076,n1077,n1078,n1079,n1080,n1081,n1082);
and (n1083,n288,n18);
and (n1084,n1020,n1085);
xor (n1085,n1086,n1621);
xor (n1086,n1087,n1618);
xor (n1087,n1088,n1617);
xor (n1088,n1089,n1609);
xor (n1089,n1090,n1608);
xor (n1090,n1091,n1594);
xor (n1091,n1092,n1593);
xor (n1092,n1093,n1573);
xor (n1093,n1094,n1572);
xor (n1094,n1095,n1546);
xor (n1095,n1096,n1545);
xor (n1096,n1097,n1513);
xor (n1097,n1098,n1512);
xor (n1098,n1099,n1473);
xor (n1099,n1100,n1472);
xor (n1100,n1101,n1428);
xor (n1101,n1102,n1427);
xor (n1102,n1103,n1377);
xor (n1103,n1104,n1376);
xor (n1104,n1105,n1320);
xor (n1105,n1106,n1319);
xor (n1106,n1107,n1258);
xor (n1107,n1108,n1257);
xor (n1108,n1109,n1189);
xor (n1109,n1110,n1188);
xor (n1110,n1111,n1114);
xor (n1111,n1112,n1113);
and (n1112,n957,n287);
and (n1113,n433,n282);
or (n1114,n1115,n1118);
and (n1115,n1116,n1117);
and (n1116,n433,n287);
and (n1117,n305,n282);
and (n1118,n1119,n1120);
xor (n1119,n1116,n1117);
or (n1120,n1121,n1124);
and (n1121,n1122,n1123);
and (n1122,n305,n287);
and (n1123,n296,n282);
and (n1124,n1125,n1126);
xor (n1125,n1122,n1123);
or (n1126,n1127,n1130);
and (n1127,n1128,n1129);
and (n1128,n296,n287);
and (n1129,n358,n282);
and (n1130,n1131,n1132);
xor (n1131,n1128,n1129);
or (n1132,n1133,n1136);
and (n1133,n1134,n1135);
and (n1134,n358,n287);
and (n1135,n346,n282);
and (n1136,n1137,n1138);
xor (n1137,n1134,n1135);
or (n1138,n1139,n1142);
and (n1139,n1140,n1141);
and (n1140,n346,n287);
and (n1141,n180,n282);
and (n1142,n1143,n1144);
xor (n1143,n1140,n1141);
or (n1144,n1145,n1147);
and (n1145,n1146,n634);
and (n1146,n180,n287);
and (n1147,n1148,n1149);
xor (n1148,n1146,n634);
or (n1149,n1150,n1153);
and (n1150,n1151,n1152);
and (n1151,n137,n287);
and (n1152,n127,n282);
and (n1153,n1154,n1155);
xor (n1154,n1151,n1152);
or (n1155,n1156,n1159);
and (n1156,n1157,n1158);
and (n1157,n127,n287);
and (n1158,n192,n282);
and (n1159,n1160,n1161);
xor (n1160,n1157,n1158);
or (n1161,n1162,n1165);
and (n1162,n1163,n1164);
and (n1163,n192,n287);
and (n1164,n258,n282);
and (n1165,n1166,n1167);
xor (n1166,n1163,n1164);
or (n1167,n1168,n1171);
and (n1168,n1169,n1170);
and (n1169,n258,n287);
and (n1170,n267,n282);
and (n1171,n1172,n1173);
xor (n1172,n1169,n1170);
or (n1173,n1174,n1177);
and (n1174,n1175,n1176);
and (n1175,n267,n287);
and (n1176,n235,n282);
and (n1177,n1178,n1179);
xor (n1178,n1175,n1176);
or (n1179,n1180,n1183);
and (n1180,n1181,n1182);
and (n1181,n235,n287);
and (n1182,n208,n282);
and (n1183,n1184,n1185);
xor (n1184,n1181,n1182);
and (n1185,n1186,n1187);
and (n1186,n208,n287);
and (n1187,n18,n282);
and (n1188,n305,n332);
or (n1189,n1190,n1193);
and (n1190,n1191,n1192);
xor (n1191,n1119,n1120);
and (n1192,n296,n332);
and (n1193,n1194,n1195);
xor (n1194,n1191,n1192);
or (n1195,n1196,n1199);
and (n1196,n1197,n1198);
xor (n1197,n1125,n1126);
and (n1198,n358,n332);
and (n1199,n1200,n1201);
xor (n1200,n1197,n1198);
or (n1201,n1202,n1205);
and (n1202,n1203,n1204);
xor (n1203,n1131,n1132);
and (n1204,n346,n332);
and (n1205,n1206,n1207);
xor (n1206,n1203,n1204);
or (n1207,n1208,n1211);
and (n1208,n1209,n1210);
xor (n1209,n1137,n1138);
and (n1210,n180,n332);
and (n1211,n1212,n1213);
xor (n1212,n1209,n1210);
or (n1213,n1214,n1217);
and (n1214,n1215,n1216);
xor (n1215,n1143,n1144);
and (n1216,n137,n332);
and (n1217,n1218,n1219);
xor (n1218,n1215,n1216);
or (n1219,n1220,n1223);
and (n1220,n1221,n1222);
xor (n1221,n1148,n1149);
and (n1222,n127,n332);
and (n1223,n1224,n1225);
xor (n1224,n1221,n1222);
or (n1225,n1226,n1229);
and (n1226,n1227,n1228);
xor (n1227,n1154,n1155);
and (n1228,n192,n332);
and (n1229,n1230,n1231);
xor (n1230,n1227,n1228);
or (n1231,n1232,n1235);
and (n1232,n1233,n1234);
xor (n1233,n1160,n1161);
and (n1234,n258,n332);
and (n1235,n1236,n1237);
xor (n1236,n1233,n1234);
or (n1237,n1238,n1241);
and (n1238,n1239,n1240);
xor (n1239,n1166,n1167);
and (n1240,n267,n332);
and (n1241,n1242,n1243);
xor (n1242,n1239,n1240);
or (n1243,n1244,n1247);
and (n1244,n1245,n1246);
xor (n1245,n1172,n1173);
and (n1246,n235,n332);
and (n1247,n1248,n1249);
xor (n1248,n1245,n1246);
or (n1249,n1250,n1253);
and (n1250,n1251,n1252);
xor (n1251,n1178,n1179);
and (n1252,n208,n332);
and (n1253,n1254,n1255);
xor (n1254,n1251,n1252);
and (n1255,n1256,n845);
xor (n1256,n1184,n1185);
and (n1257,n296,n167);
or (n1258,n1259,n1262);
and (n1259,n1260,n1261);
xor (n1260,n1194,n1195);
and (n1261,n358,n167);
and (n1262,n1263,n1264);
xor (n1263,n1260,n1261);
or (n1264,n1265,n1268);
and (n1265,n1266,n1267);
xor (n1266,n1200,n1201);
and (n1267,n346,n167);
and (n1268,n1269,n1270);
xor (n1269,n1266,n1267);
or (n1270,n1271,n1274);
and (n1271,n1272,n1273);
xor (n1272,n1206,n1207);
and (n1273,n180,n167);
and (n1274,n1275,n1276);
xor (n1275,n1272,n1273);
or (n1276,n1277,n1279);
and (n1277,n1278,n518);
xor (n1278,n1212,n1213);
and (n1279,n1280,n1281);
xor (n1280,n1278,n518);
or (n1281,n1282,n1285);
and (n1282,n1283,n1284);
xor (n1283,n1218,n1219);
and (n1284,n127,n167);
and (n1285,n1286,n1287);
xor (n1286,n1283,n1284);
or (n1287,n1288,n1291);
and (n1288,n1289,n1290);
xor (n1289,n1224,n1225);
and (n1290,n192,n167);
and (n1291,n1292,n1293);
xor (n1292,n1289,n1290);
or (n1293,n1294,n1297);
and (n1294,n1295,n1296);
xor (n1295,n1230,n1231);
and (n1296,n258,n167);
and (n1297,n1298,n1299);
xor (n1298,n1295,n1296);
or (n1299,n1300,n1303);
and (n1300,n1301,n1302);
xor (n1301,n1236,n1237);
and (n1302,n267,n167);
and (n1303,n1304,n1305);
xor (n1304,n1301,n1302);
or (n1305,n1306,n1309);
and (n1306,n1307,n1308);
xor (n1307,n1242,n1243);
and (n1308,n235,n167);
and (n1309,n1310,n1311);
xor (n1310,n1307,n1308);
or (n1311,n1312,n1315);
and (n1312,n1313,n1314);
xor (n1313,n1248,n1249);
and (n1314,n208,n167);
and (n1315,n1316,n1317);
xor (n1316,n1313,n1314);
and (n1317,n1318,n864);
xor (n1318,n1254,n1255);
and (n1319,n358,n162);
or (n1320,n1321,n1324);
and (n1321,n1322,n1323);
xor (n1322,n1263,n1264);
and (n1323,n346,n162);
and (n1324,n1325,n1326);
xor (n1325,n1322,n1323);
or (n1326,n1327,n1330);
and (n1327,n1328,n1329);
xor (n1328,n1269,n1270);
and (n1329,n180,n162);
and (n1330,n1331,n1332);
xor (n1331,n1328,n1329);
or (n1332,n1333,n1336);
and (n1333,n1334,n1335);
xor (n1334,n1275,n1276);
and (n1335,n137,n162);
and (n1336,n1337,n1338);
xor (n1337,n1334,n1335);
or (n1338,n1339,n1342);
and (n1339,n1340,n1341);
xor (n1340,n1280,n1281);
and (n1341,n127,n162);
and (n1342,n1343,n1344);
xor (n1343,n1340,n1341);
or (n1344,n1345,n1348);
and (n1345,n1346,n1347);
xor (n1346,n1286,n1287);
and (n1347,n192,n162);
and (n1348,n1349,n1350);
xor (n1349,n1346,n1347);
or (n1350,n1351,n1354);
and (n1351,n1352,n1353);
xor (n1352,n1292,n1293);
and (n1353,n258,n162);
and (n1354,n1355,n1356);
xor (n1355,n1352,n1353);
or (n1356,n1357,n1360);
and (n1357,n1358,n1359);
xor (n1358,n1298,n1299);
and (n1359,n267,n162);
and (n1360,n1361,n1362);
xor (n1361,n1358,n1359);
or (n1362,n1363,n1366);
and (n1363,n1364,n1365);
xor (n1364,n1304,n1305);
and (n1365,n235,n162);
and (n1366,n1367,n1368);
xor (n1367,n1364,n1365);
or (n1368,n1369,n1372);
and (n1369,n1370,n1371);
xor (n1370,n1310,n1311);
and (n1371,n208,n162);
and (n1372,n1373,n1374);
xor (n1373,n1370,n1371);
and (n1374,n1375,n777);
xor (n1375,n1316,n1317);
and (n1376,n346,n103);
or (n1377,n1378,n1381);
and (n1378,n1379,n1380);
xor (n1379,n1325,n1326);
and (n1380,n180,n103);
and (n1381,n1382,n1383);
xor (n1382,n1379,n1380);
or (n1383,n1384,n1387);
and (n1384,n1385,n1386);
xor (n1385,n1331,n1332);
and (n1386,n137,n103);
and (n1387,n1388,n1389);
xor (n1388,n1385,n1386);
or (n1389,n1390,n1393);
and (n1390,n1391,n1392);
xor (n1391,n1337,n1338);
and (n1392,n127,n103);
and (n1393,n1394,n1395);
xor (n1394,n1391,n1392);
or (n1395,n1396,n1399);
and (n1396,n1397,n1398);
xor (n1397,n1343,n1344);
and (n1398,n192,n103);
and (n1399,n1400,n1401);
xor (n1400,n1397,n1398);
or (n1401,n1402,n1405);
and (n1402,n1403,n1404);
xor (n1403,n1349,n1350);
and (n1404,n258,n103);
and (n1405,n1406,n1407);
xor (n1406,n1403,n1404);
or (n1407,n1408,n1411);
and (n1408,n1409,n1410);
xor (n1409,n1355,n1356);
and (n1410,n267,n103);
and (n1411,n1412,n1413);
xor (n1412,n1409,n1410);
or (n1413,n1414,n1417);
and (n1414,n1415,n1416);
xor (n1415,n1361,n1362);
and (n1416,n235,n103);
and (n1417,n1418,n1419);
xor (n1418,n1415,n1416);
or (n1419,n1420,n1423);
and (n1420,n1421,n1422);
xor (n1421,n1367,n1368);
and (n1422,n208,n103);
and (n1423,n1424,n1425);
xor (n1424,n1421,n1422);
and (n1425,n1426,n797);
xor (n1426,n1373,n1374);
and (n1427,n180,n109);
or (n1428,n1429,n1432);
and (n1429,n1430,n1431);
xor (n1430,n1382,n1383);
and (n1431,n137,n109);
and (n1432,n1433,n1434);
xor (n1433,n1430,n1431);
or (n1434,n1435,n1438);
and (n1435,n1436,n1437);
xor (n1436,n1388,n1389);
and (n1437,n127,n109);
and (n1438,n1439,n1440);
xor (n1439,n1436,n1437);
or (n1440,n1441,n1444);
and (n1441,n1442,n1443);
xor (n1442,n1394,n1395);
and (n1443,n192,n109);
and (n1444,n1445,n1446);
xor (n1445,n1442,n1443);
or (n1446,n1447,n1450);
and (n1447,n1448,n1449);
xor (n1448,n1400,n1401);
and (n1449,n258,n109);
and (n1450,n1451,n1452);
xor (n1451,n1448,n1449);
or (n1452,n1453,n1456);
and (n1453,n1454,n1455);
xor (n1454,n1406,n1407);
and (n1455,n267,n109);
and (n1456,n1457,n1458);
xor (n1457,n1454,n1455);
or (n1458,n1459,n1462);
and (n1459,n1460,n1461);
xor (n1460,n1412,n1413);
and (n1461,n235,n109);
and (n1462,n1463,n1464);
xor (n1463,n1460,n1461);
or (n1464,n1465,n1468);
and (n1465,n1466,n1467);
xor (n1466,n1418,n1419);
and (n1467,n208,n109);
and (n1468,n1469,n1470);
xor (n1469,n1466,n1467);
and (n1470,n1471,n677);
xor (n1471,n1424,n1425);
and (n1472,n137,n117);
or (n1473,n1474,n1477);
and (n1474,n1475,n1476);
xor (n1475,n1433,n1434);
and (n1476,n127,n117);
and (n1477,n1478,n1479);
xor (n1478,n1475,n1476);
or (n1479,n1480,n1483);
and (n1480,n1481,n1482);
xor (n1481,n1439,n1440);
and (n1482,n192,n117);
and (n1483,n1484,n1485);
xor (n1484,n1481,n1482);
or (n1485,n1486,n1489);
and (n1486,n1487,n1488);
xor (n1487,n1445,n1446);
and (n1488,n258,n117);
and (n1489,n1490,n1491);
xor (n1490,n1487,n1488);
or (n1491,n1492,n1495);
and (n1492,n1493,n1494);
xor (n1493,n1451,n1452);
and (n1494,n267,n117);
and (n1495,n1496,n1497);
xor (n1496,n1493,n1494);
or (n1497,n1498,n1501);
and (n1498,n1499,n1500);
xor (n1499,n1457,n1458);
and (n1500,n235,n117);
and (n1501,n1502,n1503);
xor (n1502,n1499,n1500);
or (n1503,n1504,n1507);
and (n1504,n1505,n1506);
xor (n1505,n1463,n1464);
and (n1506,n208,n117);
and (n1507,n1508,n1509);
xor (n1508,n1505,n1506);
and (n1509,n1510,n1511);
xor (n1510,n1469,n1470);
and (n1511,n18,n117);
and (n1512,n127,n248);
or (n1513,n1514,n1517);
and (n1514,n1515,n1516);
xor (n1515,n1478,n1479);
and (n1516,n192,n248);
and (n1517,n1518,n1519);
xor (n1518,n1515,n1516);
or (n1519,n1520,n1523);
and (n1520,n1521,n1522);
xor (n1521,n1484,n1485);
and (n1522,n258,n248);
and (n1523,n1524,n1525);
xor (n1524,n1521,n1522);
or (n1525,n1526,n1529);
and (n1526,n1527,n1528);
xor (n1527,n1490,n1491);
and (n1528,n267,n248);
and (n1529,n1530,n1531);
xor (n1530,n1527,n1528);
or (n1531,n1532,n1535);
and (n1532,n1533,n1534);
xor (n1533,n1496,n1497);
and (n1534,n235,n248);
and (n1535,n1536,n1537);
xor (n1536,n1533,n1534);
or (n1537,n1538,n1541);
and (n1538,n1539,n1540);
xor (n1539,n1502,n1503);
and (n1540,n208,n248);
and (n1541,n1542,n1543);
xor (n1542,n1539,n1540);
and (n1543,n1544,n560);
xor (n1544,n1508,n1509);
and (n1545,n192,n227);
or (n1546,n1547,n1550);
and (n1547,n1548,n1549);
xor (n1548,n1518,n1519);
and (n1549,n258,n227);
and (n1550,n1551,n1552);
xor (n1551,n1548,n1549);
or (n1552,n1553,n1556);
and (n1553,n1554,n1555);
xor (n1554,n1524,n1525);
and (n1555,n267,n227);
and (n1556,n1557,n1558);
xor (n1557,n1554,n1555);
or (n1558,n1559,n1562);
and (n1559,n1560,n1561);
xor (n1560,n1530,n1531);
and (n1561,n235,n227);
and (n1562,n1563,n1564);
xor (n1563,n1560,n1561);
or (n1564,n1565,n1568);
and (n1565,n1566,n1567);
xor (n1566,n1536,n1537);
and (n1567,n208,n227);
and (n1568,n1569,n1570);
xor (n1569,n1566,n1567);
and (n1570,n1571,n615);
xor (n1571,n1542,n1543);
and (n1572,n258,n219);
or (n1573,n1574,n1577);
and (n1574,n1575,n1576);
xor (n1575,n1551,n1552);
and (n1576,n267,n219);
and (n1577,n1578,n1579);
xor (n1578,n1575,n1576);
or (n1579,n1580,n1583);
and (n1580,n1581,n1582);
xor (n1581,n1557,n1558);
and (n1582,n235,n219);
and (n1583,n1584,n1585);
xor (n1584,n1581,n1582);
or (n1585,n1586,n1589);
and (n1586,n1587,n1588);
xor (n1587,n1563,n1564);
and (n1588,n208,n219);
and (n1589,n1590,n1591);
xor (n1590,n1587,n1588);
and (n1591,n1592,n375);
xor (n1592,n1569,n1570);
and (n1593,n267,n83);
or (n1594,n1595,n1598);
and (n1595,n1596,n1597);
xor (n1596,n1578,n1579);
and (n1597,n235,n83);
and (n1598,n1599,n1600);
xor (n1599,n1596,n1597);
or (n1600,n1601,n1604);
and (n1601,n1602,n1603);
xor (n1602,n1584,n1585);
and (n1603,n208,n83);
and (n1604,n1605,n1606);
xor (n1605,n1602,n1603);
and (n1606,n1607,n477);
xor (n1607,n1590,n1591);
and (n1608,n235,n68);
or (n1609,n1610,n1613);
and (n1610,n1611,n1612);
xor (n1611,n1599,n1600);
and (n1612,n208,n68);
and (n1613,n1614,n1615);
xor (n1614,n1611,n1612);
and (n1615,n1616,n17);
xor (n1616,n1605,n1606);
and (n1617,n208,n92);
and (n1618,n1619,n1620);
xor (n1619,n1614,n1615);
and (n1620,n18,n92);
and (n1621,n18,n937);
endmodule
