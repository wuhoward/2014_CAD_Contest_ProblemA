module top (out,n17,n18,n22,n24,n26,n27,n28,n32,n33
        ,n34,n41,n42,n46,n48,n50,n51,n54,n56,n58
        ,n60,n61,n62,n63,n64,n65,n66,n67,n68,n69
        ,n70,n71,n72,n73,n74,n75,n76,n77,n78,n79
        ,n80,n81,n82,n83,n84,n85,n86,n87,n88,n96
        ,n97,n98,n107,n108,n109,n113,n114,n115,n124,n125
        ,n126,n130,n131,n132,n142,n143,n144,n154,n155,n156
        ,n165,n166,n167,n170,n171,n172,n183,n184,n185,n196
        ,n197,n198,n208,n209,n210,n219,n220,n221,n240,n241
        ,n242,n261,n262,n263,n469,n470,n471,n501,n502,n503
        ,n553,n554,n558,n560,n562,n565,n566,n570,n572,n574
        ,n575,n578,n580,n582,n584,n585,n586,n587,n588,n589
        ,n590,n591,n592,n593,n594,n595,n596,n597,n598,n599
        ,n600,n601,n602,n603,n604,n605,n606,n607,n608,n609
        ,n610,n611,n612,n615,n616,n619,n620,n621,n626,n627
        ,n631,n632,n633);
output out;
input n17;
input n18;
input n22;
input n24;
input n26;
input n27;
input n28;
input n32;
input n33;
input n34;
input n41;
input n42;
input n46;
input n48;
input n50;
input n51;
input n54;
input n56;
input n58;
input n60;
input n61;
input n62;
input n63;
input n64;
input n65;
input n66;
input n67;
input n68;
input n69;
input n70;
input n71;
input n72;
input n73;
input n74;
input n75;
input n76;
input n77;
input n78;
input n79;
input n80;
input n81;
input n82;
input n83;
input n84;
input n85;
input n86;
input n87;
input n88;
input n96;
input n97;
input n98;
input n107;
input n108;
input n109;
input n113;
input n114;
input n115;
input n124;
input n125;
input n126;
input n130;
input n131;
input n132;
input n142;
input n143;
input n144;
input n154;
input n155;
input n156;
input n165;
input n166;
input n167;
input n170;
input n171;
input n172;
input n183;
input n184;
input n185;
input n196;
input n197;
input n198;
input n208;
input n209;
input n210;
input n219;
input n220;
input n221;
input n240;
input n241;
input n242;
input n261;
input n262;
input n263;
input n469;
input n470;
input n471;
input n501;
input n502;
input n503;
input n553;
input n554;
input n558;
input n560;
input n562;
input n565;
input n566;
input n570;
input n572;
input n574;
input n575;
input n578;
input n580;
input n582;
input n584;
input n585;
input n586;
input n587;
input n588;
input n589;
input n590;
input n591;
input n592;
input n593;
input n594;
input n595;
input n596;
input n597;
input n598;
input n599;
input n600;
input n601;
input n602;
input n603;
input n604;
input n605;
input n606;
input n607;
input n608;
input n609;
input n610;
input n611;
input n612;
input n615;
input n616;
input n619;
input n620;
input n621;
input n626;
input n627;
input n631;
input n632;
input n633;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n19;
wire n20;
wire n21;
wire n23;
wire n25;
wire n29;
wire n30;
wire n31;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n43;
wire n44;
wire n45;
wire n47;
wire n49;
wire n52;
wire n53;
wire n55;
wire n57;
wire n59;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n110;
wire n111;
wire n112;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n127;
wire n128;
wire n129;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n168;
wire n169;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n555;
wire n556;
wire n557;
wire n559;
wire n561;
wire n563;
wire n564;
wire n567;
wire n568;
wire n569;
wire n571;
wire n573;
wire n576;
wire n577;
wire n579;
wire n581;
wire n583;
wire n613;
wire n614;
wire n617;
wire n618;
wire n622;
wire n623;
wire n624;
wire n625;
wire n628;
wire n629;
wire n630;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
xnor (out,n0,n647);
nand (n0,n1,n535);
nand (n1,n2,n534);
or (n2,n3,n453);
nand (n3,n4,n452);
or (n4,n5,n308);
nor (n5,n6,n279);
xor (n6,n7,n244);
xor (n7,n8,n188);
or (n8,n9,n187);
and (n9,n10,n146);
xor (n10,n11,n100);
nand (n11,n12,n90);
or (n12,n13,n35);
not (n13,n14);
nor (n14,n15,n29);
wire s0n15,s1n15,notn15;
or (n15,s0n15,s1n15);
not(notn15,n28);
and (s0n15,notn15,n16);
and (s1n15,n28,n27);
wire s0n16,s1n16,notn16;
or (n16,s0n16,s1n16);
not(notn16,n19);
and (s0n16,notn16,n17);
and (s1n16,n19,n18);
and (n19,n20,n25);
and (n20,n21,n23);
not (n21,n22);
not (n23,n24);
not (n25,n26);
not (n29,n30);
wire s0n30,s1n30,notn30;
or (n30,s0n30,s1n30);
not(notn30,n28);
and (s0n30,notn30,n31);
and (s1n30,n28,n34);
wire s0n31,s1n31,notn31;
or (n31,s0n31,s1n31);
not(notn31,n19);
and (s0n31,notn31,n32);
and (s1n31,n19,n33);
not (n35,n36);
nand (n36,n37,n89);
or (n37,n30,n38);
not (n38,n39);
wire s0n39,s1n39,notn39;
or (n39,s0n39,s1n39);
not(notn39,n52);
and (s0n39,notn39,n40);
and (s1n39,n52,n51);
wire s0n40,s1n40,notn40;
or (n40,s0n40,s1n40);
not(notn40,n43);
and (s0n40,notn40,n41);
and (s1n40,n43,n42);
and (n43,n44,n49);
and (n44,n45,n47);
not (n45,n46);
not (n47,n48);
not (n49,n50);
and (n52,n53,n55);
not (n53,n54);
or (n55,n56,n57);
and (n57,n58,n59);
or (n59,n60,n61,n62,n63,n64,n65,n66,n67,n68,n69,n70,n71,n72,n73,n74,n75,n76,n77,n78,n79,n80,n81,n82,n83,n84,n85,n86,n87,n88);
nand (n89,n38,n30);
nand (n90,n91,n15);
nand (n91,n92,n99);
or (n92,n30,n93);
not (n93,n94);
wire s0n94,s1n94,notn94;
or (n94,s0n94,s1n94);
not(notn94,n52);
and (s0n94,notn94,n95);
and (s1n94,n52,n98);
wire s0n95,s1n95,notn95;
or (n95,s0n95,s1n95);
not(notn95,n43);
and (s0n95,notn95,n96);
and (s1n95,n43,n97);
nand (n99,n93,n30);
nand (n100,n101,n137);
or (n101,n102,n118);
not (n102,n103);
nand (n103,n104,n116);
or (n104,n105,n110);
wire s0n105,s1n105,notn105;
or (n105,s0n105,s1n105);
not(notn105,n28);
and (s0n105,notn105,n106);
and (s1n105,n28,n109);
wire s0n106,s1n106,notn106;
or (n106,s0n106,s1n106);
not(notn106,n19);
and (s0n106,notn106,n107);
and (s1n106,n19,n108);
not (n110,n111);
wire s0n111,s1n111,notn111;
or (n111,s0n111,s1n111);
not(notn111,n52);
and (s0n111,notn111,n112);
and (s1n111,n52,n115);
wire s0n112,s1n112,notn112;
or (n112,s0n112,s1n112);
not(notn112,n43);
and (s0n112,notn112,n113);
and (s1n112,n43,n114);
or (n116,n111,n117);
not (n117,n105);
nand (n118,n119,n134);
not (n119,n120);
nand (n120,n121,n133);
or (n121,n122,n127);
wire s0n122,s1n122,notn122;
or (n122,s0n122,s1n122);
not(notn122,n28);
and (s0n122,notn122,n123);
and (s1n122,n28,n126);
wire s0n123,s1n123,notn123;
or (n123,s0n123,s1n123);
not(notn123,n19);
and (s0n123,notn123,n124);
and (s1n123,n19,n125);
not (n127,n128);
wire s0n128,s1n128,notn128;
or (n128,s0n128,s1n128);
not(notn128,n28);
and (s0n128,notn128,n129);
and (s1n128,n28,n132);
wire s0n129,s1n129,notn129;
or (n129,s0n129,s1n129);
not(notn129,n19);
and (s0n129,notn129,n130);
and (s1n129,n19,n131);
nand (n133,n127,n122);
nand (n134,n135,n136);
or (n135,n127,n105);
nand (n136,n105,n127);
nand (n137,n138,n120);
nand (n138,n139,n145);
or (n139,n117,n140);
wire s0n140,s1n140,notn140;
or (n140,s0n140,s1n140);
not(notn140,n52);
and (s0n140,notn140,n141);
and (s1n140,n52,n144);
wire s0n141,s1n141,notn141;
or (n141,s0n141,s1n141);
not(notn141,n43);
and (s0n141,notn141,n142);
and (s1n141,n43,n143);
nand (n145,n140,n117);
nand (n146,n147,n178);
or (n147,n148,n158);
not (n148,n149);
nand (n149,n150,n157);
or (n150,n151,n152);
not (n151,n122);
wire s0n152,s1n152,notn152;
or (n152,s0n152,s1n152);
not(notn152,n52);
and (s0n152,notn152,n153);
and (s1n152,n52,n156);
wire s0n153,s1n153,notn153;
or (n153,s0n153,s1n153);
not(notn153,n43);
and (s0n153,notn153,n154);
and (s1n153,n43,n155);
nand (n157,n152,n151);
not (n158,n159);
nor (n159,n160,n174);
nand (n160,n161,n173);
or (n161,n162,n168);
not (n162,n163);
wire s0n163,s1n163,notn163;
or (n163,s0n163,s1n163);
not(notn163,n28);
and (s0n163,notn163,n164);
and (s1n163,n28,n167);
wire s0n164,s1n164,notn164;
or (n164,s0n164,s1n164);
not(notn164,n19);
and (s0n164,notn164,n165);
and (s1n164,n19,n166);
wire s0n168,s1n168,notn168;
or (n168,s0n168,s1n168);
not(notn168,n28);
and (s0n168,notn168,n169);
and (s1n168,n28,n172);
wire s0n169,s1n169,notn169;
or (n169,s0n169,s1n169);
not(notn169,n19);
and (s0n169,notn169,n170);
and (s1n169,n19,n171);
nand (n173,n168,n162);
not (n174,n175);
nand (n175,n176,n177);
or (n176,n122,n162);
nand (n177,n162,n122);
nand (n178,n179,n160);
nand (n179,n180,n186);
or (n180,n151,n181);
wire s0n181,s1n181,notn181;
or (n181,s0n181,s1n181);
not(notn181,n52);
and (s0n181,notn181,n182);
and (s1n181,n52,n185);
wire s0n182,s1n182,notn182;
or (n182,s0n182,s1n182);
not(notn182,n43);
and (s0n182,notn182,n183);
and (s1n182,n43,n184);
nand (n186,n181,n151);
and (n187,n11,n100);
xor (n188,n189,n231);
xor (n189,n190,n200);
and (n190,n191,n111);
nand (n191,n192,n199);
or (n192,n193,n105);
not (n193,n194);
wire s0n194,s1n194,notn194;
or (n194,s0n194,s1n194);
not(notn194,n28);
and (s0n194,notn194,n195);
and (s1n194,n28,n198);
wire s0n195,s1n195,notn195;
or (n195,s0n195,s1n195);
not(notn195,n19);
and (s0n195,notn195,n196);
and (s1n195,n19,n197);
nand (n199,n105,n193);
nand (n200,n201,n227);
or (n201,n202,n212);
not (n202,n203);
nand (n203,n204,n211);
or (n204,n168,n205);
not (n205,n206);
wire s0n206,s1n206,notn206;
or (n206,s0n206,s1n206);
not(notn206,n52);
and (s0n206,notn206,n207);
and (s1n206,n52,n210);
wire s0n207,s1n207,notn207;
or (n207,s0n207,s1n207);
not(notn207,n43);
and (s0n207,notn207,n208);
and (s1n207,n43,n209);
nand (n211,n205,n168);
not (n212,n213);
nor (n213,n214,n224);
nor (n214,n215,n222);
and (n215,n216,n217);
not (n216,n168);
wire s0n217,s1n217,notn217;
or (n217,s0n217,s1n217);
not(notn217,n28);
and (s0n217,notn217,n218);
and (s1n217,n28,n221);
wire s0n218,s1n218,notn218;
or (n218,s0n218,s1n218);
not(notn218,n19);
and (s0n218,notn218,n219);
and (s1n218,n19,n220);
and (n222,n168,n223);
not (n223,n217);
nand (n224,n225,n226);
or (n225,n30,n223);
nand (n226,n223,n30);
nand (n227,n228,n224);
nand (n228,n229,n230);
or (n229,n168,n38);
nand (n230,n38,n168);
nand (n231,n232,n234);
or (n232,n13,n233);
not (n233,n91);
nand (n234,n235,n15);
nand (n235,n236,n243);
or (n236,n30,n237);
not (n237,n238);
wire s0n238,s1n238,notn238;
or (n238,s0n238,s1n238);
not(notn238,n52);
and (s0n238,notn238,n239);
and (s1n238,n52,n242);
wire s0n239,s1n239,notn239;
or (n239,s0n239,s1n239);
not(notn239,n43);
and (s0n239,notn239,n240);
and (s1n239,n43,n241);
nand (n243,n237,n30);
xor (n244,n245,n265);
xor (n245,n246,n253);
nand (n246,n247,n249);
or (n247,n248,n118);
not (n248,n138);
nand (n249,n250,n120);
nand (n250,n251,n252);
or (n251,n117,n152);
nand (n252,n152,n117);
nand (n253,n254,n256);
or (n254,n255,n158);
not (n255,n179);
nand (n256,n257,n160);
nand (n257,n258,n264);
or (n258,n151,n259);
wire s0n259,s1n259,notn259;
or (n259,s0n259,s1n259);
not(notn259,n52);
and (s0n259,notn259,n260);
and (s1n259,n52,n263);
wire s0n260,s1n260,notn260;
or (n260,s0n260,s1n260);
not(notn260,n43);
and (s0n260,notn260,n261);
and (s1n260,n43,n262);
nand (n264,n259,n151);
and (n265,n266,n273);
nand (n266,n267,n272);
or (n267,n268,n212);
not (n268,n269);
nand (n269,n270,n271);
or (n270,n216,n259);
nand (n271,n259,n216);
nand (n272,n203,n224);
nor (n273,n274,n117);
and (n274,n275,n278);
nand (n275,n276,n151);
not (n276,n277);
and (n277,n111,n128);
nand (n278,n110,n127);
or (n279,n280,n307);
and (n280,n281,n306);
xor (n281,n282,n286);
nand (n282,n283,n285);
or (n283,n273,n284);
not (n284,n266);
nand (n285,n284,n273);
or (n286,n287,n305);
and (n287,n288,n298);
xor (n288,n289,n290);
and (n289,n120,n111);
nand (n290,n291,n297);
or (n291,n292,n212);
not (n292,n293);
nand (n293,n294,n296);
or (n294,n168,n295);
not (n295,n181);
nand (n296,n295,n168);
nand (n297,n269,n224);
nand (n298,n299,n304);
or (n299,n300,n158);
not (n300,n301);
nand (n301,n302,n303);
or (n302,n151,n140);
nand (n303,n140,n151);
nand (n304,n149,n160);
and (n305,n289,n290);
xor (n306,n10,n146);
and (n307,n282,n286);
not (n308,n309);
nand (n309,n310,n451);
or (n310,n311,n342);
not (n311,n312);
nand (n312,n313,n315);
not (n313,n314);
xor (n314,n281,n306);
not (n315,n316);
or (n316,n317,n341);
and (n317,n318,n340);
xor (n318,n319,n326);
nand (n319,n320,n325);
or (n320,n13,n321);
not (n321,n322);
nand (n322,n323,n324);
or (n323,n29,n206);
nand (n324,n206,n29);
nand (n325,n36,n15);
and (n326,n327,n333);
nor (n327,n328,n151);
and (n328,n329,n332);
nand (n329,n330,n216);
not (n330,n331);
and (n331,n111,n163);
nand (n332,n110,n162);
nand (n333,n334,n339);
or (n334,n335,n212);
not (n335,n336);
nand (n336,n337,n338);
or (n337,n216,n152);
nand (n338,n152,n216);
nand (n339,n293,n224);
xor (n340,n288,n298);
and (n341,n319,n326);
not (n342,n343);
nand (n343,n344,n450);
or (n344,n345,n445);
nor (n345,n346,n444);
and (n346,n347,n387);
nand (n347,n348,n367);
not (n348,n349);
xor (n349,n350,n366);
xor (n350,n351,n358);
nand (n351,n352,n357);
or (n352,n353,n158);
not (n353,n354);
nor (n354,n355,n356);
and (n355,n111,n122);
and (n356,n151,n110);
nand (n357,n160,n301);
nand (n358,n359,n361);
or (n359,n360,n321);
not (n360,n15);
nand (n361,n362,n14);
nand (n362,n363,n365);
or (n363,n30,n364);
not (n364,n259);
nand (n365,n30,n364);
xor (n366,n327,n333);
not (n367,n368);
or (n368,n369,n386);
and (n369,n370,n379);
xor (n370,n371,n372);
and (n371,n160,n111);
nand (n372,n373,n375);
or (n373,n360,n374);
not (n374,n362);
nand (n375,n376,n14);
nand (n376,n377,n378);
or (n377,n30,n295);
nand (n378,n295,n30);
nand (n379,n380,n385);
or (n380,n381,n212);
not (n381,n382);
nand (n382,n383,n384);
or (n383,n216,n140);
nand (n384,n140,n216);
nand (n385,n336,n224);
and (n386,n371,n372);
nand (n387,n388,n442);
or (n388,n389,n407);
not (n389,n390);
nand (n390,n391,n393);
not (n391,n392);
xor (n392,n370,n379);
nand (n393,n394,n401);
nand (n394,n395,n397);
or (n395,n360,n396);
not (n396,n376);
nand (n397,n398,n14);
nand (n398,n399,n400);
or (n399,n29,n152);
nand (n400,n152,n29);
nor (n401,n402,n216);
and (n402,n403,n406);
nand (n403,n404,n29);
not (n404,n405);
and (n405,n111,n217);
nand (n406,n110,n223);
not (n407,n408);
or (n408,n409,n441);
and (n409,n410,n422);
xor (n410,n411,n418);
nand (n411,n412,n417);
or (n412,n413,n212);
not (n413,n414);
nor (n414,n415,n416);
and (n415,n111,n168);
and (n416,n216,n110);
nand (n417,n224,n382);
nand (n418,n419,n421);
or (n419,n420,n394);
not (n420,n401);
nand (n421,n394,n420);
or (n422,n423,n440);
and (n423,n424,n433);
xor (n424,n425,n426);
and (n425,n111,n224);
nand (n426,n427,n429);
or (n427,n360,n428);
not (n428,n398);
nand (n429,n430,n14);
nand (n430,n431,n432);
or (n431,n29,n140);
nand (n432,n140,n29);
nor (n433,n434,n437);
nor (n434,n435,n436);
and (n435,n14,n110);
and (n436,n430,n15);
nand (n437,n438,n30);
not (n438,n439);
and (n439,n111,n15);
and (n440,n425,n426);
and (n441,n411,n418);
nand (n442,n392,n443);
not (n443,n393);
and (n444,n349,n368);
nor (n445,n446,n447);
xor (n446,n318,n340);
or (n447,n448,n449);
and (n448,n350,n366);
and (n449,n351,n358);
nand (n450,n446,n447);
nand (n451,n314,n316);
nand (n452,n6,n279);
nand (n453,n454,n533);
not (n454,n455);
nor (n455,n456,n530);
xor (n456,n457,n490);
xor (n457,n458,n487);
xor (n458,n459,n480);
xor (n459,n460,n473);
nand (n460,n461,n463);
or (n461,n13,n462);
not (n462,n235);
nand (n463,n464,n15);
nand (n464,n465,n472);
or (n465,n30,n466);
not (n466,n467);
wire s0n467,s1n467,notn467;
or (n467,s0n467,s1n467);
not(notn467,n52);
and (s0n467,notn467,n468);
and (s1n467,n52,n471);
wire s0n468,s1n468,notn468;
or (n468,s0n468,s1n468);
not(notn468,n43);
and (s0n468,notn468,n469);
and (s1n468,n43,n470);
nand (n472,n466,n30);
nand (n473,n474,n476);
or (n474,n475,n212);
not (n475,n228);
nand (n476,n477,n224);
nor (n477,n478,n479);
and (n478,n94,n168);
and (n479,n216,n93);
nand (n480,n481,n483);
or (n481,n482,n118);
not (n482,n250);
nand (n483,n484,n120);
nand (n484,n485,n486);
or (n485,n105,n295);
nand (n486,n295,n105);
or (n487,n488,n489);
and (n488,n245,n265);
and (n489,n246,n253);
xor (n490,n491,n527);
xor (n491,n492,n513);
nand (n492,n493,n509);
or (n493,n494,n505);
not (n494,n495);
nor (n495,n496,n191);
nor (n496,n497,n504);
and (n497,n498,n194);
not (n498,n499);
wire s0n499,s1n499,notn499;
or (n499,s0n499,s1n499);
not(notn499,n28);
and (s0n499,notn499,n500);
and (s1n499,n28,n503);
wire s0n500,s1n500,notn500;
or (n500,s0n500,s1n500);
not(notn500,n19);
and (s0n500,notn500,n501);
and (s1n500,n19,n502);
and (n504,n499,n193);
not (n505,n506);
nor (n506,n507,n508);
and (n507,n498,n110);
and (n508,n111,n499);
nand (n509,n191,n510);
nand (n510,n511,n512);
or (n511,n498,n140);
nand (n512,n498,n140);
xor (n513,n514,n520);
nor (n514,n515,n498);
and (n515,n516,n519);
nand (n516,n517,n117);
not (n517,n518);
and (n518,n111,n194);
nand (n519,n110,n193);
nand (n520,n521,n523);
or (n521,n158,n522);
not (n522,n257);
nand (n523,n524,n160);
nand (n524,n525,n526);
or (n525,n151,n206);
nand (n526,n206,n151);
or (n527,n528,n529);
and (n528,n189,n231);
and (n529,n190,n200);
or (n530,n531,n532);
and (n531,n7,n244);
and (n532,n8,n188);
nand (n533,n456,n530);
nand (n534,n3,n453);
not (n535,n536);
or (n536,n537,n634,n646);
and (n537,n538,n547);
xor (n538,n539,n546);
xor (n539,n540,n543);
xor (n540,n541,n542);
and (n541,n218,n111);
and (n542,n31,n140);
and (n543,n544,n545);
and (n544,n31,n111);
and (n545,n16,n140);
and (n546,n16,n152);
not (n547,n548);
xor (n548,n549,n628);
xor (n549,n550,n622);
xor (n550,n551,n613);
and (n551,n552,n563);
wire s0n552,s1n552,notn552;
or (n552,s0n552,s1n552);
not(notn552,n555);
and (s0n552,notn552,n553);
and (s1n552,n555,n554);
and (n555,n556,n561);
and (n556,n557,n559);
not (n557,n558);
not (n559,n560);
not (n561,n562);
wire s0n563,s1n563,notn563;
or (n563,s0n563,s1n563);
not(notn563,n576);
and (s0n563,notn563,n564);
and (s1n563,n576,n575);
wire s0n564,s1n564,notn564;
or (n564,s0n564,s1n564);
not(notn564,n567);
and (s0n564,notn564,n565);
and (s1n564,n567,n566);
and (n567,n568,n573);
and (n568,n569,n571);
not (n569,n570);
not (n571,n572);
not (n573,n574);
and (n576,n577,n579);
not (n577,n578);
or (n579,n580,n581);
and (n581,n582,n583);
or (n583,n584,n585,n586,n587,n588,n589,n590,n591,n592,n593,n594,n595,n596,n597,n598,n599,n600,n601,n602,n603,n604,n605,n606,n607,n608,n609,n610,n611,n612);
and (n613,n614,n617);
wire s0n614,s1n614,notn614;
or (n614,s0n614,s1n614);
not(notn614,n555);
and (s0n614,notn614,n615);
and (s1n614,n555,n616);
wire s0n617,s1n617,notn617;
or (n617,s0n617,s1n617);
not(notn617,n576);
and (s0n617,notn617,n618);
and (s1n617,n576,n621);
wire s0n618,s1n618,notn618;
or (n618,s0n618,s1n618);
not(notn618,n567);
and (s0n618,notn618,n619);
and (s1n618,n567,n620);
and (n622,n623,n624);
and (n623,n614,n563);
and (n624,n625,n617);
wire s0n625,s1n625,notn625;
or (n625,s0n625,s1n625);
not(notn625,n555);
and (s0n625,notn625,n626);
and (s1n625,n555,n627);
and (n628,n625,n629);
wire s0n629,s1n629,notn629;
or (n629,s0n629,s1n629);
not(notn629,n576);
and (s0n629,notn629,n630);
and (s1n629,n576,n633);
wire s0n630,s1n630,notn630;
or (n630,s0n630,s1n630);
not(notn630,n567);
and (s0n630,notn630,n631);
and (s1n630,n567,n632);
and (n634,n547,n635);
or (n635,n636,n640,n645);
and (n636,n637,n638);
xor (n637,n544,n545);
not (n638,n639);
xor (n639,n623,n624);
and (n640,n638,n641);
or (n641,n642,n643);
and (n642,n16,n111);
not (n643,n644);
and (n644,n625,n563);
and (n645,n637,n641);
and (n646,n538,n635);
and (n647,n535,n648);
xor (n648,n649,n508);
xor (n649,n650,n858);
xor (n650,n651,n857);
xor (n651,n652,n848);
xor (n652,n653,n847);
xor (n653,n654,n833);
xor (n654,n655,n832);
xor (n655,n656,n812);
xor (n656,n657,n811);
xor (n657,n658,n785);
xor (n658,n659,n784);
xor (n659,n660,n752);
xor (n660,n661,n751);
xor (n661,n662,n713);
xor (n662,n663,n712);
xor (n663,n664,n667);
xor (n664,n665,n666);
and (n665,n467,n15);
and (n666,n238,n30);
or (n667,n668,n671);
and (n668,n669,n670);
and (n669,n238,n15);
and (n670,n94,n30);
and (n671,n672,n673);
xor (n672,n669,n670);
or (n673,n674,n677);
and (n674,n675,n676);
and (n675,n94,n15);
and (n676,n39,n30);
and (n677,n678,n679);
xor (n678,n675,n676);
or (n679,n680,n683);
and (n680,n681,n682);
and (n681,n39,n15);
and (n682,n206,n30);
and (n683,n684,n685);
xor (n684,n681,n682);
or (n685,n686,n689);
and (n686,n687,n688);
and (n687,n206,n15);
and (n688,n259,n30);
and (n689,n690,n691);
xor (n690,n687,n688);
or (n691,n692,n695);
and (n692,n693,n694);
and (n693,n259,n15);
and (n694,n181,n30);
and (n695,n696,n697);
xor (n696,n693,n694);
or (n697,n698,n701);
and (n698,n699,n700);
and (n699,n181,n15);
and (n700,n152,n30);
and (n701,n702,n703);
xor (n702,n699,n700);
or (n703,n704,n707);
and (n704,n705,n706);
and (n705,n152,n15);
and (n706,n140,n30);
and (n707,n708,n709);
xor (n708,n705,n706);
and (n709,n710,n711);
and (n710,n140,n15);
and (n711,n111,n30);
and (n712,n94,n217);
or (n713,n714,n717);
and (n714,n715,n716);
xor (n715,n672,n673);
and (n716,n39,n217);
and (n717,n718,n719);
xor (n718,n715,n716);
or (n719,n720,n723);
and (n720,n721,n722);
xor (n721,n678,n679);
and (n722,n206,n217);
and (n723,n724,n725);
xor (n724,n721,n722);
or (n725,n726,n729);
and (n726,n727,n728);
xor (n727,n684,n685);
and (n728,n259,n217);
and (n729,n730,n731);
xor (n730,n727,n728);
or (n731,n732,n735);
and (n732,n733,n734);
xor (n733,n690,n691);
and (n734,n181,n217);
and (n735,n736,n737);
xor (n736,n733,n734);
or (n737,n738,n741);
and (n738,n739,n740);
xor (n739,n696,n697);
and (n740,n152,n217);
and (n741,n742,n743);
xor (n742,n739,n740);
or (n743,n744,n747);
and (n744,n745,n746);
xor (n745,n702,n703);
and (n746,n140,n217);
and (n747,n748,n749);
xor (n748,n745,n746);
and (n749,n750,n405);
xor (n750,n708,n709);
and (n751,n39,n168);
or (n752,n753,n756);
and (n753,n754,n755);
xor (n754,n718,n719);
and (n755,n206,n168);
and (n756,n757,n758);
xor (n757,n754,n755);
or (n758,n759,n762);
and (n759,n760,n761);
xor (n760,n724,n725);
and (n761,n259,n168);
and (n762,n763,n764);
xor (n763,n760,n761);
or (n764,n765,n768);
and (n765,n766,n767);
xor (n766,n730,n731);
and (n767,n181,n168);
and (n768,n769,n770);
xor (n769,n766,n767);
or (n770,n771,n774);
and (n771,n772,n773);
xor (n772,n736,n737);
and (n773,n152,n168);
and (n774,n775,n776);
xor (n775,n772,n773);
or (n776,n777,n780);
and (n777,n778,n779);
xor (n778,n742,n743);
and (n779,n140,n168);
and (n780,n781,n782);
xor (n781,n778,n779);
and (n782,n783,n415);
xor (n783,n748,n749);
and (n784,n206,n163);
or (n785,n786,n789);
and (n786,n787,n788);
xor (n787,n757,n758);
and (n788,n259,n163);
and (n789,n790,n791);
xor (n790,n787,n788);
or (n791,n792,n795);
and (n792,n793,n794);
xor (n793,n763,n764);
and (n794,n181,n163);
and (n795,n796,n797);
xor (n796,n793,n794);
or (n797,n798,n801);
and (n798,n799,n800);
xor (n799,n769,n770);
and (n800,n152,n163);
and (n801,n802,n803);
xor (n802,n799,n800);
or (n803,n804,n807);
and (n804,n805,n806);
xor (n805,n775,n776);
and (n806,n140,n163);
and (n807,n808,n809);
xor (n808,n805,n806);
and (n809,n810,n331);
xor (n810,n781,n782);
and (n811,n259,n122);
or (n812,n813,n816);
and (n813,n814,n815);
xor (n814,n790,n791);
and (n815,n181,n122);
and (n816,n817,n818);
xor (n817,n814,n815);
or (n818,n819,n822);
and (n819,n820,n821);
xor (n820,n796,n797);
and (n821,n152,n122);
and (n822,n823,n824);
xor (n823,n820,n821);
or (n824,n825,n828);
and (n825,n826,n827);
xor (n826,n802,n803);
and (n827,n140,n122);
and (n828,n829,n830);
xor (n829,n826,n827);
and (n830,n831,n355);
xor (n831,n808,n809);
and (n832,n181,n128);
or (n833,n834,n837);
and (n834,n835,n836);
xor (n835,n817,n818);
and (n836,n152,n128);
and (n837,n838,n839);
xor (n838,n835,n836);
or (n839,n840,n843);
and (n840,n841,n842);
xor (n841,n823,n824);
and (n842,n140,n128);
and (n843,n844,n845);
xor (n844,n841,n842);
and (n845,n846,n277);
xor (n846,n829,n830);
and (n847,n152,n105);
or (n848,n849,n852);
and (n849,n850,n851);
xor (n850,n838,n839);
and (n851,n140,n105);
and (n852,n853,n854);
xor (n853,n850,n851);
and (n854,n855,n856);
xor (n855,n844,n845);
and (n856,n111,n105);
and (n857,n140,n194);
and (n858,n859,n518);
xor (n859,n853,n854);
endmodule
