module top (out,n3,n4,n27,n28,n34,n38,n44,n53,n54
        ,n60,n64,n70,n79,n80,n92,n103,n109,n121,n122
        ,n142,n148,n157,n197,n368,n374,n381,n387,n421,n422
        ,n429,n442,n514,n534,n594);
output out;
input n3;
input n4;
input n27;
input n28;
input n34;
input n38;
input n44;
input n53;
input n54;
input n60;
input n64;
input n70;
input n79;
input n80;
input n92;
input n103;
input n109;
input n121;
input n122;
input n142;
input n148;
input n157;
input n197;
input n368;
input n374;
input n381;
input n387;
input n421;
input n422;
input n429;
input n442;
input n514;
input n534;
input n594;
wire n0;
wire n1;
wire n2;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n24;
wire n25;
wire n26;
wire n29;
wire n30;
wire n31;
wire n32;
wire n33;
wire n35;
wire n36;
wire n37;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n61;
wire n62;
wire n63;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2988;
wire n2989;
wire n2990;
wire n2991;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2996;
wire n2997;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3003;
wire n3004;
wire n3005;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3010;
wire n3011;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3038;
wire n3039;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
wire n3056;
wire n3057;
wire n3058;
wire n3059;
wire n3060;
wire n3061;
wire n3062;
wire n3063;
wire n3064;
wire n3065;
wire n3066;
wire n3067;
wire n3068;
wire n3069;
wire n3070;
wire n3071;
wire n3072;
wire n3073;
wire n3074;
wire n3075;
wire n3076;
wire n3077;
wire n3078;
wire n3079;
wire n3080;
wire n3081;
wire n3082;
wire n3083;
wire n3084;
wire n3085;
wire n3086;
wire n3087;
wire n3088;
wire n3089;
wire n3090;
wire n3091;
wire n3092;
wire n3093;
wire n3094;
wire n3095;
wire n3096;
wire n3097;
wire n3098;
wire n3099;
wire n3100;
wire n3101;
wire n3102;
wire n3103;
wire n3104;
wire n3105;
wire n3106;
wire n3107;
wire n3108;
wire n3109;
wire n3110;
wire n3111;
wire n3112;
wire n3113;
wire n3114;
wire n3115;
wire n3116;
wire n3117;
wire n3118;
wire n3119;
wire n3120;
wire n3121;
wire n3122;
wire n3123;
wire n3124;
wire n3125;
wire n3126;
wire n3127;
wire n3128;
wire n3129;
wire n3130;
wire n3131;
wire n3132;
wire n3133;
wire n3134;
wire n3135;
wire n3136;
wire n3137;
wire n3138;
wire n3139;
wire n3140;
wire n3141;
wire n3142;
wire n3143;
wire n3144;
wire n3145;
wire n3146;
wire n3147;
wire n3148;
wire n3149;
wire n3150;
wire n3151;
wire n3152;
wire n3153;
wire n3154;
wire n3155;
wire n3156;
wire n3157;
wire n3158;
wire n3159;
wire n3160;
wire n3161;
wire n3162;
wire n3163;
wire n3164;
wire n3165;
wire n3166;
wire n3167;
wire n3168;
wire n3169;
wire n3170;
wire n3171;
wire n3172;
wire n3173;
wire n3174;
wire n3175;
wire n3176;
wire n3177;
wire n3178;
wire n3179;
wire n3180;
wire n3181;
wire n3182;
wire n3183;
wire n3184;
wire n3185;
wire n3186;
wire n3187;
wire n3188;
wire n3189;
wire n3190;
wire n3191;
wire n3192;
wire n3193;
wire n3194;
wire n3195;
wire n3196;
wire n3197;
wire n3198;
wire n3199;
wire n3200;
wire n3201;
wire n3202;
wire n3203;
wire n3204;
wire n3205;
wire n3206;
wire n3207;
wire n3208;
wire n3209;
wire n3210;
wire n3211;
wire n3212;
wire n3213;
wire n3214;
wire n3215;
wire n3216;
wire n3217;
wire n3218;
wire n3219;
wire n3220;
wire n3221;
wire n3222;
wire n3223;
wire n3224;
wire n3225;
wire n3226;
wire n3227;
wire n3228;
wire n3229;
wire n3230;
wire n3231;
wire n3232;
wire n3233;
wire n3234;
wire n3235;
wire n3236;
wire n3237;
wire n3238;
wire n3239;
wire n3240;
wire n3241;
wire n3242;
wire n3243;
wire n3244;
wire n3245;
wire n3246;
wire n3247;
wire n3248;
wire n3249;
wire n3250;
wire n3251;
wire n3252;
wire n3253;
wire n3254;
wire n3255;
wire n3256;
wire n3257;
wire n3258;
wire n3259;
wire n3260;
wire n3261;
wire n3262;
wire n3263;
wire n3264;
wire n3265;
wire n3266;
wire n3267;
wire n3268;
wire n3269;
wire n3270;
wire n3271;
wire n3272;
wire n3273;
wire n3274;
wire n3275;
wire n3276;
wire n3277;
wire n3278;
wire n3279;
wire n3280;
wire n3281;
wire n3282;
wire n3283;
wire n3284;
wire n3285;
wire n3286;
wire n3287;
wire n3288;
wire n3289;
wire n3290;
wire n3291;
wire n3292;
wire n3293;
wire n3294;
wire n3295;
wire n3296;
wire n3297;
wire n3298;
wire n3299;
wire n3300;
wire n3301;
wire n3302;
wire n3303;
wire n3304;
wire n3305;
wire n3306;
wire n3307;
wire n3308;
wire n3309;
wire n3310;
wire n3311;
wire n3312;
wire n3313;
wire n3314;
wire n3315;
wire n3316;
wire n3317;
wire n3318;
wire n3319;
wire n3320;
wire n3321;
wire n3322;
wire n3323;
wire n3324;
wire n3325;
wire n3326;
wire n3327;
wire n3328;
wire n3329;
wire n3330;
wire n3331;
wire n3332;
wire n3333;
wire n3334;
wire n3335;
wire n3336;
wire n3337;
wire n3338;
wire n3339;
wire n3340;
wire n3341;
wire n3342;
wire n3343;
wire n3344;
wire n3345;
wire n3346;
wire n3347;
wire n3348;
wire n3349;
wire n3350;
wire n3351;
wire n3352;
wire n3353;
wire n3354;
wire n3355;
wire n3356;
wire n3357;
wire n3358;
wire n3359;
wire n3360;
wire n3361;
wire n3362;
wire n3363;
wire n3364;
wire n3365;
wire n3366;
wire n3367;
wire n3368;
wire n3369;
wire n3370;
wire n3371;
wire n3372;
wire n3373;
wire n3374;
wire n3375;
wire n3376;
wire n3377;
wire n3378;
wire n3379;
wire n3380;
wire n3381;
wire n3382;
wire n3383;
wire n3384;
wire n3385;
wire n3386;
wire n3387;
wire n3388;
wire n3389;
wire n3390;
wire n3391;
wire n3392;
wire n3393;
wire n3394;
wire n3395;
wire n3396;
wire n3397;
wire n3398;
wire n3399;
wire n3400;
wire n3401;
wire n3402;
wire n3403;
wire n3404;
wire n3405;
wire n3406;
wire n3407;
wire n3408;
wire n3409;
wire n3410;
wire n3411;
wire n3412;
wire n3413;
wire n3414;
wire n3415;
wire n3416;
wire n3417;
wire n3418;
wire n3419;
wire n3420;
wire n3421;
wire n3422;
wire n3423;
wire n3424;
wire n3425;
wire n3426;
wire n3427;
wire n3428;
wire n3429;
wire n3430;
wire n3431;
wire n3432;
wire n3433;
wire n3434;
wire n3435;
wire n3436;
wire n3437;
wire n3438;
wire n3439;
wire n3440;
wire n3441;
wire n3442;
wire n3443;
wire n3444;
wire n3445;
wire n3446;
wire n3447;
wire n3448;
wire n3449;
wire n3450;
wire n3451;
wire n3452;
wire n3453;
wire n3454;
wire n3455;
wire n3456;
wire n3457;
wire n3458;
wire n3459;
wire n3460;
wire n3461;
wire n3462;
wire n3463;
wire n3464;
wire n3465;
wire n3466;
wire n3467;
wire n3468;
wire n3469;
wire n3470;
wire n3471;
wire n3472;
wire n3473;
wire n3474;
wire n3475;
wire n3476;
wire n3477;
wire n3478;
wire n3479;
wire n3480;
wire n3481;
wire n3482;
wire n3483;
wire n3484;
wire n3485;
wire n3486;
wire n3487;
wire n3488;
wire n3489;
wire n3490;
wire n3491;
wire n3492;
wire n3493;
wire n3494;
wire n3495;
wire n3496;
wire n3497;
wire n3498;
wire n3499;
wire n3500;
wire n3501;
wire n3502;
wire n3503;
wire n3504;
wire n3505;
wire n3506;
wire n3507;
wire n3508;
wire n3509;
wire n3510;
wire n3511;
wire n3512;
wire n3513;
wire n3514;
wire n3515;
wire n3516;
wire n3517;
wire n3518;
wire n3519;
wire n3520;
wire n3521;
wire n3522;
wire n3523;
wire n3524;
wire n3525;
wire n3526;
wire n3527;
wire n3528;
wire n3529;
wire n3530;
wire n3531;
wire n3532;
wire n3533;
wire n3534;
wire n3535;
wire n3536;
wire n3537;
wire n3538;
wire n3539;
wire n3540;
wire n3541;
wire n3542;
wire n3543;
wire n3544;
wire n3545;
wire n3546;
wire n3547;
wire n3548;
wire n3549;
wire n3550;
wire n3551;
wire n3552;
wire n3553;
wire n3554;
wire n3555;
wire n3556;
wire n3557;
wire n3558;
wire n3559;
wire n3560;
wire n3561;
wire n3562;
wire n3563;
wire n3564;
wire n3565;
wire n3566;
wire n3567;
wire n3568;
wire n3569;
wire n3570;
wire n3571;
wire n3572;
wire n3573;
wire n3574;
wire n3575;
wire n3576;
wire n3577;
wire n3578;
wire n3579;
wire n3580;
wire n3581;
wire n3582;
wire n3583;
wire n3584;
wire n3585;
wire n3586;
wire n3587;
wire n3588;
wire n3589;
wire n3590;
wire n3591;
wire n3592;
wire n3593;
wire n3594;
wire n3595;
wire n3596;
wire n3597;
wire n3598;
wire n3599;
wire n3600;
wire n3601;
wire n3602;
wire n3603;
wire n3604;
wire n3605;
wire n3606;
wire n3607;
wire n3608;
wire n3609;
wire n3610;
wire n3611;
wire n3612;
wire n3613;
wire n3614;
wire n3615;
wire n3616;
wire n3617;
wire n3618;
wire n3619;
wire n3620;
wire n3621;
wire n3622;
wire n3623;
wire n3624;
wire n3625;
wire n3626;
wire n3627;
wire n3628;
wire n3629;
wire n3630;
wire n3631;
wire n3632;
wire n3633;
wire n3634;
wire n3635;
wire n3636;
wire n3637;
wire n3638;
wire n3639;
wire n3640;
wire n3641;
wire n3642;
wire n3643;
wire n3644;
wire n3645;
wire n3646;
wire n3647;
wire n3648;
wire n3649;
wire n3650;
wire n3651;
wire n3652;
wire n3653;
wire n3654;
wire n3655;
wire n3656;
wire n3657;
wire n3658;
wire n3659;
wire n3660;
wire n3661;
wire n3662;
wire n3663;
wire n3664;
wire n3665;
wire n3666;
wire n3667;
wire n3668;
wire n3669;
wire n3670;
wire n3671;
wire n3672;
wire n3673;
wire n3674;
wire n3675;
wire n3676;
wire n3677;
wire n3678;
wire n3679;
wire n3680;
wire n3681;
wire n3682;
wire n3683;
wire n3684;
wire n3685;
wire n3686;
wire n3687;
wire n3688;
wire n3689;
wire n3690;
wire n3691;
wire n3692;
wire n3693;
wire n3694;
wire n3695;
wire n3696;
wire n3697;
wire n3698;
wire n3699;
wire n3700;
wire n3701;
wire n3702;
wire n3703;
wire n3704;
wire n3705;
wire n3706;
wire n3707;
wire n3708;
wire n3709;
wire n3710;
wire n3711;
wire n3712;
wire n3713;
wire n3714;
wire n3715;
wire n3716;
wire n3717;
wire n3718;
wire n3719;
wire n3720;
wire n3721;
wire n3722;
wire n3723;
wire n3724;
wire n3725;
wire n3726;
wire n3727;
wire n3728;
wire n3729;
wire n3730;
wire n3731;
wire n3732;
wire n3733;
wire n3734;
wire n3735;
wire n3736;
wire n3737;
wire n3738;
wire n3739;
wire n3740;
wire n3741;
wire n3742;
wire n3743;
wire n3744;
wire n3745;
wire n3746;
wire n3747;
wire n3748;
wire n3749;
wire n3750;
wire n3751;
wire n3752;
wire n3753;
wire n3754;
wire n3755;
wire n3756;
wire n3757;
wire n3758;
wire n3759;
wire n3760;
wire n3761;
wire n3762;
wire n3763;
wire n3764;
wire n3765;
wire n3766;
wire n3767;
wire n3768;
wire n3769;
wire n3770;
wire n3771;
wire n3772;
wire n3773;
wire n3774;
wire n3775;
wire n3776;
wire n3777;
wire n3778;
wire n3779;
wire n3780;
wire n3781;
wire n3782;
wire n3783;
wire n3784;
wire n3785;
wire n3786;
wire n3787;
wire n3788;
wire n3789;
wire n3790;
wire n3791;
wire n3792;
wire n3793;
wire n3794;
wire n3795;
wire n3796;
wire n3797;
wire n3798;
wire n3799;
wire n3800;
wire n3801;
wire n3802;
wire n3803;
wire n3804;
wire n3805;
wire n3806;
wire n3807;
wire n3808;
wire n3809;
wire n3810;
wire n3811;
wire n3812;
wire n3813;
wire n3814;
wire n3815;
wire n3816;
wire n3817;
wire n3818;
wire n3819;
wire n3820;
wire n3821;
wire n3822;
wire n3823;
wire n3824;
wire n3825;
wire n3826;
wire n3827;
wire n3828;
wire n3829;
wire n3830;
wire n3831;
wire n3832;
wire n3833;
wire n3834;
wire n3835;
wire n3836;
wire n3837;
wire n3838;
wire n3839;
wire n3840;
wire n3841;
wire n3842;
wire n3843;
wire n3844;
wire n3845;
wire n3846;
wire n3847;
wire n3848;
wire n3849;
wire n3850;
wire n3851;
wire n3852;
wire n3853;
wire n3854;
wire n3855;
wire n3856;
wire n3857;
wire n3858;
wire n3859;
wire n3860;
wire n3861;
wire n3862;
wire n3863;
wire n3864;
wire n3865;
wire n3866;
wire n3867;
wire n3868;
wire n3869;
wire n3870;
wire n3871;
wire n3872;
wire n3873;
wire n3874;
wire n3875;
wire n3876;
wire n3877;
wire n3878;
wire n3879;
wire n3880;
wire n3881;
wire n3882;
wire n3883;
wire n3884;
wire n3885;
wire n3886;
wire n3887;
wire n3888;
wire n3889;
wire n3890;
wire n3891;
wire n3892;
wire n3893;
wire n3894;
wire n3895;
wire n3896;
wire n3897;
wire n3898;
wire n3899;
wire n3900;
xor (out,n0,n1621);
and (n0,n1,n5);
nor (n1,n2,n4);
not (n2,n3);
nand (n5,n6,n1619);
nand (n6,n7,n1609,n1615);
nand (n7,n8,n1582);
nand (n8,n9,n1570);
or (n9,n10,n338);
not (n10,n11);
and (n11,n12,n285,n313);
and (n12,n13,n248);
nand (n13,n14,n212);
not (n14,n15);
or (n15,n16,n211);
and (n16,n17,n181);
xor (n17,n18,n96);
or (n18,n19,n95);
and (n19,n20,n73);
xor (n20,n21,n47);
nand (n21,n22,n41);
or (n22,n23,n36);
nand (n23,n24,n31);
nor (n24,n25,n29);
and (n25,n26,n28);
not (n26,n27);
and (n29,n27,n30);
not (n30,n28);
nand (n31,n32,n35);
or (n32,n33,n28);
not (n33,n34);
nand (n35,n33,n28);
nor (n36,n37,n39);
and (n37,n33,n38);
and (n39,n34,n40);
not (n40,n38);
or (n41,n42,n24);
nor (n42,n43,n45);
and (n43,n33,n44);
and (n45,n34,n46);
not (n46,n44);
nand (n47,n48,n67);
or (n48,n49,n62);
nand (n49,n50,n57);
nor (n50,n51,n55);
and (n51,n52,n54);
not (n52,n53);
and (n55,n53,n56);
not (n56,n54);
nand (n57,n58,n61);
nand (n58,n59,n54);
not (n59,n60);
nand (n61,n60,n56);
nor (n62,n63,n65);
and (n63,n59,n64);
and (n65,n60,n66);
not (n66,n64);
or (n67,n50,n68);
nor (n68,n69,n71);
and (n69,n59,n70);
and (n71,n60,n72);
not (n72,n70);
nand (n73,n74,n89);
or (n74,n75,n86);
nand (n75,n76,n83);
nor (n76,n77,n81);
and (n77,n78,n80);
not (n78,n79);
and (n81,n79,n82);
not (n82,n80);
nand (n83,n84,n85);
or (n84,n52,n80);
nand (n85,n52,n80);
nor (n86,n87,n88);
and (n87,n52,n70);
and (n88,n53,n72);
or (n89,n76,n90);
nor (n90,n91,n93);
and (n91,n52,n92);
and (n93,n53,n94);
not (n94,n92);
and (n95,n21,n47);
xor (n96,n97,n161);
xor (n97,n98,n112);
not (n98,n99);
nand (n99,n100,n106);
or (n100,n75,n101);
nor (n101,n102,n104);
and (n102,n52,n103);
and (n104,n53,n105);
not (n105,n103);
or (n106,n76,n107);
nor (n107,n108,n110);
and (n108,n52,n109);
and (n110,n53,n111);
not (n111,n109);
or (n112,n113,n160);
and (n113,n114,n137);
xor (n114,n115,n134);
nand (n115,n116,n130);
or (n116,n117,n125);
not (n117,n118);
nor (n118,n119,n123);
and (n119,n120,n122);
not (n120,n121);
and (n123,n121,n124);
not (n124,n122);
not (n125,n126);
nand (n126,n118,n127);
nand (n127,n128,n129);
or (n128,n122,n78);
nand (n129,n78,n122);
not (n130,n131);
nor (n131,n132,n133);
and (n132,n78,n109);
and (n133,n79,n111);
nand (n134,n135,n136);
or (n135,n75,n90);
or (n136,n76,n101);
nand (n137,n138,n150);
or (n138,n139,n144);
nor (n139,n140,n143);
and (n140,n60,n141);
not (n141,n142);
and (n143,n59,n142);
not (n144,n145);
nand (n145,n146,n149);
or (n146,n27,n147);
not (n147,n148);
or (n149,n26,n148);
or (n150,n151,n155);
nand (n151,n152,n139);
or (n152,n153,n154);
and (n153,n141,n27);
and (n154,n142,n26);
nor (n155,n156,n158);
and (n156,n26,n157);
and (n158,n27,n159);
not (n159,n157);
and (n160,n115,n134);
xor (n161,n162,n175);
xor (n162,n163,n169);
nand (n163,n164,n165);
or (n164,n23,n42);
or (n165,n24,n166);
nor (n166,n167,n168);
and (n167,n33,n157);
and (n168,n34,n159);
nand (n169,n170,n171);
or (n170,n49,n68);
or (n171,n50,n172);
nor (n172,n173,n174);
and (n173,n59,n92);
and (n174,n60,n94);
nand (n175,n176,n177);
or (n176,n144,n151);
or (n177,n178,n139);
nor (n178,n179,n180);
and (n179,n26,n64);
and (n180,n27,n66);
or (n181,n182,n210);
and (n182,n183,n209);
xor (n183,n184,n208);
or (n184,n185,n207);
and (n185,n186,n201);
xor (n186,n187,n193);
nand (n187,n188,n192);
or (n188,n151,n189);
nor (n189,n190,n191);
and (n190,n44,n26);
and (n191,n27,n46);
or (n192,n155,n139);
nand (n193,n194,n200);
or (n194,n23,n195);
nor (n195,n196,n198);
and (n196,n197,n33);
and (n198,n34,n199);
not (n199,n197);
or (n200,n24,n36);
nand (n201,n202,n206);
or (n202,n126,n203);
nor (n203,n204,n205);
and (n204,n78,n103);
and (n205,n79,n105);
or (n206,n118,n131);
and (n207,n187,n193);
xor (n208,n114,n137);
xor (n209,n20,n73);
and (n210,n184,n208);
and (n211,n18,n96);
not (n212,n213);
xor (n213,n214,n245);
xor (n214,n215,n234);
xor (n215,n216,n228);
xor (n216,n217,n222);
nand (n217,n218,n221);
or (n218,n219,n220);
not (n219,n75);
not (n220,n76);
not (n221,n107);
nand (n222,n223,n224);
or (n223,n49,n172);
or (n224,n50,n225);
nor (n225,n226,n227);
and (n226,n59,n103);
and (n227,n60,n105);
nand (n228,n229,n230);
or (n229,n23,n166);
or (n230,n24,n231);
nor (n231,n232,n233);
and (n232,n33,n148);
and (n233,n34,n147);
xor (n234,n235,n242);
xor (n235,n236,n99);
nand (n236,n237,n238);
or (n237,n151,n178);
or (n238,n139,n239);
nor (n239,n240,n241);
and (n240,n26,n70);
and (n241,n27,n72);
or (n242,n243,n244);
and (n243,n162,n175);
and (n244,n163,n169);
or (n245,n246,n247);
and (n246,n97,n161);
and (n247,n98,n112);
nand (n248,n249,n253);
not (n249,n250);
or (n250,n251,n252);
and (n251,n214,n245);
and (n252,n215,n234);
not (n253,n254);
xor (n254,n255,n282);
xor (n255,n256,n259);
or (n256,n257,n258);
and (n257,n216,n228);
and (n258,n217,n222);
xor (n259,n260,n273);
xor (n260,n261,n267);
nand (n261,n262,n263);
or (n262,n151,n239);
or (n263,n264,n139);
nor (n264,n265,n266);
and (n265,n26,n92);
and (n266,n27,n94);
nand (n267,n268,n269);
or (n268,n23,n231);
or (n269,n24,n270);
nor (n270,n271,n272);
and (n271,n33,n64);
and (n272,n34,n66);
nor (n273,n274,n277);
and (n274,n275,n276);
not (n275,n49);
not (n276,n225);
and (n277,n278,n279);
not (n278,n50);
nand (n279,n280,n281);
or (n280,n60,n111);
or (n281,n59,n109);
or (n282,n283,n284);
and (n283,n235,n242);
and (n284,n236,n99);
nand (n285,n286,n290);
not (n286,n287);
or (n287,n288,n289);
and (n288,n255,n282);
and (n289,n256,n259);
not (n290,n291);
xor (n291,n292,n310);
xor (n292,n293,n294);
not (n293,n273);
xor (n294,n295,n304);
xor (n295,n296,n298);
nand (n296,n297,n279);
or (n297,n275,n278);
nand (n298,n299,n300);
or (n299,n151,n264);
or (n300,n139,n301);
nor (n301,n302,n303);
and (n302,n26,n103);
and (n303,n27,n105);
nand (n304,n305,n306);
or (n305,n23,n270);
or (n306,n24,n307);
nor (n307,n308,n309);
and (n308,n33,n70);
and (n309,n34,n72);
or (n310,n311,n312);
and (n311,n260,n273);
and (n312,n261,n267);
nand (n313,n314,n318);
not (n314,n315);
or (n315,n316,n317);
and (n316,n292,n310);
and (n317,n293,n294);
not (n318,n319);
xor (n319,n320,n335);
xor (n320,n321,n328);
nand (n321,n322,n327);
or (n322,n323,n139);
not (n323,n324);
nand (n324,n325,n326);
or (n325,n27,n111);
or (n326,n26,n109);
or (n327,n151,n301);
not (n328,n329);
nand (n329,n330,n331);
or (n330,n23,n307);
or (n331,n24,n332);
nor (n332,n333,n334);
and (n333,n33,n92);
and (n334,n34,n94);
or (n335,n336,n337);
and (n336,n295,n304);
and (n337,n296,n298);
not (n338,n339);
nand (n339,n340,n1065);
nor (n340,n341,n1053);
and (n341,n342,n956);
not (n342,n343);
nor (n343,n344,n955);
and (n344,n345,n888);
nand (n345,n346,n726);
not (n346,n347);
and (n347,n348,n658);
xor (n348,n349,n583);
xor (n349,n350,n464);
xor (n350,n351,n414);
xor (n351,n352,n391);
or (n352,n353,n390);
and (n353,n354,n377);
xor (n354,n355,n364);
nand (n355,n356,n360);
or (n356,n126,n357);
nor (n357,n358,n359);
and (n358,n78,n148);
and (n359,n79,n147);
or (n360,n118,n361);
nor (n361,n362,n363);
and (n362,n78,n64);
and (n363,n79,n66);
nand (n364,n365,n371);
or (n365,n151,n366);
nor (n366,n367,n369);
and (n367,n368,n26);
and (n369,n27,n370);
not (n370,n368);
or (n371,n372,n139);
nor (n372,n373,n375);
and (n373,n374,n26);
and (n375,n27,n376);
not (n376,n374);
nand (n377,n378,n384);
or (n378,n23,n379);
nor (n379,n380,n382);
and (n380,n381,n33);
and (n382,n34,n383);
not (n383,n381);
or (n384,n385,n24);
nor (n385,n386,n388);
and (n386,n387,n33);
and (n388,n34,n389);
not (n389,n387);
and (n390,n355,n364);
xor (n391,n392,n408);
xor (n392,n393,n402);
nand (n393,n394,n398);
or (n394,n49,n395);
nor (n395,n396,n397);
and (n396,n38,n59);
and (n397,n60,n40);
or (n398,n399,n50);
nor (n399,n400,n401);
and (n400,n44,n59);
and (n401,n60,n46);
nand (n402,n403,n404);
or (n403,n126,n361);
or (n404,n118,n405);
nor (n405,n406,n407);
and (n406,n78,n70);
and (n407,n79,n72);
nand (n408,n409,n410);
or (n409,n151,n372);
or (n410,n411,n139);
nor (n411,n412,n413);
and (n412,n197,n26);
and (n413,n27,n199);
xor (n414,n415,n454);
xor (n415,n416,n436);
nand (n416,n417,n431);
or (n417,n418,n424);
nand (n418,n419,n423);
or (n419,n420,n422);
not (n420,n421);
nand (n423,n420,n422);
not (n424,n425);
nand (n425,n426,n427);
not (n426,n418);
nand (n427,n428,n430);
or (n428,n420,n429);
nand (n430,n429,n420);
not (n431,n432);
nor (n432,n433,n435);
and (n433,n434,n109);
not (n434,n429);
and (n435,n429,n111);
nand (n436,n437,n450);
or (n437,n438,n447);
nand (n438,n439,n444);
nor (n439,n440,n443);
and (n440,n441,n429);
not (n441,n442);
and (n443,n442,n434);
nand (n444,n445,n446);
or (n445,n442,n120);
nand (n446,n120,n442);
nor (n447,n448,n449);
and (n448,n120,n92);
and (n449,n121,n94);
or (n450,n439,n451);
nor (n451,n452,n453);
and (n452,n120,n103);
and (n453,n121,n105);
nand (n454,n455,n460);
or (n455,n456,n76);
not (n456,n457);
nand (n457,n458,n459);
or (n458,n53,n147);
or (n459,n52,n148);
or (n460,n75,n461);
nor (n461,n462,n463);
and (n462,n52,n157);
and (n463,n53,n159);
xor (n464,n465,n553);
xor (n465,n466,n503);
xor (n466,n467,n480);
xor (n467,n468,n474);
nand (n468,n469,n470);
or (n469,n23,n385);
or (n470,n471,n24);
nor (n471,n472,n473);
and (n472,n33,n368);
and (n473,n34,n370);
nand (n474,n475,n479);
or (n475,n425,n476);
nor (n476,n477,n478);
and (n477,n434,n103);
and (n478,n429,n105);
or (n479,n426,n432);
or (n480,n481,n502);
and (n481,n482,n496);
xor (n482,n483,n490);
nand (n483,n484,n489);
or (n484,n485,n438);
not (n485,n486);
nand (n486,n487,n488);
or (n487,n121,n72);
or (n488,n120,n70);
or (n489,n439,n447);
nand (n490,n491,n495);
or (n491,n75,n492);
nor (n492,n493,n494);
and (n493,n52,n44);
and (n494,n53,n46);
or (n495,n76,n461);
nand (n496,n497,n501);
or (n497,n49,n498);
nor (n498,n499,n500);
and (n499,n197,n59);
and (n500,n60,n199);
or (n501,n50,n395);
and (n502,n483,n490);
or (n503,n504,n552);
and (n504,n505,n527);
xor (n505,n506,n507);
not (n506,n474);
nand (n507,n508,n520);
not (n508,n509);
nand (n509,n510,n515);
or (n510,n511,n514);
not (n511,n512);
nand (n512,n513,n422);
not (n513,n514);
not (n515,n516);
nor (n516,n517,n519);
and (n517,n518,n109);
not (n518,n422);
and (n519,n422,n111);
not (n520,n521);
nand (n521,n522,n526);
or (n522,n425,n523);
nor (n523,n524,n525);
and (n524,n434,n92);
and (n525,n429,n94);
or (n526,n426,n476);
or (n527,n528,n551);
and (n528,n529,n544);
xor (n529,n530,n538);
nand (n530,n531,n537);
or (n531,n23,n532);
nor (n532,n533,n535);
and (n533,n534,n33);
and (n535,n536,n34);
not (n536,n534);
or (n537,n379,n24);
nand (n538,n539,n543);
or (n539,n126,n540);
nor (n540,n541,n542);
and (n541,n78,n157);
and (n542,n79,n159);
or (n543,n118,n357);
nand (n544,n545,n550);
or (n545,n75,n546);
not (n546,n547);
nor (n547,n548,n549);
and (n548,n40,n52);
and (n549,n38,n53);
or (n550,n492,n76);
and (n551,n530,n538);
and (n552,n506,n507);
or (n553,n554,n582);
and (n554,n555,n581);
xor (n555,n556,n580);
or (n556,n557,n579);
and (n557,n558,n573);
xor (n558,n559,n567);
nand (n559,n560,n561);
or (n560,n439,n485);
nand (n561,n562,n566);
not (n562,n563);
nor (n563,n564,n565);
and (n564,n64,n120);
and (n565,n66,n121);
not (n566,n438);
nand (n567,n568,n572);
or (n568,n49,n569);
nor (n569,n570,n571);
and (n570,n374,n59);
and (n571,n60,n376);
or (n572,n498,n50);
nand (n573,n574,n578);
or (n574,n151,n575);
nor (n575,n576,n577);
and (n576,n387,n26);
and (n577,n27,n389);
or (n578,n366,n139);
and (n579,n559,n567);
xor (n580,n354,n377);
xor (n581,n482,n496);
and (n582,n556,n580);
or (n583,n584,n657);
and (n584,n585,n649);
xor (n585,n586,n648);
or (n586,n587,n647);
and (n587,n588,n625);
xor (n588,n589,n603);
and (n589,n590,n597);
nor (n590,n591,n33);
nor (n591,n592,n595);
and (n592,n593,n26);
nand (n593,n594,n28);
and (n595,n596,n30);
not (n596,n594);
nand (n597,n598,n602);
or (n598,n599,n512);
nor (n599,n600,n601);
and (n600,n103,n518);
and (n601,n105,n422);
or (n602,n516,n513);
or (n603,n604,n624);
and (n604,n605,n618);
xor (n605,n606,n612);
nand (n606,n607,n611);
or (n607,n425,n608);
nor (n608,n609,n610);
and (n609,n434,n70);
and (n610,n429,n72);
or (n611,n426,n523);
nand (n612,n613,n617);
or (n613,n23,n614);
nor (n614,n615,n616);
and (n615,n596,n34);
and (n616,n594,n33);
or (n617,n532,n24);
nand (n618,n619,n623);
or (n619,n126,n620);
nor (n620,n621,n622);
and (n621,n78,n44);
and (n622,n79,n46);
or (n623,n118,n540);
and (n624,n606,n612);
or (n625,n626,n646);
and (n626,n627,n640);
xor (n627,n628,n634);
nand (n628,n629,n630);
or (n629,n76,n546);
or (n630,n75,n631);
nor (n631,n632,n633);
and (n632,n52,n197);
and (n633,n53,n199);
nand (n634,n635,n639);
or (n635,n438,n636);
nor (n636,n637,n638);
and (n637,n120,n148);
and (n638,n121,n147);
or (n639,n439,n563);
nand (n640,n641,n645);
or (n641,n49,n642);
nor (n642,n643,n644);
and (n643,n59,n368);
and (n644,n60,n370);
or (n645,n50,n569);
and (n646,n628,n634);
and (n647,n589,n603);
xor (n648,n505,n527);
or (n649,n650,n656);
and (n650,n651,n655);
xor (n651,n652,n653);
xor (n652,n558,n573);
nand (n653,n654,n507);
or (n654,n508,n520);
xor (n655,n529,n544);
and (n656,n652,n653);
and (n657,n586,n648);
or (n658,n659,n725);
and (n659,n660,n724);
xor (n660,n661,n662);
xor (n661,n555,n581);
or (n662,n663,n723);
and (n663,n664,n695);
xor (n664,n665,n694);
or (n665,n666,n693);
and (n666,n667,n676);
xor (n667,n668,n675);
nand (n668,n669,n674);
or (n669,n151,n670);
not (n670,n671);
nand (n671,n672,n673);
or (n672,n383,n27);
or (n673,n26,n381);
or (n674,n575,n139);
xor (n675,n590,n597);
or (n676,n677,n692);
and (n677,n678,n686);
xor (n678,n679,n680);
nor (n679,n24,n596);
nand (n680,n681,n685);
or (n681,n682,n512);
nor (n682,n683,n684);
and (n683,n422,n94);
nor (n684,n422,n94);
or (n685,n599,n513);
nand (n686,n687,n691);
or (n687,n425,n688);
nor (n688,n689,n690);
and (n689,n434,n64);
and (n690,n429,n66);
or (n691,n426,n608);
and (n692,n679,n680);
and (n693,n668,n675);
xor (n694,n588,n625);
or (n695,n696,n722);
and (n696,n697,n721);
xor (n697,n698,n720);
or (n698,n699,n719);
and (n699,n700,n713);
xor (n700,n701,n707);
nand (n701,n702,n706);
or (n702,n126,n703);
nor (n703,n704,n705);
and (n704,n38,n78);
and (n705,n79,n40);
or (n706,n620,n118);
nand (n707,n708,n712);
or (n708,n75,n709);
nor (n709,n710,n711);
and (n710,n52,n374);
and (n711,n53,n376);
or (n712,n631,n76);
nand (n713,n714,n718);
or (n714,n438,n715);
nor (n715,n716,n717);
and (n716,n120,n157);
and (n717,n121,n159);
or (n718,n439,n636);
and (n719,n701,n707);
xor (n720,n627,n640);
xor (n721,n605,n618);
and (n722,n698,n720);
and (n723,n665,n694);
xor (n724,n585,n649);
and (n725,n661,n662);
nand (n726,n727,n887);
nand (n727,n728,n886);
or (n728,n729,n823);
nor (n729,n730,n731);
xor (n730,n660,n724);
or (n731,n732,n822);
and (n732,n733,n821);
xor (n733,n734,n735);
xor (n734,n651,n655);
or (n735,n736,n820);
and (n736,n737,n769);
xor (n737,n738,n768);
or (n738,n739,n767);
and (n739,n740,n755);
xor (n740,n741,n747);
nand (n741,n742,n746);
or (n742,n49,n743);
nor (n743,n744,n745);
and (n744,n387,n59);
and (n745,n60,n389);
or (n746,n50,n642);
nand (n747,n748,n749);
or (n748,n139,n670);
nand (n749,n750,n754);
not (n750,n751);
nor (n751,n752,n753);
and (n752,n26,n534);
and (n753,n536,n27);
not (n754,n151);
and (n755,n756,n761);
nor (n756,n757,n26);
nor (n757,n758,n760);
and (n758,n759,n59);
nand (n759,n142,n594);
and (n760,n596,n141);
nand (n761,n762,n766);
or (n762,n763,n512);
nor (n763,n764,n765);
and (n764,n518,n70);
and (n765,n422,n72);
or (n766,n682,n513);
and (n767,n741,n747);
xor (n768,n667,n676);
or (n769,n770,n819);
and (n770,n771,n818);
xor (n771,n772,n796);
or (n772,n773,n795);
and (n773,n774,n788);
xor (n774,n775,n781);
nand (n775,n776,n780);
or (n776,n425,n777);
nor (n777,n778,n779);
and (n778,n148,n434);
and (n779,n147,n429);
or (n780,n426,n688);
nand (n781,n782,n787);
or (n782,n783,n126);
not (n783,n784);
nand (n784,n785,n786);
or (n785,n79,n199);
or (n786,n78,n197);
or (n787,n703,n118);
nand (n788,n789,n794);
or (n789,n75,n790);
not (n790,n791);
nor (n791,n792,n793);
and (n792,n370,n52);
and (n793,n368,n53);
or (n794,n709,n76);
and (n795,n775,n781);
or (n796,n797,n817);
and (n797,n798,n811);
xor (n798,n799,n805);
nand (n799,n800,n804);
or (n800,n438,n801);
nor (n801,n802,n803);
and (n802,n120,n44);
and (n803,n121,n46);
or (n804,n439,n715);
nand (n805,n806,n810);
or (n806,n49,n807);
nor (n807,n808,n809);
and (n808,n381,n59);
and (n809,n60,n383);
or (n810,n743,n50);
nand (n811,n812,n816);
or (n812,n151,n813);
nor (n813,n814,n815);
and (n814,n596,n27);
and (n815,n594,n26);
or (n816,n751,n139);
and (n817,n799,n805);
xor (n818,n678,n686);
and (n819,n772,n796);
and (n820,n738,n768);
xor (n821,n664,n695);
and (n822,n734,n735);
nand (n823,n824,n825);
xor (n824,n733,n821);
or (n825,n826,n885);
and (n826,n827,n884);
xor (n827,n828,n829);
xor (n828,n697,n721);
or (n829,n830,n883);
and (n830,n831,n834);
xor (n831,n832,n833);
xor (n832,n700,n713);
xor (n833,n740,n755);
or (n834,n835,n882);
and (n835,n836,n859);
xor (n836,n837,n838);
xor (n837,n756,n761);
or (n838,n839,n858);
and (n839,n840,n851);
xor (n840,n841,n843);
and (n841,n842,n594);
not (n842,n139);
nand (n843,n844,n849);
or (n844,n845,n425);
not (n845,n846);
nand (n846,n847,n848);
or (n847,n429,n159);
or (n848,n434,n157);
nand (n849,n850,n418);
not (n850,n777);
nand (n851,n852,n857);
or (n852,n126,n853);
not (n853,n854);
nand (n854,n855,n856);
or (n855,n79,n376);
or (n856,n78,n374);
or (n857,n118,n783);
and (n858,n841,n843);
or (n859,n860,n881);
and (n860,n861,n875);
xor (n861,n862,n869);
nand (n862,n863,n868);
or (n863,n864,n75);
not (n864,n865);
nand (n865,n866,n867);
or (n866,n53,n389);
or (n867,n52,n387);
nand (n868,n791,n220);
nand (n869,n870,n871);
or (n870,n513,n763);
or (n871,n872,n512);
nor (n872,n873,n874);
and (n873,n518,n64);
and (n874,n422,n66);
nand (n875,n876,n880);
or (n876,n877,n49);
nor (n877,n878,n879);
and (n878,n534,n59);
and (n879,n60,n536);
or (n880,n807,n50);
and (n881,n862,n869);
and (n882,n837,n838);
and (n883,n832,n833);
xor (n884,n737,n769);
and (n885,n828,n829);
nand (n886,n730,n731);
or (n887,n348,n658);
or (n888,n889,n892);
or (n889,n890,n891);
and (n890,n349,n583);
and (n891,n350,n464);
xor (n892,n893,n952);
xor (n893,n894,n922);
xor (n894,n895,n902);
xor (n895,n896,n899);
or (n896,n897,n898);
and (n897,n392,n408);
and (n898,n393,n402);
or (n899,n900,n901);
and (n900,n415,n454);
and (n901,n416,n436);
xor (n902,n903,n916);
xor (n903,n904,n910);
nand (n904,n905,n906);
or (n905,n49,n399);
or (n906,n50,n907);
nor (n907,n908,n909);
and (n908,n59,n157);
and (n909,n60,n159);
nand (n910,n911,n912);
or (n911,n151,n411);
or (n912,n913,n139);
nor (n913,n914,n915);
and (n914,n26,n38);
and (n915,n27,n40);
nand (n916,n917,n918);
or (n917,n438,n451);
or (n918,n439,n919);
nor (n919,n920,n921);
and (n920,n120,n109);
and (n921,n121,n111);
xor (n922,n923,n949);
xor (n923,n924,n946);
xor (n924,n925,n939);
xor (n925,n926,n932);
nand (n926,n927,n928);
or (n927,n23,n471);
or (n928,n929,n24);
nor (n929,n930,n931);
and (n930,n374,n33);
and (n931,n34,n376);
nand (n932,n933,n934);
or (n933,n456,n75);
nand (n934,n935,n220);
not (n935,n936);
nor (n936,n937,n938);
and (n937,n52,n64);
and (n938,n53,n66);
not (n939,n940);
nand (n940,n941,n942);
or (n941,n126,n405);
or (n942,n118,n943);
nor (n943,n944,n945);
and (n944,n78,n92);
and (n945,n79,n94);
or (n946,n947,n948);
and (n947,n467,n480);
and (n948,n468,n474);
or (n949,n950,n951);
and (n950,n351,n414);
and (n951,n352,n391);
or (n952,n953,n954);
and (n953,n465,n553);
and (n954,n466,n503);
and (n955,n892,n889);
not (n956,n957);
nand (n957,n958,n1029,n1048);
not (n958,n959);
nor (n959,n960,n1007);
xor (n960,n961,n987);
xor (n961,n962,n986);
or (n962,n963,n985);
and (n963,n964,n972);
xor (n964,n965,n971);
nand (n965,n966,n970);
or (n966,n49,n967);
nor (n967,n968,n969);
and (n968,n59,n148);
and (n969,n60,n147);
or (n970,n50,n62);
not (n971,n73);
or (n972,n973,n984);
and (n973,n974,n981);
xor (n974,n975,n978);
nand (n975,n976,n977);
or (n976,n151,n913);
or (n977,n189,n139);
nand (n978,n979,n980);
or (n979,n75,n936);
or (n980,n76,n86);
nand (n981,n982,n983);
or (n982,n23,n929);
or (n983,n195,n24);
and (n984,n975,n978);
and (n985,n965,n971);
xor (n986,n183,n209);
or (n987,n988,n1006);
and (n988,n989,n1005);
xor (n989,n990,n1004);
or (n990,n991,n1003);
and (n991,n992,n1000);
xor (n992,n993,n997);
nand (n993,n994,n996);
or (n994,n566,n995);
not (n995,n439);
not (n996,n919);
nand (n997,n998,n999);
or (n998,n126,n943);
or (n999,n118,n203);
nand (n1000,n1001,n1002);
or (n1001,n49,n907);
or (n1002,n50,n967);
and (n1003,n993,n997);
xor (n1004,n186,n201);
xor (n1005,n964,n972);
and (n1006,n990,n1004);
or (n1007,n1008,n1028);
and (n1008,n1009,n1019);
xor (n1009,n1010,n1018);
or (n1010,n1011,n1017);
and (n1011,n1012,n1016);
xor (n1012,n940,n1013);
or (n1013,n1014,n1015);
and (n1014,n903,n916);
and (n1015,n904,n910);
xor (n1016,n974,n981);
and (n1017,n940,n1013);
xor (n1018,n989,n1005);
or (n1019,n1020,n1027);
and (n1020,n1021,n1026);
xor (n1021,n1022,n1023);
xor (n1022,n992,n1000);
or (n1023,n1024,n1025);
and (n1024,n925,n939);
and (n1025,n926,n932);
xor (n1026,n1012,n1016);
and (n1027,n1022,n1023);
and (n1028,n1010,n1018);
nor (n1029,n1030,n1043);
nor (n1030,n1031,n1034);
or (n1031,n1032,n1033);
and (n1032,n893,n952);
and (n1033,n894,n922);
xor (n1034,n1035,n1040);
xor (n1035,n1036,n1039);
or (n1036,n1037,n1038);
and (n1037,n895,n902);
and (n1038,n896,n899);
xor (n1039,n1021,n1026);
or (n1040,n1041,n1042);
and (n1041,n923,n949);
and (n1042,n924,n946);
nor (n1043,n1044,n1047);
or (n1044,n1045,n1046);
and (n1045,n1035,n1040);
and (n1046,n1036,n1039);
xor (n1047,n1009,n1019);
or (n1048,n1049,n1052);
or (n1049,n1050,n1051);
and (n1050,n961,n987);
and (n1051,n962,n986);
xor (n1052,n17,n181);
nand (n1053,n1054,n1064);
or (n1054,n1055,n1056);
not (n1055,n1048);
not (n1056,n1057);
nand (n1057,n1058,n1063);
nand (n1058,n958,n1059);
nand (n1059,n1060,n1062);
or (n1060,n1061,n1043);
nand (n1061,n1031,n1034);
nand (n1062,n1044,n1047);
nand (n1063,n1007,n960);
nand (n1064,n1049,n1052);
nand (n1065,n1066,n1566);
or (n1066,n1067,n1565);
and (n1067,n1068,n1131);
xor (n1068,n1069,n1130);
or (n1069,n1070,n1129);
and (n1070,n1071,n1074);
xor (n1071,n1072,n1073);
xor (n1072,n771,n818);
xor (n1073,n831,n834);
or (n1074,n1075,n1128);
and (n1075,n1076,n1079);
xor (n1076,n1077,n1078);
xor (n1077,n798,n811);
xor (n1078,n774,n788);
or (n1079,n1080,n1127);
and (n1080,n1081,n1102);
xor (n1081,n1082,n1088);
nand (n1082,n1083,n1087);
or (n1083,n438,n1084);
nor (n1084,n1085,n1086);
and (n1085,n120,n38);
and (n1086,n121,n40);
or (n1087,n439,n801);
nor (n1088,n1089,n1096);
not (n1089,n1090);
nand (n1090,n1091,n1095);
or (n1091,n1092,n425);
nor (n1092,n1093,n1094);
and (n1093,n44,n434);
and (n1094,n46,n429);
nand (n1095,n418,n846);
nand (n1096,n1097,n60);
nand (n1097,n1098,n1099);
or (n1098,n594,n54);
nand (n1099,n1100,n52);
not (n1100,n1101);
and (n1101,n594,n54);
or (n1102,n1103,n1126);
and (n1103,n1104,n1119);
xor (n1104,n1105,n1112);
nand (n1105,n1106,n1107);
or (n1106,n118,n853);
nand (n1107,n1108,n125);
not (n1108,n1109);
nor (n1109,n1110,n1111);
and (n1110,n370,n79);
and (n1111,n368,n78);
nand (n1112,n1113,n1118);
or (n1113,n1114,n75);
not (n1114,n1115);
nor (n1115,n1116,n1117);
and (n1116,n52,n383);
and (n1117,n381,n53);
nand (n1118,n220,n865);
nand (n1119,n1120,n1125);
or (n1120,n1121,n512);
not (n1121,n1122);
or (n1122,n1123,n1124);
and (n1123,n147,n422);
and (n1124,n148,n518);
or (n1125,n872,n513);
and (n1126,n1105,n1112);
and (n1127,n1082,n1088);
and (n1128,n1077,n1078);
and (n1129,n1072,n1073);
xor (n1130,n827,n884);
or (n1131,n1132,n1564);
and (n1132,n1133,n1167);
xor (n1133,n1134,n1166);
or (n1134,n1135,n1165);
and (n1135,n1136,n1164);
xor (n1136,n1137,n1138);
xor (n1137,n836,n859);
or (n1138,n1139,n1163);
and (n1139,n1140,n1143);
xor (n1140,n1141,n1142);
xor (n1141,n861,n875);
xor (n1142,n840,n851);
or (n1143,n1144,n1162);
and (n1144,n1145,n1158);
xor (n1145,n1146,n1152);
nand (n1146,n1147,n1151);
or (n1147,n49,n1148);
nor (n1148,n1149,n1150);
and (n1149,n596,n60);
and (n1150,n594,n59);
or (n1151,n877,n50);
nand (n1152,n1153,n1157);
or (n1153,n438,n1154);
nor (n1154,n1155,n1156);
and (n1155,n120,n197);
and (n1156,n121,n199);
or (n1157,n439,n1084);
nand (n1158,n1159,n1161);
or (n1159,n1160,n1089);
not (n1160,n1096);
or (n1161,n1090,n1096);
and (n1162,n1146,n1152);
and (n1163,n1141,n1142);
xor (n1164,n1076,n1079);
and (n1165,n1137,n1138);
xor (n1166,n1071,n1074);
nand (n1167,n1168,n1560);
or (n1168,n1169,n1538);
nor (n1169,n1170,n1537);
and (n1170,n1171,n1518);
or (n1171,n1172,n1517);
and (n1172,n1173,n1315);
xor (n1173,n1174,n1284);
or (n1174,n1175,n1283);
and (n1175,n1176,n1246);
xor (n1176,n1177,n1207);
xor (n1177,n1178,n1197);
xor (n1178,n1179,n1188);
nand (n1179,n1180,n1184);
or (n1180,n126,n1181);
nor (n1181,n1182,n1183);
and (n1182,n381,n78);
and (n1183,n383,n79);
or (n1184,n1185,n118);
nor (n1185,n1186,n1187);
and (n1186,n78,n387);
and (n1187,n79,n389);
nand (n1188,n1189,n1193);
or (n1189,n75,n1190);
nor (n1190,n1191,n1192);
and (n1191,n596,n53);
and (n1192,n594,n52);
or (n1193,n1194,n76);
nor (n1194,n1195,n1196);
and (n1195,n534,n52);
and (n1196,n536,n53);
nand (n1197,n1198,n1203);
or (n1198,n512,n1199);
not (n1199,n1200);
nor (n1200,n1201,n1202);
and (n1201,n44,n422);
and (n1202,n46,n518);
or (n1203,n1204,n513);
nor (n1204,n1205,n1206);
and (n1205,n157,n518);
and (n1206,n159,n422);
or (n1207,n1208,n1245);
and (n1208,n1209,n1228);
xor (n1209,n1210,n1219);
nand (n1210,n1211,n1215);
or (n1211,n425,n1212);
nor (n1212,n1213,n1214);
and (n1213,n434,n374);
and (n1214,n429,n376);
or (n1215,n426,n1216);
nor (n1216,n1217,n1218);
and (n1217,n199,n429);
and (n1218,n197,n434);
nand (n1219,n1220,n1224);
or (n1220,n438,n1221);
nor (n1221,n1222,n1223);
and (n1222,n387,n120);
and (n1223,n121,n389);
or (n1224,n439,n1225);
nor (n1225,n1226,n1227);
and (n1226,n120,n368);
and (n1227,n121,n370);
and (n1228,n1229,n1235);
nor (n1229,n1230,n78);
nor (n1230,n1231,n1234);
and (n1231,n1232,n120);
not (n1232,n1233);
and (n1233,n594,n122);
and (n1234,n596,n124);
nand (n1235,n1236,n1241);
or (n1236,n1237,n512);
not (n1237,n1238);
nor (n1238,n1239,n1240);
and (n1239,n199,n518);
and (n1240,n197,n422);
or (n1241,n1242,n513);
nor (n1242,n1243,n1244);
and (n1243,n38,n518);
and (n1244,n40,n422);
and (n1245,n1210,n1219);
xor (n1246,n1247,n1268);
xor (n1247,n1248,n1254);
nand (n1248,n1249,n1250);
or (n1249,n438,n1225);
or (n1250,n439,n1251);
nor (n1251,n1252,n1253);
and (n1252,n120,n374);
and (n1253,n121,n376);
xor (n1254,n1255,n1260);
nor (n1255,n1256,n52);
nor (n1256,n1257,n1259);
and (n1257,n1258,n78);
nand (n1258,n594,n80);
and (n1259,n596,n82);
nand (n1260,n1261,n1266);
or (n1261,n426,n1262);
not (n1262,n1263);
nand (n1263,n1264,n1265);
or (n1264,n429,n40);
or (n1265,n434,n38);
nand (n1266,n1267,n424);
not (n1267,n1216);
or (n1268,n1269,n1282);
and (n1269,n1270,n1275);
xor (n1270,n1271,n1272);
nor (n1271,n76,n596);
nand (n1272,n1273,n1274);
or (n1273,n513,n1199);
or (n1274,n1242,n512);
nand (n1275,n1276,n1277);
or (n1276,n118,n1181);
nand (n1277,n1278,n125);
not (n1278,n1279);
or (n1279,n1280,n1281);
and (n1280,n536,n78);
and (n1281,n534,n79);
and (n1282,n1271,n1272);
and (n1283,n1177,n1207);
xor (n1284,n1285,n1300);
xor (n1285,n1286,n1297);
xor (n1286,n1287,n1294);
xor (n1287,n1288,n1291);
nand (n1288,n1289,n1290);
or (n1289,n76,n1114);
or (n1290,n75,n1194);
nand (n1291,n1292,n1293);
or (n1292,n1204,n512);
nand (n1293,n1122,n514);
nand (n1294,n1295,n1296);
or (n1295,n438,n1251);
or (n1296,n439,n1154);
or (n1297,n1298,n1299);
and (n1298,n1247,n1268);
and (n1299,n1248,n1254);
xor (n1300,n1301,n1306);
xor (n1301,n1302,n1303);
and (n1302,n1255,n1260);
or (n1303,n1304,n1305);
and (n1304,n1178,n1197);
and (n1305,n1179,n1188);
xor (n1306,n1307,n1312);
xor (n1307,n1308,n1309);
nor (n1308,n50,n596);
nand (n1309,n1310,n1311);
or (n1310,n1262,n425);
or (n1311,n426,n1092);
nand (n1312,n1313,n1314);
or (n1313,n126,n1185);
or (n1314,n118,n1109);
nand (n1315,n1316,n1513,n1516);
nand (n1316,n1317,n1371,n1506);
not (n1317,n1318);
nor (n1318,n1319,n1346);
xor (n1319,n1320,n1345);
xor (n1320,n1321,n1344);
or (n1321,n1322,n1343);
and (n1322,n1323,n1337);
xor (n1323,n1324,n1330);
nand (n1324,n1325,n1329);
or (n1325,n126,n1326);
nor (n1326,n1327,n1328);
and (n1327,n596,n79);
and (n1328,n594,n78);
or (n1329,n1279,n118);
nand (n1330,n1331,n1336);
or (n1331,n1332,n425);
not (n1332,n1333);
nor (n1333,n1334,n1335);
and (n1334,n368,n429);
and (n1335,n370,n434);
or (n1336,n426,n1212);
nand (n1337,n1338,n1342);
or (n1338,n438,n1339);
nor (n1339,n1340,n1341);
and (n1340,n381,n120);
and (n1341,n121,n383);
or (n1342,n439,n1221);
and (n1343,n1324,n1330);
xor (n1344,n1270,n1275);
xor (n1345,n1209,n1228);
or (n1346,n1347,n1370);
and (n1347,n1348,n1369);
xor (n1348,n1349,n1350);
xor (n1349,n1229,n1235);
or (n1350,n1351,n1368);
and (n1351,n1352,n1361);
xor (n1352,n1353,n1354);
and (n1353,n117,n594);
nand (n1354,n1355,n1360);
or (n1355,n512,n1356);
not (n1356,n1357);
nor (n1357,n1358,n1359);
and (n1358,n376,n518);
and (n1359,n374,n422);
nand (n1360,n1238,n514);
nand (n1361,n1362,n1367);
or (n1362,n1363,n425);
not (n1363,n1364);
nor (n1364,n1365,n1366);
and (n1365,n389,n434);
and (n1366,n387,n429);
nand (n1367,n1333,n418);
and (n1368,n1353,n1354);
xor (n1369,n1323,n1337);
and (n1370,n1349,n1350);
or (n1371,n1372,n1505);
and (n1372,n1373,n1399);
xor (n1373,n1374,n1398);
or (n1374,n1375,n1397);
and (n1375,n1376,n1396);
xor (n1376,n1377,n1383);
nand (n1377,n1378,n1382);
or (n1378,n438,n1379);
nor (n1379,n1380,n1381);
and (n1380,n120,n534);
and (n1381,n121,n536);
or (n1382,n1339,n439);
and (n1383,n1384,n1390);
and (n1384,n1385,n121);
nand (n1385,n1386,n1387);
or (n1386,n594,n442);
nand (n1387,n1388,n434);
not (n1388,n1389);
and (n1389,n594,n442);
nand (n1390,n1391,n1392);
or (n1391,n513,n1356);
or (n1392,n1393,n512);
nor (n1393,n1394,n1395);
and (n1394,n518,n368);
and (n1395,n422,n370);
xor (n1396,n1352,n1361);
and (n1397,n1377,n1383);
xor (n1398,n1348,n1369);
nand (n1399,n1400,n1504);
or (n1400,n1401,n1499);
nor (n1401,n1402,n1498);
and (n1402,n1403,n1477);
nand (n1403,n1404,n1475);
or (n1404,n1405,n1459);
not (n1405,n1406);
or (n1406,n1407,n1458);
and (n1407,n1408,n1437);
xor (n1408,n1409,n1418);
nand (n1409,n1410,n1414);
or (n1410,n425,n1411);
nor (n1411,n1412,n1413);
and (n1412,n429,n596);
and (n1413,n594,n434);
or (n1414,n426,n1415);
nor (n1415,n1416,n1417);
and (n1416,n536,n429);
and (n1417,n534,n434);
nand (n1418,n1419,n1436);
or (n1419,n1420,n1426);
not (n1420,n1421);
nand (n1421,n1422,n429);
nand (n1422,n1423,n1425);
or (n1423,n1424,n422);
and (n1424,n594,n421);
nand (n1425,n596,n420);
not (n1426,n1427);
nand (n1427,n1428,n1432);
or (n1428,n1429,n512);
or (n1429,n1430,n1431);
and (n1430,n381,n422);
and (n1431,n383,n518);
or (n1432,n1433,n513);
nor (n1433,n1434,n1435);
and (n1434,n389,n422);
and (n1435,n387,n518);
or (n1436,n1427,n1421);
or (n1437,n1438,n1457);
and (n1438,n1439,n1447);
xor (n1439,n1440,n1441);
nor (n1440,n426,n596);
nand (n1441,n1442,n1446);
or (n1442,n1443,n512);
nor (n1443,n1444,n1445);
and (n1444,n536,n422);
and (n1445,n534,n518);
or (n1446,n1429,n513);
nor (n1447,n1448,n1455);
nor (n1448,n1449,n1451);
and (n1449,n1450,n514);
not (n1450,n1443);
and (n1451,n1452,n511);
nand (n1452,n1453,n1454);
or (n1453,n596,n422);
nand (n1454,n422,n596);
or (n1455,n1456,n518);
and (n1456,n594,n514);
and (n1457,n1440,n1441);
and (n1458,n1409,n1418);
not (n1459,n1460);
nand (n1460,n1461,n1474);
not (n1461,n1462);
xor (n1462,n1463,n1471);
xor (n1463,n1464,n1465);
and (n1464,n995,n594);
nand (n1465,n1466,n1467);
or (n1466,n1415,n425);
nand (n1467,n1468,n418);
nor (n1468,n1469,n1470);
and (n1469,n383,n434);
and (n1470,n381,n429);
nand (n1471,n1472,n1473);
or (n1472,n1433,n512);
or (n1473,n1393,n513);
nand (n1474,n1420,n1427);
nand (n1475,n1476,n1462);
not (n1476,n1474);
nand (n1477,n1478,n1494);
not (n1478,n1479);
xor (n1479,n1480,n1493);
xor (n1480,n1481,n1485);
nand (n1481,n1482,n1484);
or (n1482,n1483,n425);
not (n1483,n1468);
nand (n1484,n1364,n418);
nand (n1485,n1486,n1491);
or (n1486,n1487,n438);
not (n1487,n1488);
nand (n1488,n1489,n1490);
or (n1489,n594,n120);
or (n1490,n596,n121);
nand (n1491,n1492,n995);
not (n1492,n1379);
xor (n1493,n1384,n1390);
not (n1494,n1495);
or (n1495,n1496,n1497);
and (n1496,n1463,n1471);
and (n1497,n1464,n1465);
nor (n1498,n1478,n1494);
nor (n1499,n1500,n1501);
xor (n1500,n1376,n1396);
or (n1501,n1502,n1503);
and (n1502,n1480,n1493);
and (n1503,n1481,n1485);
nand (n1504,n1500,n1501);
and (n1505,n1374,n1398);
nand (n1506,n1507,n1511);
not (n1507,n1508);
or (n1508,n1509,n1510);
and (n1509,n1320,n1345);
and (n1510,n1321,n1344);
not (n1511,n1512);
xor (n1512,n1176,n1246);
nand (n1513,n1514,n1506);
not (n1514,n1515);
nand (n1515,n1319,n1346);
nand (n1516,n1512,n1508);
and (n1517,n1174,n1284);
or (n1518,n1519,n1534);
xor (n1519,n1520,n1531);
xor (n1520,n1521,n1522);
xor (n1521,n1145,n1158);
xor (n1522,n1523,n1530);
xor (n1523,n1524,n1527);
or (n1524,n1525,n1526);
and (n1525,n1307,n1312);
and (n1526,n1308,n1309);
or (n1527,n1528,n1529);
and (n1528,n1287,n1294);
and (n1529,n1288,n1291);
xor (n1530,n1104,n1119);
or (n1531,n1532,n1533);
and (n1532,n1301,n1306);
and (n1533,n1302,n1303);
or (n1534,n1535,n1536);
and (n1535,n1285,n1300);
and (n1536,n1286,n1297);
and (n1537,n1519,n1534);
nand (n1538,n1539,n1553);
not (n1539,n1540);
and (n1540,n1541,n1549);
not (n1541,n1542);
xor (n1542,n1543,n1548);
xor (n1543,n1544,n1545);
xor (n1544,n1081,n1102);
or (n1545,n1546,n1547);
and (n1546,n1523,n1530);
and (n1547,n1524,n1527);
xor (n1548,n1140,n1143);
not (n1549,n1550);
or (n1550,n1551,n1552);
and (n1551,n1520,n1531);
and (n1552,n1521,n1522);
nand (n1553,n1554,n1556);
not (n1554,n1555);
xor (n1555,n1136,n1164);
not (n1556,n1557);
or (n1557,n1558,n1559);
and (n1558,n1543,n1548);
and (n1559,n1544,n1545);
nor (n1560,n1561,n1563);
and (n1561,n1553,n1562);
nor (n1562,n1541,n1549);
nor (n1563,n1554,n1556);
and (n1564,n1134,n1166);
and (n1565,n1069,n1130);
nor (n1566,n1567,n957);
nand (n1567,n1568,n888,n887);
nor (n1568,n729,n1569);
nor (n1569,n825,n824);
nor (n1570,n1571,n1581);
and (n1571,n1572,n313);
nand (n1572,n1573,n1575);
not (n1573,n1574);
nor (n1574,n286,n290);
nand (n1575,n1576,n285);
not (n1576,n1577);
nor (n1577,n1578,n1580);
and (n1578,n1579,n248);
nor (n1579,n14,n212);
nor (n1580,n249,n253);
nor (n1581,n314,n318);
nor (n1582,n1583,n1598);
not (n1583,n1584);
or (n1584,n1585,n1588);
or (n1585,n1586,n1587);
and (n1586,n320,n335);
and (n1587,n321,n328);
xor (n1588,n1589,n329);
xor (n1589,n1590,n1592);
nand (n1590,n1591,n324);
or (n1591,n754,n842);
nand (n1592,n1593,n1594);
or (n1593,n23,n332);
or (n1594,n24,n1595);
nor (n1595,n1596,n1597);
and (n1596,n33,n103);
and (n1597,n34,n105);
and (n1598,n1599,n1603);
not (n1599,n1600);
or (n1600,n1601,n1602);
and (n1601,n1589,n329);
and (n1602,n1590,n1592);
nand (n1603,n1604,n1605);
or (n1604,n23,n1595);
or (n1605,n24,n1606);
nor (n1606,n1607,n1608);
and (n1607,n33,n109);
and (n1608,n34,n111);
nor (n1609,n1610,n1614);
and (n1610,n1611,n1613);
not (n1611,n1612);
nand (n1612,n1585,n1588);
not (n1613,n1598);
nor (n1614,n1599,n1603);
nand (n1615,n1616,n1603);
not (n1616,n1617);
nor (n1617,n1618,n1606);
and (n1618,n23,n24);
nand (n1619,n1620,n1617);
not (n1620,n1603);
and (n1621,n1622,n1);
xor (n1622,n1623,n3345);
xor (n1623,n1624,n3899);
xor (n1624,n1625,n3340);
xor (n1625,n1626,n3892);
xor (n1626,n1627,n3334);
xor (n1627,n1628,n3880);
xor (n1628,n1629,n3328);
xor (n1629,n1630,n3863);
xor (n1630,n1631,n3322);
xor (n1631,n1632,n3841);
xor (n1632,n1633,n3316);
xor (n1633,n1634,n3814);
xor (n1634,n1635,n3310);
xor (n1635,n1636,n3782);
xor (n1636,n1637,n3304);
xor (n1637,n1638,n3745);
xor (n1638,n1639,n3298);
xor (n1639,n1640,n3703);
xor (n1640,n1641,n3292);
xor (n1641,n1642,n3656);
xor (n1642,n1643,n3286);
xor (n1643,n1644,n3604);
xor (n1644,n1645,n3280);
xor (n1645,n1646,n3547);
xor (n1646,n1647,n3274);
xor (n1647,n1648,n3485);
xor (n1648,n1649,n3268);
xor (n1649,n1650,n3418);
xor (n1650,n1651,n3262);
xor (n1651,n1652,n3346);
xor (n1652,n1653,n3253);
xor (n1653,n1654,n3254);
xor (n1654,n1655,n3253);
xor (n1655,n1656,n3156);
xor (n1656,n1657,n3155);
xor (n1657,n1658,n3053);
xor (n1658,n1659,n3052);
xor (n1659,n1660,n2945);
xor (n1660,n1661,n2944);
xor (n1661,n1662,n2832);
xor (n1662,n1663,n2831);
xor (n1663,n1664,n2715);
xor (n1664,n1665,n2714);
xor (n1665,n1666,n2595);
xor (n1666,n1667,n2594);
xor (n1667,n1668,n2467);
xor (n1668,n1669,n2466);
xor (n1669,n1670,n2335);
xor (n1670,n1671,n2334);
xor (n1671,n1672,n2198);
xor (n1672,n1673,n2197);
xor (n1673,n1674,n2055);
xor (n1674,n1675,n2054);
xor (n1675,n1676,n1691);
xor (n1676,n1677,n1690);
xor (n1677,n1678,n1689);
xor (n1678,n1679,n1688);
xor (n1679,n1680,n1687);
xor (n1680,n1681,n1686);
xor (n1681,n1682,n1685);
xor (n1682,n1683,n1684);
and (n1683,n109,n514);
and (n1684,n109,n422);
and (n1685,n1683,n1684);
and (n1686,n109,n421);
and (n1687,n1681,n1686);
and (n1688,n109,n429);
and (n1689,n1679,n1688);
and (n1690,n109,n442);
or (n1691,n1692,n1693);
and (n1692,n1677,n1690);
and (n1693,n1676,n1694);
or (n1694,n1692,n1695);
and (n1695,n1676,n1696);
or (n1696,n1692,n1697);
and (n1697,n1676,n1698);
or (n1698,n1692,n1699);
and (n1699,n1676,n1700);
or (n1700,n1692,n1701);
and (n1701,n1676,n1702);
or (n1702,n1692,n1703);
and (n1703,n1676,n1704);
or (n1704,n1692,n1705);
and (n1705,n1676,n1706);
or (n1706,n1692,n1707);
and (n1707,n1676,n1708);
or (n1708,n1692,n1709);
and (n1709,n1676,n1710);
or (n1710,n1692,n1711);
and (n1711,n1676,n1712);
or (n1712,n1692,n1713);
and (n1713,n1676,n1714);
or (n1714,n1692,n1715);
and (n1715,n1676,n1716);
or (n1716,n1717,n1972);
and (n1717,n1718,n1971);
xor (n1718,n1678,n1719);
or (n1719,n1720,n1891);
and (n1720,n1721,n1890);
xor (n1721,n1680,n1722);
or (n1722,n1723,n1808);
and (n1723,n1724,n1807);
xor (n1724,n1682,n1725);
or (n1725,n1726,n1728);
and (n1726,n1683,n1727);
and (n1727,n103,n422);
and (n1728,n1729,n1730);
xor (n1729,n1683,n1727);
or (n1730,n1731,n1734);
and (n1731,n1732,n1733);
and (n1732,n103,n514);
and (n1733,n92,n422);
and (n1734,n1735,n1736);
xor (n1735,n1732,n1733);
or (n1736,n1737,n1740);
and (n1737,n1738,n1739);
and (n1738,n92,n514);
and (n1739,n70,n422);
and (n1740,n1741,n1742);
xor (n1741,n1738,n1739);
or (n1742,n1743,n1746);
and (n1743,n1744,n1745);
and (n1744,n70,n514);
and (n1745,n64,n422);
and (n1746,n1747,n1748);
xor (n1747,n1744,n1745);
or (n1748,n1749,n1752);
and (n1749,n1750,n1751);
and (n1750,n64,n514);
and (n1751,n148,n422);
and (n1752,n1753,n1754);
xor (n1753,n1750,n1751);
or (n1754,n1755,n1758);
and (n1755,n1756,n1757);
and (n1756,n148,n514);
and (n1757,n157,n422);
and (n1758,n1759,n1760);
xor (n1759,n1756,n1757);
or (n1760,n1761,n1763);
and (n1761,n1762,n1201);
and (n1762,n157,n514);
and (n1763,n1764,n1765);
xor (n1764,n1762,n1201);
or (n1765,n1766,n1769);
and (n1766,n1767,n1768);
and (n1767,n44,n514);
and (n1768,n38,n422);
and (n1769,n1770,n1771);
xor (n1770,n1767,n1768);
or (n1771,n1772,n1774);
and (n1772,n1773,n1240);
and (n1773,n38,n514);
and (n1774,n1775,n1776);
xor (n1775,n1773,n1240);
or (n1776,n1777,n1779);
and (n1777,n1778,n1359);
and (n1778,n197,n514);
and (n1779,n1780,n1781);
xor (n1780,n1778,n1359);
or (n1781,n1782,n1785);
and (n1782,n1783,n1784);
and (n1783,n374,n514);
and (n1784,n368,n422);
and (n1785,n1786,n1787);
xor (n1786,n1783,n1784);
or (n1787,n1788,n1791);
and (n1788,n1789,n1790);
and (n1789,n368,n514);
and (n1790,n387,n422);
and (n1791,n1792,n1793);
xor (n1792,n1789,n1790);
or (n1793,n1794,n1796);
and (n1794,n1795,n1430);
and (n1795,n387,n514);
and (n1796,n1797,n1798);
xor (n1797,n1795,n1430);
or (n1798,n1799,n1802);
and (n1799,n1800,n1801);
and (n1800,n381,n514);
and (n1801,n534,n422);
and (n1802,n1803,n1804);
xor (n1803,n1800,n1801);
and (n1804,n1805,n1806);
and (n1805,n534,n514);
and (n1806,n594,n422);
and (n1807,n103,n421);
and (n1808,n1809,n1810);
xor (n1809,n1724,n1807);
or (n1810,n1811,n1814);
and (n1811,n1812,n1813);
xor (n1812,n1729,n1730);
and (n1813,n92,n421);
and (n1814,n1815,n1816);
xor (n1815,n1812,n1813);
or (n1816,n1817,n1820);
and (n1817,n1818,n1819);
xor (n1818,n1735,n1736);
and (n1819,n70,n421);
and (n1820,n1821,n1822);
xor (n1821,n1818,n1819);
or (n1822,n1823,n1826);
and (n1823,n1824,n1825);
xor (n1824,n1741,n1742);
and (n1825,n64,n421);
and (n1826,n1827,n1828);
xor (n1827,n1824,n1825);
or (n1828,n1829,n1832);
and (n1829,n1830,n1831);
xor (n1830,n1747,n1748);
and (n1831,n148,n421);
and (n1832,n1833,n1834);
xor (n1833,n1830,n1831);
or (n1834,n1835,n1838);
and (n1835,n1836,n1837);
xor (n1836,n1753,n1754);
and (n1837,n157,n421);
and (n1838,n1839,n1840);
xor (n1839,n1836,n1837);
or (n1840,n1841,n1844);
and (n1841,n1842,n1843);
xor (n1842,n1759,n1760);
and (n1843,n44,n421);
and (n1844,n1845,n1846);
xor (n1845,n1842,n1843);
or (n1846,n1847,n1850);
and (n1847,n1848,n1849);
xor (n1848,n1764,n1765);
and (n1849,n38,n421);
and (n1850,n1851,n1852);
xor (n1851,n1848,n1849);
or (n1852,n1853,n1856);
and (n1853,n1854,n1855);
xor (n1854,n1770,n1771);
and (n1855,n197,n421);
and (n1856,n1857,n1858);
xor (n1857,n1854,n1855);
or (n1858,n1859,n1862);
and (n1859,n1860,n1861);
xor (n1860,n1775,n1776);
and (n1861,n374,n421);
and (n1862,n1863,n1864);
xor (n1863,n1860,n1861);
or (n1864,n1865,n1868);
and (n1865,n1866,n1867);
xor (n1866,n1780,n1781);
and (n1867,n368,n421);
and (n1868,n1869,n1870);
xor (n1869,n1866,n1867);
or (n1870,n1871,n1874);
and (n1871,n1872,n1873);
xor (n1872,n1786,n1787);
and (n1873,n387,n421);
and (n1874,n1875,n1876);
xor (n1875,n1872,n1873);
or (n1876,n1877,n1880);
and (n1877,n1878,n1879);
xor (n1878,n1792,n1793);
and (n1879,n381,n421);
and (n1880,n1881,n1882);
xor (n1881,n1878,n1879);
or (n1882,n1883,n1886);
and (n1883,n1884,n1885);
xor (n1884,n1797,n1798);
and (n1885,n534,n421);
and (n1886,n1887,n1888);
xor (n1887,n1884,n1885);
and (n1888,n1889,n1424);
xor (n1889,n1803,n1804);
and (n1890,n103,n429);
and (n1891,n1892,n1893);
xor (n1892,n1721,n1890);
or (n1893,n1894,n1897);
and (n1894,n1895,n1896);
xor (n1895,n1809,n1810);
and (n1896,n92,n429);
and (n1897,n1898,n1899);
xor (n1898,n1895,n1896);
or (n1899,n1900,n1903);
and (n1900,n1901,n1902);
xor (n1901,n1815,n1816);
and (n1902,n70,n429);
and (n1903,n1904,n1905);
xor (n1904,n1901,n1902);
or (n1905,n1906,n1909);
and (n1906,n1907,n1908);
xor (n1907,n1821,n1822);
and (n1908,n64,n429);
and (n1909,n1910,n1911);
xor (n1910,n1907,n1908);
or (n1911,n1912,n1915);
and (n1912,n1913,n1914);
xor (n1913,n1827,n1828);
and (n1914,n148,n429);
and (n1915,n1916,n1917);
xor (n1916,n1913,n1914);
or (n1917,n1918,n1921);
and (n1918,n1919,n1920);
xor (n1919,n1833,n1834);
and (n1920,n157,n429);
and (n1921,n1922,n1923);
xor (n1922,n1919,n1920);
or (n1923,n1924,n1927);
and (n1924,n1925,n1926);
xor (n1925,n1839,n1840);
and (n1926,n44,n429);
and (n1927,n1928,n1929);
xor (n1928,n1925,n1926);
or (n1929,n1930,n1933);
and (n1930,n1931,n1932);
xor (n1931,n1845,n1846);
and (n1932,n38,n429);
and (n1933,n1934,n1935);
xor (n1934,n1931,n1932);
or (n1935,n1936,n1939);
and (n1936,n1937,n1938);
xor (n1937,n1851,n1852);
and (n1938,n197,n429);
and (n1939,n1940,n1941);
xor (n1940,n1937,n1938);
or (n1941,n1942,n1945);
and (n1942,n1943,n1944);
xor (n1943,n1857,n1858);
and (n1944,n374,n429);
and (n1945,n1946,n1947);
xor (n1946,n1943,n1944);
or (n1947,n1948,n1950);
and (n1948,n1949,n1334);
xor (n1949,n1863,n1864);
and (n1950,n1951,n1952);
xor (n1951,n1949,n1334);
or (n1952,n1953,n1955);
and (n1953,n1954,n1366);
xor (n1954,n1869,n1870);
and (n1955,n1956,n1957);
xor (n1956,n1954,n1366);
or (n1957,n1958,n1960);
and (n1958,n1959,n1470);
xor (n1959,n1875,n1876);
and (n1960,n1961,n1962);
xor (n1961,n1959,n1470);
or (n1962,n1963,n1966);
and (n1963,n1964,n1965);
xor (n1964,n1881,n1882);
and (n1965,n534,n429);
and (n1966,n1967,n1968);
xor (n1967,n1964,n1965);
and (n1968,n1969,n1970);
xor (n1969,n1887,n1888);
and (n1970,n594,n429);
and (n1971,n103,n442);
and (n1972,n1973,n1974);
xor (n1973,n1718,n1971);
or (n1974,n1975,n1978);
and (n1975,n1976,n1977);
xor (n1976,n1892,n1893);
and (n1977,n92,n442);
and (n1978,n1979,n1980);
xor (n1979,n1976,n1977);
or (n1980,n1981,n1984);
and (n1981,n1982,n1983);
xor (n1982,n1898,n1899);
and (n1983,n70,n442);
and (n1984,n1985,n1986);
xor (n1985,n1982,n1983);
or (n1986,n1987,n1990);
and (n1987,n1988,n1989);
xor (n1988,n1904,n1905);
and (n1989,n64,n442);
and (n1990,n1991,n1992);
xor (n1991,n1988,n1989);
or (n1992,n1993,n1996);
and (n1993,n1994,n1995);
xor (n1994,n1910,n1911);
and (n1995,n148,n442);
and (n1996,n1997,n1998);
xor (n1997,n1994,n1995);
or (n1998,n1999,n2002);
and (n1999,n2000,n2001);
xor (n2000,n1916,n1917);
and (n2001,n157,n442);
and (n2002,n2003,n2004);
xor (n2003,n2000,n2001);
or (n2004,n2005,n2008);
and (n2005,n2006,n2007);
xor (n2006,n1922,n1923);
and (n2007,n44,n442);
and (n2008,n2009,n2010);
xor (n2009,n2006,n2007);
or (n2010,n2011,n2014);
and (n2011,n2012,n2013);
xor (n2012,n1928,n1929);
and (n2013,n38,n442);
and (n2014,n2015,n2016);
xor (n2015,n2012,n2013);
or (n2016,n2017,n2020);
and (n2017,n2018,n2019);
xor (n2018,n1934,n1935);
and (n2019,n197,n442);
and (n2020,n2021,n2022);
xor (n2021,n2018,n2019);
or (n2022,n2023,n2026);
and (n2023,n2024,n2025);
xor (n2024,n1940,n1941);
and (n2025,n374,n442);
and (n2026,n2027,n2028);
xor (n2027,n2024,n2025);
or (n2028,n2029,n2032);
and (n2029,n2030,n2031);
xor (n2030,n1946,n1947);
and (n2031,n368,n442);
and (n2032,n2033,n2034);
xor (n2033,n2030,n2031);
or (n2034,n2035,n2038);
and (n2035,n2036,n2037);
xor (n2036,n1951,n1952);
and (n2037,n387,n442);
and (n2038,n2039,n2040);
xor (n2039,n2036,n2037);
or (n2040,n2041,n2044);
and (n2041,n2042,n2043);
xor (n2042,n1956,n1957);
and (n2043,n381,n442);
and (n2044,n2045,n2046);
xor (n2045,n2042,n2043);
or (n2046,n2047,n2050);
and (n2047,n2048,n2049);
xor (n2048,n1961,n1962);
and (n2049,n534,n442);
and (n2050,n2051,n2052);
xor (n2051,n2048,n2049);
and (n2052,n2053,n1389);
xor (n2053,n1967,n1968);
and (n2054,n109,n121);
or (n2055,n2056,n2058);
and (n2056,n2057,n2054);
xor (n2057,n1676,n1694);
and (n2058,n2059,n2060);
xor (n2059,n2057,n2054);
or (n2060,n2061,n2063);
and (n2061,n2062,n2054);
xor (n2062,n1676,n1696);
and (n2063,n2064,n2065);
xor (n2064,n2062,n2054);
or (n2065,n2066,n2068);
and (n2066,n2067,n2054);
xor (n2067,n1676,n1698);
and (n2068,n2069,n2070);
xor (n2069,n2067,n2054);
or (n2070,n2071,n2073);
and (n2071,n2072,n2054);
xor (n2072,n1676,n1700);
and (n2073,n2074,n2075);
xor (n2074,n2072,n2054);
or (n2075,n2076,n2078);
and (n2076,n2077,n2054);
xor (n2077,n1676,n1702);
and (n2078,n2079,n2080);
xor (n2079,n2077,n2054);
or (n2080,n2081,n2083);
and (n2081,n2082,n2054);
xor (n2082,n1676,n1704);
and (n2083,n2084,n2085);
xor (n2084,n2082,n2054);
or (n2085,n2086,n2088);
and (n2086,n2087,n2054);
xor (n2087,n1676,n1706);
and (n2088,n2089,n2090);
xor (n2089,n2087,n2054);
or (n2090,n2091,n2093);
and (n2091,n2092,n2054);
xor (n2092,n1676,n1708);
and (n2093,n2094,n2095);
xor (n2094,n2092,n2054);
or (n2095,n2096,n2098);
and (n2096,n2097,n2054);
xor (n2097,n1676,n1710);
and (n2098,n2099,n2100);
xor (n2099,n2097,n2054);
or (n2100,n2101,n2103);
and (n2101,n2102,n2054);
xor (n2102,n1676,n1712);
and (n2103,n2104,n2105);
xor (n2104,n2102,n2054);
or (n2105,n2106,n2108);
and (n2106,n2107,n2054);
xor (n2107,n1676,n1714);
and (n2108,n2109,n2110);
xor (n2109,n2107,n2054);
or (n2110,n2111,n2114);
and (n2111,n2112,n2113);
xor (n2112,n1676,n1716);
and (n2113,n103,n121);
and (n2114,n2115,n2116);
xor (n2115,n2112,n2113);
or (n2116,n2117,n2120);
and (n2117,n2118,n2119);
xor (n2118,n1973,n1974);
and (n2119,n92,n121);
and (n2120,n2121,n2122);
xor (n2121,n2118,n2119);
or (n2122,n2123,n2126);
and (n2123,n2124,n2125);
xor (n2124,n1979,n1980);
and (n2125,n70,n121);
and (n2126,n2127,n2128);
xor (n2127,n2124,n2125);
or (n2128,n2129,n2132);
and (n2129,n2130,n2131);
xor (n2130,n1985,n1986);
and (n2131,n64,n121);
and (n2132,n2133,n2134);
xor (n2133,n2130,n2131);
or (n2134,n2135,n2138);
and (n2135,n2136,n2137);
xor (n2136,n1991,n1992);
and (n2137,n148,n121);
and (n2138,n2139,n2140);
xor (n2139,n2136,n2137);
or (n2140,n2141,n2144);
and (n2141,n2142,n2143);
xor (n2142,n1997,n1998);
and (n2143,n157,n121);
and (n2144,n2145,n2146);
xor (n2145,n2142,n2143);
or (n2146,n2147,n2150);
and (n2147,n2148,n2149);
xor (n2148,n2003,n2004);
and (n2149,n44,n121);
and (n2150,n2151,n2152);
xor (n2151,n2148,n2149);
or (n2152,n2153,n2156);
and (n2153,n2154,n2155);
xor (n2154,n2009,n2010);
and (n2155,n38,n121);
and (n2156,n2157,n2158);
xor (n2157,n2154,n2155);
or (n2158,n2159,n2162);
and (n2159,n2160,n2161);
xor (n2160,n2015,n2016);
and (n2161,n197,n121);
and (n2162,n2163,n2164);
xor (n2163,n2160,n2161);
or (n2164,n2165,n2168);
and (n2165,n2166,n2167);
xor (n2166,n2021,n2022);
and (n2167,n374,n121);
and (n2168,n2169,n2170);
xor (n2169,n2166,n2167);
or (n2170,n2171,n2174);
and (n2171,n2172,n2173);
xor (n2172,n2027,n2028);
and (n2173,n368,n121);
and (n2174,n2175,n2176);
xor (n2175,n2172,n2173);
or (n2176,n2177,n2180);
and (n2177,n2178,n2179);
xor (n2178,n2033,n2034);
and (n2179,n387,n121);
and (n2180,n2181,n2182);
xor (n2181,n2178,n2179);
or (n2182,n2183,n2186);
and (n2183,n2184,n2185);
xor (n2184,n2039,n2040);
and (n2185,n381,n121);
and (n2186,n2187,n2188);
xor (n2187,n2184,n2185);
or (n2188,n2189,n2192);
and (n2189,n2190,n2191);
xor (n2190,n2045,n2046);
and (n2191,n534,n121);
and (n2192,n2193,n2194);
xor (n2193,n2190,n2191);
and (n2194,n2195,n2196);
xor (n2195,n2051,n2052);
and (n2196,n594,n121);
and (n2197,n109,n122);
or (n2198,n2199,n2201);
and (n2199,n2200,n2197);
xor (n2200,n2059,n2060);
and (n2201,n2202,n2203);
xor (n2202,n2200,n2197);
or (n2203,n2204,n2206);
and (n2204,n2205,n2197);
xor (n2205,n2064,n2065);
and (n2206,n2207,n2208);
xor (n2207,n2205,n2197);
or (n2208,n2209,n2211);
and (n2209,n2210,n2197);
xor (n2210,n2069,n2070);
and (n2211,n2212,n2213);
xor (n2212,n2210,n2197);
or (n2213,n2214,n2216);
and (n2214,n2215,n2197);
xor (n2215,n2074,n2075);
and (n2216,n2217,n2218);
xor (n2217,n2215,n2197);
or (n2218,n2219,n2221);
and (n2219,n2220,n2197);
xor (n2220,n2079,n2080);
and (n2221,n2222,n2223);
xor (n2222,n2220,n2197);
or (n2223,n2224,n2226);
and (n2224,n2225,n2197);
xor (n2225,n2084,n2085);
and (n2226,n2227,n2228);
xor (n2227,n2225,n2197);
or (n2228,n2229,n2231);
and (n2229,n2230,n2197);
xor (n2230,n2089,n2090);
and (n2231,n2232,n2233);
xor (n2232,n2230,n2197);
or (n2233,n2234,n2236);
and (n2234,n2235,n2197);
xor (n2235,n2094,n2095);
and (n2236,n2237,n2238);
xor (n2237,n2235,n2197);
or (n2238,n2239,n2241);
and (n2239,n2240,n2197);
xor (n2240,n2099,n2100);
and (n2241,n2242,n2243);
xor (n2242,n2240,n2197);
or (n2243,n2244,n2246);
and (n2244,n2245,n2197);
xor (n2245,n2104,n2105);
and (n2246,n2247,n2248);
xor (n2247,n2245,n2197);
or (n2248,n2249,n2252);
and (n2249,n2250,n2251);
xor (n2250,n2109,n2110);
and (n2251,n103,n122);
and (n2252,n2253,n2254);
xor (n2253,n2250,n2251);
or (n2254,n2255,n2258);
and (n2255,n2256,n2257);
xor (n2256,n2115,n2116);
and (n2257,n92,n122);
and (n2258,n2259,n2260);
xor (n2259,n2256,n2257);
or (n2260,n2261,n2264);
and (n2261,n2262,n2263);
xor (n2262,n2121,n2122);
and (n2263,n70,n122);
and (n2264,n2265,n2266);
xor (n2265,n2262,n2263);
or (n2266,n2267,n2270);
and (n2267,n2268,n2269);
xor (n2268,n2127,n2128);
and (n2269,n64,n122);
and (n2270,n2271,n2272);
xor (n2271,n2268,n2269);
or (n2272,n2273,n2276);
and (n2273,n2274,n2275);
xor (n2274,n2133,n2134);
and (n2275,n148,n122);
and (n2276,n2277,n2278);
xor (n2277,n2274,n2275);
or (n2278,n2279,n2282);
and (n2279,n2280,n2281);
xor (n2280,n2139,n2140);
and (n2281,n157,n122);
and (n2282,n2283,n2284);
xor (n2283,n2280,n2281);
or (n2284,n2285,n2288);
and (n2285,n2286,n2287);
xor (n2286,n2145,n2146);
and (n2287,n44,n122);
and (n2288,n2289,n2290);
xor (n2289,n2286,n2287);
or (n2290,n2291,n2294);
and (n2291,n2292,n2293);
xor (n2292,n2151,n2152);
and (n2293,n38,n122);
and (n2294,n2295,n2296);
xor (n2295,n2292,n2293);
or (n2296,n2297,n2300);
and (n2297,n2298,n2299);
xor (n2298,n2157,n2158);
and (n2299,n197,n122);
and (n2300,n2301,n2302);
xor (n2301,n2298,n2299);
or (n2302,n2303,n2306);
and (n2303,n2304,n2305);
xor (n2304,n2163,n2164);
and (n2305,n374,n122);
and (n2306,n2307,n2308);
xor (n2307,n2304,n2305);
or (n2308,n2309,n2312);
and (n2309,n2310,n2311);
xor (n2310,n2169,n2170);
and (n2311,n368,n122);
and (n2312,n2313,n2314);
xor (n2313,n2310,n2311);
or (n2314,n2315,n2318);
and (n2315,n2316,n2317);
xor (n2316,n2175,n2176);
and (n2317,n387,n122);
and (n2318,n2319,n2320);
xor (n2319,n2316,n2317);
or (n2320,n2321,n2324);
and (n2321,n2322,n2323);
xor (n2322,n2181,n2182);
and (n2323,n381,n122);
and (n2324,n2325,n2326);
xor (n2325,n2322,n2323);
or (n2326,n2327,n2330);
and (n2327,n2328,n2329);
xor (n2328,n2187,n2188);
and (n2329,n534,n122);
and (n2330,n2331,n2332);
xor (n2331,n2328,n2329);
and (n2332,n2333,n1233);
xor (n2333,n2193,n2194);
and (n2334,n109,n79);
or (n2335,n2336,n2338);
and (n2336,n2337,n2334);
xor (n2337,n2202,n2203);
and (n2338,n2339,n2340);
xor (n2339,n2337,n2334);
or (n2340,n2341,n2343);
and (n2341,n2342,n2334);
xor (n2342,n2207,n2208);
and (n2343,n2344,n2345);
xor (n2344,n2342,n2334);
or (n2345,n2346,n2348);
and (n2346,n2347,n2334);
xor (n2347,n2212,n2213);
and (n2348,n2349,n2350);
xor (n2349,n2347,n2334);
or (n2350,n2351,n2353);
and (n2351,n2352,n2334);
xor (n2352,n2217,n2218);
and (n2353,n2354,n2355);
xor (n2354,n2352,n2334);
or (n2355,n2356,n2358);
and (n2356,n2357,n2334);
xor (n2357,n2222,n2223);
and (n2358,n2359,n2360);
xor (n2359,n2357,n2334);
or (n2360,n2361,n2363);
and (n2361,n2362,n2334);
xor (n2362,n2227,n2228);
and (n2363,n2364,n2365);
xor (n2364,n2362,n2334);
or (n2365,n2366,n2368);
and (n2366,n2367,n2334);
xor (n2367,n2232,n2233);
and (n2368,n2369,n2370);
xor (n2369,n2367,n2334);
or (n2370,n2371,n2373);
and (n2371,n2372,n2334);
xor (n2372,n2237,n2238);
and (n2373,n2374,n2375);
xor (n2374,n2372,n2334);
or (n2375,n2376,n2378);
and (n2376,n2377,n2334);
xor (n2377,n2242,n2243);
and (n2378,n2379,n2380);
xor (n2379,n2377,n2334);
or (n2380,n2381,n2384);
and (n2381,n2382,n2383);
xor (n2382,n2247,n2248);
and (n2383,n103,n79);
and (n2384,n2385,n2386);
xor (n2385,n2382,n2383);
or (n2386,n2387,n2390);
and (n2387,n2388,n2389);
xor (n2388,n2253,n2254);
and (n2389,n92,n79);
and (n2390,n2391,n2392);
xor (n2391,n2388,n2389);
or (n2392,n2393,n2396);
and (n2393,n2394,n2395);
xor (n2394,n2259,n2260);
and (n2395,n70,n79);
and (n2396,n2397,n2398);
xor (n2397,n2394,n2395);
or (n2398,n2399,n2402);
and (n2399,n2400,n2401);
xor (n2400,n2265,n2266);
and (n2401,n64,n79);
and (n2402,n2403,n2404);
xor (n2403,n2400,n2401);
or (n2404,n2405,n2408);
and (n2405,n2406,n2407);
xor (n2406,n2271,n2272);
and (n2407,n148,n79);
and (n2408,n2409,n2410);
xor (n2409,n2406,n2407);
or (n2410,n2411,n2414);
and (n2411,n2412,n2413);
xor (n2412,n2277,n2278);
and (n2413,n157,n79);
and (n2414,n2415,n2416);
xor (n2415,n2412,n2413);
or (n2416,n2417,n2420);
and (n2417,n2418,n2419);
xor (n2418,n2283,n2284);
and (n2419,n44,n79);
and (n2420,n2421,n2422);
xor (n2421,n2418,n2419);
or (n2422,n2423,n2426);
and (n2423,n2424,n2425);
xor (n2424,n2289,n2290);
and (n2425,n38,n79);
and (n2426,n2427,n2428);
xor (n2427,n2424,n2425);
or (n2428,n2429,n2432);
and (n2429,n2430,n2431);
xor (n2430,n2295,n2296);
and (n2431,n197,n79);
and (n2432,n2433,n2434);
xor (n2433,n2430,n2431);
or (n2434,n2435,n2438);
and (n2435,n2436,n2437);
xor (n2436,n2301,n2302);
and (n2437,n374,n79);
and (n2438,n2439,n2440);
xor (n2439,n2436,n2437);
or (n2440,n2441,n2444);
and (n2441,n2442,n2443);
xor (n2442,n2307,n2308);
and (n2443,n368,n79);
and (n2444,n2445,n2446);
xor (n2445,n2442,n2443);
or (n2446,n2447,n2450);
and (n2447,n2448,n2449);
xor (n2448,n2313,n2314);
and (n2449,n387,n79);
and (n2450,n2451,n2452);
xor (n2451,n2448,n2449);
or (n2452,n2453,n2456);
and (n2453,n2454,n2455);
xor (n2454,n2319,n2320);
and (n2455,n381,n79);
and (n2456,n2457,n2458);
xor (n2457,n2454,n2455);
or (n2458,n2459,n2461);
and (n2459,n2460,n1281);
xor (n2460,n2325,n2326);
and (n2461,n2462,n2463);
xor (n2462,n2460,n1281);
and (n2463,n2464,n2465);
xor (n2464,n2331,n2332);
and (n2465,n594,n79);
and (n2466,n109,n80);
or (n2467,n2468,n2470);
and (n2468,n2469,n2466);
xor (n2469,n2339,n2340);
and (n2470,n2471,n2472);
xor (n2471,n2469,n2466);
or (n2472,n2473,n2475);
and (n2473,n2474,n2466);
xor (n2474,n2344,n2345);
and (n2475,n2476,n2477);
xor (n2476,n2474,n2466);
or (n2477,n2478,n2480);
and (n2478,n2479,n2466);
xor (n2479,n2349,n2350);
and (n2480,n2481,n2482);
xor (n2481,n2479,n2466);
or (n2482,n2483,n2485);
and (n2483,n2484,n2466);
xor (n2484,n2354,n2355);
and (n2485,n2486,n2487);
xor (n2486,n2484,n2466);
or (n2487,n2488,n2490);
and (n2488,n2489,n2466);
xor (n2489,n2359,n2360);
and (n2490,n2491,n2492);
xor (n2491,n2489,n2466);
or (n2492,n2493,n2495);
and (n2493,n2494,n2466);
xor (n2494,n2364,n2365);
and (n2495,n2496,n2497);
xor (n2496,n2494,n2466);
or (n2497,n2498,n2500);
and (n2498,n2499,n2466);
xor (n2499,n2369,n2370);
and (n2500,n2501,n2502);
xor (n2501,n2499,n2466);
or (n2502,n2503,n2505);
and (n2503,n2504,n2466);
xor (n2504,n2374,n2375);
and (n2505,n2506,n2507);
xor (n2506,n2504,n2466);
or (n2507,n2508,n2511);
and (n2508,n2509,n2510);
xor (n2509,n2379,n2380);
and (n2510,n103,n80);
and (n2511,n2512,n2513);
xor (n2512,n2509,n2510);
or (n2513,n2514,n2517);
and (n2514,n2515,n2516);
xor (n2515,n2385,n2386);
and (n2516,n92,n80);
and (n2517,n2518,n2519);
xor (n2518,n2515,n2516);
or (n2519,n2520,n2523);
and (n2520,n2521,n2522);
xor (n2521,n2391,n2392);
and (n2522,n70,n80);
and (n2523,n2524,n2525);
xor (n2524,n2521,n2522);
or (n2525,n2526,n2529);
and (n2526,n2527,n2528);
xor (n2527,n2397,n2398);
and (n2528,n64,n80);
and (n2529,n2530,n2531);
xor (n2530,n2527,n2528);
or (n2531,n2532,n2535);
and (n2532,n2533,n2534);
xor (n2533,n2403,n2404);
and (n2534,n148,n80);
and (n2535,n2536,n2537);
xor (n2536,n2533,n2534);
or (n2537,n2538,n2541);
and (n2538,n2539,n2540);
xor (n2539,n2409,n2410);
and (n2540,n157,n80);
and (n2541,n2542,n2543);
xor (n2542,n2539,n2540);
or (n2543,n2544,n2547);
and (n2544,n2545,n2546);
xor (n2545,n2415,n2416);
and (n2546,n44,n80);
and (n2547,n2548,n2549);
xor (n2548,n2545,n2546);
or (n2549,n2550,n2553);
and (n2550,n2551,n2552);
xor (n2551,n2421,n2422);
and (n2552,n38,n80);
and (n2553,n2554,n2555);
xor (n2554,n2551,n2552);
or (n2555,n2556,n2559);
and (n2556,n2557,n2558);
xor (n2557,n2427,n2428);
and (n2558,n197,n80);
and (n2559,n2560,n2561);
xor (n2560,n2557,n2558);
or (n2561,n2562,n2565);
and (n2562,n2563,n2564);
xor (n2563,n2433,n2434);
and (n2564,n374,n80);
and (n2565,n2566,n2567);
xor (n2566,n2563,n2564);
or (n2567,n2568,n2571);
and (n2568,n2569,n2570);
xor (n2569,n2439,n2440);
and (n2570,n368,n80);
and (n2571,n2572,n2573);
xor (n2572,n2569,n2570);
or (n2573,n2574,n2577);
and (n2574,n2575,n2576);
xor (n2575,n2445,n2446);
and (n2576,n387,n80);
and (n2577,n2578,n2579);
xor (n2578,n2575,n2576);
or (n2579,n2580,n2583);
and (n2580,n2581,n2582);
xor (n2581,n2451,n2452);
and (n2582,n381,n80);
and (n2583,n2584,n2585);
xor (n2584,n2581,n2582);
or (n2585,n2586,n2589);
and (n2586,n2587,n2588);
xor (n2587,n2457,n2458);
and (n2588,n534,n80);
and (n2589,n2590,n2591);
xor (n2590,n2587,n2588);
and (n2591,n2592,n2593);
xor (n2592,n2462,n2463);
not (n2593,n1258);
and (n2594,n109,n53);
or (n2595,n2596,n2598);
and (n2596,n2597,n2594);
xor (n2597,n2471,n2472);
and (n2598,n2599,n2600);
xor (n2599,n2597,n2594);
or (n2600,n2601,n2603);
and (n2601,n2602,n2594);
xor (n2602,n2476,n2477);
and (n2603,n2604,n2605);
xor (n2604,n2602,n2594);
or (n2605,n2606,n2608);
and (n2606,n2607,n2594);
xor (n2607,n2481,n2482);
and (n2608,n2609,n2610);
xor (n2609,n2607,n2594);
or (n2610,n2611,n2613);
and (n2611,n2612,n2594);
xor (n2612,n2486,n2487);
and (n2613,n2614,n2615);
xor (n2614,n2612,n2594);
or (n2615,n2616,n2618);
and (n2616,n2617,n2594);
xor (n2617,n2491,n2492);
and (n2618,n2619,n2620);
xor (n2619,n2617,n2594);
or (n2620,n2621,n2623);
and (n2621,n2622,n2594);
xor (n2622,n2496,n2497);
and (n2623,n2624,n2625);
xor (n2624,n2622,n2594);
or (n2625,n2626,n2628);
and (n2626,n2627,n2594);
xor (n2627,n2501,n2502);
and (n2628,n2629,n2630);
xor (n2629,n2627,n2594);
or (n2630,n2631,n2634);
and (n2631,n2632,n2633);
xor (n2632,n2506,n2507);
and (n2633,n103,n53);
and (n2634,n2635,n2636);
xor (n2635,n2632,n2633);
or (n2636,n2637,n2640);
and (n2637,n2638,n2639);
xor (n2638,n2512,n2513);
and (n2639,n92,n53);
and (n2640,n2641,n2642);
xor (n2641,n2638,n2639);
or (n2642,n2643,n2646);
and (n2643,n2644,n2645);
xor (n2644,n2518,n2519);
and (n2645,n70,n53);
and (n2646,n2647,n2648);
xor (n2647,n2644,n2645);
or (n2648,n2649,n2652);
and (n2649,n2650,n2651);
xor (n2650,n2524,n2525);
and (n2651,n64,n53);
and (n2652,n2653,n2654);
xor (n2653,n2650,n2651);
or (n2654,n2655,n2658);
and (n2655,n2656,n2657);
xor (n2656,n2530,n2531);
and (n2657,n148,n53);
and (n2658,n2659,n2660);
xor (n2659,n2656,n2657);
or (n2660,n2661,n2664);
and (n2661,n2662,n2663);
xor (n2662,n2536,n2537);
and (n2663,n157,n53);
and (n2664,n2665,n2666);
xor (n2665,n2662,n2663);
or (n2666,n2667,n2670);
and (n2667,n2668,n2669);
xor (n2668,n2542,n2543);
and (n2669,n44,n53);
and (n2670,n2671,n2672);
xor (n2671,n2668,n2669);
or (n2672,n2673,n2675);
and (n2673,n2674,n549);
xor (n2674,n2548,n2549);
and (n2675,n2676,n2677);
xor (n2676,n2674,n549);
or (n2677,n2678,n2681);
and (n2678,n2679,n2680);
xor (n2679,n2554,n2555);
and (n2680,n197,n53);
and (n2681,n2682,n2683);
xor (n2682,n2679,n2680);
or (n2683,n2684,n2687);
and (n2684,n2685,n2686);
xor (n2685,n2560,n2561);
and (n2686,n374,n53);
and (n2687,n2688,n2689);
xor (n2688,n2685,n2686);
or (n2689,n2690,n2692);
and (n2690,n2691,n793);
xor (n2691,n2566,n2567);
and (n2692,n2693,n2694);
xor (n2693,n2691,n793);
or (n2694,n2695,n2698);
and (n2695,n2696,n2697);
xor (n2696,n2572,n2573);
and (n2697,n387,n53);
and (n2698,n2699,n2700);
xor (n2699,n2696,n2697);
or (n2700,n2701,n2703);
and (n2701,n2702,n1117);
xor (n2702,n2578,n2579);
and (n2703,n2704,n2705);
xor (n2704,n2702,n1117);
or (n2705,n2706,n2709);
and (n2706,n2707,n2708);
xor (n2707,n2584,n2585);
and (n2708,n534,n53);
and (n2709,n2710,n2711);
xor (n2710,n2707,n2708);
and (n2711,n2712,n2713);
xor (n2712,n2590,n2591);
and (n2713,n594,n53);
and (n2714,n109,n54);
or (n2715,n2716,n2718);
and (n2716,n2717,n2714);
xor (n2717,n2599,n2600);
and (n2718,n2719,n2720);
xor (n2719,n2717,n2714);
or (n2720,n2721,n2723);
and (n2721,n2722,n2714);
xor (n2722,n2604,n2605);
and (n2723,n2724,n2725);
xor (n2724,n2722,n2714);
or (n2725,n2726,n2728);
and (n2726,n2727,n2714);
xor (n2727,n2609,n2610);
and (n2728,n2729,n2730);
xor (n2729,n2727,n2714);
or (n2730,n2731,n2733);
and (n2731,n2732,n2714);
xor (n2732,n2614,n2615);
and (n2733,n2734,n2735);
xor (n2734,n2732,n2714);
or (n2735,n2736,n2738);
and (n2736,n2737,n2714);
xor (n2737,n2619,n2620);
and (n2738,n2739,n2740);
xor (n2739,n2737,n2714);
or (n2740,n2741,n2743);
and (n2741,n2742,n2714);
xor (n2742,n2624,n2625);
and (n2743,n2744,n2745);
xor (n2744,n2742,n2714);
or (n2745,n2746,n2749);
and (n2746,n2747,n2748);
xor (n2747,n2629,n2630);
and (n2748,n103,n54);
and (n2749,n2750,n2751);
xor (n2750,n2747,n2748);
or (n2751,n2752,n2755);
and (n2752,n2753,n2754);
xor (n2753,n2635,n2636);
and (n2754,n92,n54);
and (n2755,n2756,n2757);
xor (n2756,n2753,n2754);
or (n2757,n2758,n2761);
and (n2758,n2759,n2760);
xor (n2759,n2641,n2642);
and (n2760,n70,n54);
and (n2761,n2762,n2763);
xor (n2762,n2759,n2760);
or (n2763,n2764,n2767);
and (n2764,n2765,n2766);
xor (n2765,n2647,n2648);
and (n2766,n64,n54);
and (n2767,n2768,n2769);
xor (n2768,n2765,n2766);
or (n2769,n2770,n2773);
and (n2770,n2771,n2772);
xor (n2771,n2653,n2654);
and (n2772,n148,n54);
and (n2773,n2774,n2775);
xor (n2774,n2771,n2772);
or (n2775,n2776,n2779);
and (n2776,n2777,n2778);
xor (n2777,n2659,n2660);
and (n2778,n157,n54);
and (n2779,n2780,n2781);
xor (n2780,n2777,n2778);
or (n2781,n2782,n2785);
and (n2782,n2783,n2784);
xor (n2783,n2665,n2666);
and (n2784,n44,n54);
and (n2785,n2786,n2787);
xor (n2786,n2783,n2784);
or (n2787,n2788,n2791);
and (n2788,n2789,n2790);
xor (n2789,n2671,n2672);
and (n2790,n38,n54);
and (n2791,n2792,n2793);
xor (n2792,n2789,n2790);
or (n2793,n2794,n2797);
and (n2794,n2795,n2796);
xor (n2795,n2676,n2677);
and (n2796,n197,n54);
and (n2797,n2798,n2799);
xor (n2798,n2795,n2796);
or (n2799,n2800,n2803);
and (n2800,n2801,n2802);
xor (n2801,n2682,n2683);
and (n2802,n374,n54);
and (n2803,n2804,n2805);
xor (n2804,n2801,n2802);
or (n2805,n2806,n2809);
and (n2806,n2807,n2808);
xor (n2807,n2688,n2689);
and (n2808,n368,n54);
and (n2809,n2810,n2811);
xor (n2810,n2807,n2808);
or (n2811,n2812,n2815);
and (n2812,n2813,n2814);
xor (n2813,n2693,n2694);
and (n2814,n387,n54);
and (n2815,n2816,n2817);
xor (n2816,n2813,n2814);
or (n2817,n2818,n2821);
and (n2818,n2819,n2820);
xor (n2819,n2699,n2700);
and (n2820,n381,n54);
and (n2821,n2822,n2823);
xor (n2822,n2819,n2820);
or (n2823,n2824,n2827);
and (n2824,n2825,n2826);
xor (n2825,n2704,n2705);
and (n2826,n534,n54);
and (n2827,n2828,n2829);
xor (n2828,n2825,n2826);
and (n2829,n2830,n1101);
xor (n2830,n2710,n2711);
and (n2831,n109,n60);
or (n2832,n2833,n2835);
and (n2833,n2834,n2831);
xor (n2834,n2719,n2720);
and (n2835,n2836,n2837);
xor (n2836,n2834,n2831);
or (n2837,n2838,n2840);
and (n2838,n2839,n2831);
xor (n2839,n2724,n2725);
and (n2840,n2841,n2842);
xor (n2841,n2839,n2831);
or (n2842,n2843,n2845);
and (n2843,n2844,n2831);
xor (n2844,n2729,n2730);
and (n2845,n2846,n2847);
xor (n2846,n2844,n2831);
or (n2847,n2848,n2850);
and (n2848,n2849,n2831);
xor (n2849,n2734,n2735);
and (n2850,n2851,n2852);
xor (n2851,n2849,n2831);
or (n2852,n2853,n2855);
and (n2853,n2854,n2831);
xor (n2854,n2739,n2740);
and (n2855,n2856,n2857);
xor (n2856,n2854,n2831);
or (n2857,n2858,n2861);
and (n2858,n2859,n2860);
xor (n2859,n2744,n2745);
and (n2860,n103,n60);
and (n2861,n2862,n2863);
xor (n2862,n2859,n2860);
or (n2863,n2864,n2867);
and (n2864,n2865,n2866);
xor (n2865,n2750,n2751);
and (n2866,n92,n60);
and (n2867,n2868,n2869);
xor (n2868,n2865,n2866);
or (n2869,n2870,n2873);
and (n2870,n2871,n2872);
xor (n2871,n2756,n2757);
and (n2872,n70,n60);
and (n2873,n2874,n2875);
xor (n2874,n2871,n2872);
or (n2875,n2876,n2879);
and (n2876,n2877,n2878);
xor (n2877,n2762,n2763);
and (n2878,n64,n60);
and (n2879,n2880,n2881);
xor (n2880,n2877,n2878);
or (n2881,n2882,n2885);
and (n2882,n2883,n2884);
xor (n2883,n2768,n2769);
and (n2884,n148,n60);
and (n2885,n2886,n2887);
xor (n2886,n2883,n2884);
or (n2887,n2888,n2891);
and (n2888,n2889,n2890);
xor (n2889,n2774,n2775);
and (n2890,n157,n60);
and (n2891,n2892,n2893);
xor (n2892,n2889,n2890);
or (n2893,n2894,n2897);
and (n2894,n2895,n2896);
xor (n2895,n2780,n2781);
and (n2896,n44,n60);
and (n2897,n2898,n2899);
xor (n2898,n2895,n2896);
or (n2899,n2900,n2903);
and (n2900,n2901,n2902);
xor (n2901,n2786,n2787);
and (n2902,n38,n60);
and (n2903,n2904,n2905);
xor (n2904,n2901,n2902);
or (n2905,n2906,n2909);
and (n2906,n2907,n2908);
xor (n2907,n2792,n2793);
and (n2908,n197,n60);
and (n2909,n2910,n2911);
xor (n2910,n2907,n2908);
or (n2911,n2912,n2915);
and (n2912,n2913,n2914);
xor (n2913,n2798,n2799);
and (n2914,n374,n60);
and (n2915,n2916,n2917);
xor (n2916,n2913,n2914);
or (n2917,n2918,n2921);
and (n2918,n2919,n2920);
xor (n2919,n2804,n2805);
and (n2920,n368,n60);
and (n2921,n2922,n2923);
xor (n2922,n2919,n2920);
or (n2923,n2924,n2927);
and (n2924,n2925,n2926);
xor (n2925,n2810,n2811);
and (n2926,n387,n60);
and (n2927,n2928,n2929);
xor (n2928,n2925,n2926);
or (n2929,n2930,n2933);
and (n2930,n2931,n2932);
xor (n2931,n2816,n2817);
and (n2932,n381,n60);
and (n2933,n2934,n2935);
xor (n2934,n2931,n2932);
or (n2935,n2936,n2939);
and (n2936,n2937,n2938);
xor (n2937,n2822,n2823);
and (n2938,n534,n60);
and (n2939,n2940,n2941);
xor (n2940,n2937,n2938);
and (n2941,n2942,n2943);
xor (n2942,n2828,n2829);
and (n2943,n594,n60);
and (n2944,n109,n142);
or (n2945,n2946,n2948);
and (n2946,n2947,n2944);
xor (n2947,n2836,n2837);
and (n2948,n2949,n2950);
xor (n2949,n2947,n2944);
or (n2950,n2951,n2953);
and (n2951,n2952,n2944);
xor (n2952,n2841,n2842);
and (n2953,n2954,n2955);
xor (n2954,n2952,n2944);
or (n2955,n2956,n2958);
and (n2956,n2957,n2944);
xor (n2957,n2846,n2847);
and (n2958,n2959,n2960);
xor (n2959,n2957,n2944);
or (n2960,n2961,n2963);
and (n2961,n2962,n2944);
xor (n2962,n2851,n2852);
and (n2963,n2964,n2965);
xor (n2964,n2962,n2944);
or (n2965,n2966,n2969);
and (n2966,n2967,n2968);
xor (n2967,n2856,n2857);
and (n2968,n103,n142);
and (n2969,n2970,n2971);
xor (n2970,n2967,n2968);
or (n2971,n2972,n2975);
and (n2972,n2973,n2974);
xor (n2973,n2862,n2863);
and (n2974,n92,n142);
and (n2975,n2976,n2977);
xor (n2976,n2973,n2974);
or (n2977,n2978,n2981);
and (n2978,n2979,n2980);
xor (n2979,n2868,n2869);
and (n2980,n70,n142);
and (n2981,n2982,n2983);
xor (n2982,n2979,n2980);
or (n2983,n2984,n2987);
and (n2984,n2985,n2986);
xor (n2985,n2874,n2875);
and (n2986,n64,n142);
and (n2987,n2988,n2989);
xor (n2988,n2985,n2986);
or (n2989,n2990,n2993);
and (n2990,n2991,n2992);
xor (n2991,n2880,n2881);
and (n2992,n148,n142);
and (n2993,n2994,n2995);
xor (n2994,n2991,n2992);
or (n2995,n2996,n2999);
and (n2996,n2997,n2998);
xor (n2997,n2886,n2887);
and (n2998,n157,n142);
and (n2999,n3000,n3001);
xor (n3000,n2997,n2998);
or (n3001,n3002,n3005);
and (n3002,n3003,n3004);
xor (n3003,n2892,n2893);
and (n3004,n44,n142);
and (n3005,n3006,n3007);
xor (n3006,n3003,n3004);
or (n3007,n3008,n3011);
and (n3008,n3009,n3010);
xor (n3009,n2898,n2899);
and (n3010,n38,n142);
and (n3011,n3012,n3013);
xor (n3012,n3009,n3010);
or (n3013,n3014,n3017);
and (n3014,n3015,n3016);
xor (n3015,n2904,n2905);
and (n3016,n197,n142);
and (n3017,n3018,n3019);
xor (n3018,n3015,n3016);
or (n3019,n3020,n3023);
and (n3020,n3021,n3022);
xor (n3021,n2910,n2911);
and (n3022,n374,n142);
and (n3023,n3024,n3025);
xor (n3024,n3021,n3022);
or (n3025,n3026,n3029);
and (n3026,n3027,n3028);
xor (n3027,n2916,n2917);
and (n3028,n368,n142);
and (n3029,n3030,n3031);
xor (n3030,n3027,n3028);
or (n3031,n3032,n3035);
and (n3032,n3033,n3034);
xor (n3033,n2922,n2923);
and (n3034,n387,n142);
and (n3035,n3036,n3037);
xor (n3036,n3033,n3034);
or (n3037,n3038,n3041);
and (n3038,n3039,n3040);
xor (n3039,n2928,n2929);
and (n3040,n381,n142);
and (n3041,n3042,n3043);
xor (n3042,n3039,n3040);
or (n3043,n3044,n3047);
and (n3044,n3045,n3046);
xor (n3045,n2934,n2935);
and (n3046,n534,n142);
and (n3047,n3048,n3049);
xor (n3048,n3045,n3046);
and (n3049,n3050,n3051);
xor (n3050,n2940,n2941);
not (n3051,n759);
and (n3052,n109,n27);
or (n3053,n3054,n3056);
and (n3054,n3055,n3052);
xor (n3055,n2949,n2950);
and (n3056,n3057,n3058);
xor (n3057,n3055,n3052);
or (n3058,n3059,n3061);
and (n3059,n3060,n3052);
xor (n3060,n2954,n2955);
and (n3061,n3062,n3063);
xor (n3062,n3060,n3052);
or (n3063,n3064,n3066);
and (n3064,n3065,n3052);
xor (n3065,n2959,n2960);
and (n3066,n3067,n3068);
xor (n3067,n3065,n3052);
or (n3068,n3069,n3072);
and (n3069,n3070,n3071);
xor (n3070,n2964,n2965);
and (n3071,n103,n27);
and (n3072,n3073,n3074);
xor (n3073,n3070,n3071);
or (n3074,n3075,n3078);
and (n3075,n3076,n3077);
xor (n3076,n2970,n2971);
and (n3077,n92,n27);
and (n3078,n3079,n3080);
xor (n3079,n3076,n3077);
or (n3080,n3081,n3084);
and (n3081,n3082,n3083);
xor (n3082,n2976,n2977);
and (n3083,n70,n27);
and (n3084,n3085,n3086);
xor (n3085,n3082,n3083);
or (n3086,n3087,n3090);
and (n3087,n3088,n3089);
xor (n3088,n2982,n2983);
and (n3089,n64,n27);
and (n3090,n3091,n3092);
xor (n3091,n3088,n3089);
or (n3092,n3093,n3096);
and (n3093,n3094,n3095);
xor (n3094,n2988,n2989);
and (n3095,n148,n27);
and (n3096,n3097,n3098);
xor (n3097,n3094,n3095);
or (n3098,n3099,n3102);
and (n3099,n3100,n3101);
xor (n3100,n2994,n2995);
and (n3101,n157,n27);
and (n3102,n3103,n3104);
xor (n3103,n3100,n3101);
or (n3104,n3105,n3108);
and (n3105,n3106,n3107);
xor (n3106,n3000,n3001);
and (n3107,n44,n27);
and (n3108,n3109,n3110);
xor (n3109,n3106,n3107);
or (n3110,n3111,n3114);
and (n3111,n3112,n3113);
xor (n3112,n3006,n3007);
and (n3113,n38,n27);
and (n3114,n3115,n3116);
xor (n3115,n3112,n3113);
or (n3116,n3117,n3120);
and (n3117,n3118,n3119);
xor (n3118,n3012,n3013);
and (n3119,n197,n27);
and (n3120,n3121,n3122);
xor (n3121,n3118,n3119);
or (n3122,n3123,n3126);
and (n3123,n3124,n3125);
xor (n3124,n3018,n3019);
and (n3125,n374,n27);
and (n3126,n3127,n3128);
xor (n3127,n3124,n3125);
or (n3128,n3129,n3132);
and (n3129,n3130,n3131);
xor (n3130,n3024,n3025);
and (n3131,n368,n27);
and (n3132,n3133,n3134);
xor (n3133,n3130,n3131);
or (n3134,n3135,n3138);
and (n3135,n3136,n3137);
xor (n3136,n3030,n3031);
and (n3137,n387,n27);
and (n3138,n3139,n3140);
xor (n3139,n3136,n3137);
or (n3140,n3141,n3144);
and (n3141,n3142,n3143);
xor (n3142,n3036,n3037);
and (n3143,n381,n27);
and (n3144,n3145,n3146);
xor (n3145,n3142,n3143);
or (n3146,n3147,n3150);
and (n3147,n3148,n3149);
xor (n3148,n3042,n3043);
and (n3149,n534,n27);
and (n3150,n3151,n3152);
xor (n3151,n3148,n3149);
and (n3152,n3153,n3154);
xor (n3153,n3048,n3049);
and (n3154,n594,n27);
and (n3155,n109,n28);
or (n3156,n3157,n3159);
and (n3157,n3158,n3155);
xor (n3158,n3057,n3058);
and (n3159,n3160,n3161);
xor (n3160,n3158,n3155);
or (n3161,n3162,n3164);
and (n3162,n3163,n3155);
xor (n3163,n3062,n3063);
and (n3164,n3165,n3166);
xor (n3165,n3163,n3155);
or (n3166,n3167,n3170);
and (n3167,n3168,n3169);
xor (n3168,n3067,n3068);
and (n3169,n103,n28);
and (n3170,n3171,n3172);
xor (n3171,n3168,n3169);
or (n3172,n3173,n3176);
and (n3173,n3174,n3175);
xor (n3174,n3073,n3074);
and (n3175,n92,n28);
and (n3176,n3177,n3178);
xor (n3177,n3174,n3175);
or (n3178,n3179,n3182);
and (n3179,n3180,n3181);
xor (n3180,n3079,n3080);
and (n3181,n70,n28);
and (n3182,n3183,n3184);
xor (n3183,n3180,n3181);
or (n3184,n3185,n3188);
and (n3185,n3186,n3187);
xor (n3186,n3085,n3086);
and (n3187,n64,n28);
and (n3188,n3189,n3190);
xor (n3189,n3186,n3187);
or (n3190,n3191,n3194);
and (n3191,n3192,n3193);
xor (n3192,n3091,n3092);
and (n3193,n148,n28);
and (n3194,n3195,n3196);
xor (n3195,n3192,n3193);
or (n3196,n3197,n3200);
and (n3197,n3198,n3199);
xor (n3198,n3097,n3098);
and (n3199,n157,n28);
and (n3200,n3201,n3202);
xor (n3201,n3198,n3199);
or (n3202,n3203,n3206);
and (n3203,n3204,n3205);
xor (n3204,n3103,n3104);
and (n3205,n44,n28);
and (n3206,n3207,n3208);
xor (n3207,n3204,n3205);
or (n3208,n3209,n3212);
and (n3209,n3210,n3211);
xor (n3210,n3109,n3110);
and (n3211,n38,n28);
and (n3212,n3213,n3214);
xor (n3213,n3210,n3211);
or (n3214,n3215,n3218);
and (n3215,n3216,n3217);
xor (n3216,n3115,n3116);
and (n3217,n197,n28);
and (n3218,n3219,n3220);
xor (n3219,n3216,n3217);
or (n3220,n3221,n3224);
and (n3221,n3222,n3223);
xor (n3222,n3121,n3122);
and (n3223,n374,n28);
and (n3224,n3225,n3226);
xor (n3225,n3222,n3223);
or (n3226,n3227,n3230);
and (n3227,n3228,n3229);
xor (n3228,n3127,n3128);
and (n3229,n368,n28);
and (n3230,n3231,n3232);
xor (n3231,n3228,n3229);
or (n3232,n3233,n3236);
and (n3233,n3234,n3235);
xor (n3234,n3133,n3134);
and (n3235,n387,n28);
and (n3236,n3237,n3238);
xor (n3237,n3234,n3235);
or (n3238,n3239,n3242);
and (n3239,n3240,n3241);
xor (n3240,n3139,n3140);
and (n3241,n381,n28);
and (n3242,n3243,n3244);
xor (n3243,n3240,n3241);
or (n3244,n3245,n3248);
and (n3245,n3246,n3247);
xor (n3246,n3145,n3146);
and (n3247,n534,n28);
and (n3248,n3249,n3250);
xor (n3249,n3246,n3247);
and (n3250,n3251,n3252);
xor (n3251,n3151,n3152);
not (n3252,n593);
and (n3253,n109,n34);
or (n3254,n3255,n3257);
and (n3255,n3256,n3253);
xor (n3256,n3160,n3161);
and (n3257,n3258,n3259);
xor (n3258,n3256,n3253);
or (n3259,n3260,n3263);
and (n3260,n3261,n3262);
xor (n3261,n3165,n3166);
and (n3262,n103,n34);
and (n3263,n3264,n3265);
xor (n3264,n3261,n3262);
or (n3265,n3266,n3269);
and (n3266,n3267,n3268);
xor (n3267,n3171,n3172);
and (n3268,n92,n34);
and (n3269,n3270,n3271);
xor (n3270,n3267,n3268);
or (n3271,n3272,n3275);
and (n3272,n3273,n3274);
xor (n3273,n3177,n3178);
and (n3274,n70,n34);
and (n3275,n3276,n3277);
xor (n3276,n3273,n3274);
or (n3277,n3278,n3281);
and (n3278,n3279,n3280);
xor (n3279,n3183,n3184);
and (n3280,n64,n34);
and (n3281,n3282,n3283);
xor (n3282,n3279,n3280);
or (n3283,n3284,n3287);
and (n3284,n3285,n3286);
xor (n3285,n3189,n3190);
and (n3286,n148,n34);
and (n3287,n3288,n3289);
xor (n3288,n3285,n3286);
or (n3289,n3290,n3293);
and (n3290,n3291,n3292);
xor (n3291,n3195,n3196);
and (n3292,n157,n34);
and (n3293,n3294,n3295);
xor (n3294,n3291,n3292);
or (n3295,n3296,n3299);
and (n3296,n3297,n3298);
xor (n3297,n3201,n3202);
and (n3298,n44,n34);
and (n3299,n3300,n3301);
xor (n3300,n3297,n3298);
or (n3301,n3302,n3305);
and (n3302,n3303,n3304);
xor (n3303,n3207,n3208);
and (n3304,n38,n34);
and (n3305,n3306,n3307);
xor (n3306,n3303,n3304);
or (n3307,n3308,n3311);
and (n3308,n3309,n3310);
xor (n3309,n3213,n3214);
and (n3310,n197,n34);
and (n3311,n3312,n3313);
xor (n3312,n3309,n3310);
or (n3313,n3314,n3317);
and (n3314,n3315,n3316);
xor (n3315,n3219,n3220);
and (n3316,n374,n34);
and (n3317,n3318,n3319);
xor (n3318,n3315,n3316);
or (n3319,n3320,n3323);
and (n3320,n3321,n3322);
xor (n3321,n3225,n3226);
and (n3322,n368,n34);
and (n3323,n3324,n3325);
xor (n3324,n3321,n3322);
or (n3325,n3326,n3329);
and (n3326,n3327,n3328);
xor (n3327,n3231,n3232);
and (n3328,n387,n34);
and (n3329,n3330,n3331);
xor (n3330,n3327,n3328);
or (n3331,n3332,n3335);
and (n3332,n3333,n3334);
xor (n3333,n3237,n3238);
and (n3334,n381,n34);
and (n3335,n3336,n3337);
xor (n3336,n3333,n3334);
or (n3337,n3338,n3341);
and (n3338,n3339,n3340);
xor (n3339,n3243,n3244);
and (n3340,n534,n34);
and (n3341,n3342,n3343);
xor (n3342,n3339,n3340);
and (n3343,n3344,n3345);
xor (n3344,n3249,n3250);
and (n3345,n594,n34);
or (n3346,n3347,n3349);
and (n3347,n3348,n3262);
xor (n3348,n3258,n3259);
and (n3349,n3350,n3351);
xor (n3350,n3348,n3262);
or (n3351,n3352,n3354);
and (n3352,n3353,n3268);
xor (n3353,n3264,n3265);
and (n3354,n3355,n3356);
xor (n3355,n3353,n3268);
or (n3356,n3357,n3359);
and (n3357,n3358,n3274);
xor (n3358,n3270,n3271);
and (n3359,n3360,n3361);
xor (n3360,n3358,n3274);
or (n3361,n3362,n3364);
and (n3362,n3363,n3280);
xor (n3363,n3276,n3277);
and (n3364,n3365,n3366);
xor (n3365,n3363,n3280);
or (n3366,n3367,n3369);
and (n3367,n3368,n3286);
xor (n3368,n3282,n3283);
and (n3369,n3370,n3371);
xor (n3370,n3368,n3286);
or (n3371,n3372,n3374);
and (n3372,n3373,n3292);
xor (n3373,n3288,n3289);
and (n3374,n3375,n3376);
xor (n3375,n3373,n3292);
or (n3376,n3377,n3379);
and (n3377,n3378,n3298);
xor (n3378,n3294,n3295);
and (n3379,n3380,n3381);
xor (n3380,n3378,n3298);
or (n3381,n3382,n3384);
and (n3382,n3383,n3304);
xor (n3383,n3300,n3301);
and (n3384,n3385,n3386);
xor (n3385,n3383,n3304);
or (n3386,n3387,n3389);
and (n3387,n3388,n3310);
xor (n3388,n3306,n3307);
and (n3389,n3390,n3391);
xor (n3390,n3388,n3310);
or (n3391,n3392,n3394);
and (n3392,n3393,n3316);
xor (n3393,n3312,n3313);
and (n3394,n3395,n3396);
xor (n3395,n3393,n3316);
or (n3396,n3397,n3399);
and (n3397,n3398,n3322);
xor (n3398,n3318,n3319);
and (n3399,n3400,n3401);
xor (n3400,n3398,n3322);
or (n3401,n3402,n3404);
and (n3402,n3403,n3328);
xor (n3403,n3324,n3325);
and (n3404,n3405,n3406);
xor (n3405,n3403,n3328);
or (n3406,n3407,n3409);
and (n3407,n3408,n3334);
xor (n3408,n3330,n3331);
and (n3409,n3410,n3411);
xor (n3410,n3408,n3334);
or (n3411,n3412,n3414);
and (n3412,n3413,n3340);
xor (n3413,n3336,n3337);
and (n3414,n3415,n3416);
xor (n3415,n3413,n3340);
and (n3416,n3417,n3345);
xor (n3417,n3342,n3343);
or (n3418,n3419,n3421);
and (n3419,n3420,n3268);
xor (n3420,n3350,n3351);
and (n3421,n3422,n3423);
xor (n3422,n3420,n3268);
or (n3423,n3424,n3426);
and (n3424,n3425,n3274);
xor (n3425,n3355,n3356);
and (n3426,n3427,n3428);
xor (n3427,n3425,n3274);
or (n3428,n3429,n3431);
and (n3429,n3430,n3280);
xor (n3430,n3360,n3361);
and (n3431,n3432,n3433);
xor (n3432,n3430,n3280);
or (n3433,n3434,n3436);
and (n3434,n3435,n3286);
xor (n3435,n3365,n3366);
and (n3436,n3437,n3438);
xor (n3437,n3435,n3286);
or (n3438,n3439,n3441);
and (n3439,n3440,n3292);
xor (n3440,n3370,n3371);
and (n3441,n3442,n3443);
xor (n3442,n3440,n3292);
or (n3443,n3444,n3446);
and (n3444,n3445,n3298);
xor (n3445,n3375,n3376);
and (n3446,n3447,n3448);
xor (n3447,n3445,n3298);
or (n3448,n3449,n3451);
and (n3449,n3450,n3304);
xor (n3450,n3380,n3381);
and (n3451,n3452,n3453);
xor (n3452,n3450,n3304);
or (n3453,n3454,n3456);
and (n3454,n3455,n3310);
xor (n3455,n3385,n3386);
and (n3456,n3457,n3458);
xor (n3457,n3455,n3310);
or (n3458,n3459,n3461);
and (n3459,n3460,n3316);
xor (n3460,n3390,n3391);
and (n3461,n3462,n3463);
xor (n3462,n3460,n3316);
or (n3463,n3464,n3466);
and (n3464,n3465,n3322);
xor (n3465,n3395,n3396);
and (n3466,n3467,n3468);
xor (n3467,n3465,n3322);
or (n3468,n3469,n3471);
and (n3469,n3470,n3328);
xor (n3470,n3400,n3401);
and (n3471,n3472,n3473);
xor (n3472,n3470,n3328);
or (n3473,n3474,n3476);
and (n3474,n3475,n3334);
xor (n3475,n3405,n3406);
and (n3476,n3477,n3478);
xor (n3477,n3475,n3334);
or (n3478,n3479,n3481);
and (n3479,n3480,n3340);
xor (n3480,n3410,n3411);
and (n3481,n3482,n3483);
xor (n3482,n3480,n3340);
and (n3483,n3484,n3345);
xor (n3484,n3415,n3416);
or (n3485,n3486,n3488);
and (n3486,n3487,n3274);
xor (n3487,n3422,n3423);
and (n3488,n3489,n3490);
xor (n3489,n3487,n3274);
or (n3490,n3491,n3493);
and (n3491,n3492,n3280);
xor (n3492,n3427,n3428);
and (n3493,n3494,n3495);
xor (n3494,n3492,n3280);
or (n3495,n3496,n3498);
and (n3496,n3497,n3286);
xor (n3497,n3432,n3433);
and (n3498,n3499,n3500);
xor (n3499,n3497,n3286);
or (n3500,n3501,n3503);
and (n3501,n3502,n3292);
xor (n3502,n3437,n3438);
and (n3503,n3504,n3505);
xor (n3504,n3502,n3292);
or (n3505,n3506,n3508);
and (n3506,n3507,n3298);
xor (n3507,n3442,n3443);
and (n3508,n3509,n3510);
xor (n3509,n3507,n3298);
or (n3510,n3511,n3513);
and (n3511,n3512,n3304);
xor (n3512,n3447,n3448);
and (n3513,n3514,n3515);
xor (n3514,n3512,n3304);
or (n3515,n3516,n3518);
and (n3516,n3517,n3310);
xor (n3517,n3452,n3453);
and (n3518,n3519,n3520);
xor (n3519,n3517,n3310);
or (n3520,n3521,n3523);
and (n3521,n3522,n3316);
xor (n3522,n3457,n3458);
and (n3523,n3524,n3525);
xor (n3524,n3522,n3316);
or (n3525,n3526,n3528);
and (n3526,n3527,n3322);
xor (n3527,n3462,n3463);
and (n3528,n3529,n3530);
xor (n3529,n3527,n3322);
or (n3530,n3531,n3533);
and (n3531,n3532,n3328);
xor (n3532,n3467,n3468);
and (n3533,n3534,n3535);
xor (n3534,n3532,n3328);
or (n3535,n3536,n3538);
and (n3536,n3537,n3334);
xor (n3537,n3472,n3473);
and (n3538,n3539,n3540);
xor (n3539,n3537,n3334);
or (n3540,n3541,n3543);
and (n3541,n3542,n3340);
xor (n3542,n3477,n3478);
and (n3543,n3544,n3545);
xor (n3544,n3542,n3340);
and (n3545,n3546,n3345);
xor (n3546,n3482,n3483);
or (n3547,n3548,n3550);
and (n3548,n3549,n3280);
xor (n3549,n3489,n3490);
and (n3550,n3551,n3552);
xor (n3551,n3549,n3280);
or (n3552,n3553,n3555);
and (n3553,n3554,n3286);
xor (n3554,n3494,n3495);
and (n3555,n3556,n3557);
xor (n3556,n3554,n3286);
or (n3557,n3558,n3560);
and (n3558,n3559,n3292);
xor (n3559,n3499,n3500);
and (n3560,n3561,n3562);
xor (n3561,n3559,n3292);
or (n3562,n3563,n3565);
and (n3563,n3564,n3298);
xor (n3564,n3504,n3505);
and (n3565,n3566,n3567);
xor (n3566,n3564,n3298);
or (n3567,n3568,n3570);
and (n3568,n3569,n3304);
xor (n3569,n3509,n3510);
and (n3570,n3571,n3572);
xor (n3571,n3569,n3304);
or (n3572,n3573,n3575);
and (n3573,n3574,n3310);
xor (n3574,n3514,n3515);
and (n3575,n3576,n3577);
xor (n3576,n3574,n3310);
or (n3577,n3578,n3580);
and (n3578,n3579,n3316);
xor (n3579,n3519,n3520);
and (n3580,n3581,n3582);
xor (n3581,n3579,n3316);
or (n3582,n3583,n3585);
and (n3583,n3584,n3322);
xor (n3584,n3524,n3525);
and (n3585,n3586,n3587);
xor (n3586,n3584,n3322);
or (n3587,n3588,n3590);
and (n3588,n3589,n3328);
xor (n3589,n3529,n3530);
and (n3590,n3591,n3592);
xor (n3591,n3589,n3328);
or (n3592,n3593,n3595);
and (n3593,n3594,n3334);
xor (n3594,n3534,n3535);
and (n3595,n3596,n3597);
xor (n3596,n3594,n3334);
or (n3597,n3598,n3600);
and (n3598,n3599,n3340);
xor (n3599,n3539,n3540);
and (n3600,n3601,n3602);
xor (n3601,n3599,n3340);
and (n3602,n3603,n3345);
xor (n3603,n3544,n3545);
or (n3604,n3605,n3607);
and (n3605,n3606,n3286);
xor (n3606,n3551,n3552);
and (n3607,n3608,n3609);
xor (n3608,n3606,n3286);
or (n3609,n3610,n3612);
and (n3610,n3611,n3292);
xor (n3611,n3556,n3557);
and (n3612,n3613,n3614);
xor (n3613,n3611,n3292);
or (n3614,n3615,n3617);
and (n3615,n3616,n3298);
xor (n3616,n3561,n3562);
and (n3617,n3618,n3619);
xor (n3618,n3616,n3298);
or (n3619,n3620,n3622);
and (n3620,n3621,n3304);
xor (n3621,n3566,n3567);
and (n3622,n3623,n3624);
xor (n3623,n3621,n3304);
or (n3624,n3625,n3627);
and (n3625,n3626,n3310);
xor (n3626,n3571,n3572);
and (n3627,n3628,n3629);
xor (n3628,n3626,n3310);
or (n3629,n3630,n3632);
and (n3630,n3631,n3316);
xor (n3631,n3576,n3577);
and (n3632,n3633,n3634);
xor (n3633,n3631,n3316);
or (n3634,n3635,n3637);
and (n3635,n3636,n3322);
xor (n3636,n3581,n3582);
and (n3637,n3638,n3639);
xor (n3638,n3636,n3322);
or (n3639,n3640,n3642);
and (n3640,n3641,n3328);
xor (n3641,n3586,n3587);
and (n3642,n3643,n3644);
xor (n3643,n3641,n3328);
or (n3644,n3645,n3647);
and (n3645,n3646,n3334);
xor (n3646,n3591,n3592);
and (n3647,n3648,n3649);
xor (n3648,n3646,n3334);
or (n3649,n3650,n3652);
and (n3650,n3651,n3340);
xor (n3651,n3596,n3597);
and (n3652,n3653,n3654);
xor (n3653,n3651,n3340);
and (n3654,n3655,n3345);
xor (n3655,n3601,n3602);
or (n3656,n3657,n3659);
and (n3657,n3658,n3292);
xor (n3658,n3608,n3609);
and (n3659,n3660,n3661);
xor (n3660,n3658,n3292);
or (n3661,n3662,n3664);
and (n3662,n3663,n3298);
xor (n3663,n3613,n3614);
and (n3664,n3665,n3666);
xor (n3665,n3663,n3298);
or (n3666,n3667,n3669);
and (n3667,n3668,n3304);
xor (n3668,n3618,n3619);
and (n3669,n3670,n3671);
xor (n3670,n3668,n3304);
or (n3671,n3672,n3674);
and (n3672,n3673,n3310);
xor (n3673,n3623,n3624);
and (n3674,n3675,n3676);
xor (n3675,n3673,n3310);
or (n3676,n3677,n3679);
and (n3677,n3678,n3316);
xor (n3678,n3628,n3629);
and (n3679,n3680,n3681);
xor (n3680,n3678,n3316);
or (n3681,n3682,n3684);
and (n3682,n3683,n3322);
xor (n3683,n3633,n3634);
and (n3684,n3685,n3686);
xor (n3685,n3683,n3322);
or (n3686,n3687,n3689);
and (n3687,n3688,n3328);
xor (n3688,n3638,n3639);
and (n3689,n3690,n3691);
xor (n3690,n3688,n3328);
or (n3691,n3692,n3694);
and (n3692,n3693,n3334);
xor (n3693,n3643,n3644);
and (n3694,n3695,n3696);
xor (n3695,n3693,n3334);
or (n3696,n3697,n3699);
and (n3697,n3698,n3340);
xor (n3698,n3648,n3649);
and (n3699,n3700,n3701);
xor (n3700,n3698,n3340);
and (n3701,n3702,n3345);
xor (n3702,n3653,n3654);
or (n3703,n3704,n3706);
and (n3704,n3705,n3298);
xor (n3705,n3660,n3661);
and (n3706,n3707,n3708);
xor (n3707,n3705,n3298);
or (n3708,n3709,n3711);
and (n3709,n3710,n3304);
xor (n3710,n3665,n3666);
and (n3711,n3712,n3713);
xor (n3712,n3710,n3304);
or (n3713,n3714,n3716);
and (n3714,n3715,n3310);
xor (n3715,n3670,n3671);
and (n3716,n3717,n3718);
xor (n3717,n3715,n3310);
or (n3718,n3719,n3721);
and (n3719,n3720,n3316);
xor (n3720,n3675,n3676);
and (n3721,n3722,n3723);
xor (n3722,n3720,n3316);
or (n3723,n3724,n3726);
and (n3724,n3725,n3322);
xor (n3725,n3680,n3681);
and (n3726,n3727,n3728);
xor (n3727,n3725,n3322);
or (n3728,n3729,n3731);
and (n3729,n3730,n3328);
xor (n3730,n3685,n3686);
and (n3731,n3732,n3733);
xor (n3732,n3730,n3328);
or (n3733,n3734,n3736);
and (n3734,n3735,n3334);
xor (n3735,n3690,n3691);
and (n3736,n3737,n3738);
xor (n3737,n3735,n3334);
or (n3738,n3739,n3741);
and (n3739,n3740,n3340);
xor (n3740,n3695,n3696);
and (n3741,n3742,n3743);
xor (n3742,n3740,n3340);
and (n3743,n3744,n3345);
xor (n3744,n3700,n3701);
or (n3745,n3746,n3748);
and (n3746,n3747,n3304);
xor (n3747,n3707,n3708);
and (n3748,n3749,n3750);
xor (n3749,n3747,n3304);
or (n3750,n3751,n3753);
and (n3751,n3752,n3310);
xor (n3752,n3712,n3713);
and (n3753,n3754,n3755);
xor (n3754,n3752,n3310);
or (n3755,n3756,n3758);
and (n3756,n3757,n3316);
xor (n3757,n3717,n3718);
and (n3758,n3759,n3760);
xor (n3759,n3757,n3316);
or (n3760,n3761,n3763);
and (n3761,n3762,n3322);
xor (n3762,n3722,n3723);
and (n3763,n3764,n3765);
xor (n3764,n3762,n3322);
or (n3765,n3766,n3768);
and (n3766,n3767,n3328);
xor (n3767,n3727,n3728);
and (n3768,n3769,n3770);
xor (n3769,n3767,n3328);
or (n3770,n3771,n3773);
and (n3771,n3772,n3334);
xor (n3772,n3732,n3733);
and (n3773,n3774,n3775);
xor (n3774,n3772,n3334);
or (n3775,n3776,n3778);
and (n3776,n3777,n3340);
xor (n3777,n3737,n3738);
and (n3778,n3779,n3780);
xor (n3779,n3777,n3340);
and (n3780,n3781,n3345);
xor (n3781,n3742,n3743);
or (n3782,n3783,n3785);
and (n3783,n3784,n3310);
xor (n3784,n3749,n3750);
and (n3785,n3786,n3787);
xor (n3786,n3784,n3310);
or (n3787,n3788,n3790);
and (n3788,n3789,n3316);
xor (n3789,n3754,n3755);
and (n3790,n3791,n3792);
xor (n3791,n3789,n3316);
or (n3792,n3793,n3795);
and (n3793,n3794,n3322);
xor (n3794,n3759,n3760);
and (n3795,n3796,n3797);
xor (n3796,n3794,n3322);
or (n3797,n3798,n3800);
and (n3798,n3799,n3328);
xor (n3799,n3764,n3765);
and (n3800,n3801,n3802);
xor (n3801,n3799,n3328);
or (n3802,n3803,n3805);
and (n3803,n3804,n3334);
xor (n3804,n3769,n3770);
and (n3805,n3806,n3807);
xor (n3806,n3804,n3334);
or (n3807,n3808,n3810);
and (n3808,n3809,n3340);
xor (n3809,n3774,n3775);
and (n3810,n3811,n3812);
xor (n3811,n3809,n3340);
and (n3812,n3813,n3345);
xor (n3813,n3779,n3780);
or (n3814,n3815,n3817);
and (n3815,n3816,n3316);
xor (n3816,n3786,n3787);
and (n3817,n3818,n3819);
xor (n3818,n3816,n3316);
or (n3819,n3820,n3822);
and (n3820,n3821,n3322);
xor (n3821,n3791,n3792);
and (n3822,n3823,n3824);
xor (n3823,n3821,n3322);
or (n3824,n3825,n3827);
and (n3825,n3826,n3328);
xor (n3826,n3796,n3797);
and (n3827,n3828,n3829);
xor (n3828,n3826,n3328);
or (n3829,n3830,n3832);
and (n3830,n3831,n3334);
xor (n3831,n3801,n3802);
and (n3832,n3833,n3834);
xor (n3833,n3831,n3334);
or (n3834,n3835,n3837);
and (n3835,n3836,n3340);
xor (n3836,n3806,n3807);
and (n3837,n3838,n3839);
xor (n3838,n3836,n3340);
and (n3839,n3840,n3345);
xor (n3840,n3811,n3812);
or (n3841,n3842,n3844);
and (n3842,n3843,n3322);
xor (n3843,n3818,n3819);
and (n3844,n3845,n3846);
xor (n3845,n3843,n3322);
or (n3846,n3847,n3849);
and (n3847,n3848,n3328);
xor (n3848,n3823,n3824);
and (n3849,n3850,n3851);
xor (n3850,n3848,n3328);
or (n3851,n3852,n3854);
and (n3852,n3853,n3334);
xor (n3853,n3828,n3829);
and (n3854,n3855,n3856);
xor (n3855,n3853,n3334);
or (n3856,n3857,n3859);
and (n3857,n3858,n3340);
xor (n3858,n3833,n3834);
and (n3859,n3860,n3861);
xor (n3860,n3858,n3340);
and (n3861,n3862,n3345);
xor (n3862,n3838,n3839);
or (n3863,n3864,n3866);
and (n3864,n3865,n3328);
xor (n3865,n3845,n3846);
and (n3866,n3867,n3868);
xor (n3867,n3865,n3328);
or (n3868,n3869,n3871);
and (n3869,n3870,n3334);
xor (n3870,n3850,n3851);
and (n3871,n3872,n3873);
xor (n3872,n3870,n3334);
or (n3873,n3874,n3876);
and (n3874,n3875,n3340);
xor (n3875,n3855,n3856);
and (n3876,n3877,n3878);
xor (n3877,n3875,n3340);
and (n3878,n3879,n3345);
xor (n3879,n3860,n3861);
or (n3880,n3881,n3883);
and (n3881,n3882,n3334);
xor (n3882,n3867,n3868);
and (n3883,n3884,n3885);
xor (n3884,n3882,n3334);
or (n3885,n3886,n3888);
and (n3886,n3887,n3340);
xor (n3887,n3872,n3873);
and (n3888,n3889,n3890);
xor (n3889,n3887,n3340);
and (n3890,n3891,n3345);
xor (n3891,n3877,n3878);
or (n3892,n3893,n3895);
and (n3893,n3894,n3340);
xor (n3894,n3884,n3885);
and (n3895,n3896,n3897);
xor (n3896,n3894,n3340);
and (n3897,n3898,n3345);
xor (n3898,n3889,n3890);
and (n3899,n3900,n3345);
xor (n3900,n3896,n3897);
endmodule
