module top (out,n24,n29,n30,n31,n33,n34,n45,n48,n51
        ,n54,n57,n60,n63,n66,n69,n71,n74,n85,n95
        ,n100,n103,n106,n109,n112,n115,n118,n121,n124,n127
        ,n130,n132,n134,n142,n156,n161,n194,n199,n202,n205
        ,n208,n221,n266,n277,n289,n294,n297,n300,n303,n306
        ,n309,n325,n398,n408,n441,n446,n449,n636,n1083,n1119);
output out;
input n24;
input n29;
input n30;
input n31;
input n33;
input n34;
input n45;
input n48;
input n51;
input n54;
input n57;
input n60;
input n63;
input n66;
input n69;
input n71;
input n74;
input n85;
input n95;
input n100;
input n103;
input n106;
input n109;
input n112;
input n115;
input n118;
input n121;
input n124;
input n127;
input n130;
input n132;
input n134;
input n142;
input n156;
input n161;
input n194;
input n199;
input n202;
input n205;
input n208;
input n221;
input n266;
input n277;
input n289;
input n294;
input n297;
input n300;
input n303;
input n306;
input n309;
input n325;
input n398;
input n408;
input n441;
input n446;
input n449;
input n636;
input n1083;
input n1119;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n25;
wire n26;
wire n27;
wire n28;
wire n32;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n46;
wire n47;
wire n49;
wire n50;
wire n52;
wire n53;
wire n55;
wire n56;
wire n58;
wire n59;
wire n61;
wire n62;
wire n64;
wire n65;
wire n67;
wire n68;
wire n70;
wire n72;
wire n73;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n96;
wire n97;
wire n98;
wire n99;
wire n101;
wire n102;
wire n104;
wire n105;
wire n107;
wire n108;
wire n110;
wire n111;
wire n113;
wire n114;
wire n116;
wire n117;
wire n119;
wire n120;
wire n122;
wire n123;
wire n125;
wire n126;
wire n128;
wire n129;
wire n131;
wire n133;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n157;
wire n158;
wire n159;
wire n160;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n195;
wire n196;
wire n197;
wire n198;
wire n200;
wire n201;
wire n203;
wire n204;
wire n206;
wire n207;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n290;
wire n291;
wire n292;
wire n293;
wire n295;
wire n296;
wire n298;
wire n299;
wire n301;
wire n302;
wire n304;
wire n305;
wire n307;
wire n308;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n442;
wire n443;
wire n444;
wire n445;
wire n447;
wire n448;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2988;
wire n2989;
wire n2990;
wire n2991;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2996;
wire n2997;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3003;
wire n3004;
wire n3005;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3010;
wire n3011;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3038;
wire n3039;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
wire n3056;
wire n3057;
wire n3058;
wire n3059;
wire n3060;
wire n3061;
wire n3062;
wire n3063;
wire n3064;
wire n3065;
wire n3066;
wire n3067;
wire n3068;
wire n3069;
wire n3070;
wire n3071;
wire n3072;
wire n3073;
wire n3074;
wire n3075;
wire n3076;
wire n3077;
wire n3078;
wire n3079;
wire n3080;
wire n3081;
wire n3082;
wire n3083;
wire n3084;
wire n3085;
wire n3086;
wire n3087;
wire n3088;
wire n3089;
wire n3090;
wire n3091;
wire n3092;
wire n3093;
wire n3094;
wire n3095;
wire n3096;
wire n3097;
wire n3098;
wire n3099;
wire n3100;
wire n3101;
wire n3102;
wire n3103;
wire n3104;
wire n3105;
wire n3106;
wire n3107;
wire n3108;
wire n3109;
wire n3110;
wire n3111;
wire n3112;
wire n3113;
wire n3114;
wire n3115;
wire n3116;
wire n3117;
wire n3118;
wire n3119;
wire n3120;
wire n3121;
wire n3122;
wire n3123;
wire n3124;
wire n3125;
wire n3126;
wire n3127;
wire n3128;
wire n3129;
wire n3130;
wire n3131;
wire n3132;
wire n3133;
wire n3134;
wire n3135;
wire n3136;
wire n3137;
wire n3138;
wire n3139;
wire n3140;
wire n3141;
wire n3142;
wire n3143;
wire n3144;
wire n3145;
wire n3146;
wire n3147;
wire n3148;
wire n3149;
wire n3150;
wire n3151;
wire n3152;
wire n3153;
wire n3154;
wire n3155;
wire n3156;
wire n3157;
wire n3158;
wire n3159;
wire n3160;
wire n3161;
wire n3162;
wire n3163;
wire n3164;
wire n3165;
wire n3166;
wire n3167;
wire n3168;
wire n3169;
wire n3170;
wire n3171;
wire n3172;
wire n3173;
wire n3174;
wire n3175;
wire n3176;
wire n3177;
wire n3178;
wire n3179;
wire n3180;
wire n3181;
wire n3182;
wire n3183;
wire n3184;
wire n3185;
wire n3186;
wire n3187;
wire n3188;
wire n3189;
wire n3190;
wire n3191;
wire n3192;
wire n3193;
wire n3194;
wire n3195;
wire n3196;
wire n3197;
wire n3198;
wire n3199;
wire n3200;
wire n3201;
wire n3202;
wire n3203;
wire n3204;
wire n3205;
wire n3206;
wire n3207;
wire n3208;
wire n3209;
wire n3210;
wire n3211;
wire n3212;
wire n3213;
wire n3214;
wire n3215;
wire n3216;
wire n3217;
wire n3218;
wire n3219;
wire n3220;
wire n3221;
wire n3222;
wire n3223;
wire n3224;
wire n3225;
wire n3226;
wire n3227;
wire n3228;
wire n3229;
wire n3230;
wire n3231;
wire n3232;
wire n3233;
wire n3234;
wire n3235;
wire n3236;
wire n3237;
wire n3238;
wire n3239;
wire n3240;
wire n3241;
wire n3242;
wire n3243;
wire n3244;
wire n3245;
wire n3246;
wire n3247;
wire n3248;
wire n3249;
wire n3250;
wire n3251;
wire n3252;
wire n3253;
wire n3254;
wire n3255;
wire n3256;
wire n3257;
wire n3258;
wire n3259;
wire n3260;
wire n3261;
wire n3262;
wire n3263;
wire n3264;
wire n3265;
wire n3266;
wire n3267;
wire n3268;
wire n3269;
wire n3270;
wire n3271;
wire n3272;
wire n3273;
wire n3274;
wire n3275;
wire n3276;
wire n3277;
wire n3278;
wire n3279;
wire n3280;
wire n3281;
wire n3282;
wire n3283;
wire n3284;
wire n3285;
wire n3286;
wire n3287;
wire n3288;
wire n3289;
wire n3290;
wire n3291;
wire n3292;
wire n3293;
wire n3294;
wire n3295;
wire n3296;
wire n3297;
wire n3298;
wire n3299;
wire n3300;
wire n3301;
wire n3302;
wire n3303;
wire n3304;
wire n3305;
wire n3306;
wire n3307;
wire n3308;
wire n3309;
wire n3310;
wire n3311;
wire n3312;
wire n3313;
wire n3314;
wire n3315;
wire n3316;
wire n3317;
wire n3318;
wire n3319;
wire n3320;
wire n3321;
wire n3322;
wire n3323;
wire n3324;
wire n3325;
wire n3326;
wire n3327;
wire n3328;
wire n3329;
wire n3330;
wire n3331;
wire n3332;
wire n3333;
wire n3334;
wire n3335;
wire n3336;
wire n3337;
wire n3338;
wire n3339;
wire n3340;
wire n3341;
wire n3342;
wire n3343;
wire n3344;
wire n3345;
wire n3346;
wire n3347;
wire n3348;
wire n3349;
wire n3350;
wire n3351;
wire n3352;
wire n3353;
wire n3354;
wire n3355;
wire n3356;
wire n3357;
wire n3358;
wire n3359;
wire n3360;
wire n3361;
wire n3362;
wire n3363;
wire n3364;
wire n3365;
wire n3366;
wire n3367;
wire n3368;
wire n3369;
wire n3370;
wire n3371;
wire n3372;
wire n3373;
wire n3374;
wire n3375;
wire n3376;
wire n3377;
wire n3378;
wire n3379;
wire n3380;
wire n3381;
wire n3382;
wire n3383;
wire n3384;
wire n3385;
wire n3386;
wire n3387;
wire n3388;
wire n3389;
wire n3390;
wire n3391;
wire n3392;
wire n3393;
wire n3394;
wire n3395;
wire n3396;
wire n3397;
wire n3398;
wire n3399;
wire n3400;
wire n3401;
wire n3402;
wire n3403;
wire n3404;
wire n3405;
wire n3406;
wire n3407;
wire n3408;
wire n3409;
wire n3410;
wire n3411;
wire n3412;
wire n3413;
wire n3414;
wire n3415;
wire n3416;
wire n3417;
wire n3418;
wire n3419;
wire n3420;
wire n3421;
wire n3422;
wire n3423;
wire n3424;
wire n3425;
wire n3426;
wire n3427;
wire n3428;
wire n3429;
wire n3430;
wire n3431;
wire n3432;
wire n3433;
wire n3434;
wire n3435;
wire n3436;
wire n3437;
wire n3438;
wire n3439;
wire n3440;
wire n3441;
wire n3442;
wire n3443;
wire n3444;
wire n3445;
wire n3446;
wire n3447;
wire n3448;
wire n3449;
wire n3450;
wire n3451;
wire n3452;
wire n3453;
wire n3454;
wire n3455;
wire n3456;
wire n3457;
wire n3458;
wire n3459;
wire n3460;
wire n3461;
wire n3462;
wire n3463;
wire n3464;
wire n3465;
wire n3466;
wire n3467;
wire n3468;
wire n3469;
wire n3470;
wire n3471;
wire n3472;
wire n3473;
wire n3474;
wire n3475;
wire n3476;
wire n3477;
wire n3478;
wire n3479;
wire n3480;
wire n3481;
wire n3482;
wire n3483;
wire n3484;
wire n3485;
wire n3486;
wire n3487;
wire n3488;
wire n3489;
wire n3490;
wire n3491;
wire n3492;
wire n3493;
wire n3494;
wire n3495;
wire n3496;
wire n3497;
wire n3498;
wire n3499;
wire n3500;
wire n3501;
wire n3502;
wire n3503;
wire n3504;
wire n3505;
wire n3506;
wire n3507;
wire n3508;
wire n3509;
wire n3510;
wire n3511;
wire n3512;
wire n3513;
wire n3514;
wire n3515;
wire n3516;
wire n3517;
wire n3518;
wire n3519;
wire n3520;
wire n3521;
wire n3522;
wire n3523;
wire n3524;
wire n3525;
wire n3526;
wire n3527;
wire n3528;
wire n3529;
wire n3530;
wire n3531;
wire n3532;
wire n3533;
wire n3534;
wire n3535;
wire n3536;
wire n3537;
wire n3538;
wire n3539;
wire n3540;
wire n3541;
wire n3542;
wire n3543;
wire n3544;
wire n3545;
wire n3546;
wire n3547;
wire n3548;
wire n3549;
wire n3550;
wire n3551;
wire n3552;
wire n3553;
wire n3554;
wire n3555;
wire n3556;
wire n3557;
wire n3558;
wire n3559;
wire n3560;
wire n3561;
wire n3562;
wire n3563;
wire n3564;
wire n3565;
wire n3566;
wire n3567;
wire n3568;
wire n3569;
wire n3570;
wire n3571;
wire n3572;
wire n3573;
wire n3574;
wire n3575;
wire n3576;
wire n3577;
wire n3578;
wire n3579;
wire n3580;
wire n3581;
wire n3582;
wire n3583;
wire n3584;
wire n3585;
wire n3586;
wire n3587;
wire n3588;
wire n3589;
wire n3590;
wire n3591;
wire n3592;
wire n3593;
wire n3594;
wire n3595;
wire n3596;
wire n3597;
wire n3598;
wire n3599;
wire n3600;
wire n3601;
wire n3602;
wire n3603;
wire n3604;
wire n3605;
wire n3606;
wire n3607;
wire n3608;
wire n3609;
wire n3610;
wire n3611;
wire n3612;
wire n3613;
wire n3614;
wire n3615;
wire n3616;
wire n3617;
wire n3618;
wire n3619;
wire n3620;
wire n3621;
wire n3622;
wire n3623;
wire n3624;
wire n3625;
wire n3626;
wire n3627;
wire n3628;
wire n3629;
wire n3630;
wire n3631;
wire n3632;
wire n3633;
wire n3634;
wire n3635;
wire n3636;
wire n3637;
wire n3638;
wire n3639;
wire n3640;
wire n3641;
wire n3642;
wire n3643;
wire n3644;
wire n3645;
wire n3646;
wire n3647;
wire n3648;
wire n3649;
wire n3650;
wire n3651;
wire n3652;
wire n3653;
wire n3654;
wire n3655;
wire n3656;
wire n3657;
wire n3658;
wire n3659;
wire n3660;
wire n3661;
wire n3662;
wire n3663;
wire n3664;
wire n3665;
wire n3666;
wire n3667;
wire n3668;
wire n3669;
wire n3670;
wire n3671;
wire n3672;
wire n3673;
wire n3674;
wire n3675;
wire n3676;
wire n3677;
wire n3678;
wire n3679;
wire n3680;
wire n3681;
wire n3682;
wire n3683;
wire n3684;
wire n3685;
wire n3686;
wire n3687;
wire n3688;
wire n3689;
wire n3690;
wire n3691;
wire n3692;
wire n3693;
wire n3694;
wire n3695;
wire n3696;
wire n3697;
wire n3698;
wire n3699;
wire n3700;
wire n3701;
wire n3702;
wire n3703;
wire n3704;
wire n3705;
wire n3706;
wire n3707;
wire n3708;
wire n3709;
wire n3710;
wire n3711;
wire n3712;
wire n3713;
wire n3714;
wire n3715;
wire n3716;
wire n3717;
wire n3718;
wire n3719;
wire n3720;
wire n3721;
wire n3722;
wire n3723;
wire n3724;
wire n3725;
wire n3726;
wire n3727;
wire n3728;
wire n3729;
wire n3730;
wire n3731;
wire n3732;
wire n3733;
wire n3734;
wire n3735;
wire n3736;
wire n3737;
wire n3738;
wire n3739;
wire n3740;
wire n3741;
wire n3742;
wire n3743;
wire n3744;
wire n3745;
wire n3746;
wire n3747;
wire n3748;
wire n3749;
wire n3750;
wire n3751;
wire n3752;
wire n3753;
wire n3754;
wire n3755;
wire n3756;
wire n3757;
wire n3758;
wire n3759;
wire n3760;
wire n3761;
wire n3762;
wire n3763;
wire n3764;
wire n3765;
wire n3766;
wire n3767;
wire n3768;
wire n3769;
wire n3770;
wire n3771;
wire n3772;
wire n3773;
wire n3774;
wire n3775;
wire n3776;
wire n3777;
wire n3778;
wire n3779;
wire n3780;
wire n3781;
wire n3782;
wire n3783;
wire n3784;
wire n3785;
wire n3786;
wire n3787;
wire n3788;
wire n3789;
wire n3790;
wire n3791;
wire n3792;
wire n3793;
wire n3794;
wire n3795;
wire n3796;
wire n3797;
wire n3798;
wire n3799;
wire n3800;
wire n3801;
wire n3802;
wire n3803;
wire n3804;
wire n3805;
wire n3806;
wire n3807;
wire n3808;
wire n3809;
wire n3810;
wire n3811;
wire n3812;
wire n3813;
wire n3814;
wire n3815;
wire n3816;
wire n3817;
wire n3818;
wire n3819;
wire n3820;
wire n3821;
wire n3822;
wire n3823;
wire n3824;
wire n3825;
wire n3826;
wire n3827;
wire n3828;
wire n3829;
wire n3830;
wire n3831;
wire n3832;
wire n3833;
wire n3834;
wire n3835;
wire n3836;
wire n3837;
wire n3838;
wire n3839;
wire n3840;
wire n3841;
wire n3842;
wire n3843;
wire n3844;
wire n3845;
wire n3846;
wire n3847;
wire n3848;
wire n3849;
wire n3850;
wire n3851;
wire n3852;
wire n3853;
wire n3854;
wire n3855;
wire n3856;
wire n3857;
wire n3858;
wire n3859;
wire n3860;
wire n3861;
wire n3862;
wire n3863;
wire n3864;
wire n3865;
wire n3866;
wire n3867;
wire n3868;
wire n3869;
wire n3870;
wire n3871;
wire n3872;
wire n3873;
wire n3874;
wire n3875;
wire n3876;
wire n3877;
wire n3878;
wire n3879;
wire n3880;
wire n3881;
wire n3882;
wire n3883;
wire n3884;
wire n3885;
wire n3886;
wire n3887;
wire n3888;
wire n3889;
wire n3890;
wire n3891;
wire n3892;
wire n3893;
wire n3894;
wire n3895;
wire n3896;
wire n3897;
wire n3898;
wire n3899;
wire n3900;
wire n3901;
wire n3902;
wire n3903;
wire n3904;
wire n3905;
wire n3906;
wire n3907;
wire n3908;
wire n3909;
wire n3910;
wire n3911;
wire n3912;
wire n3913;
wire n3914;
wire n3915;
wire n3916;
wire n3917;
wire n3918;
wire n3919;
wire n3920;
wire n3921;
wire n3922;
wire n3923;
wire n3924;
wire n3925;
wire n3926;
wire n3927;
wire n3928;
wire n3929;
wire n3930;
wire n3931;
wire n3932;
wire n3933;
wire n3934;
wire n3935;
wire n3936;
wire n3937;
wire n3938;
wire n3939;
wire n3940;
wire n3941;
wire n3942;
wire n3943;
wire n3944;
wire n3945;
wire n3946;
wire n3947;
wire n3948;
wire n3949;
wire n3950;
wire n3951;
wire n3952;
wire n3953;
wire n3954;
wire n3955;
wire n3956;
wire n3957;
wire n3958;
wire n3959;
wire n3960;
wire n3961;
wire n3962;
wire n3963;
wire n3964;
wire n3965;
wire n3966;
wire n3967;
wire n3968;
wire n3969;
wire n3970;
wire n3971;
wire n3972;
wire n3973;
wire n3974;
wire n3975;
wire n3976;
wire n3977;
wire n3978;
wire n3979;
wire n3980;
wire n3981;
wire n3982;
wire n3983;
wire n3984;
wire n3985;
wire n3986;
wire n3987;
wire n3988;
wire n3989;
wire n3990;
wire n3991;
wire n3992;
wire n3993;
wire n3994;
wire n3995;
wire n3996;
wire n3997;
wire n3998;
wire n3999;
wire n4000;
wire n4001;
wire n4002;
wire n4003;
wire n4004;
wire n4005;
wire n4006;
wire n4007;
wire n4008;
wire n4009;
wire n4010;
wire n4011;
wire n4012;
wire n4013;
wire n4014;
wire n4015;
wire n4016;
wire n4017;
wire n4018;
wire n4019;
wire n4020;
wire n4021;
wire n4022;
wire n4023;
wire n4024;
wire n4025;
wire n4026;
wire n4027;
wire n4028;
wire n4029;
wire n4030;
wire n4031;
wire n4032;
wire n4033;
wire n4034;
wire n4035;
wire n4036;
wire n4037;
wire n4038;
wire n4039;
wire n4040;
wire n4041;
wire n4042;
wire n4043;
wire n4044;
wire n4045;
wire n4046;
wire n4047;
wire n4048;
wire n4049;
wire n4050;
wire n4051;
wire n4052;
wire n4053;
wire n4054;
wire n4055;
wire n4056;
wire n4057;
wire n4058;
wire n4059;
wire n4060;
wire n4061;
wire n4062;
wire n4063;
wire n4064;
wire n4065;
wire n4066;
wire n4067;
wire n4068;
wire n4069;
wire n4070;
wire n4071;
wire n4072;
wire n4073;
wire n4074;
wire n4075;
wire n4076;
wire n4077;
wire n4078;
wire n4079;
wire n4080;
wire n4081;
wire n4082;
wire n4083;
wire n4084;
wire n4085;
wire n4086;
wire n4087;
wire n4088;
wire n4089;
wire n4090;
wire n4091;
wire n4092;
wire n4093;
wire n4094;
wire n4095;
wire n4096;
wire n4097;
wire n4098;
wire n4099;
wire n4100;
wire n4101;
wire n4102;
wire n4103;
wire n4104;
wire n4105;
wire n4106;
wire n4107;
wire n4108;
wire n4109;
wire n4110;
wire n4111;
wire n4112;
wire n4113;
wire n4114;
wire n4115;
wire n4116;
wire n4117;
wire n4118;
wire n4119;
wire n4120;
wire n4121;
wire n4122;
wire n4123;
wire n4124;
wire n4125;
wire n4126;
wire n4127;
wire n4128;
wire n4129;
wire n4130;
wire n4131;
wire n4132;
wire n4133;
wire n4134;
wire n4135;
wire n4136;
wire n4137;
wire n4138;
wire n4139;
wire n4140;
wire n4141;
wire n4142;
wire n4143;
wire n4144;
wire n4145;
wire n4146;
wire n4147;
wire n4148;
wire n4149;
wire n4150;
wire n4151;
wire n4152;
wire n4153;
wire n4154;
wire n4155;
wire n4156;
wire n4157;
wire n4158;
wire n4159;
wire n4160;
wire n4161;
wire n4162;
wire n4163;
wire n4164;
wire n4165;
wire n4166;
wire n4167;
wire n4168;
wire n4169;
wire n4170;
wire n4171;
wire n4172;
wire n4173;
wire n4174;
wire n4175;
wire n4176;
xor (out,n0,n2388);
nand (n0,n1,n2387);
or (n1,n2,n1172);
not (n2,n3);
or (n3,n4,n1171);
and (n4,n5,n1010);
not (n5,n6);
or (n6,n7,n1009);
and (n7,n8,n881);
xor (n8,n9,n658);
xor (n9,n10,n600);
xor (n10,n11,n431);
or (n11,n12,n430);
and (n12,n13,n368);
xor (n13,n14,n242);
xor (n14,n15,n187);
xor (n15,n16,n148);
nand (n16,n17,n137);
or (n17,n18,n91);
nand (n18,n19,n81);
or (n19,n20,n78);
and (n20,n21,n75);
wire s0n21,s1n21,notn21;
or (n21,s0n21,s1n21);
not(notn21,n72);
and (s0n21,notn21,n22);
and (s1n21,n72,n41);
wire s0n22,s1n22,notn22;
or (n22,s0n22,s1n22);
not(notn22,n25);
and (s0n22,notn22,1'b0);
and (s1n22,n25,n24);
or (n25,n26,n37);
or (n26,n27,n35);
nor (n27,n28,n30,n31,n32,n34);
not (n28,n29);
not (n32,n33);
nor (n35,n29,n36,n31,n32,n34);
not (n36,n30);
or (n37,n38,n40);
and (n38,n28,n30,n31,n32,n39);
not (n39,n34);
nor (n40,n28,n36,n31,n32,n34);
xor (n41,n42,n43);
not (n42,n24);
and (n43,n44,n46);
not (n44,n45);
and (n46,n47,n49);
not (n47,n48);
and (n49,n50,n52);
not (n50,n51);
and (n52,n53,n55);
not (n53,n54);
and (n55,n56,n58);
not (n56,n57);
and (n58,n59,n61);
not (n59,n60);
and (n61,n62,n64);
not (n62,n63);
and (n64,n65,n67);
not (n65,n66);
and (n67,n68,n70);
not (n68,n69);
not (n70,n71);
and (n72,n73,n74);
or (n73,n27,n38);
wire s0n75,s1n75,notn75;
or (n75,s0n75,s1n75);
not(notn75,n72);
and (s0n75,notn75,n76);
and (s1n75,n72,n77);
wire s0n76,s1n76,notn76;
or (n76,s0n76,s1n76);
not(notn76,n25);
and (s0n76,notn76,1'b0);
and (s1n76,n25,n45);
xor (n77,n44,n46);
and (n78,n79,n80);
not (n79,n21);
not (n80,n75);
nand (n81,n82,n89);
or (n82,n79,n83);
wire s0n83,s1n83,notn83;
or (n83,s0n83,s1n83);
not(notn83,n72);
and (s0n83,notn83,n84);
and (s1n83,n72,n86);
wire s0n84,s1n84,notn84;
or (n84,s0n84,s1n84);
not(notn84,n25);
and (s0n84,notn84,1'b0);
and (s1n84,n25,n85);
xor (n86,n87,n88);
not (n87,n85);
and (n88,n42,n43);
or (n89,n90,n21);
not (n90,n83);
nor (n91,n92,n135);
and (n92,n90,n93);
wire s0n93,s1n93,notn93;
or (n93,s0n93,s1n93);
not(notn93,n133);
and (s0n93,notn93,n94);
and (s1n93,n133,n96);
wire s0n94,s1n94,notn94;
or (n94,s0n94,s1n94);
not(notn94,n25);
and (s0n94,notn94,1'b0);
and (s1n94,n25,n95);
xor (n96,n97,n98);
not (n97,n95);
and (n98,n99,n101);
not (n99,n100);
and (n101,n102,n104);
not (n102,n103);
and (n104,n105,n107);
not (n105,n106);
and (n107,n108,n110);
not (n108,n109);
and (n110,n111,n113);
not (n111,n112);
and (n113,n114,n116);
not (n114,n115);
and (n116,n117,n119);
not (n117,n118);
and (n119,n120,n122);
not (n120,n121);
and (n122,n123,n125);
not (n123,n124);
and (n125,n126,n128);
not (n126,n127);
and (n128,n129,n131);
not (n129,n130);
not (n131,n132);
and (n133,n73,n134);
and (n135,n83,n136);
not (n136,n93);
or (n137,n19,n138);
nor (n138,n139,n146);
and (n139,n90,n140);
wire s0n140,s1n140,notn140;
or (n140,s0n140,s1n140);
not(notn140,n133);
and (s0n140,notn140,n141);
and (s1n140,n133,n143);
wire s0n141,s1n141,notn141;
or (n141,s0n141,s1n141);
not(notn141,n25);
and (s0n141,notn141,1'b0);
and (s1n141,n25,n142);
xor (n143,n144,n145);
not (n144,n142);
and (n145,n97,n98);
and (n146,n83,n147);
not (n147,n140);
nand (n148,n149,n178);
or (n149,n150,n171);
or (n150,n151,n168);
nor (n151,n152,n166);
and (n152,n153,n163);
not (n153,n154);
wire s0n154,s1n154,notn154;
or (n154,s0n154,s1n154);
not(notn154,n72);
and (s0n154,notn154,n155);
and (s1n154,n72,n157);
wire s0n155,s1n155,notn155;
or (n155,s0n155,s1n155);
not(notn155,n25);
and (s0n155,notn155,1'b0);
and (s1n155,n25,n156);
xor (n157,n158,n159);
not (n158,n156);
and (n159,n160,n162);
not (n160,n161);
and (n162,n87,n88);
wire s0n163,s1n163,notn163;
or (n163,s0n163,s1n163);
not(notn163,n72);
and (s0n163,notn163,n164);
and (s1n163,n72,n165);
wire s0n164,s1n164,notn164;
or (n164,s0n164,s1n164);
not(notn164,n25);
and (s0n164,notn164,1'b0);
and (s1n164,n25,n161);
xor (n165,n160,n162);
and (n166,n167,n154);
not (n167,n163);
nor (n168,n169,n170);
and (n169,n163,n83);
and (n170,n167,n90);
nor (n171,n172,n176);
and (n172,n153,n173);
wire s0n173,s1n173,notn173;
or (n173,s0n173,s1n173);
not(notn173,n133);
and (s0n173,notn173,n174);
and (s1n173,n133,n175);
wire s0n174,s1n174,notn174;
or (n174,s0n174,s1n174);
not(notn174,n25);
and (s0n174,notn174,1'b0);
and (s1n174,n25,n103);
xor (n175,n102,n104);
and (n176,n154,n177);
not (n177,n173);
or (n178,n179,n180);
not (n179,n168);
nor (n180,n181,n185);
and (n181,n153,n182);
wire s0n182,s1n182,notn182;
or (n182,s0n182,s1n182);
not(notn182,n133);
and (s0n182,notn182,n183);
and (s1n182,n133,n184);
wire s0n183,s1n183,notn183;
or (n183,s0n183,s1n183);
not(notn183,n25);
and (s0n183,notn183,1'b0);
and (s1n183,n25,n100);
xor (n184,n99,n101);
and (n185,n154,n186);
not (n186,n182);
nand (n187,n188,n233);
or (n188,n189,n226);
or (n189,n190,n216);
nor (n190,n191,n213);
and (n191,n192,n210);
wire s0n192,s1n192,notn192;
or (n192,s0n192,s1n192);
not(notn192,n72);
and (s0n192,notn192,n193);
and (s1n192,n72,n195);
wire s0n193,s1n193,notn193;
or (n193,s0n193,s1n193);
not(notn193,n25);
and (s0n193,notn193,1'b0);
and (s1n193,n25,n194);
xor (n195,n196,n197);
not (n196,n194);
and (n197,n198,n200);
not (n198,n199);
and (n200,n201,n203);
not (n201,n202);
and (n203,n204,n206);
not (n204,n205);
and (n206,n207,n209);
not (n207,n208);
and (n209,n158,n159);
wire s0n210,s1n210,notn210;
or (n210,s0n210,s1n210);
not(notn210,n72);
and (s0n210,notn210,n211);
and (s1n210,n72,n212);
wire s0n211,s1n211,notn211;
or (n211,s0n211,s1n211);
not(notn211,n25);
and (s0n211,notn211,1'b0);
and (s1n211,n25,n199);
xor (n212,n198,n200);
and (n213,n214,n215);
not (n214,n192);
not (n215,n210);
nor (n216,n217,n225);
and (n217,n192,n218);
not (n218,n219);
wire s0n219,s1n219,notn219;
or (n219,s0n219,s1n219);
not(notn219,n72);
and (s0n219,notn219,n220);
and (s1n219,n72,n222);
wire s0n220,s1n220,notn220;
or (n220,s0n220,s1n220);
not(notn220,n25);
and (s0n220,notn220,1'b0);
and (s1n220,n25,n221);
xor (n222,n223,n224);
not (n223,n221);
and (n224,n196,n197);
and (n225,n214,n219);
nor (n226,n227,n231);
and (n227,n218,n228);
wire s0n228,s1n228,notn228;
or (n228,s0n228,s1n228);
not(notn228,n133);
and (s0n228,notn228,n229);
and (s1n228,n133,n230);
wire s0n229,s1n229,notn229;
or (n229,s0n229,s1n229);
not(notn229,n25);
and (s0n229,notn229,1'b0);
and (s1n229,n25,n121);
xor (n230,n120,n122);
and (n231,n219,n232);
not (n232,n228);
or (n233,n234,n235);
not (n234,n190);
nor (n235,n236,n240);
and (n236,n237,n218);
wire s0n237,s1n237,notn237;
or (n237,s0n237,s1n237);
not(notn237,n133);
and (s0n237,notn237,n238);
and (s1n237,n133,n239);
wire s0n238,s1n238,notn238;
or (n238,s0n238,s1n238);
not(notn238,n25);
and (s0n238,notn238,1'b0);
and (s1n238,n25,n118);
xor (n239,n117,n119);
and (n240,n241,n219);
not (n241,n237);
xor (n242,n243,n331);
xor (n243,n244,n283);
nand (n244,n245,n272);
or (n245,n246,n262);
nand (n246,n247,n254);
nor (n247,n248,n252);
and (n248,n249,n75);
wire s0n249,s1n249,notn249;
or (n249,s0n249,s1n249);
not(notn249,n72);
and (s0n249,notn249,n250);
and (s1n249,n72,n251);
wire s0n250,s1n250,notn250;
or (n250,s0n250,s1n250);
not(notn250,n25);
and (s0n250,notn250,1'b0);
and (s1n250,n25,n48);
xor (n251,n47,n49);
and (n252,n253,n80);
not (n253,n249);
not (n254,n255);
nor (n255,n256,n260);
and (n256,n257,n249);
wire s0n257,s1n257,notn257;
or (n257,s0n257,s1n257);
not(notn257,n72);
and (s0n257,notn257,n258);
and (s1n257,n72,n259);
wire s0n258,s1n258,notn258;
or (n258,s0n258,s1n258);
not(notn258,n25);
and (s0n258,notn258,1'b0);
and (s1n258,n25,n51);
xor (n259,n50,n52);
and (n260,n261,n253);
not (n261,n257);
nor (n262,n263,n270);
and (n263,n80,n264);
wire s0n264,s1n264,notn264;
or (n264,s0n264,s1n264);
not(notn264,n133);
and (s0n264,notn264,n265);
and (s1n264,n133,n267);
wire s0n265,s1n265,notn265;
or (n265,s0n265,s1n265);
not(notn265,n25);
and (s0n265,notn265,1'b0);
and (s1n265,n25,n266);
xor (n267,n268,n269);
not (n268,n266);
and (n269,n144,n145);
and (n270,n75,n271);
not (n271,n264);
or (n272,n273,n254);
nor (n273,n274,n281);
and (n274,n80,n275);
wire s0n275,s1n275,notn275;
or (n275,s0n275,s1n275);
not(notn275,n133);
and (s0n275,notn275,n276);
and (s1n275,n133,n278);
wire s0n276,s1n276,notn276;
or (n276,s0n276,s1n276);
not(notn276,n25);
and (s0n276,notn276,1'b0);
and (s1n276,n25,n277);
xor (n278,n279,n280);
not (n279,n277);
and (n280,n268,n269);
and (n281,n75,n282);
not (n282,n275);
nand (n283,n284,n320);
or (n284,n285,n317);
nor (n285,n286,n315);
and (n286,n287,n311);
wire s0n287,s1n287,notn287;
or (n287,s0n287,s1n287);
not(notn287,n133);
and (s0n287,notn287,n288);
and (s1n287,n133,n290);
wire s0n288,s1n288,notn288;
or (n288,s0n288,s1n288);
not(notn288,n25);
and (s0n288,notn288,1'b0);
and (s1n288,n25,n289);
xor (n290,n291,n292);
not (n291,n289);
and (n292,n293,n295);
not (n293,n294);
and (n295,n296,n298);
not (n296,n297);
and (n298,n299,n301);
not (n299,n300);
and (n301,n302,n304);
not (n302,n303);
and (n304,n305,n307);
not (n305,n306);
and (n307,n308,n310);
not (n308,n309);
and (n310,n279,n280);
not (n311,n312);
wire s0n312,s1n312,notn312;
or (n312,s0n312,s1n312);
not(notn312,n72);
and (s0n312,notn312,n313);
and (s1n312,n72,n314);
wire s0n313,s1n313,notn313;
or (n313,s0n313,s1n313);
not(notn313,n25);
and (s0n313,notn313,1'b0);
and (s1n313,n25,n69);
xor (n314,n68,n70);
and (n315,n316,n312);
not (n316,n287);
nand (n317,n312,n318);
not (n318,n319);
wire s0n319,s1n319,notn319;
or (n319,s0n319,s1n319);
not(notn319,n25);
and (s0n319,notn319,1'b0);
and (s1n319,n25,n71);
or (n320,n321,n318);
nor (n321,n322,n329);
and (n322,n323,n311);
wire s0n323,s1n323,notn323;
or (n323,s0n323,s1n323);
not(notn323,n133);
and (s0n323,notn323,n324);
and (s1n323,n133,n326);
wire s0n324,s1n324,notn324;
or (n324,s0n324,s1n324);
not(notn324,n25);
and (s0n324,notn324,1'b0);
and (s1n324,n25,n325);
xor (n326,n327,n328);
not (n327,n325);
and (n328,n291,n292);
and (n329,n330,n312);
not (n330,n323);
nand (n331,n332,n360);
or (n332,n333,n353);
nand (n333,n334,n345);
not (n334,n335);
nand (n335,n336,n344);
or (n336,n337,n341);
not (n337,n338);
wire s0n338,s1n338,notn338;
or (n338,s0n338,s1n338);
not(notn338,n72);
and (s0n338,notn338,n339);
and (s1n338,n72,n340);
wire s0n339,s1n339,notn339;
or (n339,s0n339,s1n339);
not(notn339,n25);
and (s0n339,notn339,1'b0);
and (s1n339,n25,n63);
xor (n340,n62,n64);
wire s0n341,s1n341,notn341;
or (n341,s0n341,s1n341);
not(notn341,n72);
and (s0n341,notn341,n342);
and (s1n341,n72,n343);
wire s0n342,s1n342,notn342;
or (n342,s0n342,s1n342);
not(notn342,n25);
and (s0n342,notn342,1'b0);
and (s1n342,n25,n60);
xor (n343,n59,n61);
nand (n344,n341,n337);
nor (n345,n346,n352);
and (n346,n347,n351);
not (n347,n348);
wire s0n348,s1n348,notn348;
or (n348,s0n348,s1n348);
not(notn348,n72);
and (s0n348,notn348,n349);
and (s1n348,n72,n350);
wire s0n349,s1n349,notn349;
or (n349,s0n349,s1n349);
not(notn349,n25);
and (s0n349,notn349,1'b0);
and (s1n349,n25,n57);
xor (n350,n56,n58);
not (n351,n341);
and (n352,n348,n341);
nor (n353,n354,n358);
and (n354,n355,n347);
wire s0n355,s1n355,notn355;
or (n355,s0n355,s1n355);
not(notn355,n133);
and (s0n355,notn355,n356);
and (s1n355,n133,n357);
wire s0n356,s1n356,notn356;
or (n356,s0n356,s1n356);
not(notn356,n25);
and (s0n356,notn356,1'b0);
and (s1n356,n25,n303);
xor (n357,n302,n304);
and (n358,n359,n348);
not (n359,n355);
or (n360,n361,n334);
nor (n361,n362,n366);
and (n362,n363,n347);
wire s0n363,s1n363,notn363;
or (n363,s0n363,s1n363);
not(notn363,n133);
and (s0n363,notn363,n364);
and (s1n363,n133,n365);
wire s0n364,s1n364,notn364;
or (n364,s0n364,s1n364);
not(notn364,n25);
and (s0n364,notn364,1'b0);
and (s1n364,n25,n300);
xor (n365,n299,n301);
and (n366,n367,n348);
not (n367,n363);
or (n368,n369,n429);
and (n369,n370,n391);
xor (n370,n371,n381);
nand (n371,n372,n380);
or (n372,n150,n373);
nor (n373,n374,n378);
and (n374,n153,n375);
wire s0n375,s1n375,notn375;
or (n375,s0n375,s1n375);
not(notn375,n133);
and (s0n375,notn375,n376);
and (s1n375,n133,n377);
wire s0n376,s1n376,notn376;
or (n376,s0n376,s1n376);
not(notn376,n25);
and (s0n376,notn376,1'b0);
and (s1n376,n25,n106);
xor (n377,n105,n107);
and (n378,n154,n379);
not (n379,n375);
or (n380,n179,n171);
nand (n381,n382,n390);
or (n382,n189,n383);
nor (n383,n384,n388);
and (n384,n385,n218);
wire s0n385,s1n385,notn385;
or (n385,s0n385,s1n385);
not(notn385,n133);
and (s0n385,notn385,n386);
and (s1n385,n133,n387);
wire s0n386,s1n386,notn386;
or (n386,s0n386,s1n386);
not(notn386,n25);
and (s0n386,notn386,1'b0);
and (s1n386,n25,n124);
xor (n387,n123,n125);
and (n388,n389,n219);
not (n389,n385);
or (n390,n234,n226);
nand (n391,n392,n421);
or (n392,n393,n414);
nand (n393,n394,n404);
nor (n394,n395,n402);
and (n395,n218,n396);
wire s0n396,s1n396,notn396;
or (n396,s0n396,s1n396);
not(notn396,n72);
and (s0n396,notn396,n397);
and (s1n396,n72,n399);
wire s0n397,s1n397,notn397;
or (n397,s0n397,s1n397);
not(notn397,n25);
and (s0n397,notn397,1'b0);
and (s1n397,n25,n398);
xor (n399,n400,n401);
not (n400,n398);
and (n401,n223,n224);
and (n402,n219,n403);
not (n403,n396);
nand (n404,n405,n412);
or (n405,n403,n406);
wire s0n406,s1n406,notn406;
or (n406,s0n406,s1n406);
not(notn406,n72);
and (s0n406,notn406,n407);
and (s1n406,n72,n409);
wire s0n407,s1n407,notn407;
or (n407,s0n407,s1n407);
not(notn407,n25);
and (s0n407,notn407,1'b0);
and (s1n407,n25,n408);
xor (n409,n410,n411);
not (n410,n408);
and (n411,n400,n401);
or (n412,n396,n413);
not (n413,n406);
nor (n414,n415,n419);
and (n415,n416,n413);
wire s0n416,s1n416,notn416;
or (n416,s0n416,s1n416);
not(notn416,n133);
and (s0n416,notn416,n417);
and (s1n416,n133,n418);
wire s0n417,s1n417,notn417;
or (n417,s0n417,s1n417);
not(notn417,n25);
and (s0n417,notn417,1'b0);
and (s1n417,n25,n130);
xor (n418,n129,n131);
and (n419,n420,n406);
not (n420,n416);
or (n421,n394,n422);
nor (n422,n423,n427);
and (n423,n424,n413);
wire s0n424,s1n424,notn424;
or (n424,s0n424,s1n424);
not(notn424,n133);
and (s0n424,notn424,n425);
and (s1n424,n133,n426);
wire s0n425,s1n425,notn425;
or (n425,s0n425,s1n425);
not(notn425,n25);
and (s0n425,notn425,1'b0);
and (s1n425,n25,n127);
xor (n426,n126,n128);
and (n427,n428,n406);
not (n428,n424);
and (n429,n371,n381);
and (n430,n14,n242);
xor (n431,n432,n573);
xor (n432,n433,n506);
xor (n433,n434,n482);
xor (n434,n435,n458);
nor (n435,n436,n456);
and (n436,n437,n454);
nand (n437,n438,n451);
not (n438,n439);
wire s0n439,s1n439,notn439;
or (n439,s0n439,s1n439);
not(notn439,n72);
and (s0n439,notn439,n440);
and (s1n439,n72,n442);
wire s0n440,s1n440,notn440;
or (n440,s0n440,s1n440);
not(notn440,n25);
and (s0n440,notn440,1'b0);
and (s1n440,n25,n441);
xor (n442,n443,n444);
not (n443,n441);
and (n444,n445,n447);
not (n445,n446);
and (n447,n448,n450);
not (n448,n449);
and (n450,n410,n411);
wire s0n451,s1n451,notn451;
or (n451,s0n451,s1n451);
not(notn451,n72);
and (s0n451,notn451,n452);
and (s1n451,n72,n453);
wire s0n452,s1n452,notn452;
or (n452,s0n452,s1n452);
not(notn452,n25);
and (s0n452,notn452,1'b0);
and (s1n452,n25,n446);
xor (n453,n445,n447);
nand (n454,n439,n455);
not (n455,n451);
not (n456,n457);
wire s0n457,s1n457,notn457;
or (n457,s0n457,s1n457);
not(notn457,n25);
and (s0n457,notn457,1'b0);
and (s1n457,n25,n132);
nand (n458,n459,n478);
or (n459,n460,n471);
nand (n460,n461,n468);
nor (n461,n462,n466);
and (n462,n311,n463);
wire s0n463,s1n463,notn463;
or (n463,s0n463,s1n463);
not(notn463,n72);
and (s0n463,notn463,n464);
and (s1n463,n72,n465);
wire s0n464,s1n464,notn464;
or (n464,s0n464,s1n464);
not(notn464,n25);
and (s0n464,notn464,1'b0);
and (s1n464,n25,n66);
xor (n465,n65,n67);
and (n466,n312,n467);
not (n467,n463);
nand (n468,n469,n470);
or (n469,n337,n463);
nand (n470,n337,n463);
nor (n471,n472,n476);
and (n472,n473,n337);
wire s0n473,s1n473,notn473;
or (n473,s0n473,s1n473);
not(notn473,n133);
and (s0n473,notn473,n474);
and (s1n473,n133,n475);
wire s0n474,s1n474,notn474;
or (n474,s0n474,s1n474);
not(notn474,n25);
and (s0n474,notn474,1'b0);
and (s1n474,n25,n294);
xor (n475,n293,n295);
and (n476,n477,n338);
not (n477,n473);
or (n478,n461,n479);
nor (n479,n480,n481);
and (n480,n287,n337);
and (n481,n316,n338);
nand (n482,n483,n502);
or (n483,n484,n495);
nand (n484,n485,n492);
or (n485,n486,n490);
and (n486,n348,n487);
wire s0n487,s1n487,notn487;
or (n487,s0n487,s1n487);
not(notn487,n72);
and (s0n487,notn487,n488);
and (s1n487,n72,n489);
wire s0n488,s1n488,notn488;
or (n488,s0n488,s1n488);
not(notn488,n25);
and (s0n488,notn488,1'b0);
and (s1n488,n25,n54);
xor (n489,n53,n55);
and (n490,n347,n491);
not (n491,n487);
nor (n492,n493,n494);
and (n493,n257,n487);
and (n494,n261,n491);
nor (n495,n496,n500);
and (n496,n497,n261);
wire s0n497,s1n497,notn497;
or (n497,s0n497,s1n497);
not(notn497,n133);
and (s0n497,notn497,n498);
and (s1n497,n133,n499);
wire s0n498,s1n498,notn498;
or (n498,s0n498,s1n498);
not(notn498,n25);
and (s0n498,notn498,1'b0);
and (s1n498,n25,n306);
xor (n499,n305,n307);
and (n500,n501,n257);
not (n501,n497);
or (n502,n503,n485);
nor (n503,n504,n505);
and (n504,n355,n261);
and (n505,n359,n257);
xor (n506,n507,n563);
xor (n507,n508,n534);
nand (n508,n509,n529);
or (n509,n510,n526);
not (n510,n511);
nor (n511,n512,n518);
nand (n512,n513,n517);
or (n513,n153,n514);
wire s0n514,s1n514,notn514;
or (n514,s0n514,s1n514);
not(notn514,n72);
and (s0n514,notn514,n515);
and (s1n514,n72,n516);
wire s0n515,s1n515,notn515;
or (n515,s0n515,s1n515);
not(notn515,n25);
and (s0n515,notn515,1'b0);
and (s1n515,n25,n208);
xor (n516,n207,n209);
nand (n517,n153,n514);
nor (n518,n519,n524);
and (n519,n520,n514);
not (n520,n521);
wire s0n521,s1n521,notn521;
or (n521,s0n521,s1n521);
not(notn521,n72);
and (s0n521,notn521,n522);
and (s1n521,n72,n523);
wire s0n522,s1n522,notn522;
or (n522,s0n522,s1n522);
not(notn522,n25);
and (s0n522,notn522,1'b0);
and (s1n522,n25,n205);
xor (n523,n204,n206);
and (n524,n525,n521);
not (n525,n514);
nor (n526,n527,n528);
and (n527,n520,n375);
and (n528,n521,n379);
or (n529,n530,n531);
not (n530,n512);
nor (n531,n532,n533);
and (n532,n520,n173);
and (n533,n521,n177);
nand (n534,n535,n555);
or (n535,n536,n548);
not (n536,n537);
and (n537,n538,n545);
nor (n538,n539,n544);
and (n539,n521,n540);
not (n540,n541);
wire s0n541,s1n541,notn541;
or (n541,s0n541,s1n541);
not(notn541,n72);
and (s0n541,notn541,n542);
and (s1n541,n72,n543);
wire s0n542,s1n542,notn542;
or (n542,s0n542,s1n542);
not(notn542,n25);
and (s0n542,notn542,1'b0);
and (s1n542,n25,n202);
xor (n543,n201,n203);
and (n544,n520,n541);
nand (n545,n546,n547);
or (n546,n540,n210);
or (n547,n215,n541);
nor (n548,n549,n553);
and (n549,n215,n550);
wire s0n550,s1n550,notn550;
or (n550,s0n550,s1n550);
not(notn550,n133);
and (s0n550,notn550,n551);
and (s1n550,n133,n552);
wire s0n551,s1n551,notn551;
or (n551,s0n551,s1n551);
not(notn551,n25);
and (s0n551,notn551,1'b0);
and (s1n551,n25,n112);
xor (n552,n111,n113);
and (n553,n210,n554);
not (n554,n550);
or (n555,n556,n538);
nor (n556,n557,n561);
and (n557,n215,n558);
wire s0n558,s1n558,notn558;
or (n558,s0n558,s1n558);
not(notn558,n133);
and (s0n558,notn558,n559);
and (s1n558,n133,n560);
wire s0n559,s1n559,notn559;
or (n559,s0n559,s1n559);
not(notn559,n25);
and (s0n559,notn559,1'b0);
and (s1n559,n25,n109);
xor (n560,n108,n110);
and (n561,n210,n562);
not (n562,n558);
nand (n563,n564,n565);
or (n564,n246,n273);
or (n565,n566,n254);
nor (n566,n567,n571);
and (n567,n80,n568);
wire s0n568,s1n568,notn568;
or (n568,s0n568,s1n568);
not(notn568,n133);
and (s0n568,notn568,n569);
and (s1n568,n133,n570);
wire s0n569,s1n569,notn569;
or (n569,s0n569,s1n569);
not(notn569,n25);
and (s0n569,notn569,1'b0);
and (s1n569,n25,n309);
xor (n570,n308,n310);
and (n571,n75,n572);
not (n572,n568);
xor (n573,n574,n591);
xor (n574,n575,n581);
nand (n575,n576,n577);
or (n576,n150,n180);
or (n577,n179,n578);
nor (n578,n579,n580);
and (n579,n153,n93);
and (n580,n154,n136);
nand (n581,n582,n583);
or (n582,n189,n235);
or (n583,n234,n584);
nor (n584,n585,n589);
and (n585,n218,n586);
wire s0n586,s1n586,notn586;
or (n586,s0n586,s1n586);
not(notn586,n133);
and (s0n586,notn586,n587);
and (s1n586,n133,n588);
wire s0n587,s1n587,notn587;
or (n587,s0n587,s1n587);
not(notn587,n25);
and (s0n587,notn587,1'b0);
and (s1n587,n25,n115);
xor (n588,n114,n116);
and (n589,n219,n590);
not (n590,n586);
nand (n591,n592,n596);
or (n592,n393,n593);
nor (n593,n594,n595);
and (n594,n385,n413);
and (n595,n389,n406);
or (n596,n394,n597);
nor (n597,n598,n599);
and (n598,n413,n228);
and (n599,n406,n232);
xor (n600,n601,n627);
xor (n601,n602,n624);
or (n602,n603,n623);
and (n603,n604,n617);
xor (n604,n605,n611);
nand (n605,n606,n610);
or (n606,n484,n607);
nor (n607,n608,n609);
and (n608,n568,n261);
and (n609,n572,n257);
or (n610,n495,n485);
nand (n611,n612,n616);
or (n612,n510,n613);
nor (n613,n614,n615);
and (n614,n520,n558);
and (n615,n521,n562);
or (n616,n530,n526);
nand (n617,n618,n622);
or (n618,n536,n619);
nor (n619,n620,n621);
and (n620,n215,n586);
and (n621,n210,n590);
or (n622,n548,n538);
and (n623,n605,n611);
or (n624,n625,n626);
and (n625,n15,n187);
and (n626,n16,n148);
xor (n627,n628,n652);
xor (n628,n629,n642);
nand (n629,n630,n631);
or (n630,n321,n317);
or (n631,n632,n318);
nor (n632,n633,n640);
and (n633,n634,n311);
wire s0n634,s1n634,notn634;
or (n634,s0n634,s1n634);
not(notn634,n133);
and (s0n634,notn634,n635);
and (s1n634,n133,n637);
wire s0n635,s1n635,notn635;
or (n635,s0n635,s1n635);
not(notn635,n25);
and (s0n635,notn635,1'b0);
and (s1n635,n25,n636);
xor (n637,n638,n639);
not (n638,n636);
and (n639,n327,n328);
and (n640,n641,n312);
not (n641,n634);
nand (n642,n643,n644);
or (n643,n333,n361);
or (n644,n334,n645);
nor (n645,n646,n650);
and (n646,n647,n347);
wire s0n647,s1n647,notn647;
or (n647,s0n647,s1n647);
not(notn647,n133);
and (s0n647,notn647,n648);
and (s1n647,n133,n649);
wire s0n648,s1n648,notn648;
or (n648,s0n648,s1n648);
not(notn648,n25);
and (s0n648,notn648,1'b0);
and (s1n648,n25,n297);
xor (n649,n296,n298);
and (n650,n651,n348);
not (n651,n647);
nand (n652,n653,n654);
or (n653,n18,n138);
or (n654,n19,n655);
nor (n655,n656,n657);
and (n656,n90,n264);
and (n657,n83,n271);
xor (n658,n659,n847);
xor (n659,n660,n786);
or (n660,n661,n785);
and (n661,n662,n703);
xor (n662,n663,n664);
xor (n663,n604,n617);
xor (n664,n665,n690);
xor (n665,n666,n669);
nand (n666,n667,n668);
or (n667,n393,n422);
or (n668,n394,n593);
nand (n669,n670,n686);
or (n670,n671,n683);
or (n671,n672,n680);
not (n672,n673);
and (n673,n674,n679);
nand (n674,n675,n406);
not (n675,n676);
wire s0n676,s1n676,notn676;
or (n676,s0n676,s1n676);
not(notn676,n72);
and (s0n676,notn676,n677);
and (s1n676,n72,n678);
wire s0n677,s1n677,notn677;
or (n677,s0n677,s1n677);
not(notn677,n25);
and (s0n677,notn677,1'b0);
and (s1n677,n25,n449);
xor (n678,n448,n450);
nand (n679,n676,n413);
nor (n680,n681,n682);
and (n681,n676,n455);
and (n682,n675,n451);
nor (n683,n684,n685);
and (n684,n451,n456);
and (n685,n455,n457);
or (n686,n673,n687);
nor (n687,n688,n689);
and (n688,n416,n455);
and (n689,n420,n451);
xor (n690,n691,n697);
nor (n691,n692,n455);
nor (n692,n693,n696);
and (n693,n694,n413);
not (n694,n695);
and (n695,n457,n676);
and (n696,n675,n456);
nand (n697,n698,n702);
or (n698,n460,n699);
nor (n699,n700,n701);
and (n700,n647,n337);
and (n701,n651,n338);
or (n702,n471,n461);
or (n703,n704,n784);
and (n704,n705,n753);
xor (n705,n706,n722);
and (n706,n707,n713);
nor (n707,n708,n413);
nor (n708,n709,n712);
and (n709,n710,n218);
not (n710,n711);
and (n711,n457,n396);
and (n712,n403,n456);
nand (n713,n714,n718);
or (n714,n460,n715);
nor (n715,n716,n717);
and (n716,n355,n337);
and (n717,n359,n338);
or (n718,n461,n719);
nor (n719,n720,n721);
and (n720,n363,n337);
and (n721,n367,n338);
or (n722,n723,n752);
and (n723,n724,n743);
xor (n724,n725,n734);
nand (n725,n726,n730);
or (n726,n246,n727);
nor (n727,n728,n729);
and (n728,n80,n93);
and (n729,n75,n136);
or (n730,n731,n254);
nor (n731,n732,n733);
and (n732,n80,n140);
and (n733,n75,n147);
nand (n734,n735,n739);
or (n735,n736,n317);
nor (n736,n737,n738);
and (n737,n647,n311);
and (n738,n651,n312);
or (n739,n740,n318);
nor (n740,n741,n742);
and (n741,n473,n311);
and (n742,n477,n312);
nand (n743,n744,n748);
or (n744,n333,n745);
nor (n745,n746,n747);
and (n746,n568,n347);
and (n747,n572,n348);
or (n748,n749,n334);
nor (n749,n750,n751);
and (n750,n497,n347);
and (n751,n501,n348);
and (n752,n725,n734);
or (n753,n754,n783);
and (n754,n755,n774);
xor (n755,n756,n765);
nand (n756,n757,n761);
or (n757,n484,n758);
nor (n758,n759,n760);
and (n759,n264,n261);
and (n760,n271,n257);
or (n761,n485,n762);
nor (n762,n763,n764);
and (n763,n275,n261);
and (n764,n282,n257);
nand (n765,n766,n770);
or (n766,n510,n767);
nor (n767,n768,n769);
and (n768,n520,n586);
and (n769,n521,n590);
or (n770,n771,n530);
nor (n771,n772,n773);
and (n772,n520,n550);
and (n773,n521,n554);
nand (n774,n775,n779);
or (n775,n536,n776);
nor (n776,n777,n778);
and (n777,n215,n228);
and (n778,n210,n232);
or (n779,n780,n538);
nor (n780,n781,n782);
and (n781,n215,n237);
and (n782,n210,n241);
and (n783,n756,n765);
and (n784,n706,n722);
and (n785,n663,n664);
xor (n786,n787,n803);
xor (n787,n788,n791);
or (n788,n789,n790);
and (n789,n665,n690);
and (n790,n666,n669);
xor (n791,n792,n800);
xor (n792,n793,n799);
nand (n793,n794,n795);
or (n794,n671,n687);
or (n795,n673,n796);
nor (n796,n797,n798);
and (n797,n424,n455);
and (n798,n428,n451);
and (n799,n691,n697);
or (n800,n801,n802);
and (n801,n243,n331);
and (n802,n244,n283);
or (n803,n804,n846);
and (n804,n805,n833);
xor (n805,n806,n822);
or (n806,n807,n821);
and (n807,n808,n815);
xor (n808,n809,n812);
nand (n809,n810,n811);
or (n810,n740,n317);
or (n811,n285,n318);
nand (n812,n813,n814);
or (n813,n333,n749);
or (n814,n353,n334);
nand (n815,n816,n820);
or (n816,n18,n817);
nor (n817,n818,n819);
and (n818,n90,n182);
and (n819,n83,n186);
or (n820,n19,n91);
and (n821,n809,n812);
or (n822,n823,n832);
and (n823,n824,n829);
xor (n824,n825,n826);
nor (n825,n673,n456);
nand (n826,n827,n828);
or (n827,n460,n719);
or (n828,n461,n699);
nand (n829,n830,n831);
or (n830,n484,n762);
or (n831,n485,n607);
and (n832,n825,n826);
or (n833,n834,n845);
and (n834,n835,n842);
xor (n835,n836,n839);
nand (n836,n837,n838);
or (n837,n510,n771);
or (n838,n530,n613);
nand (n839,n840,n841);
or (n840,n536,n780);
or (n841,n619,n538);
nand (n842,n843,n844);
or (n843,n246,n731);
or (n844,n262,n254);
and (n845,n836,n839);
and (n846,n806,n822);
or (n847,n848,n880);
and (n848,n849,n879);
xor (n849,n850,n878);
or (n850,n851,n877);
and (n851,n852,n876);
xor (n852,n853,n875);
or (n853,n854,n874);
and (n854,n855,n868);
xor (n855,n856,n862);
nand (n856,n857,n861);
or (n857,n18,n858);
nor (n858,n859,n860);
and (n859,n90,n173);
and (n860,n83,n177);
or (n861,n19,n817);
nand (n862,n863,n867);
or (n863,n150,n864);
nor (n864,n865,n866);
and (n865,n153,n558);
and (n866,n154,n562);
or (n867,n179,n373);
nand (n868,n869,n873);
or (n869,n189,n870);
nor (n870,n871,n872);
and (n871,n424,n218);
and (n872,n428,n219);
or (n873,n234,n383);
and (n874,n856,n862);
xor (n875,n808,n815);
xor (n876,n835,n842);
and (n877,n853,n875);
xor (n878,n805,n833);
xor (n879,n13,n368);
and (n880,n850,n878);
or (n881,n882,n1008);
and (n882,n883,n924);
xor (n883,n884,n885);
xor (n884,n662,n703);
or (n885,n886,n923);
and (n886,n887,n890);
xor (n887,n888,n889);
xor (n888,n824,n829);
xor (n889,n370,n391);
or (n890,n891,n922);
and (n891,n892,n900);
xor (n892,n893,n899);
nand (n893,n894,n898);
or (n894,n393,n895);
nor (n895,n896,n897);
and (n896,n406,n456);
and (n897,n413,n457);
or (n898,n394,n414);
xor (n899,n707,n713);
or (n900,n901,n921);
and (n901,n902,n915);
xor (n902,n903,n909);
nand (n903,n904,n908);
or (n904,n246,n905);
nor (n905,n906,n907);
and (n906,n80,n182);
and (n907,n75,n186);
or (n908,n727,n254);
nand (n909,n910,n914);
or (n910,n333,n911);
nor (n911,n912,n913);
and (n912,n275,n347);
and (n913,n282,n348);
or (n914,n334,n745);
nand (n915,n916,n920);
or (n916,n18,n917);
nor (n917,n918,n919);
and (n918,n90,n375);
and (n919,n83,n379);
or (n920,n19,n858);
and (n921,n903,n909);
and (n922,n893,n899);
and (n923,n888,n889);
or (n924,n925,n1007);
and (n925,n926,n972);
xor (n926,n927,n928);
xor (n927,n705,n753);
or (n928,n929,n971);
and (n929,n930,n970);
xor (n930,n931,n948);
or (n931,n932,n947);
and (n932,n933,n941);
xor (n933,n934,n935);
nor (n934,n394,n456);
nand (n935,n936,n940);
or (n936,n937,n317);
nor (n937,n938,n939);
and (n938,n363,n311);
and (n939,n367,n312);
or (n940,n736,n318);
nand (n941,n942,n946);
or (n942,n484,n943);
nor (n943,n944,n945);
and (n944,n140,n261);
and (n945,n147,n257);
or (n946,n485,n758);
and (n947,n934,n935);
or (n948,n949,n969);
and (n949,n950,n963);
xor (n950,n951,n957);
nand (n951,n952,n956);
or (n952,n510,n953);
nor (n953,n954,n955);
and (n954,n237,n520);
and (n955,n241,n521);
or (n956,n767,n530);
nand (n957,n958,n962);
or (n958,n536,n959);
nor (n959,n960,n961);
and (n960,n385,n215);
and (n961,n389,n210);
or (n962,n776,n538);
nand (n963,n964,n968);
or (n964,n460,n965);
nor (n965,n966,n967);
and (n966,n497,n337);
and (n967,n501,n338);
or (n968,n461,n715);
and (n969,n951,n957);
xor (n970,n724,n743);
and (n971,n931,n948);
or (n972,n973,n1006);
and (n973,n974,n977);
xor (n974,n975,n976);
xor (n975,n755,n774);
xor (n976,n855,n868);
or (n977,n978,n1005);
and (n978,n979,n992);
xor (n979,n980,n986);
nand (n980,n981,n985);
or (n981,n150,n982);
nor (n982,n983,n984);
and (n983,n153,n550);
and (n984,n154,n554);
or (n985,n179,n864);
nand (n986,n987,n991);
or (n987,n189,n988);
nor (n988,n989,n990);
and (n989,n416,n218);
and (n990,n420,n219);
or (n991,n234,n870);
and (n992,n993,n999);
nor (n993,n994,n218);
nor (n994,n995,n998);
and (n995,n996,n215);
not (n996,n997);
and (n997,n457,n192);
and (n998,n214,n456);
nand (n999,n1000,n1004);
or (n1000,n1001,n317);
nor (n1001,n1002,n1003);
and (n1002,n355,n311);
and (n1003,n359,n312);
or (n1004,n937,n318);
and (n1005,n980,n986);
and (n1006,n975,n976);
and (n1007,n927,n928);
and (n1008,n884,n885);
and (n1009,n9,n658);
not (n1010,n1011);
xor (n1011,n1012,n1134);
xor (n1012,n1013,n1131);
xor (n1013,n1014,n1096);
xor (n1014,n1015,n1018);
or (n1015,n1016,n1017);
and (n1016,n432,n573);
and (n1017,n433,n506);
xor (n1018,n1019,n1060);
xor (n1019,n1020,n1040);
xor (n1020,n1021,n1034);
xor (n1021,n1022,n1028);
nand (n1022,n1023,n1024);
or (n1023,n484,n503);
or (n1024,n1025,n485);
nor (n1025,n1026,n1027);
and (n1026,n363,n261);
and (n1027,n367,n257);
nand (n1028,n1029,n1030);
or (n1029,n510,n531);
or (n1030,n530,n1031);
nor (n1031,n1032,n1033);
and (n1032,n520,n182);
and (n1033,n521,n186);
nand (n1034,n1035,n1036);
or (n1035,n536,n556);
or (n1036,n1037,n538);
nor (n1037,n1038,n1039);
and (n1038,n215,n375);
and (n1039,n210,n379);
xor (n1040,n1041,n1054);
xor (n1041,n1042,n1048);
nand (n1042,n1043,n1044);
or (n1043,n333,n645);
or (n1044,n1045,n334);
nor (n1045,n1046,n1047);
and (n1046,n473,n347);
and (n1047,n477,n348);
nand (n1048,n1049,n1050);
or (n1049,n150,n578);
or (n1050,n179,n1051);
nor (n1051,n1052,n1053);
and (n1052,n153,n140);
and (n1053,n154,n147);
nand (n1054,n1055,n1056);
or (n1055,n189,n584);
or (n1056,n234,n1057);
nor (n1057,n1058,n1059);
and (n1058,n218,n550);
and (n1059,n219,n554);
xor (n1060,n1061,n1074);
xor (n1061,n1062,n1068);
nand (n1062,n1063,n1064);
or (n1063,n393,n597);
or (n1064,n394,n1065);
nor (n1065,n1066,n1067);
and (n1066,n413,n237);
and (n1067,n241,n406);
nand (n1068,n1069,n1070);
or (n1069,n671,n796);
or (n1070,n673,n1071);
nor (n1071,n1072,n1073);
and (n1072,n385,n455);
and (n1073,n389,n451);
nand (n1074,n1075,n1092);
or (n1075,n1076,n1089);
nand (n1076,n1077,n436);
or (n1077,n1078,n1087);
not (n1078,n1079);
nand (n1079,n439,n1080);
not (n1080,n1081);
wire s0n1081,s1n1081,notn1081;
or (n1081,s0n1081,s1n1081);
not(notn1081,n72);
and (s0n1081,notn1081,n1082);
and (s1n1081,n72,n1084);
wire s0n1082,s1n1082,notn1082;
or (n1082,s0n1082,s1n1082);
not(notn1082,n25);
and (s0n1082,notn1082,1'b0);
and (s1n1082,n25,n1083);
xor (n1084,n1085,n1086);
not (n1085,n1083);
and (n1086,n443,n444);
not (n1087,n1088);
nand (n1088,n438,n1081);
nor (n1089,n1090,n1091);
and (n1090,n1081,n456);
and (n1091,n1080,n457);
or (n1092,n436,n1093);
nor (n1093,n1094,n1095);
and (n1094,n416,n1080);
and (n1095,n420,n1081);
xor (n1096,n1097,n1104);
xor (n1097,n1098,n1101);
or (n1098,n1099,n1100);
and (n1099,n434,n482);
and (n1100,n435,n458);
or (n1101,n1102,n1103);
and (n1102,n574,n591);
and (n1103,n575,n581);
xor (n1104,n1105,n1125);
xor (n1105,n1106,n1112);
nand (n1106,n1107,n1108);
or (n1107,n246,n566);
or (n1108,n1109,n254);
nor (n1109,n1110,n1111);
and (n1110,n497,n80);
and (n1111,n501,n75);
nand (n1112,n1113,n1114);
or (n1113,n632,n317);
or (n1114,n1115,n318);
nor (n1115,n1116,n1123);
and (n1116,n1117,n311);
wire s0n1117,s1n1117,notn1117;
or (n1117,s0n1117,s1n1117);
not(notn1117,n133);
and (s0n1117,notn1117,n1118);
and (s1n1117,n133,n1120);
wire s0n1118,s1n1118,notn1118;
or (n1118,s0n1118,s1n1118);
not(notn1118,n25);
and (s0n1118,notn1118,1'b0);
and (s1n1118,n25,n1119);
xor (n1120,n1121,n1122);
not (n1121,n1119);
and (n1122,n638,n639);
and (n1123,n1124,n312);
not (n1124,n1117);
nand (n1125,n1126,n1127);
or (n1126,n18,n655);
or (n1127,n19,n1128);
nor (n1128,n1129,n1130);
and (n1129,n90,n275);
and (n1130,n83,n282);
or (n1131,n1132,n1133);
and (n1132,n659,n847);
and (n1133,n660,n786);
xor (n1134,n1135,n1168);
xor (n1135,n1136,n1139);
or (n1136,n1137,n1138);
and (n1137,n787,n803);
and (n1138,n788,n791);
xor (n1139,n1140,n1147);
xor (n1140,n1141,n1144);
or (n1141,n1142,n1143);
and (n1142,n792,n800);
and (n1143,n793,n799);
or (n1144,n1145,n1146);
and (n1145,n601,n627);
and (n1146,n602,n624);
xor (n1147,n1148,n1165);
xor (n1148,n1149,n1162);
xor (n1149,n1150,n1156);
nor (n1150,n1151,n1080);
nor (n1151,n1152,n1155);
and (n1152,n1153,n455);
not (n1153,n1154);
and (n1154,n457,n439);
and (n1155,n438,n456);
nand (n1156,n1157,n1158);
or (n1157,n460,n479);
or (n1158,n461,n1159);
nor (n1159,n1160,n1161);
and (n1160,n323,n337);
and (n1161,n330,n338);
or (n1162,n1163,n1164);
and (n1163,n507,n563);
and (n1164,n508,n534);
or (n1165,n1166,n1167);
and (n1166,n628,n652);
and (n1167,n629,n642);
or (n1168,n1169,n1170);
and (n1169,n10,n600);
and (n1170,n11,n431);
nor (n1171,n5,n1010);
not (n1172,n1173);
nand (n1173,n1174,n2386);
or (n1174,n1175,n2381);
nor (n1175,n1176,n2380);
and (n1176,n1177,n2367);
or (n1177,n1178,n2366);
and (n1178,n1179,n1416);
xor (n1179,n1180,n1403);
or (n1180,n1181,n1402);
and (n1181,n1182,n1317);
xor (n1182,n1183,n1236);
xor (n1183,n1184,n1235);
xor (n1184,n1185,n1186);
xor (n1185,n892,n900);
or (n1186,n1187,n1234);
and (n1187,n1188,n1233);
xor (n1188,n1189,n1211);
or (n1189,n1190,n1210);
and (n1190,n1191,n1204);
xor (n1191,n1192,n1198);
nand (n1192,n1193,n1197);
or (n1193,n484,n1194);
nor (n1194,n1195,n1196);
and (n1195,n93,n261);
and (n1196,n136,n257);
or (n1197,n485,n943);
nand (n1198,n1199,n1203);
or (n1199,n510,n1200);
nor (n1200,n1201,n1202);
and (n1201,n520,n228);
and (n1202,n232,n521);
or (n1203,n530,n953);
nand (n1204,n1205,n1209);
or (n1205,n536,n1206);
nor (n1206,n1207,n1208);
and (n1207,n424,n215);
and (n1208,n428,n210);
or (n1209,n959,n538);
and (n1210,n1192,n1198);
or (n1211,n1212,n1232);
and (n1212,n1213,n1226);
xor (n1213,n1214,n1220);
nand (n1214,n1215,n1219);
or (n1215,n460,n1216);
nor (n1216,n1217,n1218);
and (n1217,n337,n568);
and (n1218,n572,n338);
or (n1219,n965,n461);
nand (n1220,n1221,n1225);
or (n1221,n246,n1222);
nor (n1222,n1223,n1224);
and (n1223,n80,n173);
and (n1224,n75,n177);
or (n1225,n905,n254);
nand (n1226,n1227,n1231);
or (n1227,n333,n1228);
nor (n1228,n1229,n1230);
and (n1229,n264,n347);
and (n1230,n271,n348);
or (n1231,n334,n911);
and (n1232,n1214,n1220);
xor (n1233,n902,n915);
and (n1234,n1189,n1211);
xor (n1235,n930,n970);
xor (n1236,n1237,n1267);
xor (n1237,n1238,n1266);
or (n1238,n1239,n1265);
and (n1239,n1240,n1243);
xor (n1240,n1241,n1242);
xor (n1241,n933,n941);
xor (n1242,n950,n963);
or (n1243,n1244,n1264);
and (n1244,n1245,n1258);
xor (n1245,n1246,n1252);
nand (n1246,n1247,n1251);
or (n1247,n18,n1248);
nor (n1248,n1249,n1250);
and (n1249,n90,n558);
and (n1250,n83,n562);
or (n1251,n19,n917);
nand (n1252,n1253,n1257);
or (n1253,n150,n1254);
nor (n1254,n1255,n1256);
and (n1255,n153,n586);
and (n1256,n154,n590);
or (n1257,n982,n179);
nand (n1258,n1259,n1263);
or (n1259,n189,n1260);
nor (n1260,n1261,n1262);
and (n1261,n219,n456);
and (n1262,n218,n457);
or (n1263,n234,n988);
and (n1264,n1246,n1252);
and (n1265,n1241,n1242);
xor (n1266,n974,n977);
or (n1267,n1268,n1316);
and (n1268,n1269,n1315);
xor (n1269,n1270,n1271);
xor (n1270,n979,n992);
or (n1271,n1272,n1314);
and (n1272,n1273,n1292);
xor (n1273,n1274,n1275);
xor (n1274,n993,n999);
or (n1275,n1276,n1291);
and (n1276,n1277,n1285);
xor (n1277,n1278,n1279);
nor (n1278,n234,n456);
nand (n1279,n1280,n1284);
or (n1280,n1281,n317);
nor (n1281,n1282,n1283);
and (n1282,n497,n311);
and (n1283,n501,n312);
or (n1284,n1001,n318);
nand (n1285,n1286,n1287);
or (n1286,n1194,n485);
or (n1287,n484,n1288);
nor (n1288,n1289,n1290);
and (n1289,n182,n261);
and (n1290,n186,n257);
and (n1291,n1278,n1279);
or (n1292,n1293,n1313);
and (n1293,n1294,n1307);
xor (n1294,n1295,n1301);
nand (n1295,n1296,n1300);
or (n1296,n510,n1297);
nor (n1297,n1298,n1299);
and (n1298,n385,n520);
and (n1299,n389,n521);
or (n1300,n1200,n530);
nand (n1301,n1302,n1306);
or (n1302,n536,n1303);
nor (n1303,n1304,n1305);
and (n1304,n416,n215);
and (n1305,n420,n210);
or (n1306,n1206,n538);
nand (n1307,n1308,n1312);
or (n1308,n460,n1309);
nor (n1309,n1310,n1311);
and (n1310,n337,n275);
and (n1311,n282,n338);
or (n1312,n461,n1216);
and (n1313,n1295,n1301);
and (n1314,n1274,n1275);
xor (n1315,n1188,n1233);
and (n1316,n1270,n1271);
or (n1317,n1318,n1401);
and (n1318,n1319,n1349);
xor (n1319,n1320,n1348);
or (n1320,n1321,n1347);
and (n1321,n1322,n1346);
xor (n1322,n1323,n1345);
or (n1323,n1324,n1344);
and (n1324,n1325,n1338);
xor (n1325,n1326,n1332);
nand (n1326,n1327,n1331);
or (n1327,n246,n1328);
nor (n1328,n1329,n1330);
and (n1329,n80,n375);
and (n1330,n75,n379);
or (n1331,n1222,n254);
nand (n1332,n1333,n1337);
or (n1333,n333,n1334);
nor (n1334,n1335,n1336);
and (n1335,n140,n347);
and (n1336,n147,n348);
or (n1337,n334,n1228);
nand (n1338,n1339,n1343);
or (n1339,n18,n1340);
nor (n1340,n1341,n1342);
and (n1341,n90,n550);
and (n1342,n83,n554);
or (n1343,n19,n1248);
and (n1344,n1326,n1332);
xor (n1345,n1213,n1226);
xor (n1346,n1191,n1204);
and (n1347,n1323,n1345);
xor (n1348,n1240,n1243);
or (n1349,n1350,n1400);
and (n1350,n1351,n1399);
xor (n1351,n1352,n1353);
xor (n1352,n1245,n1258);
or (n1353,n1354,n1398);
and (n1354,n1355,n1375);
xor (n1355,n1356,n1362);
nand (n1356,n1357,n1361);
or (n1357,n150,n1358);
nor (n1358,n1359,n1360);
and (n1359,n153,n237);
and (n1360,n154,n241);
or (n1361,n1254,n179);
and (n1362,n1363,n1369);
nor (n1363,n1364,n215);
nor (n1364,n1365,n1368);
and (n1365,n520,n1366);
not (n1366,n1367);
and (n1367,n457,n541);
and (n1368,n540,n456);
nand (n1369,n1370,n1374);
or (n1370,n1371,n317);
nor (n1371,n1372,n1373);
and (n1372,n568,n311);
and (n1373,n572,n312);
or (n1374,n1281,n318);
or (n1375,n1376,n1397);
and (n1376,n1377,n1390);
xor (n1377,n1378,n1384);
nand (n1378,n1379,n1383);
or (n1379,n484,n1380);
nor (n1380,n1381,n1382);
and (n1381,n173,n261);
and (n1382,n177,n257);
or (n1383,n1288,n485);
nand (n1384,n1385,n1389);
or (n1385,n510,n1386);
nor (n1386,n1387,n1388);
and (n1387,n424,n520);
and (n1388,n428,n521);
or (n1389,n530,n1297);
nand (n1390,n1391,n1396);
or (n1391,n1392,n536);
not (n1392,n1393);
nand (n1393,n1394,n1395);
or (n1394,n215,n457);
or (n1395,n210,n456);
or (n1396,n1303,n538);
and (n1397,n1378,n1384);
and (n1398,n1356,n1362);
xor (n1399,n1273,n1292);
and (n1400,n1352,n1353);
and (n1401,n1320,n1348);
and (n1402,n1183,n1236);
xor (n1403,n1404,n1413);
xor (n1404,n1405,n1406);
xor (n1405,n926,n972);
xor (n1406,n1407,n1410);
xor (n1407,n1408,n1409);
xor (n1408,n852,n876);
xor (n1409,n887,n890);
or (n1410,n1411,n1412);
and (n1411,n1184,n1235);
and (n1412,n1185,n1186);
or (n1413,n1414,n1415);
and (n1414,n1237,n1267);
and (n1415,n1238,n1266);
nand (n1416,n1417,n2360);
or (n1417,n1418,n2353);
nand (n1418,n1419,n2342);
not (n1419,n1420);
nor (n1420,n1421,n2331);
nor (n1421,n1422,n2280);
nand (n1422,n1423,n2154);
or (n1423,n1424,n2153);
and (n1424,n1425,n1743);
xor (n1425,n1426,n1657);
or (n1426,n1427,n1656);
and (n1427,n1428,n1605);
xor (n1428,n1429,n1512);
xor (n1429,n1430,n1481);
xor (n1430,n1431,n1452);
xor (n1431,n1432,n1443);
xor (n1432,n1433,n1434);
nor (n1433,n530,n456);
nand (n1434,n1435,n1439);
or (n1435,n1436,n317);
nor (n1436,n1437,n1438);
and (n1437,n311,n140);
and (n1438,n147,n312);
or (n1439,n1440,n318);
nor (n1440,n1441,n1442);
and (n1441,n264,n311);
and (n1442,n271,n312);
nand (n1443,n1444,n1448);
or (n1444,n460,n1445);
nor (n1445,n1446,n1447);
and (n1446,n337,n182);
and (n1447,n186,n338);
or (n1448,n461,n1449);
nor (n1449,n1450,n1451);
and (n1450,n93,n337);
and (n1451,n136,n338);
or (n1452,n1453,n1480);
and (n1453,n1454,n1470);
xor (n1454,n1455,n1461);
nand (n1455,n1456,n1460);
or (n1456,n460,n1457);
nor (n1457,n1458,n1459);
and (n1458,n337,n173);
and (n1459,n177,n338);
or (n1460,n461,n1445);
nand (n1461,n1462,n1466);
or (n1462,n484,n1463);
nor (n1463,n1464,n1465);
and (n1464,n586,n261);
and (n1465,n590,n257);
or (n1466,n485,n1467);
nor (n1467,n1468,n1469);
and (n1468,n550,n261);
and (n1469,n554,n257);
nand (n1470,n1471,n1476);
or (n1471,n1472,n246);
not (n1472,n1473);
nand (n1473,n1474,n1475);
or (n1474,n75,n232);
or (n1475,n80,n228);
or (n1476,n1477,n254);
nor (n1477,n1478,n1479);
and (n1478,n80,n237);
and (n1479,n75,n241);
and (n1480,n1455,n1461);
or (n1481,n1482,n1511);
and (n1482,n1483,n1502);
xor (n1483,n1484,n1493);
nand (n1484,n1485,n1489);
or (n1485,n333,n1486);
nor (n1486,n1487,n1488);
and (n1487,n558,n347);
and (n1488,n562,n348);
or (n1489,n1490,n334);
nor (n1490,n1491,n1492);
and (n1491,n375,n347);
and (n1492,n379,n348);
nand (n1493,n1494,n1498);
or (n1494,n18,n1495);
nor (n1495,n1496,n1497);
and (n1496,n424,n90);
and (n1497,n428,n83);
or (n1498,n1499,n19);
nor (n1499,n1500,n1501);
and (n1500,n385,n90);
and (n1501,n389,n83);
nand (n1502,n1503,n1507);
or (n1503,n179,n1504);
nor (n1504,n1505,n1506);
and (n1505,n416,n153);
and (n1506,n420,n154);
or (n1507,n150,n1508);
nor (n1508,n1509,n1510);
and (n1509,n154,n456);
and (n1510,n153,n457);
and (n1511,n1484,n1493);
xor (n1512,n1513,n1561);
xor (n1513,n1514,n1541);
xor (n1514,n1515,n1528);
xor (n1515,n1516,n1522);
nand (n1516,n1517,n1518);
or (n1517,n18,n1499);
or (n1518,n1519,n19);
nor (n1519,n1520,n1521);
and (n1520,n90,n228);
and (n1521,n83,n232);
nand (n1522,n1523,n1524);
or (n1523,n150,n1504);
or (n1524,n1525,n179);
nor (n1525,n1526,n1527);
and (n1526,n424,n153);
and (n1527,n428,n154);
and (n1528,n1529,n1535);
nand (n1529,n1530,n1534);
or (n1530,n1531,n317);
nor (n1531,n1532,n1533);
and (n1532,n311,n93);
and (n1533,n136,n312);
or (n1534,n1436,n318);
nor (n1535,n1536,n153);
nor (n1536,n1537,n1540);
and (n1537,n90,n1538);
not (n1538,n1539);
and (n1539,n457,n163);
and (n1540,n167,n456);
xor (n1541,n1542,n1555);
xor (n1542,n1543,n1549);
nand (n1543,n1544,n1545);
or (n1544,n484,n1467);
or (n1545,n1546,n485);
nor (n1546,n1547,n1548);
and (n1547,n558,n261);
and (n1548,n562,n257);
nand (n1549,n1550,n1551);
or (n1550,n246,n1477);
or (n1551,n1552,n254);
nor (n1552,n1553,n1554);
and (n1553,n80,n586);
and (n1554,n75,n590);
nand (n1555,n1556,n1560);
or (n1556,n334,n1557);
nor (n1557,n1558,n1559);
and (n1558,n173,n347);
and (n1559,n177,n348);
or (n1560,n333,n1490);
or (n1561,n1562,n1604);
and (n1562,n1563,n1582);
xor (n1563,n1564,n1565);
xor (n1564,n1529,n1535);
or (n1565,n1566,n1581);
and (n1566,n1567,n1575);
xor (n1567,n1568,n1569);
nor (n1568,n179,n456);
nand (n1569,n1570,n1574);
or (n1570,n1571,n317);
nor (n1571,n1572,n1573);
and (n1572,n311,n182);
and (n1573,n186,n312);
or (n1574,n1531,n318);
nand (n1575,n1576,n1577);
or (n1576,n461,n1457);
or (n1577,n460,n1578);
nor (n1578,n1579,n1580);
and (n1579,n375,n337);
and (n1580,n379,n338);
and (n1581,n1568,n1569);
or (n1582,n1583,n1603);
and (n1583,n1584,n1597);
xor (n1584,n1585,n1591);
nand (n1585,n1586,n1590);
or (n1586,n484,n1587);
nor (n1587,n1588,n1589);
and (n1588,n237,n261);
and (n1589,n241,n257);
or (n1590,n1463,n485);
nand (n1591,n1592,n1593);
or (n1592,n254,n1472);
or (n1593,n246,n1594);
nor (n1594,n1595,n1596);
and (n1595,n80,n385);
and (n1596,n75,n389);
nand (n1597,n1598,n1599);
or (n1598,n19,n1495);
or (n1599,n18,n1600);
nor (n1600,n1601,n1602);
and (n1601,n416,n90);
and (n1602,n420,n83);
and (n1603,n1585,n1591);
and (n1604,n1564,n1565);
or (n1605,n1606,n1655);
and (n1606,n1607,n1610);
xor (n1607,n1608,n1609);
xor (n1608,n1483,n1502);
xor (n1609,n1454,n1470);
or (n1610,n1611,n1654);
and (n1611,n1612,n1632);
xor (n1612,n1613,n1619);
nand (n1613,n1614,n1618);
or (n1614,n333,n1615);
nor (n1615,n1616,n1617);
and (n1616,n550,n347);
and (n1617,n554,n348);
or (n1618,n334,n1486);
and (n1619,n1620,n1626);
nand (n1620,n1621,n1625);
or (n1621,n1622,n317);
nor (n1622,n1623,n1624);
and (n1623,n173,n311);
and (n1624,n177,n312);
or (n1625,n1571,n318);
nor (n1626,n1627,n90);
nor (n1627,n1628,n1631);
and (n1628,n80,n1629);
not (n1629,n1630);
and (n1630,n457,n21);
and (n1631,n79,n456);
or (n1632,n1633,n1653);
and (n1633,n1634,n1647);
xor (n1634,n1635,n1641);
nand (n1635,n1636,n1640);
or (n1636,n460,n1637);
nor (n1637,n1638,n1639);
and (n1638,n558,n337);
and (n1639,n562,n338);
or (n1640,n461,n1578);
nand (n1641,n1642,n1646);
or (n1642,n484,n1643);
nor (n1643,n1644,n1645);
and (n1644,n228,n261);
and (n1645,n232,n257);
or (n1646,n1587,n485);
nand (n1647,n1648,n1652);
or (n1648,n246,n1649);
nor (n1649,n1650,n1651);
and (n1650,n424,n80);
and (n1651,n428,n75);
or (n1652,n1594,n254);
and (n1653,n1635,n1641);
and (n1654,n1613,n1619);
and (n1655,n1608,n1609);
and (n1656,n1429,n1512);
xor (n1657,n1658,n1691);
xor (n1658,n1659,n1688);
xor (n1659,n1660,n1667);
xor (n1660,n1661,n1664);
or (n1661,n1662,n1663);
and (n1662,n1542,n1555);
and (n1663,n1543,n1549);
or (n1664,n1665,n1666);
and (n1665,n1515,n1528);
and (n1666,n1516,n1522);
xor (n1667,n1668,n1681);
xor (n1668,n1669,n1675);
nand (n1669,n1670,n1671);
or (n1670,n246,n1552);
or (n1671,n1672,n254);
nor (n1672,n1673,n1674);
and (n1673,n80,n550);
and (n1674,n75,n554);
nand (n1675,n1676,n1677);
or (n1676,n333,n1557);
or (n1677,n334,n1678);
nor (n1678,n1679,n1680);
and (n1679,n182,n347);
and (n1680,n186,n348);
nand (n1681,n1682,n1687);
or (n1682,n19,n1683);
not (n1683,n1684);
nand (n1684,n1685,n1686);
or (n1685,n241,n83);
or (n1686,n90,n237);
or (n1687,n18,n1519);
or (n1688,n1689,n1690);
and (n1689,n1513,n1561);
and (n1690,n1514,n1541);
xor (n1691,n1692,n1719);
xor (n1692,n1693,n1716);
xor (n1693,n1694,n1710);
xor (n1694,n1695,n1701);
nand (n1695,n1696,n1697);
or (n1696,n460,n1449);
or (n1697,n461,n1698);
nor (n1698,n1699,n1700);
and (n1699,n337,n140);
and (n1700,n147,n338);
nand (n1701,n1702,n1706);
or (n1702,n510,n1703);
nor (n1703,n1704,n1705);
and (n1704,n521,n456);
and (n1705,n520,n457);
or (n1706,n1707,n530);
nor (n1707,n1708,n1709);
and (n1708,n416,n520);
and (n1709,n420,n521);
nand (n1710,n1711,n1715);
or (n1711,n1712,n485);
nor (n1712,n1713,n1714);
and (n1713,n375,n261);
and (n1714,n379,n257);
or (n1715,n484,n1546);
or (n1716,n1717,n1718);
and (n1717,n1430,n1481);
and (n1718,n1431,n1452);
xor (n1719,n1720,n1740);
xor (n1720,n1721,n1727);
nand (n1721,n1722,n1723);
or (n1722,n150,n1525);
or (n1723,n1724,n179);
nor (n1724,n1725,n1726);
and (n1725,n385,n153);
and (n1726,n389,n154);
xor (n1727,n1728,n1734);
nand (n1728,n1729,n1730);
or (n1729,n1440,n317);
or (n1730,n1731,n318);
nor (n1731,n1732,n1733);
and (n1732,n275,n311);
and (n1733,n282,n312);
nor (n1734,n1735,n520);
nor (n1735,n1736,n1739);
and (n1736,n153,n1737);
not (n1737,n1738);
and (n1738,n457,n514);
and (n1739,n525,n456);
or (n1740,n1741,n1742);
and (n1741,n1432,n1443);
and (n1742,n1433,n1434);
or (n1743,n1744,n2152);
and (n1744,n1745,n1776);
xor (n1745,n1746,n1775);
or (n1746,n1747,n1774);
and (n1747,n1748,n1773);
xor (n1748,n1749,n1772);
or (n1749,n1750,n1771);
and (n1750,n1751,n1754);
xor (n1751,n1752,n1753);
xor (n1752,n1567,n1575);
xor (n1753,n1584,n1597);
or (n1754,n1755,n1770);
and (n1755,n1756,n1769);
xor (n1756,n1757,n1763);
nand (n1757,n1758,n1762);
or (n1758,n18,n1759);
nor (n1759,n1760,n1761);
and (n1760,n83,n456);
and (n1761,n90,n457);
or (n1762,n1600,n19);
nand (n1763,n1764,n1768);
or (n1764,n333,n1765);
nor (n1765,n1766,n1767);
and (n1766,n586,n347);
and (n1767,n590,n348);
or (n1768,n1615,n334);
xor (n1769,n1620,n1626);
and (n1770,n1757,n1763);
and (n1771,n1752,n1753);
xor (n1772,n1563,n1582);
xor (n1773,n1607,n1610);
and (n1774,n1749,n1772);
xor (n1775,n1428,n1605);
nand (n1776,n1777,n2149,n2151);
or (n1777,n1778,n2144);
nand (n1778,n1779,n2133);
or (n1779,n1780,n2132);
and (n1780,n1781,n1902);
xor (n1781,n1782,n1887);
or (n1782,n1783,n1886);
and (n1783,n1784,n1852);
xor (n1784,n1785,n1807);
xor (n1785,n1786,n1801);
xor (n1786,n1787,n1794);
nand (n1787,n1788,n1793);
or (n1788,n484,n1789);
not (n1789,n1790);
nor (n1790,n1791,n1792);
and (n1791,n261,n389);
and (n1792,n385,n257);
or (n1793,n1643,n485);
nand (n1794,n1795,n1800);
or (n1795,n1796,n246);
not (n1796,n1797);
nand (n1797,n1798,n1799);
or (n1798,n420,n75);
or (n1799,n416,n80);
or (n1800,n1649,n254);
nand (n1801,n1802,n1806);
or (n1802,n333,n1803);
nor (n1803,n1804,n1805);
and (n1804,n237,n347);
and (n1805,n241,n348);
or (n1806,n334,n1765);
or (n1807,n1808,n1851);
and (n1808,n1809,n1831);
xor (n1809,n1810,n1816);
nand (n1810,n1811,n1815);
or (n1811,n333,n1812);
nor (n1812,n1813,n1814);
and (n1813,n228,n347);
and (n1814,n232,n348);
or (n1815,n1803,n334);
xor (n1816,n1817,n1823);
nor (n1817,n1818,n80);
nor (n1818,n1819,n1822);
and (n1819,n1820,n261);
not (n1820,n1821);
and (n1821,n457,n249);
and (n1822,n253,n456);
nand (n1823,n1824,n1827);
or (n1824,n317,n1825);
not (n1825,n1826);
xnor (n1826,n558,n311);
or (n1827,n1828,n318);
nor (n1828,n1829,n1830);
and (n1829,n311,n375);
and (n1830,n379,n312);
or (n1831,n1832,n1850);
and (n1832,n1833,n1841);
xor (n1833,n1834,n1835);
nor (n1834,n254,n456);
nand (n1835,n1836,n1837);
or (n1836,n318,n1825);
or (n1837,n1838,n317);
nor (n1838,n1839,n1840);
and (n1839,n311,n550);
and (n1840,n554,n312);
nand (n1841,n1842,n1846);
or (n1842,n484,n1843);
nor (n1843,n1844,n1845);
and (n1844,n416,n261);
and (n1845,n420,n257);
or (n1846,n1847,n485);
nor (n1847,n1848,n1849);
and (n1848,n424,n261);
and (n1849,n428,n257);
and (n1850,n1834,n1835);
and (n1851,n1810,n1816);
xor (n1852,n1853,n1867);
xor (n1853,n1854,n1855);
and (n1854,n1817,n1823);
xor (n1855,n1856,n1861);
xor (n1856,n1857,n1858);
nor (n1857,n19,n456);
nand (n1858,n1859,n1860);
or (n1859,n1828,n317);
or (n1860,n1622,n318);
nand (n1861,n1862,n1866);
or (n1862,n460,n1863);
nor (n1863,n1864,n1865);
and (n1864,n550,n337);
and (n1865,n554,n338);
or (n1866,n461,n1637);
or (n1867,n1868,n1885);
and (n1868,n1869,n1879);
xor (n1869,n1870,n1876);
nand (n1870,n1871,n1875);
or (n1871,n460,n1872);
nor (n1872,n1873,n1874);
and (n1873,n337,n586);
and (n1874,n590,n338);
or (n1875,n1863,n461);
nand (n1876,n1877,n1878);
or (n1877,n485,n1789);
or (n1878,n1847,n484);
nand (n1879,n1880,n1881);
or (n1880,n254,n1796);
or (n1881,n246,n1882);
nor (n1882,n1883,n1884);
and (n1883,n75,n456);
and (n1884,n80,n457);
and (n1885,n1870,n1876);
and (n1886,n1785,n1807);
xor (n1887,n1888,n1893);
xor (n1888,n1889,n1890);
xor (n1889,n1634,n1647);
or (n1890,n1891,n1892);
and (n1891,n1853,n1867);
and (n1892,n1854,n1855);
xor (n1893,n1894,n1901);
xor (n1894,n1895,n1898);
or (n1895,n1896,n1897);
and (n1896,n1856,n1861);
and (n1897,n1857,n1858);
or (n1898,n1899,n1900);
and (n1899,n1786,n1801);
and (n1900,n1787,n1794);
xor (n1901,n1756,n1769);
or (n1902,n1903,n2131);
and (n1903,n1904,n1941);
xor (n1904,n1905,n1940);
or (n1905,n1906,n1939);
and (n1906,n1907,n1938);
xor (n1907,n1908,n1937);
or (n1908,n1909,n1936);
and (n1909,n1910,n1923);
xor (n1910,n1911,n1917);
nand (n1911,n1912,n1916);
or (n1912,n460,n1913);
nor (n1913,n1914,n1915);
and (n1914,n237,n337);
and (n1915,n338,n241);
or (n1916,n1872,n461);
nand (n1917,n1918,n1922);
or (n1918,n333,n1919);
nor (n1919,n1920,n1921);
and (n1920,n385,n347);
and (n1921,n389,n348);
or (n1922,n1812,n334);
and (n1923,n1924,n1930);
nor (n1924,n1925,n261);
nor (n1925,n1926,n1929);
and (n1926,n1927,n347);
not (n1927,n1928);
and (n1928,n457,n487);
and (n1929,n491,n456);
nand (n1930,n1931,n1935);
or (n1931,n1932,n317);
nor (n1932,n1933,n1934);
and (n1933,n311,n586);
and (n1934,n590,n312);
or (n1935,n1838,n318);
and (n1936,n1911,n1917);
xor (n1937,n1869,n1879);
xor (n1938,n1809,n1831);
and (n1939,n1908,n1937);
xor (n1940,n1784,n1852);
nand (n1941,n1942,n2128,n2130);
or (n1942,n1943,n2001);
nand (n1943,n1944,n1996);
not (n1944,n1945);
nor (n1945,n1946,n1972);
xor (n1946,n1947,n1971);
xor (n1947,n1948,n1970);
or (n1948,n1949,n1969);
and (n1949,n1950,n1963);
xor (n1950,n1951,n1957);
nand (n1951,n1952,n1956);
or (n1952,n484,n1953);
nor (n1953,n1954,n1955);
and (n1954,n257,n456);
and (n1955,n261,n457);
or (n1956,n1843,n485);
nand (n1957,n1958,n1962);
or (n1958,n1959,n460);
nor (n1959,n1960,n1961);
and (n1960,n338,n232);
and (n1961,n337,n228);
or (n1962,n1913,n461);
nand (n1963,n1964,n1968);
or (n1964,n333,n1965);
nor (n1965,n1966,n1967);
and (n1966,n424,n347);
and (n1967,n428,n348);
or (n1968,n1919,n334);
and (n1969,n1951,n1957);
xor (n1970,n1833,n1841);
xor (n1971,n1910,n1923);
or (n1972,n1973,n1995);
and (n1973,n1974,n1994);
xor (n1974,n1975,n1976);
xor (n1975,n1924,n1930);
or (n1976,n1977,n1993);
and (n1977,n1978,n1987);
xor (n1978,n1979,n1980);
nor (n1979,n485,n456);
nand (n1980,n1981,n1986);
or (n1981,n1982,n317);
not (n1982,n1983);
nand (n1983,n1984,n1985);
or (n1984,n312,n241);
nand (n1985,n241,n312);
or (n1986,n1932,n318);
nand (n1987,n1988,n1992);
or (n1988,n460,n1989);
nor (n1989,n1990,n1991);
and (n1990,n337,n385);
and (n1991,n338,n389);
or (n1992,n1959,n461);
and (n1993,n1979,n1980);
xor (n1994,n1950,n1963);
and (n1995,n1975,n1976);
or (n1996,n1997,n1998);
xor (n1997,n1907,n1938);
or (n1998,n1999,n2000);
and (n1999,n1947,n1971);
and (n2000,n1948,n1970);
nor (n2001,n2002,n2127);
and (n2002,n2003,n2122);
or (n2003,n2004,n2121);
and (n2004,n2005,n2046);
xor (n2005,n2006,n2039);
or (n2006,n2007,n2038);
and (n2007,n2008,n2024);
xor (n2008,n2009,n2015);
nand (n2009,n2010,n2014);
or (n2010,n460,n2011);
nor (n2011,n2012,n2013);
and (n2012,n338,n428);
and (n2013,n337,n424);
or (n2014,n1989,n461);
or (n2015,n2016,n2020);
nor (n2016,n2017,n334);
nor (n2017,n2018,n2019);
and (n2018,n347,n416);
and (n2019,n348,n420);
nor (n2020,n333,n2021);
nor (n2021,n2022,n2023);
and (n2022,n348,n456);
and (n2023,n347,n457);
xor (n2024,n2025,n2031);
nor (n2025,n2026,n347);
nor (n2026,n2027,n2030);
and (n2027,n2028,n337);
not (n2028,n2029);
and (n2029,n457,n341);
and (n2030,n351,n456);
nand (n2031,n2032,n2037);
or (n2032,n317,n2033);
not (n2033,n2034);
nand (n2034,n2035,n2036);
or (n2035,n311,n228);
nand (n2036,n228,n311);
nand (n2037,n1983,n319);
and (n2038,n2009,n2015);
xor (n2039,n2040,n2045);
xor (n2040,n2041,n2044);
nand (n2041,n2042,n2043);
or (n2042,n333,n2017);
or (n2043,n1965,n334);
and (n2044,n2025,n2031);
xor (n2045,n1978,n1987);
or (n2046,n2047,n2120);
and (n2047,n2048,n2068);
xor (n2048,n2049,n2067);
or (n2049,n2050,n2066);
and (n2050,n2051,n2060);
xor (n2051,n2052,n2053);
and (n2052,n335,n457);
nand (n2053,n2054,n2059);
or (n2054,n317,n2055);
not (n2055,n2056);
nand (n2056,n2057,n2058);
or (n2057,n312,n389);
nand (n2058,n389,n312);
nand (n2059,n2034,n319);
nand (n2060,n2061,n2065);
or (n2061,n460,n2062);
nor (n2062,n2063,n2064);
and (n2063,n337,n416);
and (n2064,n338,n420);
or (n2065,n2011,n461);
and (n2066,n2052,n2053);
xor (n2067,n2008,n2024);
or (n2068,n2069,n2119);
and (n2069,n2070,n2087);
xor (n2070,n2071,n2086);
and (n2071,n2072,n2078);
and (n2072,n2073,n338);
nand (n2073,n2074,n2077);
nand (n2074,n2075,n311);
not (n2075,n2076);
and (n2076,n457,n463);
nand (n2077,n467,n456);
nand (n2078,n2079,n2080);
or (n2079,n318,n2055);
nand (n2080,n2081,n2085);
not (n2081,n2082);
nor (n2082,n2083,n2084);
and (n2083,n428,n312);
and (n2084,n424,n311);
not (n2085,n317);
xor (n2086,n2051,n2060);
or (n2087,n2088,n2118);
and (n2088,n2089,n2097);
xor (n2089,n2090,n2096);
nand (n2090,n2091,n2095);
or (n2091,n460,n2092);
nor (n2092,n2093,n2094);
and (n2093,n338,n456);
and (n2094,n337,n457);
or (n2095,n2062,n461);
xor (n2096,n2072,n2078);
or (n2097,n2098,n2117);
and (n2098,n2099,n2107);
xor (n2099,n2100,n2101);
nor (n2100,n461,n456);
nand (n2101,n2102,n2106);
or (n2102,n2103,n317);
or (n2103,n2104,n2105);
and (n2104,n311,n420);
and (n2105,n416,n312);
or (n2106,n2082,n318);
nor (n2107,n2108,n2115);
nor (n2108,n2109,n2111);
and (n2109,n2110,n319);
not (n2110,n2103);
and (n2111,n2112,n2085);
nand (n2112,n2113,n2114);
or (n2113,n311,n457);
or (n2114,n312,n456);
or (n2115,n311,n2116);
and (n2116,n457,n319);
and (n2117,n2100,n2101);
and (n2118,n2090,n2096);
and (n2119,n2071,n2086);
and (n2120,n2049,n2067);
and (n2121,n2006,n2039);
or (n2122,n2123,n2124);
xor (n2123,n1974,n1994);
or (n2124,n2125,n2126);
and (n2125,n2040,n2045);
and (n2126,n2041,n2044);
and (n2127,n2123,n2124);
nand (n2128,n1996,n2129);
and (n2129,n1946,n1972);
nand (n2130,n1997,n1998);
and (n2131,n1905,n1940);
and (n2132,n1782,n1887);
or (n2133,n2134,n2141);
xor (n2134,n2135,n2140);
xor (n2135,n2136,n2137);
xor (n2136,n1612,n1632);
or (n2137,n2138,n2139);
and (n2138,n1894,n1901);
and (n2139,n1895,n1898);
xor (n2140,n1751,n1754);
or (n2141,n2142,n2143);
and (n2142,n1888,n1893);
and (n2143,n1889,n1890);
nor (n2144,n2145,n2146);
xor (n2145,n1748,n1773);
or (n2146,n2147,n2148);
and (n2147,n2135,n2140);
and (n2148,n2136,n2137);
or (n2149,n2144,n2150);
nand (n2150,n2134,n2141);
nand (n2151,n2145,n2146);
and (n2152,n1746,n1775);
and (n2153,n1426,n1657);
nor (n2154,n2155,n2275);
nor (n2155,n2156,n2266);
xor (n2156,n2157,n2221);
xor (n2157,n2158,n2196);
xor (n2158,n2159,n2181);
xor (n2159,n2160,n2161);
xor (n2160,n1377,n1390);
xor (n2161,n2162,n2175);
xor (n2162,n2163,n2169);
nand (n2163,n2164,n2168);
or (n2164,n460,n2165);
nor (n2165,n2166,n2167);
and (n2166,n337,n264);
and (n2167,n271,n338);
or (n2168,n461,n1309);
nand (n2169,n2170,n2174);
or (n2170,n246,n2171);
nor (n2171,n2172,n2173);
and (n2172,n80,n558);
and (n2173,n75,n562);
or (n2174,n1328,n254);
nand (n2175,n2176,n2180);
or (n2176,n2177,n333);
nor (n2177,n2178,n2179);
and (n2178,n93,n347);
and (n2179,n136,n348);
or (n2180,n334,n1334);
xor (n2181,n2182,n2195);
xor (n2182,n2183,n2189);
nand (n2183,n2184,n2188);
or (n2184,n18,n2185);
nor (n2185,n2186,n2187);
and (n2186,n90,n586);
and (n2187,n83,n590);
or (n2188,n1340,n19);
nand (n2189,n2190,n2194);
or (n2190,n150,n2191);
nor (n2191,n2192,n2193);
and (n2192,n153,n228);
and (n2193,n232,n154);
or (n2194,n179,n1358);
xor (n2195,n1363,n1369);
or (n2196,n2197,n2220);
and (n2197,n2198,n2205);
xor (n2198,n2199,n2202);
or (n2199,n2200,n2201);
and (n2200,n1720,n1740);
and (n2201,n1721,n1727);
or (n2202,n2203,n2204);
and (n2203,n1660,n1667);
and (n2204,n1661,n1664);
xor (n2205,n2206,n2217);
xor (n2206,n2207,n2208);
and (n2207,n1728,n1734);
xor (n2208,n2209,n2214);
xor (n2209,n2210,n2211);
nor (n2210,n538,n456);
nand (n2211,n2212,n2213);
or (n2212,n1731,n317);
or (n2213,n1371,n318);
nand (n2214,n2215,n2216);
or (n2215,n460,n1698);
or (n2216,n461,n2165);
or (n2217,n2218,n2219);
and (n2218,n1694,n1710);
and (n2219,n1695,n1701);
and (n2220,n2199,n2202);
xor (n2221,n2222,n2257);
xor (n2222,n2223,n2226);
or (n2223,n2224,n2225);
and (n2224,n2206,n2217);
and (n2225,n2207,n2208);
xor (n2226,n2227,n2244);
xor (n2227,n2228,n2231);
or (n2228,n2229,n2230);
and (n2229,n2209,n2214);
and (n2230,n2210,n2211);
or (n2231,n2232,n2243);
and (n2232,n2233,n2240);
xor (n2233,n2234,n2237);
nand (n2234,n2235,n2236);
or (n2235,n333,n1678);
or (n2236,n334,n2177);
nand (n2237,n2238,n2239);
or (n2238,n1683,n18);
or (n2239,n2185,n19);
nand (n2240,n2241,n2242);
or (n2241,n150,n1724);
or (n2242,n2191,n179);
and (n2243,n2234,n2237);
or (n2244,n2245,n2256);
and (n2245,n2246,n2253);
xor (n2246,n2247,n2250);
nand (n2247,n2248,n2249);
or (n2248,n510,n1707);
or (n2249,n1386,n530);
nand (n2250,n2251,n2252);
or (n2251,n484,n1712);
or (n2252,n1380,n485);
nand (n2253,n2254,n2255);
or (n2254,n246,n1672);
or (n2255,n2171,n254);
and (n2256,n2247,n2250);
or (n2257,n2258,n2265);
and (n2258,n2259,n2264);
xor (n2259,n2260,n2263);
or (n2260,n2261,n2262);
and (n2261,n1668,n1681);
and (n2262,n1669,n1675);
xor (n2263,n2233,n2240);
xor (n2264,n2246,n2253);
and (n2265,n2260,n2263);
or (n2266,n2267,n2274);
and (n2267,n2268,n2273);
xor (n2268,n2269,n2270);
xor (n2269,n2259,n2264);
or (n2270,n2271,n2272);
and (n2271,n1692,n1719);
and (n2272,n1693,n1716);
xor (n2273,n2198,n2205);
and (n2274,n2269,n2270);
nor (n2275,n2276,n2277);
xor (n2276,n2268,n2273);
or (n2277,n2278,n2279);
and (n2278,n1658,n1691);
and (n2279,n1659,n1688);
or (n2280,n2281,n2326);
nor (n2281,n2282,n2317);
xor (n2282,n2283,n2302);
xor (n2283,n2284,n2285);
xor (n2284,n1351,n1399);
or (n2285,n2286,n2301);
and (n2286,n2287,n2294);
xor (n2287,n2288,n2291);
or (n2288,n2289,n2290);
and (n2289,n2227,n2244);
and (n2290,n2228,n2231);
or (n2291,n2292,n2293);
and (n2292,n2159,n2181);
and (n2293,n2160,n2161);
xor (n2294,n2295,n2300);
xor (n2295,n2296,n2299);
or (n2296,n2297,n2298);
and (n2297,n2162,n2175);
and (n2298,n2163,n2169);
xor (n2299,n1325,n1338);
xor (n2300,n1277,n1285);
and (n2301,n2288,n2291);
xor (n2302,n2303,n2308);
xor (n2303,n2304,n2307);
or (n2304,n2305,n2306);
and (n2305,n2295,n2300);
and (n2306,n2296,n2299);
xor (n2307,n1322,n1346);
or (n2308,n2309,n2316);
and (n2309,n2310,n2315);
xor (n2310,n2311,n2312);
xor (n2311,n1294,n1307);
or (n2312,n2313,n2314);
and (n2313,n2182,n2195);
and (n2314,n2183,n2189);
xor (n2315,n1355,n1375);
and (n2316,n2311,n2312);
or (n2317,n2318,n2325);
and (n2318,n2319,n2324);
xor (n2319,n2320,n2321);
xor (n2320,n2310,n2315);
or (n2321,n2322,n2323);
and (n2322,n2222,n2257);
and (n2323,n2223,n2226);
xor (n2324,n2287,n2294);
and (n2325,n2320,n2321);
nor (n2326,n2327,n2330);
or (n2327,n2328,n2329);
and (n2328,n2157,n2221);
and (n2329,n2158,n2196);
xor (n2330,n2319,n2324);
nand (n2331,n2332,n2341);
or (n2332,n2333,n2281);
nor (n2333,n2334,n2340);
and (n2334,n2335,n2339);
nand (n2335,n2336,n2338);
or (n2336,n2155,n2337);
nand (n2337,n2276,n2277);
nand (n2338,n2156,n2266);
not (n2339,n2326);
and (n2340,n2327,n2330);
nand (n2341,n2282,n2317);
or (n2342,n2343,n2350);
xor (n2343,n2344,n2349);
xor (n2344,n2345,n2346);
xor (n2345,n1269,n1315);
or (n2346,n2347,n2348);
and (n2347,n2303,n2308);
and (n2348,n2304,n2307);
xor (n2349,n1319,n1349);
or (n2350,n2351,n2352);
and (n2351,n2283,n2302);
and (n2352,n2284,n2285);
and (n2353,n2354,n2356);
not (n2354,n2355);
xor (n2355,n1182,n1317);
not (n2356,n2357);
or (n2357,n2358,n2359);
and (n2358,n2344,n2349);
and (n2359,n2345,n2346);
nor (n2360,n2361,n2365);
and (n2361,n2362,n2363);
not (n2362,n2353);
not (n2363,n2364);
nand (n2364,n2343,n2350);
nor (n2365,n2354,n2356);
and (n2366,n1180,n1403);
nand (n2367,n2368,n2372);
not (n2368,n2369);
or (n2369,n2370,n2371);
and (n2370,n1404,n1413);
and (n2371,n1405,n1406);
not (n2372,n2373);
xor (n2373,n2374,n2379);
xor (n2374,n2375,n2376);
xor (n2375,n849,n879);
or (n2376,n2377,n2378);
and (n2377,n1407,n1410);
and (n2378,n1408,n1409);
xor (n2379,n883,n924);
nor (n2380,n2372,n2368);
nor (n2381,n2382,n2383);
xor (n2382,n8,n881);
or (n2383,n2384,n2385);
and (n2384,n2374,n2379);
and (n2385,n2375,n2376);
nand (n2386,n2382,n2383);
or (n2387,n1173,n3);
xor (n2388,n2389,n4176);
xor (n2389,n2390,n4174);
xor (n2390,n2391,n4173);
xor (n2391,n2392,n4164);
xor (n2392,n2393,n4163);
xor (n2393,n2394,n4149);
xor (n2394,n2395,n4148);
xor (n2395,n2396,n4127);
xor (n2396,n2397,n4126);
xor (n2397,n2398,n4100);
xor (n2398,n2399,n4099);
xor (n2399,n2400,n4066);
xor (n2400,n2401,n4065);
xor (n2401,n2402,n4027);
xor (n2402,n2403,n4026);
xor (n2403,n2404,n3981);
xor (n2404,n2405,n3980);
xor (n2405,n2406,n3930);
xor (n2406,n2407,n3929);
xor (n2407,n2408,n3872);
xor (n2408,n2409,n3871);
xor (n2409,n2410,n3809);
xor (n2410,n2411,n3808);
xor (n2411,n2412,n3739);
xor (n2412,n2413,n3738);
xor (n2413,n2414,n3664);
xor (n2414,n2415,n3663);
xor (n2415,n2416,n3582);
xor (n2416,n2417,n3581);
xor (n2417,n2418,n3495);
xor (n2418,n2419,n3494);
xor (n2419,n2420,n3401);
xor (n2420,n2421,n3400);
xor (n2421,n2422,n3302);
xor (n2422,n2423,n3301);
xor (n2423,n2424,n3197);
xor (n2424,n2425,n3196);
xor (n2425,n2426,n3086);
xor (n2426,n2427,n3085);
xor (n2427,n2428,n2968);
xor (n2428,n2429,n2967);
xor (n2429,n2430,n2845);
xor (n2430,n2431,n2844);
xor (n2431,n2432,n2715);
xor (n2432,n2433,n2714);
xor (n2433,n2434,n2580);
xor (n2434,n2435,n2579);
xor (n2435,n2436,n2439);
xor (n2436,n2437,n2438);
and (n2437,n1117,n319);
and (n2438,n634,n312);
or (n2439,n2440,n2443);
and (n2440,n2441,n2442);
and (n2441,n634,n319);
and (n2442,n323,n312);
and (n2443,n2444,n2445);
xor (n2444,n2441,n2442);
or (n2445,n2446,n2449);
and (n2446,n2447,n2448);
and (n2447,n323,n319);
and (n2448,n287,n312);
and (n2449,n2450,n2451);
xor (n2450,n2447,n2448);
or (n2451,n2452,n2455);
and (n2452,n2453,n2454);
and (n2453,n287,n319);
and (n2454,n473,n312);
and (n2455,n2456,n2457);
xor (n2456,n2453,n2454);
or (n2457,n2458,n2461);
and (n2458,n2459,n2460);
and (n2459,n473,n319);
and (n2460,n647,n312);
and (n2461,n2462,n2463);
xor (n2462,n2459,n2460);
or (n2463,n2464,n2467);
and (n2464,n2465,n2466);
and (n2465,n647,n319);
and (n2466,n363,n312);
and (n2467,n2468,n2469);
xor (n2468,n2465,n2466);
or (n2469,n2470,n2473);
and (n2470,n2471,n2472);
and (n2471,n363,n319);
and (n2472,n355,n312);
and (n2473,n2474,n2475);
xor (n2474,n2471,n2472);
or (n2475,n2476,n2479);
and (n2476,n2477,n2478);
and (n2477,n355,n319);
and (n2478,n497,n312);
and (n2479,n2480,n2481);
xor (n2480,n2477,n2478);
or (n2481,n2482,n2485);
and (n2482,n2483,n2484);
and (n2483,n497,n319);
and (n2484,n568,n312);
and (n2485,n2486,n2487);
xor (n2486,n2483,n2484);
or (n2487,n2488,n2491);
and (n2488,n2489,n2490);
and (n2489,n568,n319);
and (n2490,n275,n312);
and (n2491,n2492,n2493);
xor (n2492,n2489,n2490);
or (n2493,n2494,n2497);
and (n2494,n2495,n2496);
and (n2495,n275,n319);
and (n2496,n264,n312);
and (n2497,n2498,n2499);
xor (n2498,n2495,n2496);
or (n2499,n2500,n2503);
and (n2500,n2501,n2502);
and (n2501,n264,n319);
and (n2502,n140,n312);
and (n2503,n2504,n2505);
xor (n2504,n2501,n2502);
or (n2505,n2506,n2509);
and (n2506,n2507,n2508);
and (n2507,n140,n319);
and (n2508,n93,n312);
and (n2509,n2510,n2511);
xor (n2510,n2507,n2508);
or (n2511,n2512,n2515);
and (n2512,n2513,n2514);
and (n2513,n93,n319);
and (n2514,n182,n312);
and (n2515,n2516,n2517);
xor (n2516,n2513,n2514);
or (n2517,n2518,n2521);
and (n2518,n2519,n2520);
and (n2519,n182,n319);
and (n2520,n173,n312);
and (n2521,n2522,n2523);
xor (n2522,n2519,n2520);
or (n2523,n2524,n2527);
and (n2524,n2525,n2526);
and (n2525,n173,n319);
and (n2526,n375,n312);
and (n2527,n2528,n2529);
xor (n2528,n2525,n2526);
or (n2529,n2530,n2533);
and (n2530,n2531,n2532);
and (n2531,n375,n319);
and (n2532,n558,n312);
and (n2533,n2534,n2535);
xor (n2534,n2531,n2532);
or (n2535,n2536,n2539);
and (n2536,n2537,n2538);
and (n2537,n558,n319);
and (n2538,n550,n312);
and (n2539,n2540,n2541);
xor (n2540,n2537,n2538);
or (n2541,n2542,n2545);
and (n2542,n2543,n2544);
and (n2543,n550,n319);
and (n2544,n586,n312);
and (n2545,n2546,n2547);
xor (n2546,n2543,n2544);
or (n2547,n2548,n2551);
and (n2548,n2549,n2550);
and (n2549,n586,n319);
and (n2550,n237,n312);
and (n2551,n2552,n2553);
xor (n2552,n2549,n2550);
or (n2553,n2554,n2557);
and (n2554,n2555,n2556);
and (n2555,n237,n319);
and (n2556,n228,n312);
and (n2557,n2558,n2559);
xor (n2558,n2555,n2556);
or (n2559,n2560,n2563);
and (n2560,n2561,n2562);
and (n2561,n228,n319);
and (n2562,n385,n312);
and (n2563,n2564,n2565);
xor (n2564,n2561,n2562);
or (n2565,n2566,n2569);
and (n2566,n2567,n2568);
and (n2567,n385,n319);
and (n2568,n424,n312);
and (n2569,n2570,n2571);
xor (n2570,n2567,n2568);
or (n2571,n2572,n2574);
and (n2572,n2573,n2105);
and (n2573,n424,n319);
and (n2574,n2575,n2576);
xor (n2575,n2573,n2105);
and (n2576,n2577,n2578);
and (n2577,n416,n319);
and (n2578,n457,n312);
and (n2579,n323,n463);
or (n2580,n2581,n2584);
and (n2581,n2582,n2583);
xor (n2582,n2444,n2445);
and (n2583,n287,n463);
and (n2584,n2585,n2586);
xor (n2585,n2582,n2583);
or (n2586,n2587,n2590);
and (n2587,n2588,n2589);
xor (n2588,n2450,n2451);
and (n2589,n473,n463);
and (n2590,n2591,n2592);
xor (n2591,n2588,n2589);
or (n2592,n2593,n2596);
and (n2593,n2594,n2595);
xor (n2594,n2456,n2457);
and (n2595,n647,n463);
and (n2596,n2597,n2598);
xor (n2597,n2594,n2595);
or (n2598,n2599,n2602);
and (n2599,n2600,n2601);
xor (n2600,n2462,n2463);
and (n2601,n363,n463);
and (n2602,n2603,n2604);
xor (n2603,n2600,n2601);
or (n2604,n2605,n2608);
and (n2605,n2606,n2607);
xor (n2606,n2468,n2469);
and (n2607,n355,n463);
and (n2608,n2609,n2610);
xor (n2609,n2606,n2607);
or (n2610,n2611,n2614);
and (n2611,n2612,n2613);
xor (n2612,n2474,n2475);
and (n2613,n497,n463);
and (n2614,n2615,n2616);
xor (n2615,n2612,n2613);
or (n2616,n2617,n2620);
and (n2617,n2618,n2619);
xor (n2618,n2480,n2481);
and (n2619,n568,n463);
and (n2620,n2621,n2622);
xor (n2621,n2618,n2619);
or (n2622,n2623,n2626);
and (n2623,n2624,n2625);
xor (n2624,n2486,n2487);
and (n2625,n275,n463);
and (n2626,n2627,n2628);
xor (n2627,n2624,n2625);
or (n2628,n2629,n2632);
and (n2629,n2630,n2631);
xor (n2630,n2492,n2493);
and (n2631,n264,n463);
and (n2632,n2633,n2634);
xor (n2633,n2630,n2631);
or (n2634,n2635,n2638);
and (n2635,n2636,n2637);
xor (n2636,n2498,n2499);
and (n2637,n140,n463);
and (n2638,n2639,n2640);
xor (n2639,n2636,n2637);
or (n2640,n2641,n2644);
and (n2641,n2642,n2643);
xor (n2642,n2504,n2505);
and (n2643,n93,n463);
and (n2644,n2645,n2646);
xor (n2645,n2642,n2643);
or (n2646,n2647,n2650);
and (n2647,n2648,n2649);
xor (n2648,n2510,n2511);
and (n2649,n182,n463);
and (n2650,n2651,n2652);
xor (n2651,n2648,n2649);
or (n2652,n2653,n2656);
and (n2653,n2654,n2655);
xor (n2654,n2516,n2517);
and (n2655,n173,n463);
and (n2656,n2657,n2658);
xor (n2657,n2654,n2655);
or (n2658,n2659,n2662);
and (n2659,n2660,n2661);
xor (n2660,n2522,n2523);
and (n2661,n375,n463);
and (n2662,n2663,n2664);
xor (n2663,n2660,n2661);
or (n2664,n2665,n2668);
and (n2665,n2666,n2667);
xor (n2666,n2528,n2529);
and (n2667,n558,n463);
and (n2668,n2669,n2670);
xor (n2669,n2666,n2667);
or (n2670,n2671,n2674);
and (n2671,n2672,n2673);
xor (n2672,n2534,n2535);
and (n2673,n550,n463);
and (n2674,n2675,n2676);
xor (n2675,n2672,n2673);
or (n2676,n2677,n2680);
and (n2677,n2678,n2679);
xor (n2678,n2540,n2541);
and (n2679,n586,n463);
and (n2680,n2681,n2682);
xor (n2681,n2678,n2679);
or (n2682,n2683,n2686);
and (n2683,n2684,n2685);
xor (n2684,n2546,n2547);
and (n2685,n237,n463);
and (n2686,n2687,n2688);
xor (n2687,n2684,n2685);
or (n2688,n2689,n2692);
and (n2689,n2690,n2691);
xor (n2690,n2552,n2553);
and (n2691,n228,n463);
and (n2692,n2693,n2694);
xor (n2693,n2690,n2691);
or (n2694,n2695,n2698);
and (n2695,n2696,n2697);
xor (n2696,n2558,n2559);
and (n2697,n385,n463);
and (n2698,n2699,n2700);
xor (n2699,n2696,n2697);
or (n2700,n2701,n2704);
and (n2701,n2702,n2703);
xor (n2702,n2564,n2565);
and (n2703,n424,n463);
and (n2704,n2705,n2706);
xor (n2705,n2702,n2703);
or (n2706,n2707,n2710);
and (n2707,n2708,n2709);
xor (n2708,n2570,n2571);
and (n2709,n416,n463);
and (n2710,n2711,n2712);
xor (n2711,n2708,n2709);
and (n2712,n2713,n2076);
xor (n2713,n2575,n2576);
and (n2714,n287,n338);
or (n2715,n2716,n2719);
and (n2716,n2717,n2718);
xor (n2717,n2585,n2586);
and (n2718,n473,n338);
and (n2719,n2720,n2721);
xor (n2720,n2717,n2718);
or (n2721,n2722,n2725);
and (n2722,n2723,n2724);
xor (n2723,n2591,n2592);
and (n2724,n647,n338);
and (n2725,n2726,n2727);
xor (n2726,n2723,n2724);
or (n2727,n2728,n2731);
and (n2728,n2729,n2730);
xor (n2729,n2597,n2598);
and (n2730,n363,n338);
and (n2731,n2732,n2733);
xor (n2732,n2729,n2730);
or (n2733,n2734,n2737);
and (n2734,n2735,n2736);
xor (n2735,n2603,n2604);
and (n2736,n355,n338);
and (n2737,n2738,n2739);
xor (n2738,n2735,n2736);
or (n2739,n2740,n2743);
and (n2740,n2741,n2742);
xor (n2741,n2609,n2610);
and (n2742,n497,n338);
and (n2743,n2744,n2745);
xor (n2744,n2741,n2742);
or (n2745,n2746,n2749);
and (n2746,n2747,n2748);
xor (n2747,n2615,n2616);
and (n2748,n568,n338);
and (n2749,n2750,n2751);
xor (n2750,n2747,n2748);
or (n2751,n2752,n2755);
and (n2752,n2753,n2754);
xor (n2753,n2621,n2622);
and (n2754,n275,n338);
and (n2755,n2756,n2757);
xor (n2756,n2753,n2754);
or (n2757,n2758,n2761);
and (n2758,n2759,n2760);
xor (n2759,n2627,n2628);
and (n2760,n264,n338);
and (n2761,n2762,n2763);
xor (n2762,n2759,n2760);
or (n2763,n2764,n2767);
and (n2764,n2765,n2766);
xor (n2765,n2633,n2634);
and (n2766,n140,n338);
and (n2767,n2768,n2769);
xor (n2768,n2765,n2766);
or (n2769,n2770,n2773);
and (n2770,n2771,n2772);
xor (n2771,n2639,n2640);
and (n2772,n93,n338);
and (n2773,n2774,n2775);
xor (n2774,n2771,n2772);
or (n2775,n2776,n2779);
and (n2776,n2777,n2778);
xor (n2777,n2645,n2646);
and (n2778,n182,n338);
and (n2779,n2780,n2781);
xor (n2780,n2777,n2778);
or (n2781,n2782,n2785);
and (n2782,n2783,n2784);
xor (n2783,n2651,n2652);
and (n2784,n173,n338);
and (n2785,n2786,n2787);
xor (n2786,n2783,n2784);
or (n2787,n2788,n2791);
and (n2788,n2789,n2790);
xor (n2789,n2657,n2658);
and (n2790,n375,n338);
and (n2791,n2792,n2793);
xor (n2792,n2789,n2790);
or (n2793,n2794,n2797);
and (n2794,n2795,n2796);
xor (n2795,n2663,n2664);
and (n2796,n558,n338);
and (n2797,n2798,n2799);
xor (n2798,n2795,n2796);
or (n2799,n2800,n2803);
and (n2800,n2801,n2802);
xor (n2801,n2669,n2670);
and (n2802,n550,n338);
and (n2803,n2804,n2805);
xor (n2804,n2801,n2802);
or (n2805,n2806,n2809);
and (n2806,n2807,n2808);
xor (n2807,n2675,n2676);
and (n2808,n586,n338);
and (n2809,n2810,n2811);
xor (n2810,n2807,n2808);
or (n2811,n2812,n2815);
and (n2812,n2813,n2814);
xor (n2813,n2681,n2682);
and (n2814,n237,n338);
and (n2815,n2816,n2817);
xor (n2816,n2813,n2814);
or (n2817,n2818,n2821);
and (n2818,n2819,n2820);
xor (n2819,n2687,n2688);
and (n2820,n228,n338);
and (n2821,n2822,n2823);
xor (n2822,n2819,n2820);
or (n2823,n2824,n2827);
and (n2824,n2825,n2826);
xor (n2825,n2693,n2694);
and (n2826,n385,n338);
and (n2827,n2828,n2829);
xor (n2828,n2825,n2826);
or (n2829,n2830,n2833);
and (n2830,n2831,n2832);
xor (n2831,n2699,n2700);
and (n2832,n424,n338);
and (n2833,n2834,n2835);
xor (n2834,n2831,n2832);
or (n2835,n2836,n2839);
and (n2836,n2837,n2838);
xor (n2837,n2705,n2706);
and (n2838,n416,n338);
and (n2839,n2840,n2841);
xor (n2840,n2837,n2838);
and (n2841,n2842,n2843);
xor (n2842,n2711,n2712);
and (n2843,n457,n338);
and (n2844,n473,n341);
or (n2845,n2846,n2849);
and (n2846,n2847,n2848);
xor (n2847,n2720,n2721);
and (n2848,n647,n341);
and (n2849,n2850,n2851);
xor (n2850,n2847,n2848);
or (n2851,n2852,n2855);
and (n2852,n2853,n2854);
xor (n2853,n2726,n2727);
and (n2854,n363,n341);
and (n2855,n2856,n2857);
xor (n2856,n2853,n2854);
or (n2857,n2858,n2861);
and (n2858,n2859,n2860);
xor (n2859,n2732,n2733);
and (n2860,n355,n341);
and (n2861,n2862,n2863);
xor (n2862,n2859,n2860);
or (n2863,n2864,n2867);
and (n2864,n2865,n2866);
xor (n2865,n2738,n2739);
and (n2866,n497,n341);
and (n2867,n2868,n2869);
xor (n2868,n2865,n2866);
or (n2869,n2870,n2873);
and (n2870,n2871,n2872);
xor (n2871,n2744,n2745);
and (n2872,n568,n341);
and (n2873,n2874,n2875);
xor (n2874,n2871,n2872);
or (n2875,n2876,n2879);
and (n2876,n2877,n2878);
xor (n2877,n2750,n2751);
and (n2878,n275,n341);
and (n2879,n2880,n2881);
xor (n2880,n2877,n2878);
or (n2881,n2882,n2885);
and (n2882,n2883,n2884);
xor (n2883,n2756,n2757);
and (n2884,n264,n341);
and (n2885,n2886,n2887);
xor (n2886,n2883,n2884);
or (n2887,n2888,n2891);
and (n2888,n2889,n2890);
xor (n2889,n2762,n2763);
and (n2890,n140,n341);
and (n2891,n2892,n2893);
xor (n2892,n2889,n2890);
or (n2893,n2894,n2897);
and (n2894,n2895,n2896);
xor (n2895,n2768,n2769);
and (n2896,n93,n341);
and (n2897,n2898,n2899);
xor (n2898,n2895,n2896);
or (n2899,n2900,n2903);
and (n2900,n2901,n2902);
xor (n2901,n2774,n2775);
and (n2902,n182,n341);
and (n2903,n2904,n2905);
xor (n2904,n2901,n2902);
or (n2905,n2906,n2909);
and (n2906,n2907,n2908);
xor (n2907,n2780,n2781);
and (n2908,n173,n341);
and (n2909,n2910,n2911);
xor (n2910,n2907,n2908);
or (n2911,n2912,n2915);
and (n2912,n2913,n2914);
xor (n2913,n2786,n2787);
and (n2914,n375,n341);
and (n2915,n2916,n2917);
xor (n2916,n2913,n2914);
or (n2917,n2918,n2921);
and (n2918,n2919,n2920);
xor (n2919,n2792,n2793);
and (n2920,n558,n341);
and (n2921,n2922,n2923);
xor (n2922,n2919,n2920);
or (n2923,n2924,n2927);
and (n2924,n2925,n2926);
xor (n2925,n2798,n2799);
and (n2926,n550,n341);
and (n2927,n2928,n2929);
xor (n2928,n2925,n2926);
or (n2929,n2930,n2933);
and (n2930,n2931,n2932);
xor (n2931,n2804,n2805);
and (n2932,n586,n341);
and (n2933,n2934,n2935);
xor (n2934,n2931,n2932);
or (n2935,n2936,n2939);
and (n2936,n2937,n2938);
xor (n2937,n2810,n2811);
and (n2938,n237,n341);
and (n2939,n2940,n2941);
xor (n2940,n2937,n2938);
or (n2941,n2942,n2945);
and (n2942,n2943,n2944);
xor (n2943,n2816,n2817);
and (n2944,n228,n341);
and (n2945,n2946,n2947);
xor (n2946,n2943,n2944);
or (n2947,n2948,n2951);
and (n2948,n2949,n2950);
xor (n2949,n2822,n2823);
and (n2950,n385,n341);
and (n2951,n2952,n2953);
xor (n2952,n2949,n2950);
or (n2953,n2954,n2957);
and (n2954,n2955,n2956);
xor (n2955,n2828,n2829);
and (n2956,n424,n341);
and (n2957,n2958,n2959);
xor (n2958,n2955,n2956);
or (n2959,n2960,n2963);
and (n2960,n2961,n2962);
xor (n2961,n2834,n2835);
and (n2962,n416,n341);
and (n2963,n2964,n2965);
xor (n2964,n2961,n2962);
and (n2965,n2966,n2029);
xor (n2966,n2840,n2841);
and (n2967,n647,n348);
or (n2968,n2969,n2972);
and (n2969,n2970,n2971);
xor (n2970,n2850,n2851);
and (n2971,n363,n348);
and (n2972,n2973,n2974);
xor (n2973,n2970,n2971);
or (n2974,n2975,n2978);
and (n2975,n2976,n2977);
xor (n2976,n2856,n2857);
and (n2977,n355,n348);
and (n2978,n2979,n2980);
xor (n2979,n2976,n2977);
or (n2980,n2981,n2984);
and (n2981,n2982,n2983);
xor (n2982,n2862,n2863);
and (n2983,n497,n348);
and (n2984,n2985,n2986);
xor (n2985,n2982,n2983);
or (n2986,n2987,n2990);
and (n2987,n2988,n2989);
xor (n2988,n2868,n2869);
and (n2989,n568,n348);
and (n2990,n2991,n2992);
xor (n2991,n2988,n2989);
or (n2992,n2993,n2996);
and (n2993,n2994,n2995);
xor (n2994,n2874,n2875);
and (n2995,n275,n348);
and (n2996,n2997,n2998);
xor (n2997,n2994,n2995);
or (n2998,n2999,n3002);
and (n2999,n3000,n3001);
xor (n3000,n2880,n2881);
and (n3001,n264,n348);
and (n3002,n3003,n3004);
xor (n3003,n3000,n3001);
or (n3004,n3005,n3008);
and (n3005,n3006,n3007);
xor (n3006,n2886,n2887);
and (n3007,n140,n348);
and (n3008,n3009,n3010);
xor (n3009,n3006,n3007);
or (n3010,n3011,n3014);
and (n3011,n3012,n3013);
xor (n3012,n2892,n2893);
and (n3013,n93,n348);
and (n3014,n3015,n3016);
xor (n3015,n3012,n3013);
or (n3016,n3017,n3020);
and (n3017,n3018,n3019);
xor (n3018,n2898,n2899);
and (n3019,n182,n348);
and (n3020,n3021,n3022);
xor (n3021,n3018,n3019);
or (n3022,n3023,n3026);
and (n3023,n3024,n3025);
xor (n3024,n2904,n2905);
and (n3025,n173,n348);
and (n3026,n3027,n3028);
xor (n3027,n3024,n3025);
or (n3028,n3029,n3032);
and (n3029,n3030,n3031);
xor (n3030,n2910,n2911);
and (n3031,n375,n348);
and (n3032,n3033,n3034);
xor (n3033,n3030,n3031);
or (n3034,n3035,n3038);
and (n3035,n3036,n3037);
xor (n3036,n2916,n2917);
and (n3037,n558,n348);
and (n3038,n3039,n3040);
xor (n3039,n3036,n3037);
or (n3040,n3041,n3044);
and (n3041,n3042,n3043);
xor (n3042,n2922,n2923);
and (n3043,n550,n348);
and (n3044,n3045,n3046);
xor (n3045,n3042,n3043);
or (n3046,n3047,n3050);
and (n3047,n3048,n3049);
xor (n3048,n2928,n2929);
and (n3049,n586,n348);
and (n3050,n3051,n3052);
xor (n3051,n3048,n3049);
or (n3052,n3053,n3056);
and (n3053,n3054,n3055);
xor (n3054,n2934,n2935);
and (n3055,n237,n348);
and (n3056,n3057,n3058);
xor (n3057,n3054,n3055);
or (n3058,n3059,n3062);
and (n3059,n3060,n3061);
xor (n3060,n2940,n2941);
and (n3061,n228,n348);
and (n3062,n3063,n3064);
xor (n3063,n3060,n3061);
or (n3064,n3065,n3068);
and (n3065,n3066,n3067);
xor (n3066,n2946,n2947);
and (n3067,n385,n348);
and (n3068,n3069,n3070);
xor (n3069,n3066,n3067);
or (n3070,n3071,n3074);
and (n3071,n3072,n3073);
xor (n3072,n2952,n2953);
and (n3073,n424,n348);
and (n3074,n3075,n3076);
xor (n3075,n3072,n3073);
or (n3076,n3077,n3080);
and (n3077,n3078,n3079);
xor (n3078,n2958,n2959);
and (n3079,n416,n348);
and (n3080,n3081,n3082);
xor (n3081,n3078,n3079);
and (n3082,n3083,n3084);
xor (n3083,n2964,n2965);
and (n3084,n457,n348);
and (n3085,n363,n487);
or (n3086,n3087,n3090);
and (n3087,n3088,n3089);
xor (n3088,n2973,n2974);
and (n3089,n355,n487);
and (n3090,n3091,n3092);
xor (n3091,n3088,n3089);
or (n3092,n3093,n3096);
and (n3093,n3094,n3095);
xor (n3094,n2979,n2980);
and (n3095,n497,n487);
and (n3096,n3097,n3098);
xor (n3097,n3094,n3095);
or (n3098,n3099,n3102);
and (n3099,n3100,n3101);
xor (n3100,n2985,n2986);
and (n3101,n568,n487);
and (n3102,n3103,n3104);
xor (n3103,n3100,n3101);
or (n3104,n3105,n3108);
and (n3105,n3106,n3107);
xor (n3106,n2991,n2992);
and (n3107,n275,n487);
and (n3108,n3109,n3110);
xor (n3109,n3106,n3107);
or (n3110,n3111,n3114);
and (n3111,n3112,n3113);
xor (n3112,n2997,n2998);
and (n3113,n264,n487);
and (n3114,n3115,n3116);
xor (n3115,n3112,n3113);
or (n3116,n3117,n3120);
and (n3117,n3118,n3119);
xor (n3118,n3003,n3004);
and (n3119,n140,n487);
and (n3120,n3121,n3122);
xor (n3121,n3118,n3119);
or (n3122,n3123,n3126);
and (n3123,n3124,n3125);
xor (n3124,n3009,n3010);
and (n3125,n93,n487);
and (n3126,n3127,n3128);
xor (n3127,n3124,n3125);
or (n3128,n3129,n3132);
and (n3129,n3130,n3131);
xor (n3130,n3015,n3016);
and (n3131,n182,n487);
and (n3132,n3133,n3134);
xor (n3133,n3130,n3131);
or (n3134,n3135,n3138);
and (n3135,n3136,n3137);
xor (n3136,n3021,n3022);
and (n3137,n173,n487);
and (n3138,n3139,n3140);
xor (n3139,n3136,n3137);
or (n3140,n3141,n3144);
and (n3141,n3142,n3143);
xor (n3142,n3027,n3028);
and (n3143,n375,n487);
and (n3144,n3145,n3146);
xor (n3145,n3142,n3143);
or (n3146,n3147,n3150);
and (n3147,n3148,n3149);
xor (n3148,n3033,n3034);
and (n3149,n558,n487);
and (n3150,n3151,n3152);
xor (n3151,n3148,n3149);
or (n3152,n3153,n3156);
and (n3153,n3154,n3155);
xor (n3154,n3039,n3040);
and (n3155,n550,n487);
and (n3156,n3157,n3158);
xor (n3157,n3154,n3155);
or (n3158,n3159,n3162);
and (n3159,n3160,n3161);
xor (n3160,n3045,n3046);
and (n3161,n586,n487);
and (n3162,n3163,n3164);
xor (n3163,n3160,n3161);
or (n3164,n3165,n3168);
and (n3165,n3166,n3167);
xor (n3166,n3051,n3052);
and (n3167,n237,n487);
and (n3168,n3169,n3170);
xor (n3169,n3166,n3167);
or (n3170,n3171,n3174);
and (n3171,n3172,n3173);
xor (n3172,n3057,n3058);
and (n3173,n228,n487);
and (n3174,n3175,n3176);
xor (n3175,n3172,n3173);
or (n3176,n3177,n3180);
and (n3177,n3178,n3179);
xor (n3178,n3063,n3064);
and (n3179,n385,n487);
and (n3180,n3181,n3182);
xor (n3181,n3178,n3179);
or (n3182,n3183,n3186);
and (n3183,n3184,n3185);
xor (n3184,n3069,n3070);
and (n3185,n424,n487);
and (n3186,n3187,n3188);
xor (n3187,n3184,n3185);
or (n3188,n3189,n3192);
and (n3189,n3190,n3191);
xor (n3190,n3075,n3076);
and (n3191,n416,n487);
and (n3192,n3193,n3194);
xor (n3193,n3190,n3191);
and (n3194,n3195,n1928);
xor (n3195,n3081,n3082);
and (n3196,n355,n257);
or (n3197,n3198,n3201);
and (n3198,n3199,n3200);
xor (n3199,n3091,n3092);
and (n3200,n497,n257);
and (n3201,n3202,n3203);
xor (n3202,n3199,n3200);
or (n3203,n3204,n3207);
and (n3204,n3205,n3206);
xor (n3205,n3097,n3098);
and (n3206,n568,n257);
and (n3207,n3208,n3209);
xor (n3208,n3205,n3206);
or (n3209,n3210,n3213);
and (n3210,n3211,n3212);
xor (n3211,n3103,n3104);
and (n3212,n275,n257);
and (n3213,n3214,n3215);
xor (n3214,n3211,n3212);
or (n3215,n3216,n3219);
and (n3216,n3217,n3218);
xor (n3217,n3109,n3110);
and (n3218,n264,n257);
and (n3219,n3220,n3221);
xor (n3220,n3217,n3218);
or (n3221,n3222,n3225);
and (n3222,n3223,n3224);
xor (n3223,n3115,n3116);
and (n3224,n140,n257);
and (n3225,n3226,n3227);
xor (n3226,n3223,n3224);
or (n3227,n3228,n3231);
and (n3228,n3229,n3230);
xor (n3229,n3121,n3122);
and (n3230,n93,n257);
and (n3231,n3232,n3233);
xor (n3232,n3229,n3230);
or (n3233,n3234,n3237);
and (n3234,n3235,n3236);
xor (n3235,n3127,n3128);
and (n3236,n182,n257);
and (n3237,n3238,n3239);
xor (n3238,n3235,n3236);
or (n3239,n3240,n3243);
and (n3240,n3241,n3242);
xor (n3241,n3133,n3134);
and (n3242,n173,n257);
and (n3243,n3244,n3245);
xor (n3244,n3241,n3242);
or (n3245,n3246,n3249);
and (n3246,n3247,n3248);
xor (n3247,n3139,n3140);
and (n3248,n375,n257);
and (n3249,n3250,n3251);
xor (n3250,n3247,n3248);
or (n3251,n3252,n3255);
and (n3252,n3253,n3254);
xor (n3253,n3145,n3146);
and (n3254,n558,n257);
and (n3255,n3256,n3257);
xor (n3256,n3253,n3254);
or (n3257,n3258,n3261);
and (n3258,n3259,n3260);
xor (n3259,n3151,n3152);
and (n3260,n550,n257);
and (n3261,n3262,n3263);
xor (n3262,n3259,n3260);
or (n3263,n3264,n3267);
and (n3264,n3265,n3266);
xor (n3265,n3157,n3158);
and (n3266,n586,n257);
and (n3267,n3268,n3269);
xor (n3268,n3265,n3266);
or (n3269,n3270,n3273);
and (n3270,n3271,n3272);
xor (n3271,n3163,n3164);
and (n3272,n237,n257);
and (n3273,n3274,n3275);
xor (n3274,n3271,n3272);
or (n3275,n3276,n3279);
and (n3276,n3277,n3278);
xor (n3277,n3169,n3170);
and (n3278,n228,n257);
and (n3279,n3280,n3281);
xor (n3280,n3277,n3278);
or (n3281,n3282,n3284);
and (n3282,n3283,n1792);
xor (n3283,n3175,n3176);
and (n3284,n3285,n3286);
xor (n3285,n3283,n1792);
or (n3286,n3287,n3290);
and (n3287,n3288,n3289);
xor (n3288,n3181,n3182);
and (n3289,n424,n257);
and (n3290,n3291,n3292);
xor (n3291,n3288,n3289);
or (n3292,n3293,n3296);
and (n3293,n3294,n3295);
xor (n3294,n3187,n3188);
and (n3295,n416,n257);
and (n3296,n3297,n3298);
xor (n3297,n3294,n3295);
and (n3298,n3299,n3300);
xor (n3299,n3193,n3194);
and (n3300,n457,n257);
and (n3301,n497,n249);
or (n3302,n3303,n3306);
and (n3303,n3304,n3305);
xor (n3304,n3202,n3203);
and (n3305,n568,n249);
and (n3306,n3307,n3308);
xor (n3307,n3304,n3305);
or (n3308,n3309,n3312);
and (n3309,n3310,n3311);
xor (n3310,n3208,n3209);
and (n3311,n275,n249);
and (n3312,n3313,n3314);
xor (n3313,n3310,n3311);
or (n3314,n3315,n3318);
and (n3315,n3316,n3317);
xor (n3316,n3214,n3215);
and (n3317,n264,n249);
and (n3318,n3319,n3320);
xor (n3319,n3316,n3317);
or (n3320,n3321,n3324);
and (n3321,n3322,n3323);
xor (n3322,n3220,n3221);
and (n3323,n140,n249);
and (n3324,n3325,n3326);
xor (n3325,n3322,n3323);
or (n3326,n3327,n3330);
and (n3327,n3328,n3329);
xor (n3328,n3226,n3227);
and (n3329,n93,n249);
and (n3330,n3331,n3332);
xor (n3331,n3328,n3329);
or (n3332,n3333,n3336);
and (n3333,n3334,n3335);
xor (n3334,n3232,n3233);
and (n3335,n182,n249);
and (n3336,n3337,n3338);
xor (n3337,n3334,n3335);
or (n3338,n3339,n3342);
and (n3339,n3340,n3341);
xor (n3340,n3238,n3239);
and (n3341,n173,n249);
and (n3342,n3343,n3344);
xor (n3343,n3340,n3341);
or (n3344,n3345,n3348);
and (n3345,n3346,n3347);
xor (n3346,n3244,n3245);
and (n3347,n375,n249);
and (n3348,n3349,n3350);
xor (n3349,n3346,n3347);
or (n3350,n3351,n3354);
and (n3351,n3352,n3353);
xor (n3352,n3250,n3251);
and (n3353,n558,n249);
and (n3354,n3355,n3356);
xor (n3355,n3352,n3353);
or (n3356,n3357,n3360);
and (n3357,n3358,n3359);
xor (n3358,n3256,n3257);
and (n3359,n550,n249);
and (n3360,n3361,n3362);
xor (n3361,n3358,n3359);
or (n3362,n3363,n3366);
and (n3363,n3364,n3365);
xor (n3364,n3262,n3263);
and (n3365,n586,n249);
and (n3366,n3367,n3368);
xor (n3367,n3364,n3365);
or (n3368,n3369,n3372);
and (n3369,n3370,n3371);
xor (n3370,n3268,n3269);
and (n3371,n237,n249);
and (n3372,n3373,n3374);
xor (n3373,n3370,n3371);
or (n3374,n3375,n3378);
and (n3375,n3376,n3377);
xor (n3376,n3274,n3275);
and (n3377,n228,n249);
and (n3378,n3379,n3380);
xor (n3379,n3376,n3377);
or (n3380,n3381,n3384);
and (n3381,n3382,n3383);
xor (n3382,n3280,n3281);
and (n3383,n385,n249);
and (n3384,n3385,n3386);
xor (n3385,n3382,n3383);
or (n3386,n3387,n3390);
and (n3387,n3388,n3389);
xor (n3388,n3285,n3286);
and (n3389,n424,n249);
and (n3390,n3391,n3392);
xor (n3391,n3388,n3389);
or (n3392,n3393,n3396);
and (n3393,n3394,n3395);
xor (n3394,n3291,n3292);
and (n3395,n416,n249);
and (n3396,n3397,n3398);
xor (n3397,n3394,n3395);
and (n3398,n3399,n1821);
xor (n3399,n3297,n3298);
and (n3400,n568,n75);
or (n3401,n3402,n3405);
and (n3402,n3403,n3404);
xor (n3403,n3307,n3308);
and (n3404,n275,n75);
and (n3405,n3406,n3407);
xor (n3406,n3403,n3404);
or (n3407,n3408,n3411);
and (n3408,n3409,n3410);
xor (n3409,n3313,n3314);
and (n3410,n264,n75);
and (n3411,n3412,n3413);
xor (n3412,n3409,n3410);
or (n3413,n3414,n3417);
and (n3414,n3415,n3416);
xor (n3415,n3319,n3320);
and (n3416,n140,n75);
and (n3417,n3418,n3419);
xor (n3418,n3415,n3416);
or (n3419,n3420,n3423);
and (n3420,n3421,n3422);
xor (n3421,n3325,n3326);
and (n3422,n93,n75);
and (n3423,n3424,n3425);
xor (n3424,n3421,n3422);
or (n3425,n3426,n3429);
and (n3426,n3427,n3428);
xor (n3427,n3331,n3332);
and (n3428,n182,n75);
and (n3429,n3430,n3431);
xor (n3430,n3427,n3428);
or (n3431,n3432,n3435);
and (n3432,n3433,n3434);
xor (n3433,n3337,n3338);
and (n3434,n173,n75);
and (n3435,n3436,n3437);
xor (n3436,n3433,n3434);
or (n3437,n3438,n3441);
and (n3438,n3439,n3440);
xor (n3439,n3343,n3344);
and (n3440,n375,n75);
and (n3441,n3442,n3443);
xor (n3442,n3439,n3440);
or (n3443,n3444,n3447);
and (n3444,n3445,n3446);
xor (n3445,n3349,n3350);
and (n3446,n558,n75);
and (n3447,n3448,n3449);
xor (n3448,n3445,n3446);
or (n3449,n3450,n3453);
and (n3450,n3451,n3452);
xor (n3451,n3355,n3356);
and (n3452,n550,n75);
and (n3453,n3454,n3455);
xor (n3454,n3451,n3452);
or (n3455,n3456,n3459);
and (n3456,n3457,n3458);
xor (n3457,n3361,n3362);
and (n3458,n586,n75);
and (n3459,n3460,n3461);
xor (n3460,n3457,n3458);
or (n3461,n3462,n3465);
and (n3462,n3463,n3464);
xor (n3463,n3367,n3368);
and (n3464,n237,n75);
and (n3465,n3466,n3467);
xor (n3466,n3463,n3464);
or (n3467,n3468,n3471);
and (n3468,n3469,n3470);
xor (n3469,n3373,n3374);
and (n3470,n228,n75);
and (n3471,n3472,n3473);
xor (n3472,n3469,n3470);
or (n3473,n3474,n3477);
and (n3474,n3475,n3476);
xor (n3475,n3379,n3380);
and (n3476,n385,n75);
and (n3477,n3478,n3479);
xor (n3478,n3475,n3476);
or (n3479,n3480,n3483);
and (n3480,n3481,n3482);
xor (n3481,n3385,n3386);
and (n3482,n424,n75);
and (n3483,n3484,n3485);
xor (n3484,n3481,n3482);
or (n3485,n3486,n3489);
and (n3486,n3487,n3488);
xor (n3487,n3391,n3392);
and (n3488,n416,n75);
and (n3489,n3490,n3491);
xor (n3490,n3487,n3488);
and (n3491,n3492,n3493);
xor (n3492,n3397,n3398);
and (n3493,n457,n75);
and (n3494,n275,n21);
or (n3495,n3496,n3499);
and (n3496,n3497,n3498);
xor (n3497,n3406,n3407);
and (n3498,n264,n21);
and (n3499,n3500,n3501);
xor (n3500,n3497,n3498);
or (n3501,n3502,n3505);
and (n3502,n3503,n3504);
xor (n3503,n3412,n3413);
and (n3504,n140,n21);
and (n3505,n3506,n3507);
xor (n3506,n3503,n3504);
or (n3507,n3508,n3511);
and (n3508,n3509,n3510);
xor (n3509,n3418,n3419);
and (n3510,n93,n21);
and (n3511,n3512,n3513);
xor (n3512,n3509,n3510);
or (n3513,n3514,n3517);
and (n3514,n3515,n3516);
xor (n3515,n3424,n3425);
and (n3516,n182,n21);
and (n3517,n3518,n3519);
xor (n3518,n3515,n3516);
or (n3519,n3520,n3523);
and (n3520,n3521,n3522);
xor (n3521,n3430,n3431);
and (n3522,n173,n21);
and (n3523,n3524,n3525);
xor (n3524,n3521,n3522);
or (n3525,n3526,n3529);
and (n3526,n3527,n3528);
xor (n3527,n3436,n3437);
and (n3528,n375,n21);
and (n3529,n3530,n3531);
xor (n3530,n3527,n3528);
or (n3531,n3532,n3535);
and (n3532,n3533,n3534);
xor (n3533,n3442,n3443);
and (n3534,n558,n21);
and (n3535,n3536,n3537);
xor (n3536,n3533,n3534);
or (n3537,n3538,n3541);
and (n3538,n3539,n3540);
xor (n3539,n3448,n3449);
and (n3540,n550,n21);
and (n3541,n3542,n3543);
xor (n3542,n3539,n3540);
or (n3543,n3544,n3547);
and (n3544,n3545,n3546);
xor (n3545,n3454,n3455);
and (n3546,n586,n21);
and (n3547,n3548,n3549);
xor (n3548,n3545,n3546);
or (n3549,n3550,n3553);
and (n3550,n3551,n3552);
xor (n3551,n3460,n3461);
and (n3552,n237,n21);
and (n3553,n3554,n3555);
xor (n3554,n3551,n3552);
or (n3555,n3556,n3559);
and (n3556,n3557,n3558);
xor (n3557,n3466,n3467);
and (n3558,n228,n21);
and (n3559,n3560,n3561);
xor (n3560,n3557,n3558);
or (n3561,n3562,n3565);
and (n3562,n3563,n3564);
xor (n3563,n3472,n3473);
and (n3564,n385,n21);
and (n3565,n3566,n3567);
xor (n3566,n3563,n3564);
or (n3567,n3568,n3571);
and (n3568,n3569,n3570);
xor (n3569,n3478,n3479);
and (n3570,n424,n21);
and (n3571,n3572,n3573);
xor (n3572,n3569,n3570);
or (n3573,n3574,n3577);
and (n3574,n3575,n3576);
xor (n3575,n3484,n3485);
and (n3576,n416,n21);
and (n3577,n3578,n3579);
xor (n3578,n3575,n3576);
and (n3579,n3580,n1630);
xor (n3580,n3490,n3491);
and (n3581,n264,n83);
or (n3582,n3583,n3586);
and (n3583,n3584,n3585);
xor (n3584,n3500,n3501);
and (n3585,n140,n83);
and (n3586,n3587,n3588);
xor (n3587,n3584,n3585);
or (n3588,n3589,n3592);
and (n3589,n3590,n3591);
xor (n3590,n3506,n3507);
and (n3591,n93,n83);
and (n3592,n3593,n3594);
xor (n3593,n3590,n3591);
or (n3594,n3595,n3598);
and (n3595,n3596,n3597);
xor (n3596,n3512,n3513);
and (n3597,n182,n83);
and (n3598,n3599,n3600);
xor (n3599,n3596,n3597);
or (n3600,n3601,n3604);
and (n3601,n3602,n3603);
xor (n3602,n3518,n3519);
and (n3603,n173,n83);
and (n3604,n3605,n3606);
xor (n3605,n3602,n3603);
or (n3606,n3607,n3610);
and (n3607,n3608,n3609);
xor (n3608,n3524,n3525);
and (n3609,n375,n83);
and (n3610,n3611,n3612);
xor (n3611,n3608,n3609);
or (n3612,n3613,n3616);
and (n3613,n3614,n3615);
xor (n3614,n3530,n3531);
and (n3615,n558,n83);
and (n3616,n3617,n3618);
xor (n3617,n3614,n3615);
or (n3618,n3619,n3622);
and (n3619,n3620,n3621);
xor (n3620,n3536,n3537);
and (n3621,n550,n83);
and (n3622,n3623,n3624);
xor (n3623,n3620,n3621);
or (n3624,n3625,n3628);
and (n3625,n3626,n3627);
xor (n3626,n3542,n3543);
and (n3627,n586,n83);
and (n3628,n3629,n3630);
xor (n3629,n3626,n3627);
or (n3630,n3631,n3634);
and (n3631,n3632,n3633);
xor (n3632,n3548,n3549);
and (n3633,n237,n83);
and (n3634,n3635,n3636);
xor (n3635,n3632,n3633);
or (n3636,n3637,n3640);
and (n3637,n3638,n3639);
xor (n3638,n3554,n3555);
and (n3639,n228,n83);
and (n3640,n3641,n3642);
xor (n3641,n3638,n3639);
or (n3642,n3643,n3646);
and (n3643,n3644,n3645);
xor (n3644,n3560,n3561);
and (n3645,n385,n83);
and (n3646,n3647,n3648);
xor (n3647,n3644,n3645);
or (n3648,n3649,n3652);
and (n3649,n3650,n3651);
xor (n3650,n3566,n3567);
and (n3651,n424,n83);
and (n3652,n3653,n3654);
xor (n3653,n3650,n3651);
or (n3654,n3655,n3658);
and (n3655,n3656,n3657);
xor (n3656,n3572,n3573);
and (n3657,n416,n83);
and (n3658,n3659,n3660);
xor (n3659,n3656,n3657);
and (n3660,n3661,n3662);
xor (n3661,n3578,n3579);
and (n3662,n457,n83);
and (n3663,n140,n163);
or (n3664,n3665,n3668);
and (n3665,n3666,n3667);
xor (n3666,n3587,n3588);
and (n3667,n93,n163);
and (n3668,n3669,n3670);
xor (n3669,n3666,n3667);
or (n3670,n3671,n3674);
and (n3671,n3672,n3673);
xor (n3672,n3593,n3594);
and (n3673,n182,n163);
and (n3674,n3675,n3676);
xor (n3675,n3672,n3673);
or (n3676,n3677,n3680);
and (n3677,n3678,n3679);
xor (n3678,n3599,n3600);
and (n3679,n173,n163);
and (n3680,n3681,n3682);
xor (n3681,n3678,n3679);
or (n3682,n3683,n3686);
and (n3683,n3684,n3685);
xor (n3684,n3605,n3606);
and (n3685,n375,n163);
and (n3686,n3687,n3688);
xor (n3687,n3684,n3685);
or (n3688,n3689,n3692);
and (n3689,n3690,n3691);
xor (n3690,n3611,n3612);
and (n3691,n558,n163);
and (n3692,n3693,n3694);
xor (n3693,n3690,n3691);
or (n3694,n3695,n3698);
and (n3695,n3696,n3697);
xor (n3696,n3617,n3618);
and (n3697,n550,n163);
and (n3698,n3699,n3700);
xor (n3699,n3696,n3697);
or (n3700,n3701,n3704);
and (n3701,n3702,n3703);
xor (n3702,n3623,n3624);
and (n3703,n586,n163);
and (n3704,n3705,n3706);
xor (n3705,n3702,n3703);
or (n3706,n3707,n3710);
and (n3707,n3708,n3709);
xor (n3708,n3629,n3630);
and (n3709,n237,n163);
and (n3710,n3711,n3712);
xor (n3711,n3708,n3709);
or (n3712,n3713,n3716);
and (n3713,n3714,n3715);
xor (n3714,n3635,n3636);
and (n3715,n228,n163);
and (n3716,n3717,n3718);
xor (n3717,n3714,n3715);
or (n3718,n3719,n3722);
and (n3719,n3720,n3721);
xor (n3720,n3641,n3642);
and (n3721,n385,n163);
and (n3722,n3723,n3724);
xor (n3723,n3720,n3721);
or (n3724,n3725,n3728);
and (n3725,n3726,n3727);
xor (n3726,n3647,n3648);
and (n3727,n424,n163);
and (n3728,n3729,n3730);
xor (n3729,n3726,n3727);
or (n3730,n3731,n3734);
and (n3731,n3732,n3733);
xor (n3732,n3653,n3654);
and (n3733,n416,n163);
and (n3734,n3735,n3736);
xor (n3735,n3732,n3733);
and (n3736,n3737,n1539);
xor (n3737,n3659,n3660);
and (n3738,n93,n154);
or (n3739,n3740,n3743);
and (n3740,n3741,n3742);
xor (n3741,n3669,n3670);
and (n3742,n182,n154);
and (n3743,n3744,n3745);
xor (n3744,n3741,n3742);
or (n3745,n3746,n3749);
and (n3746,n3747,n3748);
xor (n3747,n3675,n3676);
and (n3748,n173,n154);
and (n3749,n3750,n3751);
xor (n3750,n3747,n3748);
or (n3751,n3752,n3755);
and (n3752,n3753,n3754);
xor (n3753,n3681,n3682);
and (n3754,n375,n154);
and (n3755,n3756,n3757);
xor (n3756,n3753,n3754);
or (n3757,n3758,n3761);
and (n3758,n3759,n3760);
xor (n3759,n3687,n3688);
and (n3760,n558,n154);
and (n3761,n3762,n3763);
xor (n3762,n3759,n3760);
or (n3763,n3764,n3767);
and (n3764,n3765,n3766);
xor (n3765,n3693,n3694);
and (n3766,n550,n154);
and (n3767,n3768,n3769);
xor (n3768,n3765,n3766);
or (n3769,n3770,n3773);
and (n3770,n3771,n3772);
xor (n3771,n3699,n3700);
and (n3772,n586,n154);
and (n3773,n3774,n3775);
xor (n3774,n3771,n3772);
or (n3775,n3776,n3779);
and (n3776,n3777,n3778);
xor (n3777,n3705,n3706);
and (n3778,n237,n154);
and (n3779,n3780,n3781);
xor (n3780,n3777,n3778);
or (n3781,n3782,n3785);
and (n3782,n3783,n3784);
xor (n3783,n3711,n3712);
and (n3784,n228,n154);
and (n3785,n3786,n3787);
xor (n3786,n3783,n3784);
or (n3787,n3788,n3791);
and (n3788,n3789,n3790);
xor (n3789,n3717,n3718);
and (n3790,n385,n154);
and (n3791,n3792,n3793);
xor (n3792,n3789,n3790);
or (n3793,n3794,n3797);
and (n3794,n3795,n3796);
xor (n3795,n3723,n3724);
and (n3796,n424,n154);
and (n3797,n3798,n3799);
xor (n3798,n3795,n3796);
or (n3799,n3800,n3803);
and (n3800,n3801,n3802);
xor (n3801,n3729,n3730);
and (n3802,n416,n154);
and (n3803,n3804,n3805);
xor (n3804,n3801,n3802);
and (n3805,n3806,n3807);
xor (n3806,n3735,n3736);
and (n3807,n457,n154);
and (n3808,n182,n514);
or (n3809,n3810,n3813);
and (n3810,n3811,n3812);
xor (n3811,n3744,n3745);
and (n3812,n173,n514);
and (n3813,n3814,n3815);
xor (n3814,n3811,n3812);
or (n3815,n3816,n3819);
and (n3816,n3817,n3818);
xor (n3817,n3750,n3751);
and (n3818,n375,n514);
and (n3819,n3820,n3821);
xor (n3820,n3817,n3818);
or (n3821,n3822,n3825);
and (n3822,n3823,n3824);
xor (n3823,n3756,n3757);
and (n3824,n558,n514);
and (n3825,n3826,n3827);
xor (n3826,n3823,n3824);
or (n3827,n3828,n3831);
and (n3828,n3829,n3830);
xor (n3829,n3762,n3763);
and (n3830,n550,n514);
and (n3831,n3832,n3833);
xor (n3832,n3829,n3830);
or (n3833,n3834,n3837);
and (n3834,n3835,n3836);
xor (n3835,n3768,n3769);
and (n3836,n586,n514);
and (n3837,n3838,n3839);
xor (n3838,n3835,n3836);
or (n3839,n3840,n3843);
and (n3840,n3841,n3842);
xor (n3841,n3774,n3775);
and (n3842,n237,n514);
and (n3843,n3844,n3845);
xor (n3844,n3841,n3842);
or (n3845,n3846,n3849);
and (n3846,n3847,n3848);
xor (n3847,n3780,n3781);
and (n3848,n228,n514);
and (n3849,n3850,n3851);
xor (n3850,n3847,n3848);
or (n3851,n3852,n3855);
and (n3852,n3853,n3854);
xor (n3853,n3786,n3787);
and (n3854,n385,n514);
and (n3855,n3856,n3857);
xor (n3856,n3853,n3854);
or (n3857,n3858,n3861);
and (n3858,n3859,n3860);
xor (n3859,n3792,n3793);
and (n3860,n424,n514);
and (n3861,n3862,n3863);
xor (n3862,n3859,n3860);
or (n3863,n3864,n3867);
and (n3864,n3865,n3866);
xor (n3865,n3798,n3799);
and (n3866,n416,n514);
and (n3867,n3868,n3869);
xor (n3868,n3865,n3866);
and (n3869,n3870,n1738);
xor (n3870,n3804,n3805);
and (n3871,n173,n521);
or (n3872,n3873,n3876);
and (n3873,n3874,n3875);
xor (n3874,n3814,n3815);
and (n3875,n375,n521);
and (n3876,n3877,n3878);
xor (n3877,n3874,n3875);
or (n3878,n3879,n3882);
and (n3879,n3880,n3881);
xor (n3880,n3820,n3821);
and (n3881,n558,n521);
and (n3882,n3883,n3884);
xor (n3883,n3880,n3881);
or (n3884,n3885,n3888);
and (n3885,n3886,n3887);
xor (n3886,n3826,n3827);
and (n3887,n550,n521);
and (n3888,n3889,n3890);
xor (n3889,n3886,n3887);
or (n3890,n3891,n3894);
and (n3891,n3892,n3893);
xor (n3892,n3832,n3833);
and (n3893,n586,n521);
and (n3894,n3895,n3896);
xor (n3895,n3892,n3893);
or (n3896,n3897,n3900);
and (n3897,n3898,n3899);
xor (n3898,n3838,n3839);
and (n3899,n237,n521);
and (n3900,n3901,n3902);
xor (n3901,n3898,n3899);
or (n3902,n3903,n3906);
and (n3903,n3904,n3905);
xor (n3904,n3844,n3845);
and (n3905,n228,n521);
and (n3906,n3907,n3908);
xor (n3907,n3904,n3905);
or (n3908,n3909,n3912);
and (n3909,n3910,n3911);
xor (n3910,n3850,n3851);
and (n3911,n385,n521);
and (n3912,n3913,n3914);
xor (n3913,n3910,n3911);
or (n3914,n3915,n3918);
and (n3915,n3916,n3917);
xor (n3916,n3856,n3857);
and (n3917,n424,n521);
and (n3918,n3919,n3920);
xor (n3919,n3916,n3917);
or (n3920,n3921,n3924);
and (n3921,n3922,n3923);
xor (n3922,n3862,n3863);
and (n3923,n416,n521);
and (n3924,n3925,n3926);
xor (n3925,n3922,n3923);
and (n3926,n3927,n3928);
xor (n3927,n3868,n3869);
and (n3928,n457,n521);
and (n3929,n375,n541);
or (n3930,n3931,n3934);
and (n3931,n3932,n3933);
xor (n3932,n3877,n3878);
and (n3933,n558,n541);
and (n3934,n3935,n3936);
xor (n3935,n3932,n3933);
or (n3936,n3937,n3940);
and (n3937,n3938,n3939);
xor (n3938,n3883,n3884);
and (n3939,n550,n541);
and (n3940,n3941,n3942);
xor (n3941,n3938,n3939);
or (n3942,n3943,n3946);
and (n3943,n3944,n3945);
xor (n3944,n3889,n3890);
and (n3945,n586,n541);
and (n3946,n3947,n3948);
xor (n3947,n3944,n3945);
or (n3948,n3949,n3952);
and (n3949,n3950,n3951);
xor (n3950,n3895,n3896);
and (n3951,n237,n541);
and (n3952,n3953,n3954);
xor (n3953,n3950,n3951);
or (n3954,n3955,n3958);
and (n3955,n3956,n3957);
xor (n3956,n3901,n3902);
and (n3957,n228,n541);
and (n3958,n3959,n3960);
xor (n3959,n3956,n3957);
or (n3960,n3961,n3964);
and (n3961,n3962,n3963);
xor (n3962,n3907,n3908);
and (n3963,n385,n541);
and (n3964,n3965,n3966);
xor (n3965,n3962,n3963);
or (n3966,n3967,n3970);
and (n3967,n3968,n3969);
xor (n3968,n3913,n3914);
and (n3969,n424,n541);
and (n3970,n3971,n3972);
xor (n3971,n3968,n3969);
or (n3972,n3973,n3976);
and (n3973,n3974,n3975);
xor (n3974,n3919,n3920);
and (n3975,n416,n541);
and (n3976,n3977,n3978);
xor (n3977,n3974,n3975);
and (n3978,n3979,n1367);
xor (n3979,n3925,n3926);
and (n3980,n558,n210);
or (n3981,n3982,n3985);
and (n3982,n3983,n3984);
xor (n3983,n3935,n3936);
and (n3984,n550,n210);
and (n3985,n3986,n3987);
xor (n3986,n3983,n3984);
or (n3987,n3988,n3991);
and (n3988,n3989,n3990);
xor (n3989,n3941,n3942);
and (n3990,n586,n210);
and (n3991,n3992,n3993);
xor (n3992,n3989,n3990);
or (n3993,n3994,n3997);
and (n3994,n3995,n3996);
xor (n3995,n3947,n3948);
and (n3996,n237,n210);
and (n3997,n3998,n3999);
xor (n3998,n3995,n3996);
or (n3999,n4000,n4003);
and (n4000,n4001,n4002);
xor (n4001,n3953,n3954);
and (n4002,n228,n210);
and (n4003,n4004,n4005);
xor (n4004,n4001,n4002);
or (n4005,n4006,n4009);
and (n4006,n4007,n4008);
xor (n4007,n3959,n3960);
and (n4008,n385,n210);
and (n4009,n4010,n4011);
xor (n4010,n4007,n4008);
or (n4011,n4012,n4015);
and (n4012,n4013,n4014);
xor (n4013,n3965,n3966);
and (n4014,n424,n210);
and (n4015,n4016,n4017);
xor (n4016,n4013,n4014);
or (n4017,n4018,n4021);
and (n4018,n4019,n4020);
xor (n4019,n3971,n3972);
and (n4020,n416,n210);
and (n4021,n4022,n4023);
xor (n4022,n4019,n4020);
and (n4023,n4024,n4025);
xor (n4024,n3977,n3978);
and (n4025,n457,n210);
and (n4026,n550,n192);
or (n4027,n4028,n4031);
and (n4028,n4029,n4030);
xor (n4029,n3986,n3987);
and (n4030,n586,n192);
and (n4031,n4032,n4033);
xor (n4032,n4029,n4030);
or (n4033,n4034,n4037);
and (n4034,n4035,n4036);
xor (n4035,n3992,n3993);
and (n4036,n237,n192);
and (n4037,n4038,n4039);
xor (n4038,n4035,n4036);
or (n4039,n4040,n4043);
and (n4040,n4041,n4042);
xor (n4041,n3998,n3999);
and (n4042,n228,n192);
and (n4043,n4044,n4045);
xor (n4044,n4041,n4042);
or (n4045,n4046,n4049);
and (n4046,n4047,n4048);
xor (n4047,n4004,n4005);
and (n4048,n385,n192);
and (n4049,n4050,n4051);
xor (n4050,n4047,n4048);
or (n4051,n4052,n4055);
and (n4052,n4053,n4054);
xor (n4053,n4010,n4011);
and (n4054,n424,n192);
and (n4055,n4056,n4057);
xor (n4056,n4053,n4054);
or (n4057,n4058,n4061);
and (n4058,n4059,n4060);
xor (n4059,n4016,n4017);
and (n4060,n416,n192);
and (n4061,n4062,n4063);
xor (n4062,n4059,n4060);
and (n4063,n4064,n997);
xor (n4064,n4022,n4023);
and (n4065,n586,n219);
or (n4066,n4067,n4070);
and (n4067,n4068,n4069);
xor (n4068,n4032,n4033);
and (n4069,n237,n219);
and (n4070,n4071,n4072);
xor (n4071,n4068,n4069);
or (n4072,n4073,n4076);
and (n4073,n4074,n4075);
xor (n4074,n4038,n4039);
and (n4075,n228,n219);
and (n4076,n4077,n4078);
xor (n4077,n4074,n4075);
or (n4078,n4079,n4082);
and (n4079,n4080,n4081);
xor (n4080,n4044,n4045);
and (n4081,n385,n219);
and (n4082,n4083,n4084);
xor (n4083,n4080,n4081);
or (n4084,n4085,n4088);
and (n4085,n4086,n4087);
xor (n4086,n4050,n4051);
and (n4087,n424,n219);
and (n4088,n4089,n4090);
xor (n4089,n4086,n4087);
or (n4090,n4091,n4094);
and (n4091,n4092,n4093);
xor (n4092,n4056,n4057);
and (n4093,n416,n219);
and (n4094,n4095,n4096);
xor (n4095,n4092,n4093);
and (n4096,n4097,n4098);
xor (n4097,n4062,n4063);
and (n4098,n457,n219);
and (n4099,n237,n396);
or (n4100,n4101,n4104);
and (n4101,n4102,n4103);
xor (n4102,n4071,n4072);
and (n4103,n228,n396);
and (n4104,n4105,n4106);
xor (n4105,n4102,n4103);
or (n4106,n4107,n4110);
and (n4107,n4108,n4109);
xor (n4108,n4077,n4078);
and (n4109,n385,n396);
and (n4110,n4111,n4112);
xor (n4111,n4108,n4109);
or (n4112,n4113,n4116);
and (n4113,n4114,n4115);
xor (n4114,n4083,n4084);
and (n4115,n424,n396);
and (n4116,n4117,n4118);
xor (n4117,n4114,n4115);
or (n4118,n4119,n4122);
and (n4119,n4120,n4121);
xor (n4120,n4089,n4090);
and (n4121,n416,n396);
and (n4122,n4123,n4124);
xor (n4123,n4120,n4121);
and (n4124,n4125,n711);
xor (n4125,n4095,n4096);
and (n4126,n228,n406);
or (n4127,n4128,n4131);
and (n4128,n4129,n4130);
xor (n4129,n4105,n4106);
and (n4130,n385,n406);
and (n4131,n4132,n4133);
xor (n4132,n4129,n4130);
or (n4133,n4134,n4137);
and (n4134,n4135,n4136);
xor (n4135,n4111,n4112);
and (n4136,n424,n406);
and (n4137,n4138,n4139);
xor (n4138,n4135,n4136);
or (n4139,n4140,n4143);
and (n4140,n4141,n4142);
xor (n4141,n4117,n4118);
and (n4142,n416,n406);
and (n4143,n4144,n4145);
xor (n4144,n4141,n4142);
and (n4145,n4146,n4147);
xor (n4146,n4123,n4124);
and (n4147,n457,n406);
and (n4148,n385,n676);
or (n4149,n4150,n4153);
and (n4150,n4151,n4152);
xor (n4151,n4132,n4133);
and (n4152,n424,n676);
and (n4153,n4154,n4155);
xor (n4154,n4151,n4152);
or (n4155,n4156,n4159);
and (n4156,n4157,n4158);
xor (n4157,n4138,n4139);
and (n4158,n416,n676);
and (n4159,n4160,n4161);
xor (n4160,n4157,n4158);
and (n4161,n4162,n695);
xor (n4162,n4144,n4145);
and (n4163,n424,n451);
or (n4164,n4165,n4168);
and (n4165,n4166,n4167);
xor (n4166,n4154,n4155);
and (n4167,n416,n451);
and (n4168,n4169,n4170);
xor (n4169,n4166,n4167);
and (n4170,n4171,n4172);
xor (n4171,n4160,n4161);
and (n4172,n457,n451);
and (n4173,n416,n439);
and (n4174,n4175,n1154);
xor (n4175,n4169,n4170);
and (n4176,n457,n1081);
endmodule
