module top (out,n17,n20,n21,n22,n30,n31,n37,n38,n43
        ,n51,n53,n54,n63,n64,n74,n89,n90,n93,n99
        ,n121,n122,n129,n237,n238,n246,n303,n309);
output out;
input n17;
input n20;
input n21;
input n22;
input n30;
input n31;
input n37;
input n38;
input n43;
input n51;
input n53;
input n54;
input n63;
input n64;
input n74;
input n89;
input n90;
input n93;
input n99;
input n121;
input n122;
input n129;
input n237;
input n238;
input n246;
input n303;
input n309;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n18;
wire n19;
wire n23;
wire n24;
wire n25;
wire n26;
wire n27;
wire n28;
wire n29;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n39;
wire n40;
wire n41;
wire n42;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n52;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n91;
wire n92;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n302;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
xor (out,n0,n339);
nand (n0,n1,n338);
or (n1,n2,n285);
not (n2,n3);
nor (n3,n4,n283);
and (n4,n5,n226);
or (n5,n6,n225);
and (n6,n7,n141);
xor (n7,n8,n104);
or (n8,n9,n103);
and (n9,n10,n77);
xor (n10,n11,n46);
nand (n11,n12,n40);
or (n12,n13,n24);
not (n13,n14);
nor (n14,n15,n23);
and (n15,n16,n18);
not (n16,n17);
not (n18,n19);
wire s0n19,s1n19,notn19;
or (n19,s0n19,s1n19);
not(notn19,n22);
and (s0n19,notn19,n20);
and (s1n19,n22,n21);
and (n23,n17,n19);
not (n24,n25);
and (n25,n26,n33);
nand (n26,n27,n32);
or (n27,n28,n19);
not (n28,n29);
wire s0n29,s1n29,notn29;
or (n29,s0n29,s1n29);
not(notn29,n22);
and (s0n29,notn29,n30);
and (s1n29,n22,n31);
nand (n32,n19,n28);
not (n33,n34);
nand (n34,n35,n39);
or (n35,n28,n36);
wire s0n36,s1n36,notn36;
or (n36,s0n36,s1n36);
not(notn36,n22);
and (s0n36,notn36,n37);
and (s1n36,n22,n38);
nand (n39,n36,n28);
nand (n40,n34,n41);
nor (n41,n42,n44);
and (n42,n43,n19);
and (n44,n18,n45);
not (n45,n43);
nand (n46,n47,n66);
or (n47,n48,n58);
not (n48,n49);
nor (n49,n50,n55);
and (n50,n51,n52);
wire s0n52,s1n52,notn52;
or (n52,s0n52,s1n52);
not(notn52,n22);
and (s0n52,notn52,n53);
and (s1n52,n22,n54);
and (n55,n56,n57);
not (n56,n51);
not (n57,n52);
not (n58,n59);
nand (n59,n60,n65);
or (n60,n61,n19);
not (n61,n62);
wire s0n62,s1n62,notn62;
or (n62,s0n62,s1n62);
not(notn62,n22);
and (s0n62,notn62,n63);
and (s1n62,n22,n64);
nand (n65,n19,n61);
nand (n66,n67,n72);
not (n67,n68);
nand (n68,n58,n69);
nand (n69,n70,n71);
or (n70,n61,n52);
nand (n71,n52,n61);
nand (n72,n73,n75);
or (n73,n57,n74);
or (n75,n52,n76);
not (n76,n74);
xor (n77,n78,n83);
and (n78,n79,n52);
nand (n79,n80,n82);
or (n80,n19,n81);
and (n81,n74,n62);
or (n82,n62,n74);
nand (n83,n84,n96);
or (n84,n85,n91);
not (n85,n86);
nor (n86,n87,n88);
not (n87,n36);
wire s0n88,s1n88,notn88;
or (n88,s0n88,s1n88);
not(notn88,n22);
and (s0n88,notn88,n89);
and (s1n88,n22,n90);
nor (n91,n92,n94);
and (n92,n87,n93);
and (n94,n36,n95);
not (n95,n93);
or (n96,n97,n102);
nor (n97,n98,n100);
and (n98,n99,n87);
and (n100,n101,n36);
not (n101,n99);
not (n102,n88);
and (n103,n11,n46);
xor (n104,n105,n113);
xor (n105,n106,n112);
nand (n106,n107,n108);
or (n107,n48,n68);
or (n108,n58,n109);
nor (n109,n110,n111);
and (n110,n57,n17);
and (n111,n52,n16);
and (n112,n78,n83);
xor (n113,n114,n134);
xor (n114,n115,n124);
and (n115,n116,n74);
not (n116,n117);
nor (n117,n118,n123);
and (n118,n119,n52);
not (n119,n120);
wire s0n120,s1n120,notn120;
or (n120,s0n120,s1n120);
not(notn120,n22);
and (s0n120,notn120,n121);
and (s1n120,n22,n122);
and (n123,n120,n57);
nand (n124,n125,n132);
or (n125,n102,n126);
not (n126,n127);
nor (n127,n128,n130);
and (n128,n129,n36);
and (n130,n131,n87);
not (n131,n129);
nand (n132,n133,n86);
not (n133,n97);
nand (n134,n135,n137);
or (n135,n136,n24);
not (n136,n41);
nand (n137,n34,n138);
nand (n138,n139,n140);
or (n139,n19,n95);
or (n140,n18,n93);
or (n141,n142,n224);
and (n142,n143,n164);
xor (n143,n144,n163);
or (n144,n145,n162);
and (n145,n146,n155);
xor (n146,n147,n148);
and (n147,n59,n74);
nand (n148,n149,n154);
or (n149,n150,n24);
not (n150,n151);
nor (n151,n152,n153);
and (n152,n51,n19);
and (n153,n56,n18);
nand (n154,n14,n34);
nand (n155,n156,n161);
or (n156,n85,n157);
not (n157,n158);
nor (n158,n159,n160);
and (n159,n45,n87);
and (n160,n43,n36);
or (n161,n91,n102);
and (n162,n147,n148);
xor (n163,n10,n77);
or (n164,n165,n223);
and (n165,n166,n222);
xor (n166,n167,n181);
nor (n167,n168,n176);
not (n168,n169);
nand (n169,n170,n175);
or (n170,n171,n85);
not (n171,n172);
nand (n172,n173,n174);
or (n173,n16,n36);
nand (n174,n36,n16);
nand (n175,n158,n88);
nand (n176,n177,n19);
nand (n177,n178,n180);
or (n178,n36,n179);
and (n179,n74,n29);
or (n180,n29,n74);
nand (n181,n182,n220);
or (n182,n183,n206);
not (n183,n184);
nand (n184,n185,n205);
or (n185,n186,n195);
nor (n186,n187,n194);
nand (n187,n188,n193);
or (n188,n189,n85);
not (n189,n190);
nand (n190,n191,n192);
or (n191,n56,n36);
nand (n192,n36,n56);
nand (n193,n172,n88);
nor (n194,n33,n76);
nand (n195,n196,n203);
nand (n196,n197,n202);
or (n197,n198,n85);
not (n198,n199);
nand (n199,n200,n201);
or (n200,n87,n74);
or (n201,n36,n76);
nand (n202,n190,n88);
nor (n203,n204,n87);
and (n204,n74,n88);
nand (n205,n187,n194);
not (n206,n207);
nand (n207,n208,n216);
not (n208,n209);
nand (n209,n210,n215);
or (n210,n211,n24);
not (n211,n212);
nand (n212,n213,n214);
or (n213,n18,n74);
or (n214,n19,n76);
nand (n215,n34,n151);
nor (n216,n217,n219);
and (n217,n168,n218);
not (n218,n176);
and (n219,n169,n176);
nand (n220,n221,n209);
not (n221,n216);
xor (n222,n146,n155);
and (n223,n167,n181);
and (n224,n144,n163);
and (n225,n8,n104);
or (n226,n227,n280);
xor (n227,n228,n251);
xor (n228,n229,n248);
xor (n229,n230,n239);
nor (n230,n231,n235);
nor (n231,n232,n234);
and (n232,n57,n233);
nand (n233,n120,n74);
and (n234,n119,n76);
not (n235,n236);
wire s0n236,s1n236,notn236;
or (n236,s0n236,s1n236);
not(notn236,n22);
and (s0n236,notn236,n237);
and (s1n236,n22,n238);
nand (n239,n240,n241);
or (n240,n126,n85);
nand (n241,n242,n88);
not (n242,n243);
nor (n243,n244,n247);
and (n244,n245,n36);
not (n245,n246);
and (n247,n246,n87);
or (n248,n249,n250);
and (n249,n114,n134);
and (n250,n115,n124);
xor (n251,n252,n274);
xor (n252,n253,n267);
nand (n253,n254,n263);
or (n254,n255,n259);
not (n255,n256);
nand (n256,n257,n258);
or (n257,n235,n74);
or (n258,n236,n76);
nand (n259,n117,n260);
nand (n260,n261,n262);
or (n261,n119,n236);
nand (n262,n236,n119);
or (n263,n117,n264);
nor (n264,n265,n266);
and (n265,n51,n235);
and (n266,n56,n236);
nand (n267,n268,n270);
or (n268,n269,n24);
not (n269,n138);
nand (n270,n34,n271);
nor (n271,n272,n273);
and (n272,n99,n19);
and (n273,n101,n18);
nand (n274,n275,n276);
or (n275,n68,n109);
or (n276,n58,n277);
nor (n277,n278,n279);
and (n278,n57,n43);
and (n279,n52,n45);
or (n280,n281,n282);
and (n281,n105,n113);
and (n282,n106,n112);
not (n283,n284);
nand (n284,n227,n280);
not (n285,n286);
nor (n286,n287,n337);
not (n287,n288);
nand (n288,n289,n334);
xor (n289,n290,n318);
xor (n290,n291,n294);
or (n291,n292,n293);
and (n292,n252,n274);
and (n293,n253,n267);
xor (n294,n295,n312);
xor (n295,n296,n304);
and (n296,n297,n74);
not (n297,n298);
nand (n298,n236,n299);
not (n299,n300);
wire s0n300,s1n300,notn300;
or (n300,s0n300,s1n300);
not(notn300,n22);
and (s0n300,notn300,1'b0);
and (s1n300,n22,n302);
and (n302,n303,n238);
nand (n304,n305,n306);
or (n305,n85,n243);
or (n306,n307,n102);
nor (n307,n308,n310);
and (n308,n87,n309);
and (n310,n36,n311);
not (n311,n309);
nand (n312,n313,n314);
or (n313,n259,n264);
or (n314,n117,n315);
nor (n315,n316,n317);
and (n316,n17,n235);
and (n317,n16,n236);
xor (n318,n319,n333);
xor (n319,n320,n327);
nand (n320,n321,n323);
or (n321,n24,n322);
not (n322,n271);
or (n323,n33,n324);
nor (n324,n325,n326);
and (n325,n18,n129);
and (n326,n19,n131);
nand (n327,n328,n329);
or (n328,n68,n277);
or (n329,n58,n330);
nor (n330,n331,n332);
and (n331,n57,n93);
and (n332,n52,n95);
and (n333,n230,n239);
or (n334,n335,n336);
and (n335,n228,n251);
and (n336,n229,n248);
nor (n337,n289,n334);
or (n338,n286,n3);
xor (n339,n340,n500);
xor (n340,n341,n497);
xor (n341,n342,n496);
xor (n342,n343,n487);
xor (n343,n344,n486);
xor (n344,n345,n472);
xor (n345,n346,n471);
xor (n346,n347,n451);
xor (n347,n348,n450);
xor (n348,n349,n426);
xor (n349,n350,n272);
xor (n350,n351,n394);
xor (n351,n352,n393);
xor (n352,n353,n356);
xor (n353,n354,n355);
and (n354,n309,n88);
and (n355,n246,n36);
or (n356,n357,n359);
and (n357,n358,n128);
and (n358,n246,n88);
and (n359,n360,n361);
xor (n360,n358,n128);
or (n361,n362,n365);
and (n362,n363,n364);
and (n363,n129,n88);
and (n364,n99,n36);
and (n365,n366,n367);
xor (n366,n363,n364);
or (n367,n368,n371);
and (n368,n369,n370);
and (n369,n99,n88);
and (n370,n93,n36);
and (n371,n372,n373);
xor (n372,n369,n370);
or (n373,n374,n376);
and (n374,n375,n160);
and (n375,n93,n88);
and (n376,n377,n378);
xor (n377,n375,n160);
or (n378,n379,n382);
and (n379,n380,n381);
and (n380,n43,n88);
and (n381,n17,n36);
and (n382,n383,n384);
xor (n383,n380,n381);
or (n384,n385,n388);
and (n385,n386,n387);
and (n386,n17,n88);
and (n387,n51,n36);
and (n388,n389,n390);
xor (n389,n386,n387);
and (n390,n391,n392);
and (n391,n51,n88);
and (n392,n74,n36);
and (n393,n129,n29);
or (n394,n395,n398);
and (n395,n396,n397);
xor (n396,n360,n361);
and (n397,n99,n29);
and (n398,n399,n400);
xor (n399,n396,n397);
or (n400,n401,n404);
and (n401,n402,n403);
xor (n402,n366,n367);
and (n403,n93,n29);
and (n404,n405,n406);
xor (n405,n402,n403);
or (n406,n407,n410);
and (n407,n408,n409);
xor (n408,n372,n373);
and (n409,n43,n29);
and (n410,n411,n412);
xor (n411,n408,n409);
or (n412,n413,n416);
and (n413,n414,n415);
xor (n414,n377,n378);
and (n415,n17,n29);
and (n416,n417,n418);
xor (n417,n414,n415);
or (n418,n419,n422);
and (n419,n420,n421);
xor (n420,n383,n384);
and (n421,n51,n29);
and (n422,n423,n424);
xor (n423,n420,n421);
and (n424,n425,n179);
xor (n425,n389,n390);
or (n426,n427,n430);
and (n427,n428,n429);
xor (n428,n399,n400);
and (n429,n93,n19);
and (n430,n431,n432);
xor (n431,n428,n429);
or (n432,n433,n435);
and (n433,n434,n42);
xor (n434,n405,n406);
and (n435,n436,n437);
xor (n436,n434,n42);
or (n437,n438,n440);
and (n438,n439,n23);
xor (n439,n411,n412);
and (n440,n441,n442);
xor (n441,n439,n23);
or (n442,n443,n445);
and (n443,n444,n152);
xor (n444,n417,n418);
and (n445,n446,n447);
xor (n446,n444,n152);
and (n447,n448,n449);
xor (n448,n423,n424);
and (n449,n74,n19);
and (n450,n93,n62);
or (n451,n452,n455);
and (n452,n453,n454);
xor (n453,n431,n432);
and (n454,n43,n62);
and (n455,n456,n457);
xor (n456,n453,n454);
or (n457,n458,n461);
and (n458,n459,n460);
xor (n459,n436,n437);
and (n460,n17,n62);
and (n461,n462,n463);
xor (n462,n459,n460);
or (n463,n464,n467);
and (n464,n465,n466);
xor (n465,n441,n442);
and (n466,n51,n62);
and (n467,n468,n469);
xor (n468,n465,n466);
and (n469,n470,n81);
xor (n470,n446,n447);
and (n471,n43,n52);
or (n472,n473,n476);
and (n473,n474,n475);
xor (n474,n456,n457);
and (n475,n17,n52);
and (n476,n477,n478);
xor (n477,n474,n475);
or (n478,n479,n481);
and (n479,n480,n50);
xor (n480,n462,n463);
and (n481,n482,n483);
xor (n482,n480,n50);
and (n483,n484,n485);
xor (n484,n468,n469);
and (n485,n74,n52);
and (n486,n17,n120);
or (n487,n488,n491);
and (n488,n489,n490);
xor (n489,n477,n478);
and (n490,n51,n120);
and (n491,n492,n493);
xor (n492,n489,n490);
and (n493,n494,n495);
xor (n494,n482,n483);
not (n495,n233);
and (n496,n51,n236);
and (n497,n498,n499);
xor (n498,n492,n493);
and (n499,n74,n236);
and (n500,n74,n300);
endmodule
