module top (out,n5,n6,n7,n33,n35,n39,n49,n51,n58
        ,n63,n69,n76,n77,n85,n86,n96,n106,n108,n115
        ,n120,n126,n133,n134,n142,n143,n152,n160,n161,n167
        ,n171,n177,n188,n189,n195,n206,n214,n220,n223,n229
        ,n238,n245,n246,n265,n266,n270,n272,n284,n286,n292
        ,n298,n303,n312,n313,n323,n338,n344,n368,n380,n388
        ,n396,n417,n423,n432,n444,n445,n450,n456,n461,n473
        ,n478,n496,n502,n535,n553,n565,n583,n615,n640,n646
        ,n653,n660,n667,n679,n735,n761,n794,n847,n853,n1241
        ,n1260,n1266,n1317,n1559,n1590,n1633,n1734,n1780,n1822,n1829
        ,n1835);
output out;
input n5;
input n6;
input n7;
input n33;
input n35;
input n39;
input n49;
input n51;
input n58;
input n63;
input n69;
input n76;
input n77;
input n85;
input n86;
input n96;
input n106;
input n108;
input n115;
input n120;
input n126;
input n133;
input n134;
input n142;
input n143;
input n152;
input n160;
input n161;
input n167;
input n171;
input n177;
input n188;
input n189;
input n195;
input n206;
input n214;
input n220;
input n223;
input n229;
input n238;
input n245;
input n246;
input n265;
input n266;
input n270;
input n272;
input n284;
input n286;
input n292;
input n298;
input n303;
input n312;
input n313;
input n323;
input n338;
input n344;
input n368;
input n380;
input n388;
input n396;
input n417;
input n423;
input n432;
input n444;
input n445;
input n450;
input n456;
input n461;
input n473;
input n478;
input n496;
input n502;
input n535;
input n553;
input n565;
input n583;
input n615;
input n640;
input n646;
input n653;
input n660;
input n667;
input n679;
input n735;
input n761;
input n794;
input n847;
input n853;
input n1241;
input n1260;
input n1266;
input n1317;
input n1559;
input n1590;
input n1633;
input n1734;
input n1780;
input n1822;
input n1829;
input n1835;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n24;
wire n25;
wire n26;
wire n27;
wire n28;
wire n29;
wire n30;
wire n31;
wire n32;
wire n34;
wire n36;
wire n37;
wire n38;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n50;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n59;
wire n60;
wire n61;
wire n62;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n107;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n116;
wire n117;
wire n118;
wire n119;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n168;
wire n169;
wire n170;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n221;
wire n222;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n267;
wire n268;
wire n269;
wire n271;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n285;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n299;
wire n300;
wire n301;
wire n302;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n446;
wire n447;
wire n448;
wire n449;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n457;
wire n458;
wire n459;
wire n460;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n474;
wire n475;
wire n476;
wire n477;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2988;
wire n2989;
wire n2990;
wire n2991;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2996;
wire n2997;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3003;
wire n3004;
wire n3005;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3010;
wire n3011;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3038;
wire n3039;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
wire n3056;
wire n3057;
wire n3058;
wire n3059;
wire n3060;
wire n3061;
wire n3062;
wire n3063;
wire n3064;
wire n3065;
wire n3066;
wire n3067;
wire n3068;
wire n3069;
wire n3070;
wire n3071;
wire n3072;
wire n3073;
wire n3074;
wire n3075;
wire n3076;
wire n3077;
wire n3078;
wire n3079;
wire n3080;
wire n3081;
wire n3082;
wire n3083;
wire n3084;
wire n3085;
wire n3086;
wire n3087;
wire n3088;
wire n3089;
wire n3090;
wire n3091;
wire n3092;
wire n3093;
wire n3094;
wire n3095;
wire n3096;
wire n3097;
wire n3098;
wire n3099;
wire n3100;
wire n3101;
wire n3102;
wire n3103;
wire n3104;
wire n3105;
wire n3106;
wire n3107;
wire n3108;
wire n3109;
wire n3110;
wire n3111;
wire n3112;
wire n3113;
wire n3114;
wire n3115;
wire n3116;
wire n3117;
wire n3118;
wire n3119;
wire n3120;
wire n3121;
wire n3122;
wire n3123;
wire n3124;
wire n3125;
wire n3126;
wire n3127;
wire n3128;
wire n3129;
wire n3130;
wire n3131;
wire n3132;
wire n3133;
wire n3134;
wire n3135;
wire n3136;
wire n3137;
wire n3138;
wire n3139;
wire n3140;
wire n3141;
wire n3142;
wire n3143;
wire n3144;
wire n3145;
wire n3146;
wire n3147;
wire n3148;
wire n3149;
wire n3150;
wire n3151;
wire n3152;
wire n3153;
wire n3154;
wire n3155;
wire n3156;
wire n3157;
wire n3158;
wire n3159;
wire n3160;
wire n3161;
wire n3162;
wire n3163;
wire n3164;
wire n3165;
wire n3166;
wire n3167;
wire n3168;
wire n3169;
wire n3170;
wire n3171;
wire n3172;
wire n3173;
wire n3174;
wire n3175;
wire n3176;
wire n3177;
wire n3178;
wire n3179;
wire n3180;
wire n3181;
wire n3182;
wire n3183;
wire n3184;
wire n3185;
wire n3186;
wire n3187;
wire n3188;
wire n3189;
wire n3190;
wire n3191;
wire n3192;
wire n3193;
wire n3194;
wire n3195;
wire n3196;
wire n3197;
wire n3198;
wire n3199;
wire n3200;
wire n3201;
wire n3202;
wire n3203;
wire n3204;
wire n3205;
wire n3206;
wire n3207;
wire n3208;
wire n3209;
wire n3210;
wire n3211;
wire n3212;
wire n3213;
wire n3214;
wire n3215;
wire n3216;
wire n3217;
wire n3218;
wire n3219;
wire n3220;
wire n3221;
wire n3222;
wire n3223;
wire n3224;
wire n3225;
wire n3226;
wire n3227;
wire n3228;
wire n3229;
wire n3230;
wire n3231;
wire n3232;
wire n3233;
wire n3234;
wire n3235;
wire n3236;
wire n3237;
wire n3238;
wire n3239;
wire n3240;
wire n3241;
wire n3242;
wire n3243;
wire n3244;
wire n3245;
wire n3246;
wire n3247;
wire n3248;
wire n3249;
wire n3250;
wire n3251;
wire n3252;
wire n3253;
wire n3254;
wire n3255;
wire n3256;
wire n3257;
wire n3258;
wire n3259;
wire n3260;
wire n3261;
wire n3262;
wire n3263;
wire n3264;
wire n3265;
wire n3266;
wire n3267;
wire n3268;
wire n3269;
wire n3270;
wire n3271;
wire n3272;
wire n3273;
wire n3274;
wire n3275;
wire n3276;
wire n3277;
wire n3278;
wire n3279;
wire n3280;
wire n3281;
wire n3282;
wire n3283;
wire n3284;
wire n3285;
wire n3286;
wire n3287;
wire n3288;
wire n3289;
wire n3290;
wire n3291;
wire n3292;
wire n3293;
wire n3294;
wire n3295;
wire n3296;
wire n3297;
wire n3298;
wire n3299;
wire n3300;
wire n3301;
wire n3302;
wire n3303;
wire n3304;
wire n3305;
wire n3306;
wire n3307;
wire n3308;
wire n3309;
wire n3310;
wire n3311;
wire n3312;
wire n3313;
wire n3314;
wire n3315;
wire n3316;
wire n3317;
wire n3318;
wire n3319;
wire n3320;
wire n3321;
wire n3322;
wire n3323;
wire n3324;
wire n3325;
wire n3326;
wire n3327;
wire n3328;
wire n3329;
wire n3330;
wire n3331;
wire n3332;
wire n3333;
wire n3334;
wire n3335;
wire n3336;
wire n3337;
wire n3338;
wire n3339;
wire n3340;
wire n3341;
wire n3342;
wire n3343;
wire n3344;
wire n3345;
wire n3346;
wire n3347;
wire n3348;
wire n3349;
wire n3350;
wire n3351;
wire n3352;
wire n3353;
wire n3354;
wire n3355;
wire n3356;
wire n3357;
wire n3358;
wire n3359;
wire n3360;
wire n3361;
wire n3362;
wire n3363;
wire n3364;
wire n3365;
wire n3366;
wire n3367;
wire n3368;
wire n3369;
wire n3370;
wire n3371;
wire n3372;
wire n3373;
wire n3374;
wire n3375;
wire n3376;
wire n3377;
wire n3378;
wire n3379;
wire n3380;
wire n3381;
wire n3382;
wire n3383;
wire n3384;
wire n3385;
wire n3386;
wire n3387;
wire n3388;
wire n3389;
wire n3390;
wire n3391;
wire n3392;
wire n3393;
wire n3394;
wire n3395;
wire n3396;
wire n3397;
wire n3398;
wire n3399;
wire n3400;
wire n3401;
wire n3402;
wire n3403;
wire n3404;
wire n3405;
wire n3406;
wire n3407;
wire n3408;
wire n3409;
wire n3410;
wire n3411;
wire n3412;
wire n3413;
wire n3414;
wire n3415;
wire n3416;
wire n3417;
wire n3418;
wire n3419;
wire n3420;
wire n3421;
wire n3422;
wire n3423;
wire n3424;
wire n3425;
wire n3426;
wire n3427;
wire n3428;
wire n3429;
wire n3430;
wire n3431;
wire n3432;
wire n3433;
wire n3434;
wire n3435;
wire n3436;
wire n3437;
wire n3438;
wire n3439;
wire n3440;
wire n3441;
wire n3442;
wire n3443;
wire n3444;
wire n3445;
wire n3446;
wire n3447;
wire n3448;
wire n3449;
wire n3450;
wire n3451;
wire n3452;
wire n3453;
wire n3454;
wire n3455;
wire n3456;
wire n3457;
wire n3458;
wire n3459;
wire n3460;
wire n3461;
wire n3462;
wire n3463;
wire n3464;
wire n3465;
wire n3466;
wire n3467;
wire n3468;
wire n3469;
wire n3470;
wire n3471;
wire n3472;
wire n3473;
wire n3474;
wire n3475;
wire n3476;
wire n3477;
wire n3478;
wire n3479;
wire n3480;
wire n3481;
wire n3482;
wire n3483;
wire n3484;
wire n3485;
wire n3486;
wire n3487;
wire n3488;
wire n3489;
wire n3490;
wire n3491;
wire n3492;
wire n3493;
wire n3494;
wire n3495;
wire n3496;
wire n3497;
wire n3498;
wire n3499;
wire n3500;
wire n3501;
wire n3502;
wire n3503;
wire n3504;
wire n3505;
wire n3506;
wire n3507;
wire n3508;
wire n3509;
wire n3510;
wire n3511;
wire n3512;
wire n3513;
wire n3514;
wire n3515;
wire n3516;
wire n3517;
wire n3518;
wire n3519;
wire n3520;
wire n3521;
wire n3522;
wire n3523;
wire n3524;
wire n3525;
wire n3526;
wire n3527;
wire n3528;
wire n3529;
wire n3530;
wire n3531;
wire n3532;
wire n3533;
wire n3534;
wire n3535;
wire n3536;
wire n3537;
wire n3538;
wire n3539;
wire n3540;
wire n3541;
wire n3542;
wire n3543;
wire n3544;
wire n3545;
wire n3546;
wire n3547;
wire n3548;
wire n3549;
wire n3550;
wire n3551;
wire n3552;
wire n3553;
wire n3554;
wire n3555;
wire n3556;
wire n3557;
wire n3558;
wire n3559;
wire n3560;
wire n3561;
wire n3562;
wire n3563;
wire n3564;
wire n3565;
wire n3566;
wire n3567;
wire n3568;
wire n3569;
wire n3570;
wire n3571;
wire n3572;
wire n3573;
wire n3574;
wire n3575;
wire n3576;
wire n3577;
wire n3578;
wire n3579;
wire n3580;
wire n3581;
wire n3582;
wire n3583;
wire n3584;
wire n3585;
wire n3586;
wire n3587;
wire n3588;
wire n3589;
wire n3590;
wire n3591;
wire n3592;
wire n3593;
wire n3594;
wire n3595;
wire n3596;
wire n3597;
wire n3598;
wire n3599;
wire n3600;
wire n3601;
wire n3602;
wire n3603;
wire n3604;
wire n3605;
wire n3606;
wire n3607;
wire n3608;
wire n3609;
wire n3610;
wire n3611;
wire n3612;
wire n3613;
wire n3614;
wire n3615;
wire n3616;
wire n3617;
wire n3618;
wire n3619;
wire n3620;
wire n3621;
wire n3622;
wire n3623;
wire n3624;
wire n3625;
wire n3626;
wire n3627;
wire n3628;
wire n3629;
wire n3630;
wire n3631;
wire n3632;
wire n3633;
wire n3634;
wire n3635;
wire n3636;
wire n3637;
wire n3638;
wire n3639;
wire n3640;
wire n3641;
wire n3642;
wire n3643;
wire n3644;
wire n3645;
wire n3646;
wire n3647;
wire n3648;
wire n3649;
wire n3650;
wire n3651;
wire n3652;
wire n3653;
wire n3654;
wire n3655;
wire n3656;
wire n3657;
wire n3658;
wire n3659;
wire n3660;
wire n3661;
wire n3662;
wire n3663;
wire n3664;
wire n3665;
wire n3666;
wire n3667;
wire n3668;
wire n3669;
wire n3670;
wire n3671;
wire n3672;
wire n3673;
wire n3674;
wire n3675;
wire n3676;
wire n3677;
wire n3678;
wire n3679;
wire n3680;
wire n3681;
wire n3682;
wire n3683;
wire n3684;
wire n3685;
wire n3686;
wire n3687;
wire n3688;
wire n3689;
wire n3690;
wire n3691;
wire n3692;
wire n3693;
wire n3694;
wire n3695;
wire n3696;
wire n3697;
wire n3698;
wire n3699;
wire n3700;
wire n3701;
wire n3702;
wire n3703;
wire n3704;
wire n3705;
wire n3706;
wire n3707;
wire n3708;
wire n3709;
wire n3710;
wire n3711;
wire n3712;
wire n3713;
wire n3714;
wire n3715;
wire n3716;
wire n3717;
wire n3718;
wire n3719;
wire n3720;
wire n3721;
wire n3722;
wire n3723;
wire n3724;
wire n3725;
wire n3726;
wire n3727;
wire n3728;
wire n3729;
wire n3730;
wire n3731;
wire n3732;
wire n3733;
wire n3734;
wire n3735;
wire n3736;
wire n3737;
wire n3738;
wire n3739;
wire n3740;
wire n3741;
wire n3742;
wire n3743;
wire n3744;
wire n3745;
wire n3746;
wire n3747;
wire n3748;
wire n3749;
wire n3750;
wire n3751;
wire n3752;
wire n3753;
wire n3754;
wire n3755;
wire n3756;
wire n3757;
wire n3758;
wire n3759;
wire n3760;
wire n3761;
wire n3762;
wire n3763;
wire n3764;
wire n3765;
wire n3766;
wire n3767;
wire n3768;
wire n3769;
wire n3770;
wire n3771;
wire n3772;
wire n3773;
wire n3774;
wire n3775;
wire n3776;
wire n3777;
wire n3778;
wire n3779;
wire n3780;
wire n3781;
wire n3782;
wire n3783;
wire n3784;
wire n3785;
wire n3786;
wire n3787;
wire n3788;
wire n3789;
wire n3790;
wire n3791;
wire n3792;
wire n3793;
wire n3794;
wire n3795;
wire n3796;
wire n3797;
wire n3798;
wire n3799;
wire n3800;
wire n3801;
wire n3802;
wire n3803;
wire n3804;
wire n3805;
wire n3806;
wire n3807;
wire n3808;
wire n3809;
wire n3810;
wire n3811;
wire n3812;
wire n3813;
wire n3814;
wire n3815;
wire n3816;
wire n3817;
wire n3818;
wire n3819;
wire n3820;
wire n3821;
wire n3822;
wire n3823;
wire n3824;
wire n3825;
wire n3826;
wire n3827;
wire n3828;
wire n3829;
wire n3830;
wire n3831;
wire n3832;
wire n3833;
wire n3834;
wire n3835;
wire n3836;
wire n3837;
wire n3838;
wire n3839;
wire n3840;
wire n3841;
wire n3842;
wire n3843;
wire n3844;
wire n3845;
wire n3846;
wire n3847;
wire n3848;
wire n3849;
wire n3850;
wire n3851;
wire n3852;
wire n3853;
wire n3854;
wire n3855;
wire n3856;
wire n3857;
wire n3858;
wire n3859;
wire n3860;
wire n3861;
wire n3862;
wire n3863;
wire n3864;
wire n3865;
wire n3866;
wire n3867;
wire n3868;
wire n3869;
wire n3870;
wire n3871;
wire n3872;
wire n3873;
wire n3874;
wire n3875;
wire n3876;
wire n3877;
wire n3878;
wire n3879;
wire n3880;
wire n3881;
wire n3882;
wire n3883;
wire n3884;
wire n3885;
wire n3886;
wire n3887;
wire n3888;
wire n3889;
wire n3890;
wire n3891;
wire n3892;
wire n3893;
wire n3894;
wire n3895;
wire n3896;
wire n3897;
wire n3898;
wire n3899;
wire n3900;
wire n3901;
wire n3902;
wire n3903;
wire n3904;
wire n3905;
wire n3906;
wire n3907;
wire n3908;
wire n3909;
wire n3910;
wire n3911;
wire n3912;
wire n3913;
wire n3914;
wire n3915;
wire n3916;
wire n3917;
wire n3918;
wire n3919;
wire n3920;
wire n3921;
wire n3922;
wire n3923;
wire n3924;
wire n3925;
wire n3926;
wire n3927;
wire n3928;
wire n3929;
wire n3930;
wire n3931;
wire n3932;
wire n3933;
wire n3934;
wire n3935;
wire n3936;
wire n3937;
wire n3938;
wire n3939;
wire n3940;
wire n3941;
wire n3942;
wire n3943;
wire n3944;
wire n3945;
wire n3946;
wire n3947;
wire n3948;
wire n3949;
wire n3950;
wire n3951;
wire n3952;
wire n3953;
wire n3954;
wire n3955;
wire n3956;
wire n3957;
wire n3958;
wire n3959;
wire n3960;
wire n3961;
wire n3962;
wire n3963;
wire n3964;
wire n3965;
wire n3966;
wire n3967;
wire n3968;
wire n3969;
wire n3970;
wire n3971;
wire n3972;
wire n3973;
wire n3974;
wire n3975;
wire n3976;
wire n3977;
wire n3978;
wire n3979;
wire n3980;
wire n3981;
wire n3982;
wire n3983;
wire n3984;
wire n3985;
wire n3986;
wire n3987;
wire n3988;
wire n3989;
wire n3990;
wire n3991;
wire n3992;
wire n3993;
wire n3994;
wire n3995;
wire n3996;
wire n3997;
wire n3998;
wire n3999;
wire n4000;
wire n4001;
wire n4002;
wire n4003;
wire n4004;
wire n4005;
wire n4006;
wire n4007;
wire n4008;
wire n4009;
wire n4010;
wire n4011;
wire n4012;
wire n4013;
wire n4014;
wire n4015;
wire n4016;
wire n4017;
wire n4018;
wire n4019;
wire n4020;
wire n4021;
wire n4022;
wire n4023;
wire n4024;
wire n4025;
wire n4026;
wire n4027;
wire n4028;
wire n4029;
wire n4030;
wire n4031;
wire n4032;
wire n4033;
wire n4034;
wire n4035;
wire n4036;
wire n4037;
wire n4038;
wire n4039;
wire n4040;
wire n4041;
wire n4042;
wire n4043;
wire n4044;
wire n4045;
wire n4046;
wire n4047;
wire n4048;
wire n4049;
wire n4050;
wire n4051;
wire n4052;
wire n4053;
wire n4054;
wire n4055;
wire n4056;
wire n4057;
wire n4058;
wire n4059;
wire n4060;
wire n4061;
wire n4062;
wire n4063;
wire n4064;
wire n4065;
wire n4066;
wire n4067;
wire n4068;
wire n4069;
wire n4070;
wire n4071;
wire n4072;
wire n4073;
wire n4074;
wire n4075;
wire n4076;
wire n4077;
wire n4078;
wire n4079;
wire n4080;
wire n4081;
wire n4082;
wire n4083;
wire n4084;
wire n4085;
wire n4086;
wire n4087;
wire n4088;
wire n4089;
wire n4090;
wire n4091;
wire n4092;
wire n4093;
wire n4094;
wire n4095;
wire n4096;
wire n4097;
wire n4098;
wire n4099;
wire n4100;
wire n4101;
wire n4102;
wire n4103;
wire n4104;
wire n4105;
wire n4106;
wire n4107;
wire n4108;
wire n4109;
wire n4110;
wire n4111;
wire n4112;
wire n4113;
wire n4114;
wire n4115;
wire n4116;
wire n4117;
wire n4118;
wire n4119;
wire n4120;
wire n4121;
wire n4122;
wire n4123;
wire n4124;
wire n4125;
wire n4126;
wire n4127;
wire n4128;
wire n4129;
wire n4130;
wire n4131;
wire n4132;
wire n4133;
wire n4134;
wire n4135;
wire n4136;
wire n4137;
wire n4138;
wire n4139;
wire n4140;
wire n4141;
wire n4142;
wire n4143;
wire n4144;
wire n4145;
wire n4146;
wire n4147;
wire n4148;
wire n4149;
wire n4150;
wire n4151;
wire n4152;
wire n4153;
wire n4154;
wire n4155;
wire n4156;
wire n4157;
wire n4158;
wire n4159;
wire n4160;
wire n4161;
wire n4162;
wire n4163;
wire n4164;
wire n4165;
wire n4166;
wire n4167;
wire n4168;
wire n4169;
wire n4170;
wire n4171;
wire n4172;
wire n4173;
wire n4174;
wire n4175;
wire n4176;
wire n4177;
wire n4178;
wire n4179;
wire n4180;
wire n4181;
wire n4182;
wire n4183;
wire n4184;
wire n4185;
wire n4186;
wire n4187;
wire n4188;
wire n4189;
wire n4190;
wire n4191;
wire n4192;
wire n4193;
wire n4194;
wire n4195;
wire n4196;
wire n4197;
wire n4198;
wire n4199;
wire n4200;
wire n4201;
wire n4202;
wire n4203;
wire n4204;
wire n4205;
wire n4206;
wire n4207;
wire n4208;
wire n4209;
wire n4210;
wire n4211;
wire n4212;
wire n4213;
wire n4214;
wire n4215;
wire n4216;
wire n4217;
wire n4218;
wire n4219;
wire n4220;
wire n4221;
wire n4222;
wire n4223;
wire n4224;
wire n4225;
wire n4226;
wire n4227;
wire n4228;
wire n4229;
wire n4230;
wire n4231;
wire n4232;
wire n4233;
wire n4234;
wire n4235;
wire n4236;
wire n4237;
wire n4238;
wire n4239;
wire n4240;
wire n4241;
wire n4242;
wire n4243;
wire n4244;
wire n4245;
wire n4246;
wire n4247;
wire n4248;
wire n4249;
wire n4250;
wire n4251;
wire n4252;
wire n4253;
wire n4254;
wire n4255;
wire n4256;
wire n4257;
wire n4258;
wire n4259;
wire n4260;
wire n4261;
wire n4262;
wire n4263;
wire n4264;
wire n4265;
wire n4266;
wire n4267;
wire n4268;
wire n4269;
wire n4270;
wire n4271;
wire n4272;
wire n4273;
wire n4274;
wire n4275;
wire n4276;
wire n4277;
wire n4278;
wire n4279;
wire n4280;
wire n4281;
wire n4282;
wire n4283;
wire n4284;
wire n4285;
wire n4286;
wire n4287;
wire n4288;
wire n4289;
wire n4290;
wire n4291;
wire n4292;
wire n4293;
wire n4294;
wire n4295;
wire n4296;
wire n4297;
wire n4298;
wire n4299;
wire n4300;
wire n4301;
wire n4302;
wire n4303;
wire n4304;
wire n4305;
wire n4306;
wire n4307;
wire n4308;
wire n4309;
wire n4310;
wire n4311;
wire n4312;
wire n4313;
wire n4314;
wire n4315;
wire n4316;
wire n4317;
wire n4318;
wire n4319;
wire n4320;
wire n4321;
wire n4322;
wire n4323;
wire n4324;
wire n4325;
wire n4326;
wire n4327;
wire n4328;
wire n4329;
wire n4330;
wire n4331;
wire n4332;
wire n4333;
wire n4334;
wire n4335;
wire n4336;
wire n4337;
wire n4338;
wire n4339;
wire n4340;
wire n4341;
wire n4342;
wire n4343;
wire n4344;
wire n4345;
wire n4346;
wire n4347;
wire n4348;
wire n4349;
wire n4350;
wire n4351;
wire n4352;
wire n4353;
wire n4354;
wire n4355;
wire n4356;
wire n4357;
wire n4358;
wire n4359;
wire n4360;
wire n4361;
wire n4362;
wire n4363;
wire n4364;
wire n4365;
wire n4366;
wire n4367;
wire n4368;
wire n4369;
wire n4370;
wire n4371;
wire n4372;
wire n4373;
wire n4374;
wire n4375;
wire n4376;
wire n4377;
wire n4378;
wire n4379;
wire n4380;
wire n4381;
wire n4382;
wire n4383;
wire n4384;
wire n4385;
wire n4386;
wire n4387;
wire n4388;
wire n4389;
wire n4390;
wire n4391;
wire n4392;
wire n4393;
wire n4394;
wire n4395;
wire n4396;
wire n4397;
wire n4398;
wire n4399;
wire n4400;
wire n4401;
wire n4402;
wire n4403;
wire n4404;
wire n4405;
wire n4406;
wire n4407;
wire n4408;
wire n4409;
wire n4410;
wire n4411;
wire n4412;
wire n4413;
wire n4414;
wire n4415;
wire n4416;
wire n4417;
wire n4418;
wire n4419;
wire n4420;
wire n4421;
wire n4422;
wire n4423;
wire n4424;
wire n4425;
wire n4426;
wire n4427;
wire n4428;
wire n4429;
wire n4430;
wire n4431;
wire n4432;
wire n4433;
wire n4434;
wire n4435;
wire n4436;
wire n4437;
wire n4438;
wire n4439;
wire n4440;
wire n4441;
wire n4442;
wire n4443;
wire n4444;
wire n4445;
wire n4446;
wire n4447;
wire n4448;
wire n4449;
wire n4450;
wire n4451;
wire n4452;
wire n4453;
wire n4454;
wire n4455;
wire n4456;
wire n4457;
wire n4458;
wire n4459;
wire n4460;
wire n4461;
wire n4462;
wire n4463;
wire n4464;
wire n4465;
wire n4466;
wire n4467;
wire n4468;
wire n4469;
wire n4470;
wire n4471;
wire n4472;
wire n4473;
wire n4474;
wire n4475;
wire n4476;
wire n4477;
wire n4478;
wire n4479;
wire n4480;
wire n4481;
wire n4482;
wire n4483;
wire n4484;
wire n4485;
wire n4486;
wire n4487;
wire n4488;
wire n4489;
wire n4490;
wire n4491;
wire n4492;
wire n4493;
wire n4494;
wire n4495;
wire n4496;
wire n4497;
wire n4498;
wire n4499;
wire n4500;
wire n4501;
wire n4502;
wire n4503;
wire n4504;
wire n4505;
wire n4506;
wire n4507;
wire n4508;
wire n4509;
wire n4510;
wire n4511;
wire n4512;
wire n4513;
wire n4514;
wire n4515;
wire n4516;
wire n4517;
wire n4518;
wire n4519;
wire n4520;
wire n4521;
wire n4522;
wire n4523;
wire n4524;
wire n4525;
wire n4526;
wire n4527;
wire n4528;
wire n4529;
wire n4530;
wire n4531;
wire n4532;
wire n4533;
wire n4534;
wire n4535;
wire n4536;
wire n4537;
wire n4538;
wire n4539;
wire n4540;
wire n4541;
wire n4542;
wire n4543;
wire n4544;
wire n4545;
wire n4546;
wire n4547;
wire n4548;
wire n4549;
wire n4550;
wire n4551;
wire n4552;
wire n4553;
wire n4554;
wire n4555;
wire n4556;
wire n4557;
wire n4558;
wire n4559;
wire n4560;
wire n4561;
wire n4562;
wire n4563;
wire n4564;
wire n4565;
wire n4566;
wire n4567;
wire n4568;
wire n4569;
wire n4570;
wire n4571;
wire n4572;
wire n4573;
wire n4574;
wire n4575;
wire n4576;
wire n4577;
wire n4578;
wire n4579;
wire n4580;
wire n4581;
wire n4582;
wire n4583;
wire n4584;
wire n4585;
wire n4586;
wire n4587;
wire n4588;
wire n4589;
wire n4590;
wire n4591;
wire n4592;
wire n4593;
wire n4594;
wire n4595;
wire n4596;
wire n4597;
wire n4598;
wire n4599;
wire n4600;
wire n4601;
wire n4602;
wire n4603;
wire n4604;
wire n4605;
wire n4606;
wire n4607;
wire n4608;
wire n4609;
wire n4610;
wire n4611;
wire n4612;
wire n4613;
wire n4614;
wire n4615;
wire n4616;
wire n4617;
wire n4618;
wire n4619;
wire n4620;
wire n4621;
wire n4622;
wire n4623;
wire n4624;
wire n4625;
wire n4626;
wire n4627;
wire n4628;
wire n4629;
wire n4630;
wire n4631;
wire n4632;
wire n4633;
wire n4634;
wire n4635;
wire n4636;
wire n4637;
wire n4638;
wire n4639;
wire n4640;
wire n4641;
wire n4642;
wire n4643;
wire n4644;
wire n4645;
wire n4646;
wire n4647;
wire n4648;
wire n4649;
wire n4650;
wire n4651;
wire n4652;
wire n4653;
wire n4654;
wire n4655;
wire n4656;
wire n4657;
wire n4658;
wire n4659;
wire n4660;
wire n4661;
wire n4662;
wire n4663;
wire n4664;
wire n4665;
wire n4666;
wire n4667;
wire n4668;
wire n4669;
wire n4670;
wire n4671;
wire n4672;
wire n4673;
wire n4674;
wire n4675;
wire n4676;
wire n4677;
wire n4678;
wire n4679;
wire n4680;
wire n4681;
wire n4682;
wire n4683;
wire n4684;
wire n4685;
wire n4686;
wire n4687;
wire n4688;
wire n4689;
wire n4690;
wire n4691;
wire n4692;
wire n4693;
wire n4694;
wire n4695;
wire n4696;
wire n4697;
wire n4698;
wire n4699;
wire n4700;
wire n4701;
wire n4702;
wire n4703;
wire n4704;
wire n4705;
wire n4706;
wire n4707;
wire n4708;
wire n4709;
wire n4710;
wire n4711;
wire n4712;
wire n4713;
wire n4714;
wire n4715;
wire n4716;
wire n4717;
wire n4718;
wire n4719;
wire n4720;
wire n4721;
wire n4722;
wire n4723;
wire n4724;
wire n4725;
wire n4726;
wire n4727;
wire n4728;
wire n4729;
wire n4730;
wire n4731;
wire n4732;
wire n4733;
wire n4734;
wire n4735;
wire n4736;
wire n4737;
wire n4738;
wire n4739;
wire n4740;
wire n4741;
wire n4742;
wire n4743;
wire n4744;
wire n4745;
wire n4746;
wire n4747;
wire n4748;
wire n4749;
wire n4750;
wire n4751;
wire n4752;
wire n4753;
wire n4754;
wire n4755;
wire n4756;
wire n4757;
wire n4758;
wire n4759;
wire n4760;
wire n4761;
wire n4762;
wire n4763;
wire n4764;
wire n4765;
wire n4766;
wire n4767;
wire n4768;
wire n4769;
wire n4770;
wire n4771;
wire n4772;
wire n4773;
wire n4774;
wire n4775;
wire n4776;
wire n4777;
wire n4778;
wire n4779;
wire n4780;
wire n4781;
wire n4782;
wire n4783;
wire n4784;
wire n4785;
wire n4786;
wire n4787;
wire n4788;
wire n4789;
wire n4790;
wire n4791;
wire n4792;
wire n4793;
wire n4794;
wire n4795;
wire n4796;
wire n4797;
wire n4798;
wire n4799;
wire n4800;
wire n4801;
wire n4802;
wire n4803;
wire n4804;
wire n4805;
wire n4806;
wire n4807;
wire n4808;
wire n4809;
wire n4810;
wire n4811;
wire n4812;
wire n4813;
wire n4814;
wire n4815;
wire n4816;
wire n4817;
wire n4818;
wire n4819;
wire n4820;
wire n4821;
wire n4822;
wire n4823;
wire n4824;
wire n4825;
wire n4826;
wire n4827;
wire n4828;
wire n4829;
wire n4830;
wire n4831;
wire n4832;
wire n4833;
wire n4834;
wire n4835;
wire n4836;
wire n4837;
wire n4838;
wire n4839;
wire n4840;
wire n4841;
wire n4842;
wire n4843;
wire n4844;
wire n4845;
wire n4846;
wire n4847;
wire n4848;
wire n4849;
wire n4850;
wire n4851;
wire n4852;
wire n4853;
wire n4854;
wire n4855;
wire n4856;
wire n4857;
wire n4858;
wire n4859;
wire n4860;
wire n4861;
wire n4862;
wire n4863;
wire n4864;
wire n4865;
wire n4866;
wire n4867;
wire n4868;
wire n4869;
wire n4870;
wire n4871;
wire n4872;
wire n4873;
wire n4874;
wire n4875;
wire n4876;
wire n4877;
wire n4878;
wire n4879;
wire n4880;
wire n4881;
wire n4882;
wire n4883;
wire n4884;
wire n4885;
wire n4886;
wire n4887;
wire n4888;
wire n4889;
wire n4890;
wire n4891;
wire n4892;
wire n4893;
wire n4894;
wire n4895;
wire n4896;
wire n4897;
wire n4898;
wire n4899;
wire n4900;
wire n4901;
wire n4902;
wire n4903;
wire n4904;
wire n4905;
wire n4906;
wire n4907;
wire n4908;
wire n4909;
wire n4910;
wire n4911;
wire n4912;
wire n4913;
wire n4914;
wire n4915;
wire n4916;
wire n4917;
wire n4918;
wire n4919;
wire n4920;
wire n4921;
wire n4922;
wire n4923;
wire n4924;
wire n4925;
wire n4926;
wire n4927;
wire n4928;
wire n4929;
wire n4930;
wire n4931;
wire n4932;
wire n4933;
wire n4934;
wire n4935;
wire n4936;
wire n4937;
wire n4938;
wire n4939;
wire n4940;
wire n4941;
wire n4942;
wire n4943;
wire n4944;
wire n4945;
wire n4946;
wire n4947;
wire n4948;
wire n4949;
wire n4950;
wire n4951;
wire n4952;
wire n4953;
wire n4954;
wire n4955;
wire n4956;
wire n4957;
wire n4958;
wire n4959;
wire n4960;
wire n4961;
wire n4962;
wire n4963;
wire n4964;
wire n4965;
wire n4966;
wire n4967;
wire n4968;
wire n4969;
wire n4970;
wire n4971;
wire n4972;
wire n4973;
wire n4974;
wire n4975;
wire n4976;
wire n4977;
wire n4978;
wire n4979;
wire n4980;
wire n4981;
wire n4982;
wire n4983;
wire n4984;
wire n4985;
wire n4986;
wire n4987;
wire n4988;
wire n4989;
wire n4990;
wire n4991;
wire n4992;
wire n4993;
wire n4994;
wire n4995;
wire n4996;
wire n4997;
wire n4998;
wire n4999;
wire n5000;
wire n5001;
wire n5002;
wire n5003;
wire n5004;
wire n5005;
wire n5006;
wire n5007;
wire n5008;
wire n5009;
wire n5010;
wire n5011;
wire n5012;
wire n5013;
wire n5014;
wire n5015;
wire n5016;
wire n5017;
wire n5018;
wire n5019;
wire n5020;
wire n5021;
wire n5022;
wire n5023;
wire n5024;
wire n5025;
wire n5026;
wire n5027;
wire n5028;
wire n5029;
wire n5030;
wire n5031;
wire n5032;
wire n5033;
wire n5034;
wire n5035;
wire n5036;
wire n5037;
wire n5038;
wire n5039;
wire n5040;
wire n5041;
wire n5042;
wire n5043;
wire n5044;
wire n5045;
wire n5046;
wire n5047;
wire n5048;
wire n5049;
wire n5050;
wire n5051;
wire n5052;
wire n5053;
wire n5054;
wire n5055;
wire n5056;
wire n5057;
wire n5058;
wire n5059;
wire n5060;
wire n5061;
wire n5062;
wire n5063;
wire n5064;
wire n5065;
wire n5066;
wire n5067;
wire n5068;
wire n5069;
wire n5070;
wire n5071;
wire n5072;
wire n5073;
wire n5074;
wire n5075;
wire n5076;
wire n5077;
wire n5078;
wire n5079;
wire n5080;
wire n5081;
wire n5082;
wire n5083;
wire n5084;
wire n5085;
wire n5086;
wire n5087;
wire n5088;
wire n5089;
wire n5090;
wire n5091;
wire n5092;
wire n5093;
wire n5094;
wire n5095;
wire n5096;
wire n5097;
wire n5098;
wire n5099;
wire n5100;
wire n5101;
wire n5102;
wire n5103;
wire n5104;
wire n5105;
wire n5106;
wire n5107;
wire n5108;
wire n5109;
wire n5110;
wire n5111;
wire n5112;
wire n5113;
wire n5114;
wire n5115;
wire n5116;
wire n5117;
wire n5118;
wire n5119;
wire n5120;
wire n5121;
wire n5122;
wire n5123;
wire n5124;
wire n5125;
wire n5126;
wire n5127;
wire n5128;
wire n5129;
wire n5130;
wire n5131;
wire n5132;
wire n5133;
wire n5134;
wire n5135;
wire n5136;
wire n5137;
wire n5138;
wire n5139;
wire n5140;
wire n5141;
wire n5142;
wire n5143;
wire n5144;
wire n5145;
wire n5146;
wire n5147;
wire n5148;
wire n5149;
wire n5150;
wire n5151;
wire n5152;
wire n5153;
wire n5154;
wire n5155;
wire n5156;
wire n5157;
wire n5158;
wire n5159;
wire n5160;
wire n5161;
wire n5162;
wire n5163;
wire n5164;
wire n5165;
wire n5166;
wire n5167;
wire n5168;
wire n5169;
wire n5170;
wire n5171;
wire n5172;
wire n5173;
wire n5174;
wire n5175;
wire n5176;
wire n5177;
wire n5178;
wire n5179;
wire n5180;
wire n5181;
wire n5182;
wire n5183;
wire n5184;
wire n5185;
wire n5186;
wire n5187;
wire n5188;
wire n5189;
wire n5190;
wire n5191;
wire n5192;
wire n5193;
wire n5194;
wire n5195;
wire n5196;
wire n5197;
wire n5198;
wire n5199;
wire n5200;
wire n5201;
wire n5202;
wire n5203;
wire n5204;
wire n5205;
wire n5206;
wire n5207;
wire n5208;
wire n5209;
wire n5210;
wire n5211;
wire n5212;
wire n5213;
wire n5214;
wire n5215;
wire n5216;
wire n5217;
wire n5218;
wire n5219;
wire n5220;
wire n5221;
wire n5222;
wire n5223;
wire n5224;
wire n5225;
wire n5226;
wire n5227;
wire n5228;
wire n5229;
wire n5230;
wire n5231;
wire n5232;
wire n5233;
wire n5234;
wire n5235;
wire n5236;
wire n5237;
wire n5238;
wire n5239;
wire n5240;
wire n5241;
wire n5242;
wire n5243;
wire n5244;
wire n5245;
wire n5246;
wire n5247;
wire n5248;
wire n5249;
wire n5250;
wire n5251;
wire n5252;
wire n5253;
wire n5254;
wire n5255;
wire n5256;
wire n5257;
wire n5258;
wire n5259;
wire n5260;
wire n5261;
wire n5262;
wire n5263;
wire n5264;
wire n5265;
wire n5266;
wire n5267;
wire n5268;
wire n5269;
wire n5270;
wire n5271;
wire n5272;
wire n5273;
wire n5274;
wire n5275;
wire n5276;
wire n5277;
wire n5278;
wire n5279;
wire n5280;
wire n5281;
wire n5282;
wire n5283;
wire n5284;
wire n5285;
wire n5286;
wire n5287;
wire n5288;
wire n5289;
wire n5290;
wire n5291;
wire n5292;
wire n5293;
wire n5294;
wire n5295;
wire n5296;
wire n5297;
wire n5298;
wire n5299;
wire n5300;
wire n5301;
wire n5302;
wire n5303;
wire n5304;
wire n5305;
wire n5306;
wire n5307;
wire n5308;
wire n5309;
wire n5310;
wire n5311;
wire n5312;
wire n5313;
wire n5314;
wire n5315;
wire n5316;
wire n5317;
wire n5318;
wire n5319;
wire n5320;
wire n5321;
wire n5322;
wire n5323;
wire n5324;
wire n5325;
wire n5326;
wire n5327;
wire n5328;
wire n5329;
wire n5330;
wire n5331;
wire n5332;
wire n5333;
wire n5334;
wire n5335;
wire n5336;
wire n5337;
wire n5338;
wire n5339;
wire n5340;
wire n5341;
wire n5342;
wire n5343;
wire n5344;
wire n5345;
wire n5346;
wire n5347;
wire n5348;
wire n5349;
wire n5350;
wire n5351;
wire n5352;
wire n5353;
wire n5354;
wire n5355;
wire n5356;
wire n5357;
wire n5358;
wire n5359;
wire n5360;
wire n5361;
wire n5362;
wire n5363;
wire n5364;
wire n5365;
wire n5366;
wire n5367;
wire n5368;
wire n5369;
wire n5370;
wire n5371;
wire n5372;
wire n5373;
wire n5374;
wire n5375;
wire n5376;
wire n5377;
wire n5378;
wire n5379;
wire n5380;
wire n5381;
wire n5382;
wire n5383;
wire n5384;
wire n5385;
wire n5386;
wire n5387;
wire n5388;
wire n5389;
wire n5390;
wire n5391;
wire n5392;
wire n5393;
wire n5394;
wire n5395;
wire n5396;
wire n5397;
wire n5398;
wire n5399;
wire n5400;
wire n5401;
wire n5402;
wire n5403;
wire n5404;
wire n5405;
wire n5406;
wire n5407;
wire n5408;
wire n5409;
wire n5410;
wire n5411;
wire n5412;
wire n5413;
wire n5414;
wire n5415;
wire n5416;
wire n5417;
wire n5418;
wire n5419;
wire n5420;
wire n5421;
wire n5422;
wire n5423;
wire n5424;
wire n5425;
wire n5426;
wire n5427;
wire n5428;
wire n5429;
wire n5430;
wire n5431;
wire n5432;
wire n5433;
wire n5434;
wire n5435;
wire n5436;
wire n5437;
wire n5438;
wire n5439;
wire n5440;
wire n5441;
wire n5442;
wire n5443;
wire n5444;
wire n5445;
wire n5446;
wire n5447;
wire n5448;
wire n5449;
wire n5450;
wire n5451;
wire n5452;
wire n5453;
wire n5454;
wire n5455;
wire n5456;
wire n5457;
wire n5458;
wire n5459;
wire n5460;
wire n5461;
wire n5462;
wire n5463;
wire n5464;
wire n5465;
wire n5466;
wire n5467;
wire n5468;
wire n5469;
wire n5470;
wire n5471;
wire n5472;
wire n5473;
wire n5474;
wire n5475;
wire n5476;
wire n5477;
wire n5478;
wire n5479;
wire n5480;
wire n5481;
wire n5482;
wire n5483;
wire n5484;
wire n5485;
wire n5486;
wire n5487;
wire n5488;
wire n5489;
wire n5490;
wire n5491;
wire n5492;
wire n5493;
wire n5494;
wire n5495;
wire n5496;
wire n5497;
wire n5498;
wire n5499;
wire n5500;
wire n5501;
wire n5502;
wire n5503;
wire n5504;
wire n5505;
wire n5506;
wire n5507;
wire n5508;
wire n5509;
wire n5510;
wire n5511;
wire n5512;
wire n5513;
wire n5514;
wire n5515;
wire n5516;
wire n5517;
wire n5518;
wire n5519;
wire n5520;
wire n5521;
wire n5522;
wire n5523;
wire n5524;
wire n5525;
wire n5526;
wire n5527;
wire n5528;
wire n5529;
wire n5530;
wire n5531;
wire n5532;
wire n5533;
wire n5534;
wire n5535;
wire n5536;
wire n5537;
wire n5538;
wire n5539;
wire n5540;
wire n5541;
wire n5542;
wire n5543;
wire n5544;
wire n5545;
wire n5546;
wire n5547;
wire n5548;
wire n5549;
wire n5550;
wire n5551;
wire n5552;
wire n5553;
wire n5554;
wire n5555;
wire n5556;
wire n5557;
wire n5558;
wire n5559;
wire n5560;
wire n5561;
wire n5562;
wire n5563;
wire n5564;
wire n5565;
wire n5566;
wire n5567;
wire n5568;
wire n5569;
wire n5570;
wire n5571;
wire n5572;
wire n5573;
wire n5574;
wire n5575;
wire n5576;
wire n5577;
wire n5578;
wire n5579;
wire n5580;
wire n5581;
wire n5582;
wire n5583;
wire n5584;
wire n5585;
wire n5586;
wire n5587;
wire n5588;
wire n5589;
wire n5590;
wire n5591;
wire n5592;
wire n5593;
wire n5594;
wire n5595;
wire n5596;
wire n5597;
wire n5598;
wire n5599;
wire n5600;
wire n5601;
wire n5602;
wire n5603;
wire n5604;
wire n5605;
wire n5606;
wire n5607;
wire n5608;
wire n5609;
wire n5610;
wire n5611;
wire n5612;
wire n5613;
wire n5614;
wire n5615;
wire n5616;
wire n5617;
wire n5618;
wire n5619;
wire n5620;
wire n5621;
wire n5622;
wire n5623;
wire n5624;
wire n5625;
wire n5626;
wire n5627;
wire n5628;
wire n5629;
wire n5630;
wire n5631;
wire n5632;
wire n5633;
wire n5634;
wire n5635;
wire n5636;
wire n5637;
wire n5638;
wire n5639;
wire n5640;
wire n5641;
wire n5642;
wire n5643;
wire n5644;
wire n5645;
wire n5646;
wire n5647;
wire n5648;
wire n5649;
wire n5650;
wire n5651;
wire n5652;
wire n5653;
wire n5654;
wire n5655;
wire n5656;
wire n5657;
wire n5658;
wire n5659;
wire n5660;
wire n5661;
wire n5662;
wire n5663;
wire n5664;
wire n5665;
wire n5666;
wire n5667;
wire n5668;
wire n5669;
wire n5670;
wire n5671;
wire n5672;
wire n5673;
wire n5674;
wire n5675;
wire n5676;
wire n5677;
wire n5678;
wire n5679;
wire n5680;
wire n5681;
wire n5682;
wire n5683;
wire n5684;
wire n5685;
wire n5686;
wire n5687;
wire n5688;
wire n5689;
wire n5690;
wire n5691;
wire n5692;
wire n5693;
wire n5694;
wire n5695;
wire n5696;
wire n5697;
wire n5698;
wire n5699;
wire n5700;
wire n5701;
wire n5702;
wire n5703;
wire n5704;
wire n5705;
wire n5706;
wire n5707;
wire n5708;
wire n5709;
wire n5710;
wire n5711;
wire n5712;
wire n5713;
wire n5714;
wire n5715;
wire n5716;
wire n5717;
wire n5718;
wire n5719;
wire n5720;
wire n5721;
wire n5722;
wire n5723;
wire n5724;
wire n5725;
wire n5726;
wire n5727;
wire n5728;
wire n5729;
wire n5730;
wire n5731;
wire n5732;
wire n5733;
wire n5734;
wire n5735;
wire n5736;
wire n5737;
wire n5738;
wire n5739;
wire n5740;
wire n5741;
wire n5742;
wire n5743;
wire n5744;
wire n5745;
wire n5746;
wire n5747;
wire n5748;
wire n5749;
wire n5750;
wire n5751;
wire n5752;
wire n5753;
wire n5754;
wire n5755;
wire n5756;
wire n5757;
wire n5758;
wire n5759;
wire n5760;
wire n5761;
wire n5762;
wire n5763;
wire n5764;
wire n5765;
wire n5766;
wire n5767;
wire n5768;
wire n5769;
wire n5770;
wire n5771;
wire n5772;
wire n5773;
wire n5774;
wire n5775;
wire n5776;
wire n5777;
wire n5778;
wire n5779;
wire n5780;
wire n5781;
wire n5782;
wire n5783;
wire n5784;
wire n5785;
wire n5786;
wire n5787;
wire n5788;
wire n5789;
wire n5790;
wire n5791;
wire n5792;
wire n5793;
wire n5794;
wire n5795;
wire n5796;
wire n5797;
wire n5798;
wire n5799;
wire n5800;
wire n5801;
wire n5802;
wire n5803;
wire n5804;
wire n5805;
wire n5806;
wire n5807;
wire n5808;
wire n5809;
wire n5810;
wire n5811;
wire n5812;
wire n5813;
wire n5814;
wire n5815;
wire n5816;
wire n5817;
wire n5818;
wire n5819;
wire n5820;
wire n5821;
wire n5822;
wire n5823;
wire n5824;
wire n5825;
wire n5826;
wire n5827;
wire n5828;
wire n5829;
wire n5830;
wire n5831;
wire n5832;
wire n5833;
wire n5834;
wire n5835;
wire n5836;
wire n5837;
wire n5838;
wire n5839;
wire n5840;
wire n5841;
wire n5842;
wire n5843;
wire n5844;
wire n5845;
wire n5846;
wire n5847;
wire n5848;
wire n5849;
wire n5850;
wire n5851;
wire n5852;
wire n5853;
wire n5854;
wire n5855;
wire n5856;
wire n5857;
wire n5858;
wire n5859;
wire n5860;
wire n5861;
wire n5862;
wire n5863;
wire n5864;
wire n5865;
wire n5866;
wire n5867;
wire n5868;
wire n5869;
wire n5870;
wire n5871;
wire n5872;
wire n5873;
wire n5874;
wire n5875;
wire n5876;
wire n5877;
wire n5878;
wire n5879;
wire n5880;
wire n5881;
wire n5882;
wire n5883;
wire n5884;
wire n5885;
wire n5886;
wire n5887;
wire n5888;
wire n5889;
wire n5890;
wire n5891;
wire n5892;
wire n5893;
wire n5894;
wire n5895;
wire n5896;
wire n5897;
wire n5898;
wire n5899;
wire n5900;
wire n5901;
wire n5902;
wire n5903;
wire n5904;
wire n5905;
wire n5906;
wire n5907;
wire n5908;
wire n5909;
wire n5910;
wire n5911;
wire n5912;
wire n5913;
wire n5914;
wire n5915;
wire n5916;
wire n5917;
wire n5918;
wire n5919;
wire n5920;
wire n5921;
wire n5922;
wire n5923;
wire n5924;
wire n5925;
wire n5926;
wire n5927;
wire n5928;
wire n5929;
wire n5930;
wire n5931;
wire n5932;
wire n5933;
wire n5934;
wire n5935;
wire n5936;
wire n5937;
wire n5938;
wire n5939;
wire n5940;
wire n5941;
wire n5942;
wire n5943;
wire n5944;
wire n5945;
wire n5946;
wire n5947;
wire n5948;
wire n5949;
wire n5950;
wire n5951;
wire n5952;
wire n5953;
wire n5954;
wire n5955;
wire n5956;
wire n5957;
wire n5958;
wire n5959;
wire n5960;
wire n5961;
wire n5962;
wire n5963;
wire n5964;
wire n5965;
wire n5966;
wire n5967;
wire n5968;
wire n5969;
wire n5970;
wire n5971;
wire n5972;
wire n5973;
wire n5974;
wire n5975;
wire n5976;
wire n5977;
wire n5978;
wire n5979;
wire n5980;
wire n5981;
wire n5982;
wire n5983;
wire n5984;
wire n5985;
wire n5986;
wire n5987;
wire n5988;
wire n5989;
wire n5990;
wire n5991;
wire n5992;
wire n5993;
wire n5994;
wire n5995;
wire n5996;
wire n5997;
wire n5998;
wire n5999;
wire n6000;
wire n6001;
wire n6002;
wire n6003;
wire n6004;
wire n6005;
wire n6006;
wire n6007;
wire n6008;
wire n6009;
wire n6010;
wire n6011;
wire n6012;
wire n6013;
wire n6014;
wire n6015;
wire n6016;
wire n6017;
wire n6018;
wire n6019;
wire n6020;
wire n6021;
wire n6022;
wire n6023;
wire n6024;
wire n6025;
wire n6026;
wire n6027;
wire n6028;
wire n6029;
wire n6030;
wire n6031;
wire n6032;
wire n6033;
wire n6034;
wire n6035;
wire n6036;
wire n6037;
wire n6038;
wire n6039;
wire n6040;
wire n6041;
wire n6042;
wire n6043;
wire n6044;
wire n6045;
wire n6046;
wire n6047;
wire n6048;
wire n6049;
wire n6050;
wire n6051;
wire n6052;
wire n6053;
wire n6054;
wire n6055;
wire n6056;
wire n6057;
wire n6058;
wire n6059;
wire n6060;
wire n6061;
wire n6062;
wire n6063;
wire n6064;
wire n6065;
wire n6066;
wire n6067;
wire n6068;
wire n6069;
wire n6070;
wire n6071;
wire n6072;
wire n6073;
wire n6074;
wire n6075;
wire n6076;
wire n6077;
wire n6078;
wire n6079;
wire n6080;
wire n6081;
wire n6082;
wire n6083;
wire n6084;
wire n6085;
wire n6086;
wire n6087;
wire n6088;
wire n6089;
wire n6090;
wire n6091;
wire n6092;
wire n6093;
wire n6094;
wire n6095;
wire n6096;
wire n6097;
wire n6098;
wire n6099;
wire n6100;
wire n6101;
wire n6102;
wire n6103;
wire n6104;
wire n6105;
wire n6106;
wire n6107;
wire n6108;
wire n6109;
wire n6110;
wire n6111;
wire n6112;
wire n6113;
wire n6114;
wire n6115;
wire n6116;
wire n6117;
wire n6118;
wire n6119;
wire n6120;
wire n6121;
wire n6122;
wire n6123;
wire n6124;
wire n6125;
wire n6126;
wire n6127;
wire n6128;
wire n6129;
wire n6130;
wire n6131;
wire n6132;
wire n6133;
wire n6134;
wire n6135;
wire n6136;
wire n6137;
wire n6138;
wire n6139;
wire n6140;
wire n6141;
wire n6142;
wire n6143;
wire n6144;
wire n6145;
wire n6146;
wire n6147;
wire n6148;
wire n6149;
wire n6150;
wire n6151;
wire n6152;
wire n6153;
wire n6154;
wire n6155;
wire n6156;
wire n6157;
wire n6158;
wire n6159;
wire n6160;
wire n6161;
wire n6162;
wire n6163;
wire n6164;
wire n6165;
wire n6166;
wire n6167;
wire n6168;
wire n6169;
wire n6170;
wire n6171;
wire n6172;
wire n6173;
wire n6174;
wire n6175;
wire n6176;
wire n6177;
wire n6178;
wire n6179;
wire n6180;
wire n6181;
wire n6182;
wire n6183;
wire n6184;
wire n6185;
wire n6186;
wire n6187;
wire n6188;
wire n6189;
wire n6190;
wire n6191;
wire n6192;
wire n6193;
wire n6194;
wire n6195;
wire n6196;
wire n6197;
wire n6198;
wire n6199;
wire n6200;
wire n6201;
wire n6202;
wire n6203;
wire n6204;
wire n6205;
wire n6206;
wire n6207;
wire n6208;
wire n6209;
wire n6210;
wire n6211;
wire n6212;
wire n6213;
wire n6214;
wire n6215;
wire n6216;
wire n6217;
wire n6218;
wire n6219;
wire n6220;
wire n6221;
wire n6222;
wire n6223;
wire n6224;
wire n6225;
wire n6226;
wire n6227;
wire n6228;
wire n6229;
wire n6230;
wire n6231;
wire n6232;
wire n6233;
wire n6234;
wire n6235;
wire n6236;
wire n6237;
wire n6238;
wire n6239;
wire n6240;
wire n6241;
wire n6242;
wire n6243;
wire n6244;
wire n6245;
wire n6246;
wire n6247;
wire n6248;
wire n6249;
wire n6250;
wire n6251;
wire n6252;
wire n6253;
wire n6254;
wire n6255;
wire n6256;
wire n6257;
wire n6258;
wire n6259;
wire n6260;
wire n6261;
wire n6262;
wire n6263;
wire n6264;
wire n6265;
wire n6266;
wire n6267;
wire n6268;
wire n6269;
wire n6270;
wire n6271;
wire n6272;
wire n6273;
wire n6274;
wire n6275;
wire n6276;
wire n6277;
wire n6278;
wire n6279;
wire n6280;
wire n6281;
wire n6282;
wire n6283;
wire n6284;
wire n6285;
wire n6286;
wire n6287;
wire n6288;
wire n6289;
wire n6290;
wire n6291;
wire n6292;
wire n6293;
wire n6294;
wire n6295;
wire n6296;
wire n6297;
wire n6298;
wire n6299;
wire n6300;
wire n6301;
wire n6302;
wire n6303;
wire n6304;
wire n6305;
wire n6306;
wire n6307;
wire n6308;
wire n6309;
wire n6310;
wire n6311;
wire n6312;
wire n6313;
wire n6314;
wire n6315;
wire n6316;
wire n6317;
wire n6318;
wire n6319;
wire n6320;
wire n6321;
wire n6322;
wire n6323;
wire n6324;
wire n6325;
wire n6326;
wire n6327;
wire n6328;
wire n6329;
wire n6330;
wire n6331;
wire n6332;
wire n6333;
wire n6334;
wire n6335;
wire n6336;
wire n6337;
wire n6338;
wire n6339;
wire n6340;
wire n6341;
wire n6342;
wire n6343;
wire n6344;
wire n6345;
wire n6346;
wire n6347;
wire n6348;
wire n6349;
wire n6350;
wire n6351;
wire n6352;
wire n6353;
wire n6354;
wire n6355;
wire n6356;
wire n6357;
wire n6358;
wire n6359;
wire n6360;
wire n6361;
wire n6362;
wire n6363;
wire n6364;
wire n6365;
wire n6366;
wire n6367;
wire n6368;
wire n6369;
wire n6370;
wire n6371;
wire n6372;
wire n6373;
wire n6374;
wire n6375;
wire n6376;
wire n6377;
wire n6378;
wire n6379;
wire n6380;
wire n6381;
wire n6382;
wire n6383;
wire n6384;
wire n6385;
wire n6386;
wire n6387;
wire n6388;
wire n6389;
wire n6390;
wire n6391;
wire n6392;
wire n6393;
wire n6394;
wire n6395;
wire n6396;
wire n6397;
wire n6398;
wire n6399;
wire n6400;
wire n6401;
wire n6402;
wire n6403;
wire n6404;
wire n6405;
wire n6406;
wire n6407;
wire n6408;
wire n6409;
wire n6410;
wire n6411;
wire n6412;
wire n6413;
wire n6414;
wire n6415;
wire n6416;
wire n6417;
wire n6418;
wire n6419;
wire n6420;
wire n6421;
wire n6422;
wire n6423;
wire n6424;
wire n6425;
wire n6426;
wire n6427;
wire n6428;
wire n6429;
wire n6430;
wire n6431;
wire n6432;
wire n6433;
wire n6434;
wire n6435;
wire n6436;
wire n6437;
wire n6438;
wire n6439;
wire n6440;
wire n6441;
wire n6442;
wire n6443;
wire n6444;
wire n6445;
wire n6446;
wire n6447;
wire n6448;
wire n6449;
wire n6450;
wire n6451;
wire n6452;
wire n6453;
wire n6454;
wire n6455;
wire n6456;
wire n6457;
wire n6458;
wire n6459;
wire n6460;
wire n6461;
wire n6462;
wire n6463;
wire n6464;
wire n6465;
wire n6466;
wire n6467;
wire n6468;
wire n6469;
wire n6470;
wire n6471;
wire n6472;
wire n6473;
wire n6474;
wire n6475;
wire n6476;
wire n6477;
wire n6478;
wire n6479;
wire n6480;
wire n6481;
wire n6482;
wire n6483;
wire n6484;
wire n6485;
wire n6486;
wire n6487;
wire n6488;
wire n6489;
wire n6490;
wire n6491;
wire n6492;
wire n6493;
wire n6494;
wire n6495;
wire n6496;
wire n6497;
wire n6498;
wire n6499;
wire n6500;
wire n6501;
wire n6502;
wire n6503;
wire n6504;
wire n6505;
wire n6506;
wire n6507;
wire n6508;
wire n6509;
wire n6510;
wire n6511;
wire n6512;
wire n6513;
wire n6514;
wire n6515;
wire n6516;
wire n6517;
wire n6518;
wire n6519;
wire n6520;
wire n6521;
wire n6522;
wire n6523;
wire n6524;
wire n6525;
wire n6526;
wire n6527;
wire n6528;
wire n6529;
wire n6530;
wire n6531;
wire n6532;
wire n6533;
wire n6534;
wire n6535;
wire n6536;
wire n6537;
wire n6538;
wire n6539;
wire n6540;
wire n6541;
wire n6542;
wire n6543;
wire n6544;
wire n6545;
wire n6546;
wire n6547;
wire n6548;
wire n6549;
wire n6550;
wire n6551;
wire n6552;
wire n6553;
wire n6554;
wire n6555;
wire n6556;
wire n6557;
wire n6558;
wire n6559;
wire n6560;
wire n6561;
wire n6562;
wire n6563;
wire n6564;
wire n6565;
wire n6566;
wire n6567;
wire n6568;
wire n6569;
wire n6570;
wire n6571;
wire n6572;
wire n6573;
wire n6574;
wire n6575;
wire n6576;
wire n6577;
wire n6578;
wire n6579;
wire n6580;
wire n6581;
wire n6582;
wire n6583;
wire n6584;
wire n6585;
wire n6586;
wire n6587;
wire n6588;
wire n6589;
wire n6590;
wire n6591;
wire n6592;
wire n6593;
wire n6594;
wire n6595;
wire n6596;
wire n6597;
wire n6598;
wire n6599;
wire n6600;
wire n6601;
wire n6602;
wire n6603;
wire n6604;
wire n6605;
wire n6606;
wire n6607;
wire n6608;
wire n6609;
wire n6610;
wire n6611;
wire n6612;
wire n6613;
wire n6614;
wire n6615;
wire n6616;
wire n6617;
wire n6618;
wire n6619;
wire n6620;
wire n6621;
wire n6622;
wire n6623;
wire n6624;
wire n6625;
wire n6626;
wire n6627;
wire n6628;
wire n6629;
wire n6630;
wire n6631;
wire n6632;
wire n6633;
wire n6634;
wire n6635;
wire n6636;
wire n6637;
wire n6638;
wire n6639;
wire n6640;
wire n6641;
wire n6642;
wire n6643;
wire n6644;
wire n6645;
wire n6646;
wire n6647;
wire n6648;
wire n6649;
wire n6650;
wire n6651;
wire n6652;
wire n6653;
wire n6654;
wire n6655;
wire n6656;
wire n6657;
wire n6658;
wire n6659;
wire n6660;
wire n6661;
wire n6662;
wire n6663;
wire n6664;
wire n6665;
wire n6666;
wire n6667;
wire n6668;
wire n6669;
wire n6670;
wire n6671;
wire n6672;
wire n6673;
wire n6674;
wire n6675;
wire n6676;
wire n6677;
wire n6678;
wire n6679;
wire n6680;
wire n6681;
wire n6682;
wire n6683;
wire n6684;
wire n6685;
wire n6686;
wire n6687;
wire n6688;
wire n6689;
wire n6690;
wire n6691;
wire n6692;
wire n6693;
wire n6694;
wire n6695;
wire n6696;
wire n6697;
wire n6698;
wire n6699;
wire n6700;
wire n6701;
wire n6702;
wire n6703;
wire n6704;
wire n6705;
wire n6706;
wire n6707;
wire n6708;
wire n6709;
wire n6710;
wire n6711;
wire n6712;
wire n6713;
wire n6714;
wire n6715;
wire n6716;
wire n6717;
wire n6718;
wire n6719;
wire n6720;
wire n6721;
wire n6722;
wire n6723;
wire n6724;
wire n6725;
wire n6726;
wire n6727;
wire n6728;
wire n6729;
wire n6730;
wire n6731;
wire n6732;
wire n6733;
wire n6734;
wire n6735;
wire n6736;
wire n6737;
wire n6738;
wire n6739;
wire n6740;
wire n6741;
wire n6742;
wire n6743;
wire n6744;
wire n6745;
wire n6746;
wire n6747;
wire n6748;
wire n6749;
wire n6750;
wire n6751;
wire n6752;
wire n6753;
wire n6754;
wire n6755;
wire n6756;
wire n6757;
wire n6758;
wire n6759;
wire n6760;
wire n6761;
wire n6762;
wire n6763;
wire n6764;
wire n6765;
wire n6766;
wire n6767;
wire n6768;
wire n6769;
wire n6770;
wire n6771;
wire n6772;
wire n6773;
wire n6774;
wire n6775;
wire n6776;
wire n6777;
wire n6778;
wire n6779;
wire n6780;
wire n6781;
wire n6782;
wire n6783;
wire n6784;
wire n6785;
wire n6786;
wire n6787;
wire n6788;
wire n6789;
wire n6790;
wire n6791;
wire n6792;
wire n6793;
wire n6794;
wire n6795;
wire n6796;
wire n6797;
wire n6798;
wire n6799;
wire n6800;
wire n6801;
wire n6802;
wire n6803;
wire n6804;
wire n6805;
wire n6806;
wire n6807;
wire n6808;
wire n6809;
wire n6810;
wire n6811;
wire n6812;
wire n6813;
wire n6814;
wire n6815;
wire n6816;
wire n6817;
wire n6818;
wire n6819;
wire n6820;
wire n6821;
wire n6822;
wire n6823;
wire n6824;
wire n6825;
wire n6826;
wire n6827;
wire n6828;
wire n6829;
wire n6830;
wire n6831;
wire n6832;
wire n6833;
wire n6834;
wire n6835;
wire n6836;
wire n6837;
wire n6838;
wire n6839;
wire n6840;
wire n6841;
wire n6842;
wire n6843;
wire n6844;
wire n6845;
wire n6846;
wire n6847;
wire n6848;
wire n6849;
wire n6850;
wire n6851;
wire n6852;
wire n6853;
wire n6854;
wire n6855;
wire n6856;
wire n6857;
wire n6858;
wire n6859;
wire n6860;
wire n6861;
wire n6862;
wire n6863;
wire n6864;
wire n6865;
wire n6866;
wire n6867;
wire n6868;
wire n6869;
wire n6870;
wire n6871;
wire n6872;
wire n6873;
wire n6874;
wire n6875;
wire n6876;
wire n6877;
wire n6878;
wire n6879;
wire n6880;
wire n6881;
wire n6882;
wire n6883;
wire n6884;
wire n6885;
wire n6886;
wire n6887;
wire n6888;
wire n6889;
wire n6890;
wire n6891;
wire n6892;
wire n6893;
wire n6894;
wire n6895;
wire n6896;
wire n6897;
wire n6898;
wire n6899;
wire n6900;
wire n6901;
wire n6902;
wire n6903;
wire n6904;
wire n6905;
wire n6906;
wire n6907;
wire n6908;
wire n6909;
wire n6910;
wire n6911;
wire n6912;
wire n6913;
wire n6914;
wire n6915;
wire n6916;
wire n6917;
wire n6918;
wire n6919;
wire n6920;
wire n6921;
wire n6922;
wire n6923;
wire n6924;
wire n6925;
wire n6926;
wire n6927;
wire n6928;
wire n6929;
wire n6930;
wire n6931;
wire n6932;
wire n6933;
wire n6934;
wire n6935;
wire n6936;
wire n6937;
wire n6938;
wire n6939;
wire n6940;
wire n6941;
wire n6942;
wire n6943;
wire n6944;
wire n6945;
wire n6946;
wire n6947;
wire n6948;
wire n6949;
wire n6950;
wire n6951;
wire n6952;
wire n6953;
wire n6954;
wire n6955;
wire n6956;
wire n6957;
wire n6958;
wire n6959;
wire n6960;
wire n6961;
wire n6962;
wire n6963;
wire n6964;
wire n6965;
wire n6966;
wire n6967;
wire n6968;
wire n6969;
wire n6970;
wire n6971;
wire n6972;
wire n6973;
wire n6974;
wire n6975;
wire n6976;
wire n6977;
wire n6978;
wire n6979;
wire n6980;
wire n6981;
wire n6982;
wire n6983;
wire n6984;
wire n6985;
wire n6986;
wire n6987;
wire n6988;
wire n6989;
wire n6990;
wire n6991;
wire n6992;
wire n6993;
wire n6994;
wire n6995;
wire n6996;
wire n6997;
wire n6998;
wire n6999;
wire n7000;
wire n7001;
wire n7002;
wire n7003;
wire n7004;
wire n7005;
wire n7006;
wire n7007;
wire n7008;
wire n7009;
wire n7010;
wire n7011;
wire n7012;
wire n7013;
wire n7014;
wire n7015;
wire n7016;
wire n7017;
wire n7018;
wire n7019;
wire n7020;
wire n7021;
wire n7022;
wire n7023;
wire n7024;
wire n7025;
wire n7026;
wire n7027;
wire n7028;
wire n7029;
wire n7030;
wire n7031;
wire n7032;
wire n7033;
wire n7034;
wire n7035;
wire n7036;
wire n7037;
wire n7038;
wire n7039;
wire n7040;
wire n7041;
wire n7042;
wire n7043;
wire n7044;
wire n7045;
wire n7046;
wire n7047;
wire n7048;
wire n7049;
wire n7050;
wire n7051;
wire n7052;
wire n7053;
wire n7054;
wire n7055;
wire n7056;
wire n7057;
wire n7058;
wire n7059;
wire n7060;
wire n7061;
wire n7062;
wire n7063;
wire n7064;
wire n7065;
wire n7066;
wire n7067;
wire n7068;
wire n7069;
wire n7070;
wire n7071;
wire n7072;
wire n7073;
wire n7074;
wire n7075;
wire n7076;
wire n7077;
wire n7078;
wire n7079;
wire n7080;
wire n7081;
wire n7082;
wire n7083;
wire n7084;
wire n7085;
wire n7086;
wire n7087;
wire n7088;
wire n7089;
wire n7090;
wire n7091;
wire n7092;
wire n7093;
wire n7094;
wire n7095;
wire n7096;
wire n7097;
wire n7098;
wire n7099;
wire n7100;
wire n7101;
wire n7102;
wire n7103;
wire n7104;
wire n7105;
wire n7106;
wire n7107;
wire n7108;
wire n7109;
wire n7110;
wire n7111;
wire n7112;
wire n7113;
wire n7114;
wire n7115;
wire n7116;
wire n7117;
wire n7118;
wire n7119;
wire n7120;
wire n7121;
wire n7122;
wire n7123;
wire n7124;
wire n7125;
wire n7126;
wire n7127;
wire n7128;
wire n7129;
wire n7130;
wire n7131;
wire n7132;
wire n7133;
wire n7134;
wire n7135;
wire n7136;
wire n7137;
wire n7138;
wire n7139;
wire n7140;
wire n7141;
wire n7142;
wire n7143;
wire n7144;
wire n7145;
wire n7146;
wire n7147;
wire n7148;
wire n7149;
wire n7150;
wire n7151;
wire n7152;
wire n7153;
wire n7154;
wire n7155;
wire n7156;
wire n7157;
wire n7158;
wire n7159;
wire n7160;
wire n7161;
wire n7162;
wire n7163;
wire n7164;
wire n7165;
wire n7166;
wire n7167;
wire n7168;
wire n7169;
wire n7170;
wire n7171;
wire n7172;
wire n7173;
wire n7174;
wire n7175;
wire n7176;
wire n7177;
wire n7178;
wire n7179;
wire n7180;
wire n7181;
wire n7182;
wire n7183;
wire n7184;
wire n7185;
wire n7186;
wire n7187;
wire n7188;
wire n7189;
wire n7190;
wire n7191;
wire n7192;
wire n7193;
wire n7194;
wire n7195;
wire n7196;
wire n7197;
wire n7198;
wire n7199;
wire n7200;
wire n7201;
wire n7202;
wire n7203;
wire n7204;
wire n7205;
wire n7206;
wire n7207;
wire n7208;
wire n7209;
wire n7210;
wire n7211;
wire n7212;
wire n7213;
wire n7214;
wire n7215;
wire n7216;
wire n7217;
wire n7218;
wire n7219;
wire n7220;
wire n7221;
wire n7222;
wire n7223;
wire n7224;
wire n7225;
wire n7226;
wire n7227;
wire n7228;
wire n7229;
wire n7230;
wire n7231;
wire n7232;
wire n7233;
wire n7234;
wire n7235;
wire n7236;
wire n7237;
wire n7238;
wire n7239;
wire n7240;
wire n7241;
wire n7242;
wire n7243;
wire n7244;
wire n7245;
wire n7246;
wire n7247;
wire n7248;
wire n7249;
wire n7250;
wire n7251;
wire n7252;
wire n7253;
wire n7254;
wire n7255;
wire n7256;
wire n7257;
wire n7258;
wire n7259;
wire n7260;
wire n7261;
wire n7262;
wire n7263;
wire n7264;
wire n7265;
wire n7266;
wire n7267;
wire n7268;
wire n7269;
wire n7270;
wire n7271;
wire n7272;
wire n7273;
wire n7274;
wire n7275;
wire n7276;
wire n7277;
wire n7278;
wire n7279;
wire n7280;
wire n7281;
wire n7282;
wire n7283;
wire n7284;
wire n7285;
wire n7286;
wire n7287;
wire n7288;
wire n7289;
wire n7290;
wire n7291;
wire n7292;
wire n7293;
wire n7294;
wire n7295;
wire n7296;
wire n7297;
wire n7298;
wire n7299;
wire n7300;
wire n7301;
wire n7302;
wire n7303;
wire n7304;
wire n7305;
wire n7306;
wire n7307;
wire n7308;
wire n7309;
wire n7310;
wire n7311;
wire n7312;
wire n7313;
wire n7314;
wire n7315;
wire n7316;
wire n7317;
wire n7318;
wire n7319;
wire n7320;
wire n7321;
wire n7322;
wire n7323;
wire n7324;
wire n7325;
wire n7326;
wire n7327;
wire n7328;
wire n7329;
wire n7330;
wire n7331;
wire n7332;
wire n7333;
wire n7334;
wire n7335;
wire n7336;
wire n7337;
wire n7338;
wire n7339;
wire n7340;
wire n7341;
wire n7342;
wire n7343;
wire n7344;
wire n7345;
wire n7346;
wire n7347;
wire n7348;
wire n7349;
wire n7350;
wire n7351;
wire n7352;
wire n7353;
wire n7354;
wire n7355;
wire n7356;
wire n7357;
wire n7358;
wire n7359;
wire n7360;
wire n7361;
wire n7362;
wire n7363;
wire n7364;
wire n7365;
wire n7366;
wire n7367;
wire n7368;
wire n7369;
wire n7370;
wire n7371;
wire n7372;
wire n7373;
wire n7374;
wire n7375;
wire n7376;
wire n7377;
wire n7378;
wire n7379;
wire n7380;
wire n7381;
wire n7382;
wire n7383;
wire n7384;
wire n7385;
wire n7386;
wire n7387;
wire n7388;
wire n7389;
wire n7390;
wire n7391;
wire n7392;
wire n7393;
wire n7394;
wire n7395;
wire n7396;
wire n7397;
wire n7398;
wire n7399;
wire n7400;
wire n7401;
wire n7402;
wire n7403;
wire n7404;
wire n7405;
wire n7406;
wire n7407;
wire n7408;
wire n7409;
wire n7410;
wire n7411;
wire n7412;
wire n7413;
wire n7414;
wire n7415;
wire n7416;
wire n7417;
wire n7418;
wire n7419;
wire n7420;
wire n7421;
wire n7422;
wire n7423;
wire n7424;
wire n7425;
wire n7426;
wire n7427;
wire n7428;
wire n7429;
wire n7430;
wire n7431;
wire n7432;
wire n7433;
wire n7434;
wire n7435;
wire n7436;
wire n7437;
wire n7438;
wire n7439;
wire n7440;
wire n7441;
wire n7442;
wire n7443;
wire n7444;
wire n7445;
wire n7446;
wire n7447;
wire n7448;
wire n7449;
wire n7450;
wire n7451;
wire n7452;
wire n7453;
wire n7454;
wire n7455;
wire n7456;
wire n7457;
wire n7458;
wire n7459;
wire n7460;
wire n7461;
wire n7462;
wire n7463;
wire n7464;
wire n7465;
wire n7466;
wire n7467;
wire n7468;
wire n7469;
wire n7470;
wire n7471;
wire n7472;
wire n7473;
wire n7474;
wire n7475;
wire n7476;
wire n7477;
wire n7478;
wire n7479;
wire n7480;
wire n7481;
wire n7482;
wire n7483;
wire n7484;
wire n7485;
wire n7486;
wire n7487;
wire n7488;
wire n7489;
wire n7490;
wire n7491;
wire n7492;
wire n7493;
wire n7494;
wire n7495;
wire n7496;
wire n7497;
wire n7498;
wire n7499;
wire n7500;
wire n7501;
wire n7502;
wire n7503;
wire n7504;
wire n7505;
wire n7506;
wire n7507;
wire n7508;
wire n7509;
wire n7510;
wire n7511;
wire n7512;
wire n7513;
wire n7514;
wire n7515;
wire n7516;
wire n7517;
wire n7518;
wire n7519;
wire n7520;
wire n7521;
wire n7522;
wire n7523;
wire n7524;
wire n7525;
wire n7526;
wire n7527;
wire n7528;
wire n7529;
wire n7530;
wire n7531;
wire n7532;
wire n7533;
wire n7534;
wire n7535;
wire n7536;
wire n7537;
wire n7538;
wire n7539;
wire n7540;
wire n7541;
wire n7542;
wire n7543;
wire n7544;
wire n7545;
wire n7546;
wire n7547;
wire n7548;
wire n7549;
wire n7550;
wire n7551;
wire n7552;
wire n7553;
wire n7554;
wire n7555;
wire n7556;
wire n7557;
wire n7558;
wire n7559;
wire n7560;
wire n7561;
wire n7562;
wire n7563;
wire n7564;
wire n7565;
wire n7566;
wire n7567;
wire n7568;
wire n7569;
wire n7570;
wire n7571;
wire n7572;
wire n7573;
wire n7574;
wire n7575;
wire n7576;
wire n7577;
wire n7578;
wire n7579;
wire n7580;
wire n7581;
wire n7582;
wire n7583;
wire n7584;
wire n7585;
wire n7586;
wire n7587;
wire n7588;
wire n7589;
wire n7590;
wire n7591;
wire n7592;
wire n7593;
wire n7594;
wire n7595;
wire n7596;
wire n7597;
wire n7598;
wire n7599;
wire n7600;
wire n7601;
wire n7602;
wire n7603;
wire n7604;
wire n7605;
wire n7606;
wire n7607;
wire n7608;
wire n7609;
wire n7610;
wire n7611;
wire n7612;
wire n7613;
wire n7614;
wire n7615;
wire n7616;
wire n7617;
wire n7618;
wire n7619;
wire n7620;
wire n7621;
wire n7622;
wire n7623;
wire n7624;
wire n7625;
wire n7626;
wire n7627;
wire n7628;
wire n7629;
wire n7630;
wire n7631;
wire n7632;
wire n7633;
wire n7634;
wire n7635;
wire n7636;
wire n7637;
wire n7638;
wire n7639;
wire n7640;
wire n7641;
wire n7642;
wire n7643;
wire n7644;
wire n7645;
wire n7646;
wire n7647;
wire n7648;
wire n7649;
wire n7650;
wire n7651;
wire n7652;
wire n7653;
wire n7654;
wire n7655;
wire n7656;
wire n7657;
wire n7658;
wire n7659;
wire n7660;
wire n7661;
wire n7662;
wire n7663;
wire n7664;
wire n7665;
wire n7666;
wire n7667;
wire n7668;
wire n7669;
wire n7670;
wire n7671;
wire n7672;
wire n7673;
wire n7674;
wire n7675;
wire n7676;
wire n7677;
wire n7678;
wire n7679;
wire n7680;
wire n7681;
wire n7682;
wire n7683;
wire n7684;
wire n7685;
wire n7686;
wire n7687;
wire n7688;
wire n7689;
wire n7690;
wire n7691;
wire n7692;
wire n7693;
wire n7694;
wire n7695;
wire n7696;
wire n7697;
wire n7698;
wire n7699;
wire n7700;
wire n7701;
wire n7702;
wire n7703;
wire n7704;
wire n7705;
wire n7706;
wire n7707;
wire n7708;
wire n7709;
wire n7710;
wire n7711;
wire n7712;
wire n7713;
wire n7714;
wire n7715;
wire n7716;
wire n7717;
wire n7718;
wire n7719;
wire n7720;
wire n7721;
wire n7722;
wire n7723;
wire n7724;
wire n7725;
wire n7726;
wire n7727;
wire n7728;
wire n7729;
wire n7730;
wire n7731;
wire n7732;
wire n7733;
wire n7734;
wire n7735;
wire n7736;
wire n7737;
wire n7738;
wire n7739;
wire n7740;
wire n7741;
wire n7742;
wire n7743;
wire n7744;
wire n7745;
wire n7746;
wire n7747;
wire n7748;
wire n7749;
wire n7750;
wire n7751;
wire n7752;
wire n7753;
wire n7754;
wire n7755;
wire n7756;
wire n7757;
wire n7758;
wire n7759;
wire n7760;
wire n7761;
wire n7762;
wire n7763;
wire n7764;
wire n7765;
wire n7766;
wire n7767;
wire n7768;
wire n7769;
wire n7770;
wire n7771;
wire n7772;
wire n7773;
wire n7774;
wire n7775;
wire n7776;
wire n7777;
wire n7778;
wire n7779;
wire n7780;
wire n7781;
wire n7782;
wire n7783;
wire n7784;
wire n7785;
wire n7786;
wire n7787;
wire n7788;
wire n7789;
wire n7790;
wire n7791;
wire n7792;
wire n7793;
wire n7794;
wire n7795;
wire n7796;
wire n7797;
wire n7798;
wire n7799;
wire n7800;
wire n7801;
wire n7802;
wire n7803;
wire n7804;
wire n7805;
wire n7806;
wire n7807;
wire n7808;
wire n7809;
wire n7810;
wire n7811;
wire n7812;
wire n7813;
wire n7814;
wire n7815;
wire n7816;
wire n7817;
wire n7818;
wire n7819;
wire n7820;
wire n7821;
wire n7822;
wire n7823;
wire n7824;
wire n7825;
wire n7826;
wire n7827;
wire n7828;
wire n7829;
wire n7830;
wire n7831;
wire n7832;
wire n7833;
wire n7834;
wire n7835;
wire n7836;
wire n7837;
wire n7838;
wire n7839;
wire n7840;
wire n7841;
wire n7842;
wire n7843;
wire n7844;
wire n7845;
wire n7846;
wire n7847;
wire n7848;
wire n7849;
wire n7850;
wire n7851;
wire n7852;
wire n7853;
wire n7854;
wire n7855;
wire n7856;
wire n7857;
wire n7858;
wire n7859;
wire n7860;
wire n7861;
wire n7862;
wire n7863;
wire n7864;
wire n7865;
wire n7866;
wire n7867;
wire n7868;
wire n7869;
wire n7870;
wire n7871;
wire n7872;
wire n7873;
wire n7874;
wire n7875;
wire n7876;
wire n7877;
wire n7878;
wire n7879;
wire n7880;
wire n7881;
wire n7882;
wire n7883;
wire n7884;
wire n7885;
wire n7886;
wire n7887;
wire n7888;
wire n7889;
wire n7890;
wire n7891;
wire n7892;
wire n7893;
wire n7894;
wire n7895;
wire n7896;
wire n7897;
wire n7898;
wire n7899;
wire n7900;
wire n7901;
wire n7902;
wire n7903;
wire n7904;
wire n7905;
wire n7906;
wire n7907;
wire n7908;
wire n7909;
wire n7910;
wire n7911;
wire n7912;
wire n7913;
wire n7914;
wire n7915;
wire n7916;
wire n7917;
wire n7918;
wire n7919;
wire n7920;
wire n7921;
wire n7922;
wire n7923;
wire n7924;
wire n7925;
wire n7926;
wire n7927;
wire n7928;
wire n7929;
wire n7930;
wire n7931;
wire n7932;
wire n7933;
wire n7934;
wire n7935;
wire n7936;
wire n7937;
wire n7938;
wire n7939;
wire n7940;
wire n7941;
wire n7942;
wire n7943;
wire n7944;
wire n7945;
wire n7946;
wire n7947;
wire n7948;
wire n7949;
wire n7950;
wire n7951;
wire n7952;
wire n7953;
wire n7954;
wire n7955;
wire n7956;
wire n7957;
wire n7958;
wire n7959;
wire n7960;
wire n7961;
wire n7962;
wire n7963;
wire n7964;
wire n7965;
wire n7966;
wire n7967;
wire n7968;
wire n7969;
wire n7970;
wire n7971;
wire n7972;
wire n7973;
wire n7974;
wire n7975;
wire n7976;
wire n7977;
wire n7978;
wire n7979;
wire n7980;
wire n7981;
wire n7982;
wire n7983;
wire n7984;
wire n7985;
wire n7986;
wire n7987;
wire n7988;
wire n7989;
wire n7990;
wire n7991;
wire n7992;
wire n7993;
wire n7994;
wire n7995;
wire n7996;
wire n7997;
wire n7998;
wire n7999;
wire n8000;
wire n8001;
wire n8002;
wire n8003;
wire n8004;
wire n8005;
wire n8006;
wire n8007;
wire n8008;
wire n8009;
wire n8010;
wire n8011;
wire n8012;
wire n8013;
wire n8014;
wire n8015;
wire n8016;
wire n8017;
wire n8018;
wire n8019;
wire n8020;
wire n8021;
wire n8022;
wire n8023;
wire n8024;
wire n8025;
wire n8026;
wire n8027;
wire n8028;
wire n8029;
wire n8030;
wire n8031;
wire n8032;
wire n8033;
wire n8034;
wire n8035;
wire n8036;
wire n8037;
wire n8038;
wire n8039;
wire n8040;
wire n8041;
wire n8042;
wire n8043;
wire n8044;
wire n8045;
wire n8046;
wire n8047;
wire n8048;
wire n8049;
wire n8050;
wire n8051;
wire n8052;
wire n8053;
wire n8054;
wire n8055;
wire n8056;
wire n8057;
wire n8058;
wire n8059;
wire n8060;
wire n8061;
wire n8062;
wire n8063;
wire n8064;
wire n8065;
wire n8066;
wire n8067;
wire n8068;
wire n8069;
wire n8070;
wire n8071;
wire n8072;
wire n8073;
wire n8074;
wire n8075;
wire n8076;
wire n8077;
wire n8078;
wire n8079;
wire n8080;
wire n8081;
wire n8082;
wire n8083;
wire n8084;
wire n8085;
wire n8086;
wire n8087;
wire n8088;
wire n8089;
wire n8090;
wire n8091;
wire n8092;
wire n8093;
wire n8094;
wire n8095;
wire n8096;
wire n8097;
wire n8098;
wire n8099;
wire n8100;
wire n8101;
wire n8102;
wire n8103;
wire n8104;
wire n8105;
wire n8106;
wire n8107;
wire n8108;
wire n8109;
wire n8110;
wire n8111;
wire n8112;
wire n8113;
wire n8114;
wire n8115;
wire n8116;
wire n8117;
wire n8118;
wire n8119;
wire n8120;
wire n8121;
wire n8122;
wire n8123;
wire n8124;
wire n8125;
wire n8126;
wire n8127;
wire n8128;
wire n8129;
wire n8130;
wire n8131;
wire n8132;
wire n8133;
wire n8134;
wire n8135;
wire n8136;
wire n8137;
wire n8138;
wire n8139;
wire n8140;
wire n8141;
wire n8142;
wire n8143;
wire n8144;
wire n8145;
wire n8146;
wire n8147;
wire n8148;
wire n8149;
wire n8150;
wire n8151;
wire n8152;
wire n8153;
wire n8154;
wire n8155;
wire n8156;
wire n8157;
wire n8158;
wire n8159;
wire n8160;
wire n8161;
wire n8162;
wire n8163;
wire n8164;
wire n8165;
wire n8166;
wire n8167;
wire n8168;
wire n8169;
wire n8170;
wire n8171;
wire n8172;
wire n8173;
wire n8174;
wire n8175;
wire n8176;
wire n8177;
wire n8178;
wire n8179;
wire n8180;
wire n8181;
wire n8182;
wire n8183;
wire n8184;
wire n8185;
wire n8186;
wire n8187;
wire n8188;
wire n8189;
wire n8190;
wire n8191;
wire n8192;
wire n8193;
wire n8194;
wire n8195;
wire n8196;
wire n8197;
wire n8198;
wire n8199;
wire n8200;
wire n8201;
wire n8202;
wire n8203;
wire n8204;
wire n8205;
wire n8206;
wire n8207;
wire n8208;
wire n8209;
wire n8210;
wire n8211;
wire n8212;
wire n8213;
wire n8214;
wire n8215;
wire n8216;
wire n8217;
wire n8218;
wire n8219;
wire n8220;
wire n8221;
wire n8222;
wire n8223;
wire n8224;
wire n8225;
wire n8226;
wire n8227;
wire n8228;
wire n8229;
wire n8230;
wire n8231;
wire n8232;
wire n8233;
wire n8234;
wire n8235;
wire n8236;
wire n8237;
wire n8238;
wire n8239;
wire n8240;
wire n8241;
wire n8242;
wire n8243;
wire n8244;
wire n8245;
wire n8246;
wire n8247;
wire n8248;
wire n8249;
wire n8250;
wire n8251;
wire n8252;
wire n8253;
wire n8254;
wire n8255;
wire n8256;
wire n8257;
wire n8258;
wire n8259;
wire n8260;
wire n8261;
wire n8262;
wire n8263;
wire n8264;
wire n8265;
wire n8266;
wire n8267;
wire n8268;
wire n8269;
wire n8270;
wire n8271;
wire n8272;
wire n8273;
wire n8274;
wire n8275;
wire n8276;
wire n8277;
wire n8278;
wire n8279;
wire n8280;
wire n8281;
wire n8282;
wire n8283;
wire n8284;
wire n8285;
wire n8286;
wire n8287;
wire n8288;
wire n8289;
wire n8290;
wire n8291;
wire n8292;
wire n8293;
wire n8294;
wire n8295;
wire n8296;
wire n8297;
wire n8298;
wire n8299;
wire n8300;
wire n8301;
wire n8302;
wire n8303;
wire n8304;
wire n8305;
wire n8306;
wire n8307;
wire n8308;
wire n8309;
wire n8310;
wire n8311;
wire n8312;
wire n8313;
wire n8314;
wire n8315;
wire n8316;
wire n8317;
wire n8318;
wire n8319;
wire n8320;
wire n8321;
wire n8322;
wire n8323;
wire n8324;
wire n8325;
wire n8326;
wire n8327;
wire n8328;
wire n8329;
wire n8330;
wire n8331;
wire n8332;
wire n8333;
wire n8334;
wire n8335;
wire n8336;
wire n8337;
wire n8338;
wire n8339;
wire n8340;
wire n8341;
wire n8342;
wire n8343;
wire n8344;
wire n8345;
wire n8346;
wire n8347;
wire n8348;
wire n8349;
wire n8350;
wire n8351;
wire n8352;
wire n8353;
wire n8354;
wire n8355;
wire n8356;
wire n8357;
wire n8358;
wire n8359;
wire n8360;
wire n8361;
wire n8362;
wire n8363;
wire n8364;
wire n8365;
wire n8366;
wire n8367;
wire n8368;
wire n8369;
wire n8370;
wire n8371;
wire n8372;
wire n8373;
wire n8374;
wire n8375;
wire n8376;
wire n8377;
wire n8378;
wire n8379;
wire n8380;
wire n8381;
wire n8382;
wire n8383;
wire n8384;
wire n8385;
wire n8386;
wire n8387;
wire n8388;
wire n8389;
wire n8390;
wire n8391;
wire n8392;
wire n8393;
wire n8394;
wire n8395;
wire n8396;
wire n8397;
wire n8398;
wire n8399;
wire n8400;
wire n8401;
wire n8402;
wire n8403;
wire n8404;
wire n8405;
wire n8406;
wire n8407;
wire n8408;
wire n8409;
wire n8410;
wire n8411;
wire n8412;
wire n8413;
wire n8414;
wire n8415;
wire n8416;
wire n8417;
wire n8418;
wire n8419;
wire n8420;
wire n8421;
wire n8422;
wire n8423;
wire n8424;
wire n8425;
wire n8426;
wire n8427;
wire n8428;
wire n8429;
wire n8430;
wire n8431;
wire n8432;
wire n8433;
wire n8434;
wire n8435;
wire n8436;
wire n8437;
wire n8438;
wire n8439;
wire n8440;
wire n8441;
wire n8442;
wire n8443;
wire n8444;
wire n8445;
wire n8446;
wire n8447;
wire n8448;
wire n8449;
wire n8450;
wire n8451;
wire n8452;
wire n8453;
wire n8454;
wire n8455;
wire n8456;
wire n8457;
wire n8458;
wire n8459;
wire n8460;
wire n8461;
wire n8462;
wire n8463;
wire n8464;
wire n8465;
wire n8466;
wire n8467;
wire n8468;
wire n8469;
wire n8470;
wire n8471;
wire n8472;
wire n8473;
wire n8474;
wire n8475;
wire n8476;
wire n8477;
wire n8478;
wire n8479;
wire n8480;
wire n8481;
wire n8482;
wire n8483;
wire n8484;
wire n8485;
wire n8486;
wire n8487;
wire n8488;
wire n8489;
wire n8490;
wire n8491;
wire n8492;
wire n8493;
wire n8494;
wire n8495;
wire n8496;
wire n8497;
wire n8498;
wire n8499;
wire n8500;
wire n8501;
wire n8502;
wire n8503;
wire n8504;
wire n8505;
wire n8506;
wire n8507;
wire n8508;
wire n8509;
wire n8510;
wire n8511;
wire n8512;
wire n8513;
wire n8514;
wire n8515;
wire n8516;
wire n8517;
wire n8518;
wire n8519;
wire n8520;
wire n8521;
wire n8522;
wire n8523;
wire n8524;
wire n8525;
wire n8526;
wire n8527;
wire n8528;
wire n8529;
wire n8530;
wire n8531;
wire n8532;
wire n8533;
wire n8534;
wire n8535;
wire n8536;
wire n8537;
wire n8538;
wire n8539;
wire n8540;
wire n8541;
wire n8542;
wire n8543;
wire n8544;
wire n8545;
wire n8546;
wire n8547;
wire n8548;
wire n8549;
wire n8550;
wire n8551;
wire n8552;
wire n8553;
wire n8554;
wire n8555;
wire n8556;
wire n8557;
wire n8558;
wire n8559;
wire n8560;
wire n8561;
wire n8562;
wire n8563;
wire n8564;
wire n8565;
wire n8566;
wire n8567;
wire n8568;
wire n8569;
wire n8570;
wire n8571;
wire n8572;
wire n8573;
wire n8574;
wire n8575;
wire n8576;
wire n8577;
wire n8578;
wire n8579;
wire n8580;
wire n8581;
wire n8582;
wire n8583;
wire n8584;
wire n8585;
wire n8586;
wire n8587;
wire n8588;
wire n8589;
wire n8590;
wire n8591;
wire n8592;
wire n8593;
wire n8594;
wire n8595;
wire n8596;
wire n8597;
wire n8598;
wire n8599;
wire n8600;
wire n8601;
wire n8602;
wire n8603;
wire n8604;
wire n8605;
wire n8606;
wire n8607;
wire n8608;
wire n8609;
wire n8610;
wire n8611;
wire n8612;
wire n8613;
wire n8614;
wire n8615;
wire n8616;
wire n8617;
wire n8618;
wire n8619;
wire n8620;
wire n8621;
wire n8622;
wire n8623;
wire n8624;
wire n8625;
wire n8626;
wire n8627;
wire n8628;
wire n8629;
wire n8630;
wire n8631;
wire n8632;
wire n8633;
wire n8634;
wire n8635;
wire n8636;
wire n8637;
wire n8638;
wire n8639;
wire n8640;
wire n8641;
wire n8642;
wire n8643;
wire n8644;
wire n8645;
wire n8646;
wire n8647;
wire n8648;
wire n8649;
wire n8650;
wire n8651;
wire n8652;
wire n8653;
wire n8654;
wire n8655;
wire n8656;
wire n8657;
wire n8658;
wire n8659;
wire n8660;
wire n8661;
wire n8662;
wire n8663;
wire n8664;
wire n8665;
wire n8666;
wire n8667;
wire n8668;
wire n8669;
wire n8670;
wire n8671;
wire n8672;
wire n8673;
wire n8674;
wire n8675;
wire n8676;
wire n8677;
wire n8678;
wire n8679;
wire n8680;
wire n8681;
wire n8682;
wire n8683;
wire n8684;
wire n8685;
wire n8686;
wire n8687;
wire n8688;
wire n8689;
wire n8690;
wire n8691;
wire n8692;
wire n8693;
wire n8694;
wire n8695;
wire n8696;
wire n8697;
wire n8698;
wire n8699;
wire n8700;
wire n8701;
wire n8702;
wire n8703;
wire n8704;
wire n8705;
wire n8706;
wire n8707;
wire n8708;
wire n8709;
wire n8710;
wire n8711;
wire n8712;
wire n8713;
wire n8714;
wire n8715;
wire n8716;
wire n8717;
wire n8718;
wire n8719;
wire n8720;
wire n8721;
wire n8722;
wire n8723;
wire n8724;
wire n8725;
wire n8726;
wire n8727;
wire n8728;
wire n8729;
wire n8730;
wire n8731;
wire n8732;
wire n8733;
wire n8734;
wire n8735;
wire n8736;
wire n8737;
wire n8738;
wire n8739;
wire n8740;
wire n8741;
wire n8742;
wire n8743;
wire n8744;
wire n8745;
wire n8746;
wire n8747;
wire n8748;
wire n8749;
wire n8750;
wire n8751;
wire n8752;
wire n8753;
wire n8754;
wire n8755;
wire n8756;
wire n8757;
wire n8758;
wire n8759;
wire n8760;
wire n8761;
wire n8762;
wire n8763;
wire n8764;
wire n8765;
wire n8766;
wire n8767;
wire n8768;
wire n8769;
wire n8770;
wire n8771;
wire n8772;
wire n8773;
wire n8774;
wire n8775;
wire n8776;
wire n8777;
wire n8778;
wire n8779;
wire n8780;
wire n8781;
wire n8782;
wire n8783;
wire n8784;
wire n8785;
wire n8786;
wire n8787;
wire n8788;
wire n8789;
wire n8790;
wire n8791;
wire n8792;
wire n8793;
wire n8794;
wire n8795;
wire n8796;
wire n8797;
wire n8798;
wire n8799;
wire n8800;
wire n8801;
wire n8802;
wire n8803;
wire n8804;
wire n8805;
wire n8806;
wire n8807;
wire n8808;
wire n8809;
wire n8810;
wire n8811;
wire n8812;
wire n8813;
wire n8814;
wire n8815;
wire n8816;
wire n8817;
wire n8818;
wire n8819;
wire n8820;
wire n8821;
wire n8822;
wire n8823;
wire n8824;
wire n8825;
wire n8826;
wire n8827;
wire n8828;
wire n8829;
wire n8830;
wire n8831;
wire n8832;
wire n8833;
wire n8834;
wire n8835;
wire n8836;
wire n8837;
wire n8838;
wire n8839;
wire n8840;
wire n8841;
wire n8842;
wire n8843;
wire n8844;
wire n8845;
wire n8846;
wire n8847;
wire n8848;
wire n8849;
wire n8850;
wire n8851;
wire n8852;
wire n8853;
wire n8854;
wire n8855;
xor (out,n0,n4671);
or (n0,n1,n8);
and (n1,n2,n7);
not (n2,n3);
nor (n3,n4,n6);
not (n4,n5);
and (n8,n3,n9);
nand (n9,n10,n4670);
or (n10,n11,n2014);
nand (n11,n12,n2013);
not (n12,n13);
nor (n13,n14,n1848);
or (n14,n15,n1847);
and (n15,n16,n1509);
xor (n16,n17,n1059);
or (n17,n18,n1058);
and (n18,n19,n985);
xor (n19,n20,n524);
xor (n20,n21,n404);
xor (n21,n22,n255);
or (n22,n23,n254);
and (n23,n24,n180);
xor (n24,n25,n99);
xor (n25,n26,n71);
xor (n26,n27,n43);
not (n27,n28);
nor (n28,n29,n34);
and (n29,n30,n37);
not (n30,n31);
nand (n31,n32,n36);
or (n32,n33,n34);
not (n34,n35);
nand (n36,n34,n33);
nor (n37,n38,n41);
and (n38,n39,n40);
not (n40,n33);
and (n41,n42,n33);
not (n42,n39);
nand (n43,n44,n65);
or (n44,n45,n53);
not (n45,n46);
nor (n46,n47,n52);
and (n47,n48,n50);
not (n48,n49);
not (n50,n51);
and (n52,n49,n51);
not (n53,n54);
nor (n54,n55,n60);
nor (n55,n56,n59);
and (n56,n49,n57);
not (n57,n58);
nor (n59,n49,n57);
nand (n60,n61,n64);
or (n61,n62,n58);
not (n62,n63);
nand (n64,n62,n58);
nand (n65,n66,n60);
nor (n66,n67,n70);
and (n67,n48,n68);
not (n68,n69);
and (n70,n49,n69);
nand (n71,n72,n92);
or (n72,n73,n81);
not (n73,n74);
nor (n74,n75,n78);
and (n75,n76,n77);
and (n78,n79,n80);
not (n79,n76);
not (n80,n77);
nand (n81,n82,n89);
nor (n82,n83,n87);
and (n83,n84,n86);
not (n84,n85);
and (n87,n85,n88);
not (n88,n86);
nand (n89,n90,n91);
or (n90,n86,n79);
nand (n91,n79,n86);
nand (n92,n93,n98);
nand (n93,n94,n97);
or (n94,n95,n76);
not (n95,n96);
or (n97,n79,n96);
not (n98,n82);
xor (n99,n100,n154);
xor (n100,n101,n128);
nand (n101,n102,n122);
or (n102,n103,n110);
not (n103,n104);
nand (n104,n105,n109);
or (n105,n106,n107);
not (n107,n108);
nand (n109,n106,n107);
not (n110,n111);
nor (n111,n112,n117);
nor (n112,n113,n116);
and (n113,n108,n114);
not (n114,n115);
and (n116,n107,n115);
nand (n117,n118,n121);
or (n118,n119,n115);
not (n119,n120);
nand (n121,n119,n115);
nand (n122,n123,n117);
nor (n123,n124,n127);
and (n124,n125,n107);
not (n125,n126);
and (n127,n126,n108);
nand (n128,n129,n148);
or (n129,n130,n137);
nor (n130,n131,n135);
and (n131,n132,n134);
not (n132,n133);
and (n135,n133,n136);
not (n136,n134);
nand (n137,n138,n145);
not (n138,n139);
nand (n139,n140,n144);
or (n140,n141,n143);
not (n141,n142);
nand (n144,n141,n143);
nand (n145,n146,n147);
or (n146,n142,n132);
nand (n147,n132,n142);
nand (n148,n149,n139);
nor (n149,n150,n153);
and (n150,n132,n151);
not (n151,n152);
and (n153,n133,n152);
nand (n154,n155,n174);
or (n155,n156,n169);
nand (n156,n157,n164);
nor (n157,n158,n162);
and (n158,n159,n161);
not (n159,n160);
and (n162,n160,n163);
not (n163,n161);
nand (n164,n165,n168);
or (n165,n161,n166);
not (n166,n167);
nand (n168,n166,n161);
nor (n169,n170,n172);
and (n170,n166,n171);
and (n172,n167,n173);
not (n173,n171);
or (n174,n175,n157);
nor (n175,n176,n178);
and (n176,n177,n166);
and (n178,n179,n167);
not (n179,n177);
xor (n180,n181,n233);
xor (n181,n182,n208);
nand (n182,n183,n197);
or (n183,n184,n191);
not (n184,n185);
nand (n185,n186,n190);
or (n186,n187,n189);
not (n187,n188);
nand (n190,n187,n189);
not (n191,n192);
nor (n192,n193,n196);
and (n193,n119,n194);
not (n194,n195);
and (n196,n120,n195);
or (n197,n198,n202);
nand (n198,n184,n199);
nand (n199,n200,n201);
or (n200,n189,n119);
nand (n201,n119,n189);
not (n202,n203);
nand (n203,n204,n207);
or (n204,n120,n205);
not (n205,n206);
nand (n207,n120,n205);
nand (n208,n209,n226);
or (n209,n210,n216);
not (n210,n211);
nor (n211,n212,n215);
and (n212,n213,n159);
not (n213,n214);
and (n215,n214,n160);
not (n216,n217);
nor (n217,n218,n221);
xnor (n218,n159,n219);
not (n219,n220);
nor (n221,n222,n224);
and (n222,n223,n220);
and (n224,n225,n219);
not (n225,n223);
or (n226,n227,n232);
nor (n227,n228,n230);
and (n228,n159,n229);
and (n230,n231,n160);
not (n231,n229);
not (n232,n221);
nand (n233,n234,n252);
or (n234,n235,n241);
nor (n235,n236,n239);
and (n236,n237,n143);
not (n237,n238);
and (n239,n238,n240);
not (n240,n143);
nand (n241,n242,n249);
nor (n242,n243,n247);
and (n243,n244,n246);
not (n244,n245);
and (n247,n245,n248);
not (n248,n246);
nand (n249,n250,n251);
or (n250,n246,n240);
nand (n251,n240,n246);
nand (n252,n253,n143);
not (n253,n242);
and (n254,n25,n99);
xor (n255,n256,n371);
xor (n256,n257,n330);
xor (n257,n258,n305);
xor (n258,n259,n278);
nand (n259,n260,n277);
nand (n260,n261,n268,n274);
not (n261,n262);
nand (n262,n263,n267);
or (n263,n264,n266);
not (n264,n265);
nand (n267,n264,n266);
nand (n268,n269,n273);
or (n269,n270,n271);
not (n271,n272);
nand (n273,n270,n271);
nand (n274,n275,n276);
or (n275,n264,n272);
nand (n276,n264,n272);
nand (n277,n262,n272);
nand (n278,n279,n300);
or (n279,n280,n288);
not (n280,n281);
nor (n281,n282,n287);
and (n282,n283,n285);
not (n283,n284);
not (n285,n286);
and (n287,n284,n286);
not (n288,n289);
nor (n289,n290,n295);
nor (n290,n291,n293);
and (n291,n283,n292);
and (n293,n294,n284);
not (n294,n292);
nand (n295,n296,n299);
or (n296,n297,n292);
not (n297,n298);
nand (n299,n297,n292);
nand (n300,n301,n295);
nand (n301,n302,n304);
or (n302,n303,n283);
nand (n304,n303,n283);
nand (n305,n306,n326);
or (n306,n307,n321);
not (n307,n308);
nor (n308,n309,n317);
not (n309,n310);
nor (n310,n311,n314);
and (n311,n312,n313);
and (n314,n315,n316);
not (n315,n312);
not (n316,n313);
not (n317,n318);
or (n318,n319,n320);
and (n319,n312,n49);
and (n320,n315,n48);
nor (n321,n322,n324);
and (n322,n323,n316);
and (n324,n325,n313);
not (n325,n323);
or (n326,n327,n318);
nor (n327,n328,n329);
and (n328,n316,n51);
and (n329,n313,n50);
xor (n330,n331,n362);
xor (n331,n332,n355);
nand (n332,n333,n350);
or (n333,n334,n340);
not (n334,n335);
nor (n335,n336,n339);
and (n336,n337,n62);
not (n337,n338);
and (n339,n338,n63);
not (n340,n341);
and (n341,n342,n347);
nor (n342,n343,n345);
and (n343,n166,n344);
and (n345,n167,n346);
not (n346,n344);
nand (n347,n348,n349);
or (n348,n344,n62);
nand (n349,n62,n344);
nand (n350,n351,n354);
nand (n351,n352,n353);
or (n352,n171,n62);
nand (n353,n171,n62);
not (n354,n342);
nand (n355,n356,n357);
or (n356,n175,n156);
nand (n357,n358,n359);
not (n358,n157);
nor (n359,n360,n361);
and (n360,n213,n166);
and (n361,n214,n167);
nand (n362,n363,n365);
or (n363,n81,n364);
not (n364,n93);
or (n365,n366,n82);
nor (n366,n367,n369);
and (n367,n368,n79);
and (n369,n370,n76);
not (n370,n368);
xor (n371,n372,n391);
xor (n372,n373,n383);
nand (n373,n374,n376);
or (n374,n53,n375);
not (n375,n66);
or (n376,n377,n382);
nor (n377,n378,n381);
and (n378,n379,n49);
not (n379,n380);
and (n381,n48,n380);
not (n382,n60);
nand (n383,n384,n385);
or (n384,n216,n227);
or (n385,n386,n232);
nor (n386,n387,n389);
and (n387,n159,n388);
and (n389,n390,n160);
not (n390,n388);
not (n391,n392);
nand (n392,n393,n223);
or (n393,n394,n398);
nand (n394,n395,n397);
or (n395,n34,n396);
nand (n397,n34,n396);
not (n398,n399);
nand (n399,n400,n403);
nand (n400,n401,n402);
or (n401,n396,n225);
nand (n402,n225,n396);
not (n403,n394);
xor (n404,n405,n465);
xor (n405,n406,n409);
or (n406,n407,n408);
and (n407,n26,n71);
and (n408,n27,n43);
xor (n409,n410,n437);
xor (n410,n411,n435);
nand (n411,n412,n428);
or (n412,n413,n419);
not (n413,n414);
nor (n414,n415,n418);
and (n415,n187,n416);
not (n416,n417);
and (n418,n188,n417);
nand (n419,n420,n425);
nor (n420,n421,n424);
and (n421,n272,n422);
not (n422,n423);
and (n424,n271,n423);
nand (n425,n426,n427);
or (n426,n422,n188);
nand (n427,n188,n422);
nand (n428,n429,n434);
nand (n429,n430,n433);
or (n430,n188,n431);
not (n431,n432);
nand (n433,n188,n431);
not (n434,n420);
nor (n435,n436,n240);
and (n436,n241,n242);
nand (n437,n438,n458);
or (n438,n439,n452);
not (n439,n440);
nor (n440,n441,n448);
nor (n441,n442,n446);
and (n442,n443,n445);
not (n443,n444);
and (n446,n447,n444);
not (n447,n445);
nand (n448,n449,n451);
or (n449,n447,n450);
nand (n451,n447,n450);
not (n452,n453);
nor (n453,n454,n457);
and (n454,n443,n455);
not (n455,n456);
and (n457,n444,n456);
or (n458,n459,n464);
nor (n459,n460,n462);
and (n460,n461,n443);
and (n462,n444,n463);
not (n463,n461);
not (n464,n448);
xor (n465,n466,n515);
xor (n466,n467,n489);
nand (n467,n468,n484);
or (n468,n469,n475);
not (n469,n470);
nor (n470,n471,n474);
and (n471,n84,n472);
not (n472,n473);
and (n474,n85,n473);
nand (n475,n476,n481);
nor (n476,n477,n479);
and (n477,n132,n478);
and (n479,n133,n480);
not (n480,n478);
nand (n481,n482,n483);
or (n482,n480,n85);
nand (n483,n85,n480);
nand (n484,n485,n488);
nor (n485,n486,n487);
and (n486,n84,n136);
and (n487,n85,n134);
not (n488,n476);
nand (n489,n490,n509);
or (n490,n491,n498);
not (n491,n492);
nor (n492,n493,n497);
and (n493,n494,n495);
not (n494,n450);
not (n495,n496);
and (n497,n450,n496);
nand (n498,n499,n506);
or (n499,n500,n503);
not (n500,n501);
nand (n501,n494,n502);
not (n503,n504);
nand (n504,n450,n505);
not (n505,n502);
nor (n506,n507,n508);
and (n507,n107,n502);
and (n508,n108,n505);
nand (n509,n510,n511);
not (n510,n506);
nor (n511,n512,n514);
and (n512,n494,n513);
not (n513,n106);
and (n514,n450,n106);
nand (n515,n516,n518);
or (n516,n110,n517);
not (n517,n123);
or (n518,n519,n523);
not (n519,n520);
nor (n520,n521,n522);
and (n521,n107,n205);
and (n522,n108,n206);
not (n523,n117);
or (n524,n525,n984);
and (n525,n526,n833);
xor (n526,n527,n682);
xor (n527,n528,n595);
xor (n528,n529,n568);
xor (n529,n530,n546);
xor (n530,n531,n539);
nand (n531,n532,n538);
or (n532,n307,n533);
nor (n533,n534,n536);
and (n534,n316,n535);
and (n536,n313,n537);
not (n537,n535);
or (n538,n321,n318);
nand (n539,n540,n545);
or (n540,n340,n541);
not (n541,n542);
nor (n542,n543,n544);
and (n543,n380,n63);
and (n544,n379,n62);
or (n545,n342,n334);
nand (n546,n547,n562);
or (n547,n548,n558);
not (n548,n549);
and (n549,n550,n555);
not (n550,n551);
nand (n551,n552,n554);
or (n552,n79,n553);
nand (n554,n79,n553);
nand (n555,n556,n557);
or (n556,n553,n297);
nand (n557,n297,n553);
nor (n558,n559,n560);
and (n559,n297,n303);
and (n560,n298,n561);
not (n561,n303);
or (n562,n563,n550);
nor (n563,n564,n566);
and (n564,n297,n565);
and (n566,n567,n298);
not (n567,n565);
xor (n568,n569,n586);
xor (n569,n570,n577);
nand (n570,n571,n572);
or (n571,n506,n491);
or (n572,n498,n573);
not (n573,n574);
nand (n574,n575,n576);
or (n575,n450,n463);
nand (n576,n463,n450);
nand (n577,n578,n585);
or (n578,n579,n419);
not (n579,n580);
nor (n580,n581,n584);
and (n581,n582,n187);
not (n582,n583);
and (n584,n583,n188);
nand (n585,n434,n414);
nand (n586,n587,n593);
or (n587,n588,n589);
nand (n588,n261,n274);
not (n589,n590);
nand (n590,n591,n592);
or (n591,n272,n431);
or (n592,n271,n432);
or (n593,n261,n594);
not (n594,n268);
or (n595,n596,n681);
and (n596,n597,n663);
xor (n597,n598,n621);
or (n598,n599,n610);
nand (n599,n600,n605);
or (n600,n110,n601);
not (n601,n602);
nand (n602,n603,n604);
or (n603,n463,n108);
nand (n604,n463,n108);
nand (n605,n606,n117);
not (n606,n607);
nor (n607,n608,n609);
and (n608,n496,n107);
and (n609,n495,n108);
nand (n610,n611,n617);
or (n611,n612,n548);
not (n612,n613);
nand (n613,n614,n616);
or (n614,n615,n297);
nand (n616,n297,n615);
nand (n617,n618,n551);
nand (n618,n619,n620);
or (n619,n285,n298);
or (n620,n297,n286);
or (n621,n622,n662);
and (n622,n623,n648);
xor (n623,n624,n634);
nand (n624,n625,n630);
or (n625,n626,n399);
not (n626,n627);
nand (n627,n628,n629);
or (n628,n214,n225);
nand (n629,n225,n214);
nand (n630,n631,n394);
nand (n631,n632,n633);
or (n632,n229,n225);
nand (n633,n225,n229);
nand (n634,n635,n642);
or (n635,n636,n439);
not (n636,n637);
nand (n637,n638,n641);
or (n638,n444,n639);
not (n639,n640);
nand (n641,n444,n639);
nand (n642,n448,n643);
nor (n643,n644,n647);
and (n644,n645,n443);
not (n645,n646);
and (n647,n646,n444);
nand (n648,n649,n656);
or (n649,n650,n288);
not (n650,n651);
nor (n651,n652,n654);
and (n652,n284,n653);
and (n654,n283,n655);
not (n655,n653);
nand (n656,n295,n657);
nor (n657,n658,n661);
and (n658,n283,n659);
not (n659,n660);
and (n661,n284,n660);
and (n662,n624,n634);
or (n663,n664,n680);
and (n664,n665,n678);
xor (n665,n666,n668);
not (n666,n667);
nand (n668,n669,n676);
or (n669,n670,n674);
not (n670,n671);
nand (n671,n672,n673);
or (n672,n388,n34);
nand (n673,n388,n34);
not (n674,n675);
and (n675,n31,n37);
nand (n676,n677,n35);
not (n677,n37);
not (n678,n679);
and (n680,n666,n668);
and (n681,n598,n621);
or (n682,n683,n832);
and (n683,n684,n831);
xor (n684,n685,n769);
or (n685,n686,n768);
and (n686,n687,n721);
xor (n687,n688,n689);
xor (n688,n623,n648);
xor (n689,n690,n711);
xor (n690,n691,n701);
nand (n691,n692,n697);
or (n692,n693,n137);
not (n693,n694);
nor (n694,n695,n696);
and (n695,n133,n368);
and (n696,n132,n370);
nand (n697,n139,n698);
nand (n698,n699,n700);
or (n699,n473,n132);
nand (n700,n473,n132);
nand (n701,n702,n707);
or (n702,n703,n156);
not (n703,n704);
nand (n704,n705,n706);
or (n705,n380,n166);
nand (n706,n166,n380);
nand (n707,n358,n708);
nand (n708,n709,n710);
or (n709,n338,n166);
nand (n710,n166,n338);
nand (n711,n712,n717);
or (n712,n216,n713);
not (n713,n714);
nand (n714,n715,n716);
or (n715,n171,n159);
nand (n716,n159,n171);
or (n717,n718,n232);
nor (n718,n719,n720);
and (n719,n177,n159);
and (n720,n179,n160);
xor (n721,n722,n756);
xor (n722,n723,n746);
nand (n723,n724,n740);
or (n724,n725,n730);
not (n725,n726);
nand (n726,n727,n729);
or (n727,n432,n728);
not (n728,n266);
nand (n729,n728,n432);
not (n730,n731);
and (n731,n732,n737);
nand (n732,n733,n736);
or (n733,n734,n266);
not (n734,n735);
nand (n736,n266,n734);
nor (n737,n738,n739);
and (n738,n666,n735);
and (n739,n667,n734);
nand (n740,n741,n742);
not (n741,n737);
nor (n742,n743,n745);
and (n743,n744,n728);
not (n744,n270);
and (n745,n270,n266);
nand (n746,n747,n752);
or (n747,n340,n748);
not (n748,n749);
nand (n749,n750,n751);
or (n750,n51,n62);
nand (n751,n62,n51);
nand (n752,n354,n753);
nand (n753,n754,n755);
or (n754,n68,n63);
or (n755,n62,n69);
nand (n756,n757,n763);
or (n757,n498,n758);
not (n758,n759);
nand (n759,n760,n762);
or (n760,n761,n494);
nand (n762,n761,n494);
or (n763,n506,n764);
not (n764,n765);
nand (n765,n766,n767);
or (n766,n450,n455);
nand (n767,n455,n450);
and (n768,n688,n689);
xor (n769,n770,n818);
xor (n770,n771,n815);
or (n771,n772,n814);
and (n772,n773,n803);
xor (n773,n774,n784);
nand (n774,n775,n780);
or (n775,n776,n241);
not (n776,n777);
nand (n777,n778,n779);
or (n778,n134,n240);
nand (n779,n240,n134);
nand (n780,n253,n781);
nand (n781,n782,n783);
or (n782,n152,n240);
or (n783,n151,n143);
nand (n784,n785,n801);
or (n785,n786,n790);
not (n786,n787);
nand (n787,n788,n789);
or (n788,n238,n244);
nand (n789,n244,n238);
nand (n790,n791,n798);
or (n791,n792,n795);
not (n792,n793);
nand (n793,n244,n794);
not (n795,n796);
nand (n796,n245,n797);
not (n797,n794);
nor (n798,n799,n800);
and (n799,n678,n794);
and (n800,n679,n797);
nand (n801,n802,n245);
not (n802,n798);
nand (n803,n804,n809);
or (n804,n805,n261);
not (n805,n806);
nand (n806,n807,n808);
or (n807,n416,n272);
or (n808,n271,n417);
or (n809,n588,n810);
not (n810,n811);
nand (n811,n812,n813);
or (n812,n272,n582);
nand (n813,n582,n272);
and (n814,n774,n784);
or (n815,n816,n817);
and (n816,n690,n711);
and (n817,n691,n701);
xor (n818,n819,n827);
xor (n819,n820,n823);
nand (n820,n821,n822);
or (n821,n110,n607);
nand (n822,n117,n104);
nand (n823,n824,n826);
or (n824,n137,n825);
not (n825,n698);
or (n826,n130,n138);
nand (n827,n828,n830);
or (n828,n156,n829);
not (n829,n708);
or (n830,n169,n157);
xor (n831,n597,n663);
and (n832,n685,n769);
xor (n833,n834,n954);
xor (n834,n835,n904);
or (n835,n836,n903);
and (n836,n837,n900);
xor (n837,n838,n866);
or (n838,n839,n865);
and (n839,n840,n855);
xor (n840,n841,n42);
nand (n841,n842,n849);
or (n842,n843,n307);
not (n843,n844);
nor (n844,n845,n848);
and (n845,n316,n846);
not (n846,n847);
and (n848,n313,n847);
nand (n849,n850,n317);
nor (n850,n851,n854);
and (n851,n316,n852);
not (n852,n853);
and (n854,n313,n853);
nand (n855,n856,n861);
or (n856,n198,n857);
not (n857,n858);
nand (n858,n859,n860);
or (n859,n106,n119);
nand (n860,n119,n106);
or (n861,n862,n184);
nor (n862,n863,n864);
and (n863,n119,n126);
and (n864,n120,n125);
and (n865,n841,n42);
or (n866,n867,n899);
and (n867,n868,n889);
xor (n868,n869,n879);
nand (n869,n870,n875);
or (n870,n871,n475);
not (n871,n872);
nand (n872,n873,n874);
or (n873,n77,n84);
or (n874,n80,n85);
nand (n875,n876,n488);
nand (n876,n877,n878);
or (n877,n96,n84);
nand (n878,n96,n84);
nand (n879,n880,n885);
or (n880,n881,n81);
not (n881,n882);
nor (n882,n883,n884);
and (n883,n561,n79);
and (n884,n303,n76);
nand (n885,n886,n98);
nor (n886,n887,n888);
and (n887,n79,n567);
and (n888,n76,n565);
nand (n889,n890,n894);
or (n890,n53,n891);
nor (n891,n892,n893);
and (n892,n48,n535);
and (n893,n49,n537);
or (n894,n895,n382);
not (n895,n896);
nor (n896,n897,n898);
and (n897,n48,n325);
and (n898,n49,n323);
and (n899,n869,n879);
or (n900,n901,n902);
and (n901,n722,n756);
and (n902,n723,n746);
and (n903,n838,n866);
xor (n904,n905,n937);
xor (n905,n906,n923);
or (n906,n907,n922);
and (n907,n908,n919);
xor (n908,n909,n912);
nand (n909,n910,n911);
or (n910,n764,n498);
nand (n911,n574,n510);
nand (n912,n913,n918);
or (n913,n914,n419);
not (n914,n915);
nor (n915,n916,n917);
and (n916,n187,n194);
and (n917,n188,n195);
nand (n918,n580,n434);
nand (n919,n920,n921);
or (n920,n805,n588);
nand (n921,n262,n590);
and (n922,n909,n912);
or (n923,n924,n936);
and (n924,n925,n932);
xor (n925,n926,n929);
nand (n926,n927,n928);
or (n927,n862,n198);
nand (n928,n203,n185);
nand (n929,n930,n931);
or (n930,n718,n216);
nand (n931,n211,n221);
nand (n932,n933,n935);
or (n933,n241,n934);
not (n934,n781);
or (n935,n235,n242);
and (n936,n926,n929);
or (n937,n938,n953);
and (n938,n939,n949);
xor (n939,n940,n945);
nand (n940,n941,n943);
or (n941,n942,n307);
not (n942,n850);
nand (n943,n944,n317);
not (n944,n533);
nand (n945,n946,n948);
or (n946,n947,n340);
not (n947,n753);
nand (n948,n354,n542);
nand (n949,n950,n952);
or (n950,n548,n951);
not (n951,n618);
or (n952,n558,n550);
and (n953,n940,n945);
or (n954,n955,n983);
and (n955,n956,n982);
xor (n956,n957,n981);
xor (n957,n958,n974);
xor (n958,n959,n967);
nand (n959,n960,n962);
or (n960,n961,n439);
not (n961,n643);
nand (n962,n448,n963);
nor (n963,n964,n966);
and (n964,n443,n965);
not (n965,n761);
and (n966,n444,n761);
nand (n967,n968,n970);
or (n968,n969,n475);
not (n969,n876);
nand (n970,n971,n488);
nor (n971,n972,n973);
and (n972,n84,n370);
and (n973,n85,n368);
nand (n974,n975,n977);
or (n975,n399,n976);
not (n976,n631);
or (n977,n978,n403);
nor (n978,n979,n980);
and (n979,n225,n388);
and (n980,n223,n390);
xor (n981,n925,n932);
xor (n982,n939,n949);
and (n983,n957,n981);
and (n984,n527,n682);
xor (n985,n986,n993);
xor (n986,n987,n990);
or (n987,n988,n989);
and (n988,n528,n595);
and (n989,n529,n568);
or (n990,n991,n992);
and (n991,n834,n954);
and (n992,n835,n904);
xor (n993,n994,n1055);
xor (n994,n995,n1017);
xor (n995,n996,n1010);
xor (n996,n997,n1004);
nand (n997,n998,n999);
or (n998,n198,n191);
or (n999,n1000,n184);
not (n1000,n1001);
nor (n1001,n1002,n1003);
and (n1002,n119,n582);
and (n1003,n120,n583);
nand (n1004,n1005,n1006);
or (n1005,n548,n563);
or (n1006,n1007,n550);
nor (n1007,n1008,n1009);
and (n1008,n298,n80);
and (n1009,n297,n77);
nand (n1010,n1011,n1015);
or (n1011,n1012,n138);
nor (n1012,n1013,n1014);
and (n1013,n132,n238);
and (n1014,n133,n237);
or (n1015,n137,n1016);
not (n1016,n149);
or (n1017,n1018,n1054);
and (n1018,n1019,n1043);
xor (n1019,n1020,n1040);
or (n1020,n1021,n1039);
and (n1021,n1022,n1035);
xor (n1022,n1023,n1027);
nand (n1023,n1024,n1026);
or (n1024,n1025,n730);
not (n1025,n742);
nand (n1026,n741,n266);
nand (n1027,n1028,n1030);
or (n1028,n1029,n288);
not (n1029,n657);
nand (n1030,n1031,n295);
nor (n1031,n1032,n1034);
and (n1032,n283,n1033);
not (n1033,n615);
and (n1034,n284,n615);
not (n1035,n1036);
nand (n1036,n1037,n245);
or (n1037,n802,n1038);
not (n1038,n790);
and (n1039,n1023,n1027);
or (n1040,n1041,n1042);
and (n1041,n819,n827);
and (n1042,n820,n823);
or (n1043,n1044,n1053);
and (n1044,n1045,n1049);
xor (n1045,n28,n1046);
nand (n1046,n1047,n1048);
or (n1047,n895,n53);
nand (n1048,n46,n60);
nand (n1049,n1050,n1052);
or (n1050,n1051,n81);
not (n1051,n886);
nand (n1052,n74,n98);
and (n1053,n28,n1046);
and (n1054,n1020,n1040);
or (n1055,n1056,n1057);
and (n1056,n905,n937);
and (n1057,n906,n923);
and (n1058,n20,n524);
xor (n1059,n1060,n1367);
xor (n1060,n1061,n1139);
xor (n1061,n1062,n1136);
xor (n1062,n1063,n1117);
or (n1063,n1064,n1116);
and (n1064,n1065,n1107);
xor (n1065,n1066,n1084);
xor (n1066,n1067,n1081);
xor (n1067,n1068,n1078);
or (n1068,n1069,n1077);
and (n1069,n1070,n1036);
xor (n1070,n1071,n1073);
nand (n1071,n1072,n266);
or (n1072,n734,n666);
nand (n1073,n1074,n1076);
or (n1074,n1075,n288);
not (n1075,n1031);
nand (n1076,n281,n295);
and (n1077,n1071,n1073);
or (n1078,n1079,n1080);
and (n1079,n100,n154);
and (n1080,n101,n128);
or (n1081,n1082,n1083);
and (n1082,n181,n233);
and (n1083,n182,n208);
xor (n1084,n1085,n1104);
xor (n1085,n1086,n1101);
or (n1086,n1087,n1100);
and (n1087,n1088,n1097);
xor (n1088,n1089,n1093);
nand (n1089,n1090,n1092);
or (n1090,n1091,n439);
not (n1091,n963);
nand (n1092,n453,n448);
nand (n1093,n1094,n1096);
or (n1094,n1095,n475);
not (n1095,n971);
nand (n1096,n470,n488);
nand (n1097,n1098,n1099);
or (n1098,n399,n978);
or (n1099,n403,n225);
and (n1100,n1089,n1093);
or (n1101,n1102,n1103);
and (n1102,n569,n586);
and (n1103,n570,n577);
or (n1104,n1105,n1106);
and (n1105,n530,n546);
and (n1106,n531,n539);
or (n1107,n1108,n1115);
and (n1108,n1109,n1114);
xor (n1109,n1110,n1113);
or (n1110,n1111,n1112);
and (n1111,n958,n974);
and (n1112,n959,n967);
xor (n1113,n1070,n1036);
xor (n1114,n1088,n1097);
and (n1115,n1110,n1113);
and (n1116,n1066,n1084);
xor (n1117,n1118,n1125);
xor (n1118,n1119,n1122);
or (n1119,n1120,n1121);
and (n1120,n1085,n1104);
and (n1121,n1086,n1101);
or (n1122,n1123,n1124);
and (n1123,n1067,n1081);
and (n1124,n1068,n1078);
xor (n1125,n1126,n1133);
xor (n1126,n1127,n1130);
or (n1127,n1128,n1129);
and (n1128,n331,n362);
and (n1129,n332,n355);
or (n1130,n1131,n1132);
and (n1131,n372,n391);
and (n1132,n373,n383);
or (n1133,n1134,n1135);
and (n1134,n996,n1010);
and (n1135,n997,n1004);
or (n1136,n1137,n1138);
and (n1137,n21,n404);
and (n1138,n22,n255);
or (n1139,n1140,n1366);
and (n1140,n1141,n1158);
xor (n1141,n1142,n1157);
or (n1142,n1143,n1156);
and (n1143,n1144,n1155);
xor (n1144,n1145,n1152);
or (n1145,n1146,n1151);
and (n1146,n1147,n1150);
xor (n1147,n1148,n1149);
xor (n1148,n1045,n1049);
xor (n1149,n908,n919);
xor (n1150,n1022,n1035);
and (n1151,n1148,n1149);
or (n1152,n1153,n1154);
and (n1153,n770,n818);
and (n1154,n771,n815);
xor (n1155,n1019,n1043);
and (n1156,n1145,n1152);
xor (n1157,n1065,n1107);
or (n1158,n1159,n1365);
and (n1159,n1160,n1163);
xor (n1160,n1161,n1162);
xor (n1161,n24,n180);
xor (n1162,n1109,n1114);
or (n1163,n1164,n1364);
and (n1164,n1165,n1299);
xor (n1165,n1166,n1245);
or (n1166,n1167,n1244);
and (n1167,n1168,n1217);
xor (n1168,n1169,n1193);
or (n1169,n1170,n1192);
and (n1170,n1171,n1185);
xor (n1171,n1172,n1178);
nand (n1172,n1173,n1177);
nand (n1173,n1174,n242,n249);
nand (n1174,n1175,n1176);
or (n1175,n143,n472);
nand (n1176,n472,n143);
nand (n1177,n777,n253);
nand (n1178,n1179,n1184);
or (n1179,n1180,n216);
not (n1180,n1181);
nand (n1181,n1182,n1183);
or (n1182,n160,n337);
nand (n1183,n337,n160);
nand (n1184,n714,n221);
nand (n1185,n1186,n1191);
or (n1186,n1187,n81);
not (n1187,n1188);
nor (n1188,n1189,n1190);
and (n1189,n285,n79);
and (n1190,n286,n76);
nand (n1191,n882,n98);
and (n1192,n1172,n1178);
or (n1193,n1194,n1216);
and (n1194,n1195,n1210);
xor (n1195,n1196,n1203);
nand (n1196,n1197,n1202);
or (n1197,n1198,n340);
not (n1198,n1199);
nand (n1199,n1200,n1201);
or (n1200,n323,n62);
nand (n1201,n62,n323);
nand (n1202,n749,n354);
nand (n1203,n1204,n1209);
or (n1204,n1205,n674);
not (n1205,n1206);
nand (n1206,n1207,n1208);
or (n1207,n35,n231);
nand (n1208,n231,n35);
nand (n1209,n671,n677);
nand (n1210,n1211,n1212);
or (n1211,n871,n476);
or (n1212,n475,n1213);
nor (n1213,n1214,n1215);
and (n1214,n565,n84);
and (n1215,n567,n85);
and (n1216,n1196,n1203);
or (n1217,n1218,n1243);
and (n1218,n1219,n1234);
xor (n1219,n1220,n1227);
nand (n1220,n1221,n1226);
or (n1221,n1222,n730);
not (n1222,n1223);
nand (n1223,n1224,n1225);
or (n1224,n266,n416);
nand (n1225,n416,n266);
nand (n1226,n726,n741);
nand (n1227,n1228,n1233);
or (n1228,n1229,n156);
not (n1229,n1230);
nor (n1230,n1231,n1232);
and (n1231,n166,n68);
and (n1232,n167,n69);
nand (n1233,n358,n704);
nand (n1234,n1235,n1236);
or (n1235,n318,n843);
or (n1236,n307,n1237);
not (n1237,n1238);
nor (n1238,n1239,n1242);
and (n1239,n316,n1240);
not (n1240,n1241);
and (n1242,n313,n1241);
and (n1243,n1220,n1227);
and (n1244,n1169,n1193);
or (n1245,n1246,n1298);
and (n1246,n1247,n1273);
xor (n1247,n1248,n1254);
nand (n1248,n1249,n1253);
or (n1249,n419,n1250);
nor (n1250,n1251,n1252);
and (n1251,n187,n206);
and (n1252,n188,n205);
or (n1253,n420,n914);
nor (n1254,n1255,n1264);
not (n1255,n1256);
nand (n1256,n1257,n1263);
or (n1257,n1258,n288);
nor (n1258,n1259,n1261);
and (n1259,n283,n1260);
and (n1261,n1262,n284);
not (n1262,n1260);
nand (n1263,n651,n295);
nor (n1264,n1265,n1267);
and (n1265,n667,n1266);
and (n1267,n1268,n1271);
nor (n1268,n1269,n1270);
and (n1269,n666,n744);
and (n1270,n667,n270);
and (n1271,n667,n1272);
not (n1272,n1266);
or (n1273,n1274,n1297);
and (n1274,n1275,n1290);
xor (n1275,n1276,n1283);
nand (n1276,n1277,n1282);
or (n1277,n1278,n548);
not (n1278,n1279);
nand (n1279,n1280,n1281);
or (n1280,n660,n297);
nand (n1281,n297,n660);
nand (n1282,n613,n551);
nand (n1283,n1284,n1289);
or (n1284,n1285,n498);
not (n1285,n1286);
nand (n1286,n1287,n1288);
or (n1287,n646,n494);
nand (n1288,n494,n646);
nand (n1289,n759,n510);
nand (n1290,n1291,n1296);
or (n1291,n137,n1292);
not (n1292,n1293);
nor (n1293,n1294,n1295);
and (n1294,n133,n96);
and (n1295,n132,n95);
or (n1296,n693,n138);
and (n1297,n1276,n1283);
and (n1298,n1248,n1254);
or (n1299,n1300,n1363);
and (n1300,n1301,n1346);
xor (n1301,n1302,n1328);
or (n1302,n1303,n1327);
and (n1303,n1304,n1320);
xor (n1304,n1305,n1312);
nand (n1305,n1306,n1311);
or (n1306,n1307,n790);
not (n1307,n1308);
nand (n1308,n1309,n1310);
or (n1309,n152,n244);
nand (n1310,n244,n152);
nand (n1311,n787,n802);
nand (n1312,n1313,n1319);
or (n1313,n1314,n439);
not (n1314,n1315);
nand (n1315,n1316,n1318);
or (n1316,n1317,n443);
nand (n1318,n443,n1317);
nand (n1319,n637,n448);
nand (n1320,n1321,n1326);
or (n1321,n1322,n588);
not (n1322,n1323);
nand (n1323,n1324,n1325);
or (n1324,n195,n271);
nand (n1325,n195,n271);
nand (n1326,n262,n811);
and (n1327,n1305,n1312);
or (n1328,n1329,n1345);
and (n1329,n1330,n1338);
xor (n1330,n39,n1331);
nand (n1331,n1332,n1337);
or (n1332,n1333,n110);
not (n1333,n1334);
nand (n1334,n1335,n1336);
or (n1335,n456,n107);
nand (n1336,n456,n107);
nand (n1337,n117,n602);
nand (n1338,n1339,n1344);
or (n1339,n399,n1340);
not (n1340,n1341);
nor (n1341,n1342,n1343);
and (n1342,n179,n225);
and (n1343,n177,n223);
or (n1344,n626,n403);
and (n1345,n39,n1331);
or (n1346,n1347,n1362);
and (n1347,n1348,n1356);
xor (n1348,n1349,n679);
nand (n1349,n1350,n1355);
or (n1350,n1351,n198);
not (n1351,n1352);
nand (n1352,n1353,n1354);
or (n1353,n119,n496);
nand (n1354,n119,n496);
nand (n1355,n185,n858);
nand (n1356,n1357,n1361);
or (n1357,n53,n1358);
nor (n1358,n1359,n1360);
and (n1359,n48,n853);
and (n1360,n49,n852);
or (n1361,n382,n891);
and (n1362,n1349,n679);
and (n1363,n1302,n1328);
and (n1364,n1166,n1245);
and (n1365,n1161,n1162);
and (n1366,n1142,n1157);
xor (n1367,n1368,n1506);
xor (n1368,n1369,n1388);
xor (n1369,n1370,n1385);
xor (n1370,n1371,n1382);
xor (n1371,n1372,n1379);
xor (n1372,n1373,n1376);
or (n1373,n1374,n1375);
and (n1374,n258,n305);
and (n1375,n259,n278);
or (n1376,n1377,n1378);
and (n1377,n410,n437);
and (n1378,n411,n435);
or (n1379,n1380,n1381);
and (n1380,n466,n515);
and (n1381,n467,n489);
or (n1382,n1383,n1384);
and (n1383,n405,n465);
and (n1384,n406,n409);
or (n1385,n1386,n1387);
and (n1386,n256,n371);
and (n1387,n257,n330);
xor (n1388,n1389,n1503);
xor (n1389,n1390,n1448);
xor (n1390,n1391,n1432);
xor (n1391,n1392,n1414);
xor (n1392,n1393,n1408);
xor (n1393,n1394,n1401);
nand (n1394,n1395,n1397);
or (n1395,n1396,n475);
not (n1396,n485);
nand (n1397,n1398,n488);
nor (n1398,n1399,n1400);
and (n1399,n84,n151);
and (n1400,n85,n152);
nand (n1401,n1402,n1404);
or (n1402,n1403,n498);
not (n1403,n511);
nand (n1404,n1405,n510);
nor (n1405,n1406,n1407);
and (n1406,n494,n125);
and (n1407,n450,n126);
nand (n1408,n1409,n1410);
or (n1409,n519,n110);
nand (n1410,n117,n1411);
nor (n1411,n1412,n1413);
and (n1412,n194,n107);
and (n1413,n195,n108);
xor (n1414,n1415,n1426);
xor (n1415,n1416,n1419);
nand (n1416,n1417,n272);
or (n1417,n262,n1418);
not (n1418,n588);
nand (n1419,n1420,n1422);
or (n1420,n1421,n288);
not (n1421,n301);
nand (n1422,n1423,n295);
nor (n1423,n1424,n1425);
and (n1424,n283,n567);
and (n1425,n284,n565);
nand (n1426,n1427,n1428);
or (n1427,n307,n327);
or (n1428,n1429,n318);
nor (n1429,n1430,n1431);
and (n1430,n69,n316);
and (n1431,n68,n313);
xor (n1432,n1433,n1442);
xor (n1433,n1434,n1441);
nand (n1434,n1435,n1437);
or (n1435,n419,n1436);
not (n1436,n429);
nand (n1437,n434,n1438);
nand (n1438,n1439,n1440);
or (n1439,n744,n188);
or (n1440,n187,n270);
not (n1441,n435);
nand (n1442,n1443,n1444);
or (n1443,n439,n459);
or (n1444,n1445,n464);
nor (n1445,n1446,n1447);
and (n1446,n444,n495);
and (n1447,n443,n496);
xor (n1448,n1449,n1484);
xor (n1449,n1450,n1473);
xor (n1450,n1451,n1467);
xor (n1451,n1452,n1459);
nand (n1452,n1453,n1455);
or (n1453,n1454,n340);
not (n1454,n351);
nand (n1455,n354,n1456);
nor (n1456,n1457,n1458);
and (n1457,n179,n62);
and (n1458,n177,n63);
nand (n1459,n1460,n1465);
or (n1460,n157,n1461);
not (n1461,n1462);
nor (n1462,n1463,n1464);
and (n1463,n231,n166);
and (n1464,n229,n167);
nand (n1465,n1466,n359);
not (n1466,n156);
nand (n1467,n1468,n1469);
or (n1468,n81,n366);
or (n1469,n1470,n82);
nor (n1470,n1471,n1472);
and (n1471,n473,n79);
and (n1472,n472,n76);
xor (n1473,n1474,n392);
xor (n1474,n1475,n1481);
nand (n1475,n1476,n1477);
or (n1476,n377,n53);
nand (n1477,n1478,n60);
nor (n1478,n1479,n1480);
and (n1479,n48,n337);
and (n1480,n49,n338);
nand (n1481,n1482,n1483);
or (n1482,n386,n216);
nand (n1483,n221,n160);
xor (n1484,n1485,n1500);
xor (n1485,n1486,n1492);
nand (n1486,n1487,n1488);
or (n1487,n1000,n198);
nand (n1488,n1489,n185);
nor (n1489,n1490,n1491);
and (n1490,n119,n416);
and (n1491,n120,n417);
nand (n1492,n1493,n1498);
or (n1493,n550,n1494);
not (n1494,n1495);
nand (n1495,n1496,n1497);
or (n1496,n95,n298);
or (n1497,n297,n96);
nand (n1498,n1499,n549);
not (n1499,n1007);
nand (n1500,n1501,n1502);
or (n1501,n137,n1012);
or (n1502,n138,n132);
or (n1503,n1504,n1505);
and (n1504,n994,n1055);
and (n1505,n995,n1017);
or (n1506,n1507,n1508);
and (n1507,n986,n993);
and (n1508,n987,n990);
or (n1509,n1510,n1846);
and (n1510,n1511,n1569);
xor (n1511,n1512,n1513);
xor (n1512,n1141,n1158);
or (n1513,n1514,n1568);
and (n1514,n1515,n1567);
xor (n1515,n1516,n1566);
or (n1516,n1517,n1565);
and (n1517,n1518,n1528);
xor (n1518,n1519,n1527);
or (n1519,n1520,n1526);
and (n1520,n1521,n1525);
xor (n1521,n1522,n1524);
nand (n1522,n598,n1523);
nand (n1523,n599,n610);
xor (n1524,n773,n803);
xor (n1525,n840,n855);
and (n1526,n1522,n1524);
xor (n1527,n837,n900);
or (n1528,n1529,n1564);
and (n1529,n1530,n1533);
xor (n1530,n1531,n1532);
xor (n1531,n868,n889);
xor (n1532,n665,n678);
or (n1533,n1534,n1563);
and (n1534,n1535,n1543);
xor (n1535,n1536,n1542);
nand (n1536,n1537,n1541);
or (n1537,n419,n1538);
nor (n1538,n1539,n1540);
and (n1539,n187,n126);
and (n1540,n188,n125);
or (n1541,n420,n1250);
xor (n1542,n1264,n1255);
and (n1543,n1544,n1553);
nand (n1544,n1545,n1547);
or (n1545,n1272,n1546);
not (n1546,n1268);
or (n1547,n1548,n1552);
not (n1548,n1549);
nor (n1549,n1550,n1551);
and (n1550,n666,n431);
and (n1551,n432,n667);
not (n1552,n1271);
nand (n1553,n1554,n1561);
or (n1554,n288,n1555);
not (n1555,n1556);
nor (n1556,n1557,n1560);
and (n1557,n283,n1558);
not (n1558,n1559);
and (n1560,n1559,n284);
or (n1561,n1258,n1562);
not (n1562,n295);
and (n1563,n1536,n1542);
and (n1564,n1531,n1532);
and (n1565,n1519,n1527);
xor (n1566,n1144,n1155);
xor (n1567,n1160,n1163);
and (n1568,n1516,n1566);
or (n1569,n1570,n1845);
and (n1570,n1571,n1844);
xor (n1571,n1572,n1747);
or (n1572,n1573,n1746);
and (n1573,n1574,n1577);
xor (n1574,n1575,n1576);
xor (n1575,n1147,n1150);
xor (n1576,n956,n982);
or (n1577,n1578,n1745);
and (n1578,n1579,n1664);
xor (n1579,n1580,n1663);
or (n1580,n1581,n1662);
and (n1581,n1582,n1637);
xor (n1582,n1583,n1611);
or (n1583,n1584,n1610);
and (n1584,n1585,n1603);
xor (n1585,n1586,n1596);
nand (n1586,n1587,n1595);
or (n1587,n1588,n1591);
not (n1588,n1589);
nor (n1589,n42,n1590);
not (n1591,n1592);
nor (n1592,n1593,n1594);
and (n1593,n42,n390);
and (n1594,n388,n39);
nand (n1595,n39,n1590);
nand (n1596,n1597,n1602);
or (n1597,n1598,n110);
not (n1598,n1599);
nand (n1599,n1600,n1601);
or (n1600,n761,n107);
nand (n1601,n107,n761);
nand (n1602,n1334,n117);
nand (n1603,n1604,n1609);
or (n1604,n1605,n399);
not (n1605,n1606);
nor (n1606,n1607,n1608);
and (n1607,n225,n173);
and (n1608,n171,n223);
nand (n1609,n1341,n394);
and (n1610,n1586,n1596);
or (n1611,n1612,n1636);
and (n1612,n1613,n1628);
xor (n1613,n1614,n1621);
nand (n1614,n1615,n1620);
or (n1615,n1616,n730);
not (n1616,n1617);
nand (n1617,n1618,n1619);
or (n1618,n583,n728);
nand (n1619,n583,n728);
nand (n1620,n1223,n741);
nand (n1621,n1622,n1627);
or (n1622,n1623,n156);
not (n1623,n1624);
nand (n1624,n1625,n1626);
or (n1625,n167,n50);
nand (n1626,n50,n167);
nand (n1627,n1230,n358);
nand (n1628,n1629,n1635);
or (n1629,n1630,n307);
not (n1630,n1631);
nand (n1631,n1632,n1634);
or (n1632,n316,n1633);
nand (n1634,n1633,n316);
nand (n1635,n1238,n317);
and (n1636,n1614,n1621);
or (n1637,n1638,n1661);
and (n1638,n1639,n1654);
xor (n1639,n1640,n1647);
nand (n1640,n1641,n1646);
or (n1641,n1642,n241);
not (n1642,n1643);
nand (n1643,n1644,n1645);
or (n1644,n143,n370);
nand (n1645,n143,n370);
nand (n1646,n253,n1174);
nand (n1647,n1648,n1653);
or (n1648,n216,n1649);
not (n1649,n1650);
nand (n1650,n1651,n1652);
or (n1651,n160,n379);
nand (n1652,n160,n379);
nand (n1653,n1181,n221);
nand (n1654,n1655,n1660);
or (n1655,n81,n1656);
not (n1656,n1657);
nor (n1657,n1658,n1659);
and (n1658,n79,n1033);
and (n1659,n615,n76);
or (n1660,n82,n1187);
and (n1661,n1640,n1647);
and (n1662,n1583,n1611);
xor (n1663,n1247,n1273);
or (n1664,n1665,n1744);
and (n1665,n1666,n1715);
xor (n1666,n1667,n1691);
or (n1667,n1668,n1690);
and (n1668,n1669,n1683);
xor (n1669,n1670,n1677);
nand (n1670,n1671,n1676);
or (n1671,n1672,n548);
not (n1672,n1673);
nand (n1673,n1674,n1675);
or (n1674,n653,n297);
nand (n1675,n653,n297);
nand (n1676,n1279,n551);
nand (n1677,n1678,n1682);
or (n1678,n1679,n498);
nor (n1679,n1680,n1681);
and (n1680,n494,n640);
and (n1681,n450,n639);
nand (n1682,n1286,n510);
nand (n1683,n1684,n1689);
or (n1684,n1685,n137);
not (n1685,n1686);
nor (n1686,n1687,n1688);
and (n1687,n132,n80);
and (n1688,n77,n133);
nand (n1689,n1293,n139);
and (n1690,n1670,n1677);
or (n1691,n1692,n1714);
and (n1692,n1693,n1708);
xor (n1693,n1694,n1701);
nand (n1694,n1695,n1700);
or (n1695,n1696,n340);
not (n1696,n1697);
nand (n1697,n1698,n1699);
or (n1698,n535,n62);
nand (n1699,n535,n62);
nand (n1700,n354,n1199);
nand (n1701,n1702,n1707);
or (n1702,n1703,n674);
not (n1703,n1704);
nand (n1704,n1705,n1706);
or (n1705,n35,n213);
or (n1706,n214,n34);
nand (n1707,n1206,n677);
nand (n1708,n1709,n1713);
or (n1709,n475,n1710);
nor (n1710,n1711,n1712);
and (n1711,n561,n85);
and (n1712,n303,n84);
or (n1713,n476,n1213);
and (n1714,n1694,n1701);
or (n1715,n1716,n1743);
and (n1716,n1717,n1736);
xor (n1717,n1718,n1725);
nand (n1718,n1719,n1720);
or (n1719,n184,n1351);
or (n1720,n198,n1721);
not (n1721,n1722);
nor (n1722,n1723,n1724);
and (n1723,n119,n463);
and (n1724,n461,n120);
nand (n1725,n1726,n1735);
or (n1726,n1727,n1731);
not (n1727,n1728);
nor (n1728,n1729,n1730);
and (n1729,n678,n237);
and (n1730,n238,n679);
not (n1731,n1732);
and (n1732,n679,n1733);
not (n1733,n1734);
or (n1735,n678,n1733);
nand (n1736,n1737,n1742);
or (n1737,n53,n1738);
not (n1738,n1739);
nor (n1739,n1740,n1741);
and (n1740,n847,n49);
and (n1741,n48,n846);
or (n1742,n1358,n382);
and (n1743,n1718,n1725);
and (n1744,n1667,n1691);
and (n1745,n1580,n1663);
and (n1746,n1575,n1576);
or (n1747,n1748,n1843);
and (n1748,n1749,n1796);
xor (n1749,n1750,n1795);
or (n1750,n1751,n1794);
and (n1751,n1752,n1761);
xor (n1752,n1753,n1754);
xor (n1753,n1168,n1217);
or (n1754,n1755,n1760);
and (n1755,n1756,n1759);
xor (n1756,n1757,n1758);
xor (n1757,n1304,n1320);
xor (n1758,n1171,n1185);
xor (n1759,n1219,n1234);
and (n1760,n1757,n1758);
or (n1761,n1762,n1793);
and (n1762,n1763,n1792);
xor (n1763,n1764,n1791);
or (n1764,n1765,n1790);
and (n1765,n1766,n1783);
xor (n1766,n1767,n1774);
nand (n1767,n1768,n1773);
or (n1768,n1769,n790);
not (n1769,n1770);
nand (n1770,n1771,n1772);
or (n1771,n134,n244);
nand (n1772,n244,n134);
nand (n1773,n1308,n802);
nand (n1774,n1775,n1782);
or (n1775,n1776,n439);
not (n1776,n1777);
nand (n1777,n1778,n1781);
or (n1778,n444,n1779);
not (n1779,n1780);
nand (n1781,n1779,n444);
nand (n1782,n448,n1315);
nand (n1783,n1784,n1789);
or (n1784,n588,n1785);
not (n1785,n1786);
nand (n1786,n1787,n1788);
or (n1787,n271,n206);
nand (n1788,n206,n271);
or (n1789,n1322,n261);
and (n1790,n1767,n1774);
xor (n1791,n1330,n1338);
xor (n1792,n1348,n1356);
and (n1793,n1764,n1791);
and (n1794,n1753,n1754);
xor (n1795,n1165,n1299);
or (n1796,n1797,n1842);
and (n1797,n1798,n1801);
xor (n1798,n1799,n1800);
xor (n1799,n1301,n1346);
xor (n1800,n1521,n1525);
or (n1801,n1802,n1841);
and (n1802,n1803,n1806);
xor (n1803,n1804,n1805);
xor (n1804,n1275,n1290);
xor (n1805,n1195,n1210);
or (n1806,n1807,n1840);
and (n1807,n1808,n1839);
xor (n1808,n1809,n1815);
nand (n1809,n1810,n1814);
or (n1810,n419,n1811);
nor (n1811,n1812,n1813);
and (n1812,n187,n106);
and (n1813,n513,n188);
or (n1814,n420,n1538);
or (n1815,n1816,n1838);
and (n1816,n1817,n1831);
xor (n1817,n1818,n1825);
nor (n1818,n1819,n443);
nor (n1819,n1820,n1823);
and (n1820,n1821,n447);
not (n1821,n1822);
nor (n1823,n1824,n450);
and (n1824,n1822,n445);
and (n1825,n1826,n313);
nand (n1826,n1827,n1830);
or (n1827,n1828,n49);
and (n1828,n1829,n312);
or (n1830,n1829,n312);
nor (n1831,n1832,n283);
nor (n1832,n1833,n1836);
and (n1833,n1834,n297);
nand (n1834,n1835,n292);
and (n1836,n1837,n294);
not (n1837,n1835);
and (n1838,n1818,n1825);
xor (n1839,n1544,n1553);
and (n1840,n1809,n1815);
and (n1841,n1804,n1805);
and (n1842,n1799,n1800);
and (n1843,n1750,n1795);
xor (n1844,n526,n833);
and (n1845,n1572,n1747);
and (n1846,n1512,n1513);
and (n1847,n17,n1059);
xor (n1848,n1849,n2010);
xor (n1849,n1850,n1853);
or (n1850,n1851,n1852);
and (n1851,n1368,n1506);
and (n1852,n1369,n1388);
xor (n1853,n1854,n1909);
xor (n1854,n1855,n1906);
xor (n1855,n1856,n1903);
xor (n1856,n1857,n1900);
xor (n1857,n1858,n1897);
xor (n1858,n1859,n1875);
xor (n1859,n1860,n1869);
xor (n1860,n1861,n1863);
nor (n1861,n1862,n132);
and (n1862,n137,n138);
nand (n1863,n1864,n1865);
or (n1864,n439,n1445);
or (n1865,n1866,n464);
nor (n1866,n1867,n1868);
and (n1867,n444,n513);
and (n1868,n443,n106);
nand (n1869,n1870,n1871);
or (n1870,n81,n1470);
or (n1871,n1872,n82);
nor (n1872,n1873,n1874);
and (n1873,n79,n134);
and (n1874,n76,n136);
xor (n1875,n1876,n1891);
xor (n1876,n1877,n1884);
nand (n1877,n1878,n1880);
or (n1878,n1879,n475);
not (n1879,n1398);
nand (n1880,n1881,n488);
nor (n1881,n1882,n1883);
and (n1882,n237,n84);
and (n1883,n238,n85);
nand (n1884,n1885,n1887);
or (n1885,n1886,n498);
not (n1886,n1405);
nand (n1887,n1888,n510);
nor (n1888,n1889,n1890);
and (n1889,n494,n205);
and (n1890,n450,n206);
nand (n1891,n1892,n1893);
or (n1892,n307,n1429);
or (n1893,n1894,n318);
nor (n1894,n1895,n1896);
and (n1895,n380,n316);
and (n1896,n379,n313);
or (n1897,n1898,n1899);
and (n1898,n1372,n1379);
and (n1899,n1373,n1376);
or (n1900,n1901,n1902);
and (n1901,n1370,n1385);
and (n1902,n1371,n1382);
or (n1903,n1904,n1905);
and (n1904,n1118,n1125);
and (n1905,n1119,n1122);
or (n1906,n1907,n1908);
and (n1907,n1062,n1136);
and (n1908,n1063,n1117);
xor (n1909,n1910,n2007);
xor (n1910,n1911,n1980);
xor (n1911,n1912,n1919);
xor (n1912,n1913,n1916);
or (n1913,n1914,n1915);
and (n1914,n1391,n1432);
and (n1915,n1392,n1414);
or (n1916,n1917,n1918);
and (n1917,n1449,n1484);
and (n1918,n1450,n1473);
xor (n1919,n1920,n1958);
xor (n1920,n1921,n1938);
xor (n1921,n1922,n1931);
xor (n1922,n1923,n1925);
nor (n1923,n1924,n159);
and (n1924,n216,n232);
nand (n1925,n1926,n1927);
or (n1926,n1494,n548);
nand (n1927,n1928,n551);
nor (n1928,n1929,n1930);
and (n1929,n297,n370);
and (n1930,n298,n368);
nand (n1931,n1932,n1934);
or (n1932,n340,n1933);
not (n1933,n1456);
or (n1934,n342,n1935);
nor (n1935,n1936,n1937);
and (n1936,n62,n214);
and (n1937,n63,n213);
xor (n1938,n1939,n1951);
xor (n1939,n1940,n1944);
nand (n1940,n1941,n1943);
or (n1941,n1942,n419);
not (n1942,n1438);
nand (n1943,n434,n188);
nand (n1944,n1945,n1947);
or (n1945,n1946,n288);
not (n1946,n1423);
nand (n1947,n1948,n295);
nor (n1948,n1949,n1950);
and (n1949,n283,n80);
and (n1950,n284,n77);
nand (n1951,n1952,n1954);
or (n1952,n53,n1953);
not (n1953,n1478);
or (n1954,n1955,n382);
nor (n1955,n1956,n1957);
and (n1956,n171,n48);
and (n1957,n173,n49);
xor (n1958,n1959,n1973);
xor (n1959,n1960,n1966);
nand (n1960,n1961,n1962);
or (n1961,n1461,n156);
nand (n1962,n1963,n358);
nor (n1963,n1964,n1965);
and (n1964,n390,n166);
and (n1965,n388,n167);
nand (n1966,n1967,n1969);
or (n1967,n1968,n110);
not (n1968,n1411);
nand (n1969,n117,n1970);
nand (n1970,n1971,n1972);
or (n1971,n108,n582);
or (n1972,n107,n583);
nand (n1973,n1974,n1976);
or (n1974,n198,n1975);
not (n1975,n1489);
or (n1976,n1977,n184);
nor (n1977,n1978,n1979);
and (n1978,n119,n432);
and (n1979,n120,n431);
xor (n1980,n1981,n1996);
xor (n1981,n1982,n1985);
or (n1982,n1983,n1984);
and (n1983,n1126,n1133);
and (n1984,n1127,n1130);
xor (n1985,n1986,n1993);
xor (n1986,n1987,n1990);
or (n1987,n1988,n1989);
and (n1988,n1485,n1500);
and (n1989,n1486,n1492);
or (n1990,n1991,n1992);
and (n1991,n1474,n392);
and (n1992,n1475,n1481);
or (n1993,n1994,n1995);
and (n1994,n1451,n1467);
and (n1995,n1452,n1459);
xor (n1996,n1997,n2004);
xor (n1997,n1998,n2001);
or (n1998,n1999,n2000);
and (n1999,n1415,n1426);
and (n2000,n1416,n1419);
or (n2001,n2002,n2003);
and (n2002,n1433,n1442);
and (n2003,n1434,n1441);
or (n2004,n2005,n2006);
and (n2005,n1393,n1408);
and (n2006,n1394,n1401);
or (n2007,n2008,n2009);
and (n2008,n1389,n1503);
and (n2009,n1390,n1448);
or (n2010,n2011,n2012);
and (n2011,n1060,n1367);
and (n2012,n1061,n1139);
nand (n2013,n14,n1848);
not (n2014,n2015);
nor (n2015,n2016,n4668);
and (n2016,n2017,n4662);
nand (n2017,n2018,n4655);
or (n2018,n2019,n4623);
nor (n2019,n2020,n4608);
and (n2020,n2021,n3182,n4591);
nor (n2021,n2022,n3151);
nor (n2022,n2023,n2998);
xor (n2023,n2024,n2782);
xor (n2024,n2025,n2709);
or (n2025,n2026,n2708);
and (n2026,n2027,n2542);
xor (n2027,n2028,n2134);
or (n2028,n2029,n2133);
and (n2029,n2030,n2041);
xor (n2030,n2031,n2036);
xor (n2031,n2032,n2035);
xor (n2032,n2033,n2034);
xor (n2033,n1585,n1603);
xor (n2034,n1766,n1783);
xor (n2035,n1639,n1654);
xor (n2036,n2037,n2040);
xor (n2037,n2038,n2039);
xor (n2038,n1613,n1628);
xor (n2039,n1669,n1683);
xor (n2040,n1693,n1708);
or (n2041,n2042,n2132);
and (n2042,n2043,n2090);
xor (n2043,n2044,n2068);
xor (n2044,n2045,n2060);
xor (n2045,n2046,n2053);
nand (n2046,n2047,n2048);
or (n2047,n318,n1630);
or (n2048,n307,n2049);
nor (n2049,n2050,n2052);
and (n2050,n313,n2051);
not (n2051,n1829);
and (n2052,n1829,n316);
nand (n2053,n2054,n2059);
or (n2054,n2055,n241);
not (n2055,n2056);
nand (n2056,n2057,n2058);
or (n2057,n96,n240);
nand (n2058,n240,n96);
nand (n2059,n1643,n253);
nand (n2060,n2061,n2066);
or (n2061,n2062,n1588);
not (n2062,n2063);
nor (n2063,n2064,n2065);
and (n2064,n42,n231);
and (n2065,n229,n39);
or (n2066,n1591,n2067);
not (n2067,n1590);
xor (n2068,n2069,n2084);
xor (n2069,n2070,n2077);
nand (n2070,n2071,n2076);
or (n2071,n1731,n2072);
not (n2072,n2073);
nor (n2073,n2074,n2075);
and (n2074,n678,n151);
and (n2075,n152,n679);
nand (n2076,n1728,n1734);
nand (n2077,n2078,n2083);
or (n2078,n2079,n216);
not (n2079,n2080);
nand (n2080,n2081,n2082);
or (n2081,n69,n159);
nand (n2082,n69,n159);
nand (n2083,n1650,n221);
nand (n2084,n2085,n2086);
or (n2085,n138,n1685);
or (n2086,n137,n2087);
nor (n2087,n2088,n2089);
and (n2088,n565,n132);
and (n2089,n567,n133);
xor (n2090,n2091,n2100);
xor (n2091,n2092,n2099);
or (n2092,n2093,n2098);
and (n2093,n2094,n2097);
xor (n2094,n2095,n2096);
and (n2095,n448,n1822);
and (n2096,n317,n1829);
nor (n2097,n1562,n1837);
and (n2098,n2095,n2096);
xor (n2099,n1817,n1831);
or (n2100,n2101,n2131);
and (n2101,n2102,n2119);
xor (n2102,n2103,n2109);
nand (n2103,n2104,n2105);
or (n2104,n2067,n2062);
nand (n2105,n2106,n1589);
nor (n2106,n2107,n2108);
and (n2107,n42,n213);
and (n2108,n214,n39);
nand (n2109,n2110,n2115);
or (n2110,n2111,n198);
not (n2111,n2112);
nor (n2112,n2113,n2114);
and (n2113,n119,n965);
and (n2114,n761,n120);
nand (n2115,n185,n2116);
nand (n2116,n2117,n2118);
or (n2117,n120,n455);
nand (n2118,n120,n455);
nand (n2119,n2120,n2125);
or (n2120,n2121,n382);
not (n2121,n2122);
nand (n2122,n2123,n2124);
or (n2123,n49,n1240);
nand (n2124,n1240,n49);
nand (n2125,n2126,n54);
not (n2126,n2127);
nor (n2127,n2128,n2129);
and (n2128,n1633,n48);
and (n2129,n2130,n49);
not (n2130,n1633);
and (n2131,n2103,n2109);
and (n2132,n2044,n2068);
and (n2133,n2031,n2036);
or (n2134,n2135,n2541);
and (n2135,n2136,n2532);
xor (n2136,n2137,n2405);
or (n2137,n2138,n2404);
and (n2138,n2139,n2343);
xor (n2139,n2140,n2246);
or (n2140,n2141,n2245);
and (n2141,n2142,n2211);
xor (n2142,n2143,n2176);
or (n2143,n2144,n2175);
and (n2144,n2145,n2166);
xor (n2145,n2146,n2156);
nand (n2146,n2147,n2152);
or (n2147,n2148,n548);
not (n2148,n2149);
nor (n2149,n2150,n2151);
and (n2150,n1837,n297);
and (n2151,n1835,n298);
nand (n2152,n2153,n551);
nor (n2153,n2154,n2155);
and (n2154,n1558,n297);
and (n2155,n1559,n298);
nand (n2156,n2157,n2162);
or (n2157,n2158,n730);
not (n2158,n2159);
nor (n2159,n2160,n2161);
and (n2160,n125,n728);
and (n2161,n126,n266);
nand (n2162,n2163,n741);
nor (n2163,n2164,n2165);
and (n2164,n205,n728);
and (n2165,n206,n266);
nand (n2166,n2167,n2171);
or (n2167,n137,n2168);
nor (n2168,n2169,n2170);
and (n2169,n132,n286);
and (n2170,n133,n285);
nand (n2171,n2172,n139);
or (n2172,n2173,n2174);
and (n2173,n303,n132);
and (n2174,n561,n133);
and (n2175,n2146,n2156);
or (n2176,n2177,n2210);
and (n2177,n2178,n2200);
xor (n2178,n2179,n2189);
nand (n2179,n2180,n2185);
or (n2180,n2181,n241);
not (n2181,n2182);
nand (n2182,n2183,n2184);
or (n2183,n565,n240);
or (n2184,n143,n567);
nand (n2185,n253,n2186);
nand (n2186,n2187,n2188);
or (n2187,n80,n143);
nand (n2188,n143,n80);
nand (n2189,n2190,n2196);
or (n2190,n110,n2191);
not (n2191,n2192);
nor (n2192,n2193,n2195);
and (n2193,n2194,n107);
not (n2194,n1317);
and (n2195,n1317,n108);
nand (n2196,n117,n2197);
nor (n2197,n2198,n2199);
and (n2198,n639,n107);
and (n2199,n640,n108);
nand (n2200,n2201,n2206);
or (n2201,n674,n2202);
not (n2202,n2203);
nor (n2203,n2204,n2205);
and (n2204,n34,n337);
and (n2205,n338,n35);
or (n2206,n2207,n37);
nor (n2207,n2208,n2209);
and (n2208,n34,n171);
and (n2209,n35,n173);
and (n2210,n2179,n2189);
or (n2211,n2212,n2244);
and (n2212,n2213,n2234);
xor (n2213,n2214,n2224);
nand (n2214,n2215,n2220);
or (n2215,n2216,n81);
not (n2216,n2217);
nand (n2217,n2218,n2219);
or (n2218,n76,n1262);
or (n2219,n1260,n79);
nand (n2220,n2221,n98);
nor (n2221,n2222,n2223);
and (n2222,n79,n655);
and (n2223,n653,n76);
nand (n2224,n2225,n2230);
or (n2225,n1733,n2226);
not (n2226,n2227);
nor (n2227,n2228,n2229);
and (n2228,n678,n136);
and (n2229,n134,n679);
nand (n2230,n2231,n1732);
nor (n2231,n2232,n2233);
and (n2232,n678,n472);
and (n2233,n473,n679);
nand (n2234,n2235,n2240);
or (n2235,n1552,n2236);
not (n2236,n2237);
nor (n2237,n2238,n2239);
and (n2238,n194,n666);
and (n2239,n195,n667);
or (n2240,n2241,n1272);
nor (n2241,n2242,n2243);
and (n2242,n583,n666);
and (n2243,n667,n582);
and (n2244,n2214,n2224);
and (n2245,n2143,n2176);
or (n2246,n2247,n2342);
and (n2247,n2248,n2317);
xor (n2248,n2249,n2283);
or (n2249,n2250,n2282);
and (n2250,n2251,n2272);
xor (n2251,n2252,n2262);
nand (n2252,n2253,n2258);
or (n2253,n2254,n419);
not (n2254,n2255);
nor (n2255,n2256,n2257);
and (n2256,n187,n455);
and (n2257,n456,n188);
nand (n2258,n2259,n434);
nor (n2259,n2260,n2261);
and (n2260,n187,n463);
and (n2261,n461,n188);
nand (n2262,n2263,n2268);
or (n2263,n2264,n399);
not (n2264,n2265);
nor (n2265,n2266,n2267);
and (n2266,n69,n223);
and (n2267,n68,n225);
nand (n2268,n2269,n394);
nor (n2269,n2270,n2271);
and (n2270,n379,n225);
and (n2271,n380,n223);
nand (n2272,n2273,n2278);
or (n2273,n588,n2274);
not (n2274,n2275);
nor (n2275,n2276,n2277);
and (n2276,n496,n272);
and (n2277,n495,n271);
or (n2278,n2279,n261);
nor (n2279,n2280,n2281);
and (n2280,n272,n513);
and (n2281,n271,n106);
and (n2282,n2252,n2262);
or (n2283,n2284,n2316);
and (n2284,n2285,n2306);
xor (n2285,n2286,n2296);
nand (n2286,n2287,n2292);
or (n2287,n2288,n216);
not (n2288,n2289);
nand (n2289,n2290,n2291);
or (n2290,n323,n159);
nand (n2291,n323,n159);
nand (n2292,n2293,n221);
nand (n2293,n2294,n2295);
or (n2294,n51,n159);
nand (n2295,n159,n51);
nand (n2296,n2297,n2302);
or (n2297,n2298,n156);
not (n2298,n2299);
nor (n2299,n2300,n2301);
and (n2300,n166,n852);
and (n2301,n853,n167);
nand (n2302,n2303,n358);
nand (n2303,n2304,n2305);
or (n2304,n535,n166);
nand (n2305,n535,n166);
nand (n2306,n2307,n2312);
or (n2307,n2308,n475);
not (n2308,n2309);
nor (n2309,n2310,n2311);
and (n2310,n84,n659);
and (n2311,n660,n85);
nand (n2312,n2313,n488);
nor (n2313,n2314,n2315);
and (n2314,n1033,n84);
and (n2315,n615,n85);
and (n2316,n2286,n2296);
or (n2317,n2318,n2341);
and (n2318,n2319,n2335);
xor (n2319,n2320,n2327);
nand (n2320,n2321,n2323);
or (n2321,n2067,n2322);
not (n2322,n2106);
or (n2323,n2324,n1588);
nor (n2324,n2325,n2326);
and (n2325,n177,n42);
and (n2326,n179,n39);
nand (n2327,n2328,n2329);
or (n2328,n184,n2111);
nand (n2329,n2330,n2334);
not (n2330,n2331);
nor (n2331,n2332,n2333);
and (n2332,n119,n646);
and (n2333,n645,n120);
not (n2334,n198);
nand (n2335,n2336,n2340);
or (n2336,n53,n2337);
nor (n2337,n2338,n2339);
and (n2338,n2051,n49);
and (n2339,n1829,n48);
or (n2340,n2127,n382);
and (n2341,n2320,n2327);
and (n2342,n2249,n2283);
or (n2343,n2344,n2403);
and (n2344,n2345,n2369);
xor (n2345,n2346,n2368);
or (n2346,n2347,n2367);
and (n2347,n2348,n2361);
xor (n2348,n2349,n2355);
and (n2349,n2350,n450);
nand (n2350,n2351,n2352);
or (n2351,n502,n1822);
nand (n2352,n2353,n107);
not (n2353,n2354);
and (n2354,n1822,n502);
nor (n2355,n2356,n48);
not (n2356,n2357);
nand (n2357,n2358,n2359);
or (n2358,n1829,n58);
nand (n2359,n2360,n62);
nand (n2360,n1829,n58);
nor (n2361,n2362,n297);
nor (n2362,n2363,n2365);
and (n2363,n2364,n79);
nand (n2364,n1835,n553);
and (n2365,n1837,n2366);
not (n2366,n553);
and (n2367,n2349,n2355);
xor (n2368,n2094,n2097);
or (n2369,n2370,n2402);
and (n2370,n2371,n2392);
xor (n2371,n2372,n2382);
nand (n2372,n2373,n2378);
or (n2373,n2374,n340);
not (n2374,n2375);
nand (n2375,n2376,n2377);
or (n2376,n1241,n62);
nand (n2377,n62,n1241);
nand (n2378,n2379,n354);
nand (n2379,n2380,n2381);
or (n2380,n847,n62);
nand (n2381,n62,n847);
nand (n2382,n2383,n2388);
or (n2383,n2384,n790);
not (n2384,n2385);
nor (n2385,n2386,n2387);
and (n2386,n244,n95);
and (n2387,n96,n245);
nand (n2388,n2389,n802);
nand (n2389,n2390,n2391);
or (n2390,n368,n244);
nand (n2391,n244,n368);
nand (n2392,n2393,n2398);
or (n2393,n2394,n498);
not (n2394,n2395);
nand (n2395,n2396,n2397);
or (n2396,n1822,n494);
or (n2397,n1821,n450);
nand (n2398,n2399,n510);
nand (n2399,n2400,n2401);
or (n2400,n1780,n494);
nand (n2401,n494,n1780);
and (n2402,n2372,n2382);
and (n2403,n2346,n2368);
and (n2404,n2140,n2246);
or (n2405,n2406,n2531);
and (n2406,n2407,n2520);
xor (n2407,n2408,n2473);
or (n2408,n2409,n2472);
and (n2409,n2410,n2449);
xor (n2410,n2411,n2430);
xor (n2411,n2412,n2424);
xor (n2412,n2413,n2417);
nand (n2413,n2414,n2416);
or (n2414,n2415,n241);
not (n2415,n2186);
nand (n2416,n2056,n253);
nand (n2417,n2418,n2420);
or (n2418,n2419,n110);
not (n2419,n2197);
nand (n2420,n117,n2421);
nand (n2421,n2422,n2423);
or (n2422,n108,n645);
nand (n2423,n108,n645);
nand (n2424,n2425,n2426);
or (n2425,n2207,n674);
nand (n2426,n2427,n677);
nor (n2427,n2428,n2429);
and (n2428,n177,n35);
and (n2429,n179,n34);
xor (n2430,n2431,n2442);
xor (n2431,n2432,n2439);
nand (n2432,n2433,n2435);
or (n2433,n2434,n81);
not (n2434,n2221);
nand (n2435,n2436,n98);
nand (n2436,n2437,n2438);
or (n2437,n76,n659);
nand (n2438,n76,n659);
nand (n2439,n2440,n2441);
or (n2440,n1731,n2226);
nand (n2441,n2073,n1734);
nand (n2442,n2443,n2444);
or (n2443,n2241,n1552);
or (n2444,n2445,n1272);
not (n2445,n2446);
nor (n2446,n2447,n2448);
and (n2447,n666,n416);
and (n2448,n417,n667);
xor (n2449,n2450,n2465);
xor (n2450,n2451,n2458);
nand (n2451,n2452,n2454);
or (n2452,n2453,n340);
not (n2453,n2379);
nand (n2454,n354,n2455);
nand (n2455,n2456,n2457);
or (n2456,n853,n62);
nand (n2457,n853,n62);
nand (n2458,n2459,n2461);
or (n2459,n2460,n790);
not (n2460,n2389);
nand (n2461,n2462,n802);
nand (n2462,n2463,n2464);
or (n2463,n245,n472);
nand (n2464,n245,n472);
nand (n2465,n2466,n2468);
or (n2466,n498,n2467);
not (n2467,n2399);
or (n2468,n2469,n506);
nor (n2469,n2470,n2471);
and (n2470,n2194,n450);
and (n2471,n1317,n494);
and (n2472,n2411,n2430);
or (n2473,n2474,n2519);
and (n2474,n2475,n2498);
xor (n2475,n2476,n2497);
xor (n2476,n2477,n2490);
xor (n2477,n2478,n2485);
nand (n2478,n2479,n2481);
or (n2479,n2480,n419);
not (n2480,n2259);
nand (n2481,n2482,n434);
nand (n2482,n2483,n2484);
or (n2483,n496,n187);
nand (n2484,n496,n187);
nand (n2485,n2486,n2488);
or (n2486,n2487,n399);
not (n2487,n2269);
nand (n2488,n2489,n394);
xnor (n2489,n225,n338);
nand (n2490,n2491,n2492);
or (n2491,n588,n2279);
or (n2492,n261,n2493);
not (n2493,n2494);
nor (n2494,n2495,n2496);
and (n2495,n271,n125);
and (n2496,n126,n272);
xor (n2497,n2102,n2119);
xor (n2498,n2499,n2512);
xor (n2499,n2500,n2504);
nand (n2500,n2501,n2503);
or (n2501,n216,n2502);
not (n2502,n2293);
or (n2503,n2079,n232);
nand (n2504,n2505,n2507);
or (n2505,n156,n2506);
not (n2506,n2303);
or (n2507,n157,n2508);
not (n2508,n2509);
nor (n2509,n2510,n2511);
and (n2510,n166,n325);
and (n2511,n323,n167);
nand (n2512,n2513,n2515);
or (n2513,n475,n2514);
not (n2514,n2313);
or (n2515,n2516,n476);
nor (n2516,n2517,n2518);
and (n2517,n84,n286);
and (n2518,n85,n285);
and (n2519,n2476,n2497);
xor (n2520,n2521,n2528);
xor (n2521,n2522,n2525);
or (n2522,n2523,n2524);
and (n2523,n2477,n2490);
and (n2524,n2478,n2485);
or (n2525,n2526,n2527);
and (n2526,n2499,n2512);
and (n2527,n2500,n2504);
or (n2528,n2529,n2530);
and (n2529,n2412,n2424);
and (n2530,n2413,n2417);
and (n2531,n2408,n2473);
xor (n2532,n2533,n2538);
xor (n2533,n2534,n2535);
xor (n2534,n1808,n1839);
or (n2535,n2536,n2537);
and (n2536,n2091,n2100);
and (n2537,n2092,n2099);
or (n2538,n2539,n2540);
and (n2539,n2521,n2528);
and (n2540,n2522,n2525);
and (n2541,n2137,n2405);
or (n2542,n2543,n2707);
and (n2543,n2544,n2700);
xor (n2544,n2545,n2655);
xor (n2545,n2546,n2630);
xor (n2546,n2547,n2586);
xor (n2547,n2548,n2583);
xor (n2548,n2549,n2565);
or (n2549,n2550,n2564);
and (n2550,n2551,n2561);
xor (n2551,n2552,n2558);
nand (n2552,n2553,n2557);
nand (n2553,n2554,n737,n732);
nand (n2554,n2555,n2556);
or (n2555,n266,n194);
nand (n2556,n266,n194);
nand (n2557,n741,n1617);
nand (n2558,n2559,n2560);
nand (n2559,n2455,n342,n347);
nand (n2560,n1697,n354);
nand (n2561,n2562,n2563);
or (n2562,n2508,n156);
nand (n2563,n1624,n358);
and (n2564,n2552,n2558);
or (n2565,n2566,n2582);
and (n2566,n2567,n2578);
xor (n2567,n2568,n2571);
nand (n2568,n2569,n2570);
or (n2569,n403,n1605);
nand (n2570,n2489,n400,n403);
nand (n2571,n2572,n2577);
or (n2572,n2573,n439);
not (n2573,n2574);
nor (n2574,n2575,n2576);
and (n2575,n443,n1821);
and (n2576,n1822,n444);
nand (n2577,n1777,n448);
nand (n2578,n2579,n2581);
or (n2579,n419,n2580);
not (n2580,n2482);
or (n2581,n1811,n420);
and (n2582,n2568,n2571);
or (n2583,n2584,n2585);
and (n2584,n2069,n2084);
and (n2585,n2070,n2077);
or (n2586,n2587,n2629);
and (n2587,n2588,n2618);
xor (n2588,n2589,n2605);
xor (n2589,n2590,n2601);
xor (n2590,n2591,n2594);
nand (n2591,n2592,n2593);
or (n2592,n2121,n53);
nand (n2593,n1739,n60);
nand (n2594,n2595,n2600);
or (n2595,n2596,n288);
not (n2596,n2597);
nor (n2597,n2598,n2599);
and (n2598,n283,n1837);
and (n2599,n1835,n284);
nand (n2600,n1556,n295);
nand (n2601,n2602,n2604);
or (n2602,n2603,n110);
not (n2603,n2421);
nand (n2604,n117,n1599);
xor (n2605,n2606,n2614);
xor (n2606,n2607,n2611);
nand (n2607,n2608,n2610);
or (n2608,n2609,n198);
not (n2609,n2116);
nand (n2610,n1722,n185);
nand (n2611,n2612,n2613);
nand (n2612,n1549,n1266);
nand (n2613,n2446,n1271);
nand (n2614,n2615,n2617);
or (n2615,n2616,n81);
not (n2616,n2436);
nand (n2617,n1657,n98);
xor (n2618,n2619,n2626);
xor (n2619,n2620,n2623);
nand (n2620,n2621,n2622);
or (n2621,n2493,n588);
nand (n2622,n1786,n262);
nand (n2623,n2624,n2625);
or (n2624,n37,n1703);
nand (n2625,n675,n2427);
nand (n2626,n2627,n2628);
or (n2627,n475,n2516);
or (n2628,n476,n1710);
and (n2629,n2589,n2605);
xor (n2630,n2631,n2652);
xor (n2631,n2632,n2649);
or (n2632,n2633,n2648);
and (n2633,n2634,n2645);
xor (n2634,n2635,n2641);
nand (n2635,n2636,n2640);
or (n2636,n548,n2637);
nor (n2637,n2638,n2639);
and (n2638,n297,n1260);
and (n2639,n1262,n298);
nand (n2640,n1673,n551);
nand (n2641,n2642,n2644);
or (n2642,n2643,n790);
not (n2643,n2462);
nand (n2644,n1770,n802);
nand (n2645,n2646,n2647);
or (n2646,n498,n2469);
or (n2647,n1679,n506);
and (n2648,n2635,n2641);
or (n2649,n2650,n2651);
and (n2650,n2045,n2060);
and (n2651,n2046,n2053);
or (n2652,n2653,n2654);
and (n2653,n2619,n2626);
and (n2654,n2620,n2623);
xor (n2655,n2656,n2693);
xor (n2656,n2657,n2684);
or (n2657,n2658,n2683);
and (n2658,n2659,n2666);
xor (n2659,n2660,n2663);
or (n2660,n2661,n2662);
and (n2661,n2450,n2465);
and (n2662,n2451,n2458);
or (n2663,n2664,n2665);
and (n2664,n2431,n2442);
and (n2665,n2432,n2439);
or (n2666,n2667,n2682);
and (n2667,n2668,n2678);
xor (n2668,n2669,n2673);
nand (n2669,n2670,n2672);
or (n2670,n548,n2671);
not (n2671,n2153);
or (n2672,n550,n2637);
nand (n2673,n2674,n2676);
or (n2674,n730,n2675);
not (n2675,n2163);
or (n2676,n737,n2677);
not (n2677,n2554);
nand (n2678,n2679,n2681);
or (n2679,n137,n2680);
not (n2680,n2172);
or (n2681,n2087,n138);
and (n2682,n2669,n2673);
and (n2683,n2660,n2663);
xor (n2684,n2685,n2692);
xor (n2685,n2686,n2689);
or (n2686,n2687,n2688);
and (n2687,n2606,n2614);
and (n2688,n2607,n2611);
or (n2689,n2690,n2691);
and (n2690,n2590,n2601);
and (n2691,n2591,n2594);
xor (n2692,n1717,n1736);
or (n2693,n2694,n2699);
and (n2694,n2695,n2698);
xor (n2695,n2696,n2697);
xor (n2696,n2551,n2561);
xor (n2697,n2567,n2578);
xor (n2698,n2634,n2645);
and (n2699,n2696,n2697);
or (n2700,n2701,n2706);
and (n2701,n2702,n2705);
xor (n2702,n2703,n2704);
xor (n2703,n2659,n2666);
xor (n2704,n2695,n2698);
xor (n2705,n2588,n2618);
and (n2706,n2703,n2704);
and (n2707,n2545,n2655);
and (n2708,n2028,n2134);
xor (n2709,n2710,n2761);
xor (n2710,n2711,n2738);
or (n2711,n2712,n2737);
and (n2712,n2713,n2730);
xor (n2713,n2714,n2723);
xor (n2714,n2715,n2720);
xor (n2715,n2716,n2719);
or (n2716,n2717,n2718);
and (n2717,n2037,n2040);
and (n2718,n2038,n2039);
xor (n2719,n1582,n1637);
or (n2720,n2721,n2722);
and (n2721,n2032,n2035);
and (n2722,n2033,n2034);
xor (n2723,n2724,n2729);
xor (n2724,n2725,n2728);
or (n2725,n2726,n2727);
and (n2726,n2685,n2692);
and (n2727,n2686,n2689);
xor (n2728,n1666,n1715);
xor (n2729,n1763,n1792);
xor (n2730,n2731,n2734);
xor (n2731,n2732,n2733);
xor (n2732,n1756,n1759);
xor (n2733,n1803,n1806);
or (n2734,n2735,n2736);
and (n2735,n2533,n2538);
and (n2736,n2534,n2535);
and (n2737,n2714,n2723);
xor (n2738,n2739,n2746);
xor (n2739,n2740,n2743);
or (n2740,n2741,n2742);
and (n2741,n2724,n2729);
and (n2742,n2725,n2728);
or (n2743,n2744,n2745);
and (n2744,n2731,n2734);
and (n2745,n2732,n2733);
xor (n2746,n2747,n2750);
xor (n2747,n2748,n2749);
xor (n2748,n687,n721);
xor (n2749,n1530,n1533);
or (n2750,n2751,n2760);
and (n2751,n2752,n2759);
xor (n2752,n2753,n2756);
or (n2753,n2754,n2755);
and (n2754,n2631,n2652);
and (n2755,n2632,n2649);
or (n2756,n2757,n2758);
and (n2757,n2548,n2583);
and (n2758,n2549,n2565);
xor (n2759,n1535,n1543);
and (n2760,n2753,n2756);
xor (n2761,n2762,n2775);
xor (n2762,n2763,n2764);
xor (n2763,n1798,n1801);
or (n2764,n2765,n2774);
and (n2765,n2766,n2771);
xor (n2766,n2767,n2770);
or (n2767,n2768,n2769);
and (n2768,n2546,n2630);
and (n2769,n2547,n2586);
xor (n2770,n2752,n2759);
or (n2771,n2772,n2773);
and (n2772,n2656,n2693);
and (n2773,n2657,n2684);
and (n2774,n2767,n2770);
xor (n2775,n2776,n2781);
xor (n2776,n2777,n2778);
xor (n2777,n1579,n1664);
or (n2778,n2779,n2780);
and (n2779,n2715,n2720);
and (n2780,n2716,n2719);
xor (n2781,n1752,n1761);
or (n2782,n2783,n2997);
and (n2783,n2784,n2787);
xor (n2784,n2785,n2786);
xor (n2785,n2766,n2771);
xor (n2786,n2713,n2730);
or (n2787,n2788,n2996);
and (n2788,n2789,n2971);
xor (n2789,n2790,n2791);
xor (n2790,n2030,n2041);
or (n2791,n2792,n2970);
and (n2792,n2793,n2912);
xor (n2793,n2794,n2795);
xor (n2794,n2043,n2090);
or (n2795,n2796,n2911);
and (n2796,n2797,n2875);
xor (n2797,n2798,n2799);
xor (n2798,n2668,n2678);
or (n2799,n2800,n2874);
and (n2800,n2801,n2849);
xor (n2801,n2802,n2826);
or (n2802,n2803,n2825);
and (n2803,n2804,n2819);
xor (n2804,n2805,n2812);
nand (n2805,n2806,n2811);
or (n2806,n2807,n790);
not (n2807,n2808);
nand (n2808,n2809,n2810);
or (n2809,n77,n244);
nand (n2810,n77,n244);
nand (n2811,n2385,n802);
nand (n2812,n2813,n2815);
or (n2813,n1733,n2814);
not (n2814,n2231);
nand (n2815,n2816,n1732);
nor (n2816,n2817,n2818);
and (n2817,n678,n370);
and (n2818,n368,n679);
nand (n2819,n2820,n2821);
or (n2820,n420,n2254);
or (n2821,n419,n2822);
nor (n2822,n2823,n2824);
and (n2823,n761,n187);
and (n2824,n188,n965);
and (n2825,n2805,n2812);
or (n2826,n2827,n2848);
and (n2827,n2828,n2842);
xor (n2828,n2829,n2835);
nand (n2829,n2830,n2831);
or (n2830,n1272,n2236);
or (n2831,n2832,n1552);
nor (n2832,n2833,n2834);
and (n2833,n666,n206);
and (n2834,n667,n205);
nand (n2835,n2836,n2841);
or (n2836,n2837,n340);
not (n2837,n2838);
nand (n2838,n2839,n2840);
or (n2839,n63,n2130);
or (n2840,n62,n1633);
nand (n2841,n354,n2375);
nand (n2842,n2843,n2847);
or (n2843,n81,n2844);
nor (n2844,n2845,n2846);
and (n2845,n79,n1559);
and (n2846,n76,n1558);
or (n2847,n2216,n82);
and (n2848,n2829,n2835);
or (n2849,n2850,n2873);
and (n2850,n2851,n2866);
xor (n2851,n2852,n2859);
nand (n2852,n2853,n2858);
or (n2853,n2854,n475);
not (n2854,n2855);
nand (n2855,n2856,n2857);
or (n2856,n653,n84);
nand (n2857,n653,n84);
nand (n2858,n2309,n488);
nand (n2859,n2860,n2865);
or (n2860,n2861,n588);
not (n2861,n2862);
nor (n2862,n2863,n2864);
and (n2863,n271,n463);
and (n2864,n461,n272);
nand (n2865,n2275,n262);
nand (n2866,n2867,n2872);
or (n2867,n2868,n241);
not (n2868,n2869);
nand (n2869,n2870,n2871);
or (n2870,n143,n561);
or (n2871,n240,n303);
nand (n2872,n253,n2182);
and (n2873,n2852,n2859);
and (n2874,n2802,n2826);
or (n2875,n2876,n2910);
and (n2876,n2877,n2886);
xor (n2877,n2878,n2885);
or (n2878,n2879,n2884);
and (n2879,n2880,n2883);
xor (n2880,n2881,n2882);
and (n2881,n510,n1822);
and (n2882,n551,n1835);
nor (n2883,n382,n2051);
and (n2884,n2881,n2882);
xor (n2885,n2348,n2361);
or (n2886,n2887,n2909);
and (n2887,n2888,n2903);
xor (n2888,n2889,n2896);
nand (n2889,n2890,n2895);
or (n2890,n216,n2891);
not (n2891,n2892);
nor (n2892,n2893,n2894);
and (n2893,n159,n537);
and (n2894,n535,n160);
or (n2895,n2288,n232);
nand (n2896,n2897,n2902);
or (n2897,n2898,n730);
not (n2898,n2899);
nand (n2899,n2900,n2901);
or (n2900,n106,n728);
nand (n2901,n106,n728);
nand (n2902,n741,n2159);
nand (n2903,n2904,n2908);
or (n2904,n198,n2905);
nor (n2905,n2906,n2907);
and (n2906,n640,n119);
and (n2907,n120,n639);
or (n2908,n2331,n184);
and (n2909,n2889,n2896);
and (n2910,n2878,n2885);
and (n2911,n2798,n2799);
or (n2912,n2913,n2969);
and (n2913,n2914,n2917);
xor (n2914,n2915,n2916);
xor (n2915,n2345,n2369);
xor (n2916,n2142,n2211);
or (n2917,n2918,n2968);
and (n2918,n2919,n2967);
xor (n2919,n2920,n2944);
or (n2920,n2921,n2943);
and (n2921,n2922,n2936);
xor (n2922,n2923,n2930);
nand (n2923,n2924,n2929);
or (n2924,n2925,n110);
not (n2925,n2926);
nand (n2926,n2927,n2928);
or (n2927,n1780,n107);
nand (n2928,n1780,n107);
nand (n2929,n2192,n117);
nand (n2930,n2931,n2932);
or (n2931,n403,n2264);
nand (n2932,n398,n2933);
nand (n2933,n2934,n2935);
or (n2934,n51,n225);
nand (n2935,n51,n225);
nand (n2936,n2937,n2942);
or (n2937,n156,n2938);
not (n2938,n2939);
nand (n2939,n2940,n2941);
or (n2940,n846,n167);
or (n2941,n166,n847);
or (n2942,n2298,n157);
and (n2943,n2923,n2930);
or (n2944,n2945,n2966);
and (n2945,n2946,n2960);
xor (n2946,n2947,n2954);
nand (n2947,n2948,n2953);
or (n2948,n2949,n674);
not (n2949,n2950);
nand (n2950,n2951,n2952);
or (n2951,n34,n380);
nand (n2952,n380,n34);
nand (n2953,n2203,n677);
nand (n2954,n2955,n2959);
or (n2955,n2956,n1588);
nor (n2956,n2957,n2958);
and (n2957,n42,n171);
and (n2958,n39,n173);
or (n2959,n2324,n2067);
nand (n2960,n2961,n2965);
or (n2961,n137,n2962);
nor (n2962,n2963,n2964);
and (n2963,n615,n132);
and (n2964,n133,n1033);
or (n2965,n2168,n138);
and (n2966,n2947,n2954);
xor (n2967,n2319,n2335);
and (n2968,n2920,n2944);
and (n2969,n2915,n2916);
and (n2970,n2794,n2795);
or (n2971,n2972,n2995);
and (n2972,n2973,n2994);
xor (n2973,n2974,n2993);
or (n2974,n2975,n2992);
and (n2975,n2976,n2985);
xor (n2976,n2977,n2984);
or (n2977,n2978,n2983);
and (n2978,n2979,n2982);
xor (n2979,n2980,n2981);
xor (n2980,n2371,n2392);
xor (n2981,n2285,n2306);
xor (n2982,n2213,n2234);
and (n2983,n2980,n2981);
xor (n2984,n2248,n2317);
or (n2985,n2986,n2991);
and (n2986,n2987,n2990);
xor (n2987,n2988,n2989);
xor (n2988,n2145,n2166);
xor (n2989,n2178,n2200);
xor (n2990,n2251,n2272);
and (n2991,n2988,n2989);
and (n2992,n2977,n2984);
xor (n2993,n2139,n2343);
xor (n2994,n2407,n2520);
and (n2995,n2974,n2993);
and (n2996,n2790,n2791);
and (n2997,n2785,n2786);
or (n2998,n2999,n3150);
and (n2999,n3000,n3149);
xor (n3000,n3001,n3002);
xor (n3001,n2027,n2542);
or (n3002,n3003,n3148);
and (n3003,n3004,n3007);
xor (n3004,n3005,n3006);
xor (n3005,n2136,n2532);
xor (n3006,n2544,n2700);
or (n3007,n3008,n3147);
and (n3008,n3009,n3146);
xor (n3009,n3010,n3145);
or (n3010,n3011,n3144);
and (n3011,n3012,n3015);
xor (n3012,n3013,n3014);
xor (n3013,n2410,n2449);
xor (n3014,n2475,n2498);
or (n3015,n3016,n3143);
and (n3016,n3017,n3142);
xor (n3017,n3018,n3092);
or (n3018,n3019,n3091);
and (n3019,n3020,n3068);
xor (n3020,n3021,n3045);
or (n3021,n3022,n3044);
and (n3022,n3023,n3038);
xor (n3023,n3024,n3031);
nand (n3024,n3025,n3030);
or (n3025,n3026,n110);
not (n3026,n3027);
nand (n3027,n3028,n3029);
or (n3028,n1822,n107);
or (n3029,n108,n1821);
nand (n3030,n2926,n117);
nand (n3031,n3032,n3037);
or (n3032,n399,n3033);
not (n3033,n3034);
nor (n3034,n3035,n3036);
and (n3035,n225,n325);
and (n3036,n323,n223);
nand (n3037,n2933,n394);
nand (n3038,n3039,n3040);
or (n3039,n157,n2938);
or (n3040,n156,n3041);
nor (n3041,n3042,n3043);
and (n3042,n166,n1241);
and (n3043,n167,n1240);
and (n3044,n3024,n3031);
or (n3045,n3046,n3067);
and (n3046,n3047,n3060);
xor (n3047,n3048,n3054);
nand (n3048,n3049,n3050);
or (n3049,n37,n2949);
or (n3050,n674,n3051);
nor (n3051,n3052,n3053);
and (n3052,n34,n69);
and (n3053,n35,n68);
nand (n3054,n3055,n3059);
or (n3055,n3056,n1588);
nor (n3056,n3057,n3058);
and (n3057,n42,n338);
and (n3058,n39,n337);
or (n3059,n2956,n2067);
nand (n3060,n3061,n3066);
or (n3061,n137,n3062);
not (n3062,n3063);
nor (n3063,n3064,n3065);
and (n3064,n132,n659);
and (n3065,n660,n133);
or (n3066,n2962,n138);
and (n3067,n3048,n3054);
or (n3068,n3069,n3090);
and (n3069,n3070,n3084);
xor (n3070,n3071,n3078);
nand (n3071,n3072,n3077);
or (n3072,n3073,n1552);
not (n3073,n3074);
nand (n3074,n3075,n3076);
or (n3075,n666,n126);
nand (n3076,n126,n666);
or (n3077,n2832,n1272);
nand (n3078,n3079,n3080);
or (n3079,n342,n2837);
or (n3080,n340,n3081);
nor (n3081,n3082,n3083);
and (n3082,n63,n2051);
and (n3083,n62,n1829);
nand (n3084,n3085,n3089);
or (n3085,n81,n3086);
nor (n3086,n3087,n3088);
and (n3087,n1837,n76);
and (n3088,n1835,n79);
or (n3089,n2844,n82);
and (n3090,n3071,n3078);
and (n3091,n3021,n3045);
or (n3092,n3093,n3141);
and (n3093,n3094,n3116);
xor (n3094,n3095,n3115);
or (n3095,n3096,n3114);
and (n3096,n3097,n3109);
xor (n3097,n3098,n3103);
nor (n3098,n3099,n107);
nor (n3099,n3100,n3102);
nor (n3100,n3101,n120);
and (n3101,n1822,n115);
nor (n3102,n1822,n115);
and (n3103,n3104,n76);
nand (n3104,n3105,n3106);
or (n3105,n86,n1835);
nand (n3106,n3107,n84);
not (n3107,n3108);
and (n3108,n1835,n86);
nor (n3109,n3110,n62);
nor (n3110,n3111,n3113);
and (n3111,n3112,n166);
nand (n3112,n1829,n344);
and (n3113,n2051,n346);
and (n3114,n3098,n3103);
xor (n3115,n2880,n2883);
or (n3116,n3117,n3140);
and (n3117,n3118,n3133);
xor (n3118,n3119,n3126);
nand (n3119,n3120,n3125);
or (n3120,n3121,n790);
not (n3121,n3122);
nand (n3122,n3123,n3124);
or (n3123,n567,n245);
or (n3124,n244,n565);
nand (n3125,n802,n2808);
nand (n3126,n3127,n3131);
or (n3127,n3128,n1731);
nor (n3128,n3129,n3130);
and (n3129,n96,n678);
and (n3130,n95,n679);
or (n3131,n3132,n1733);
not (n3132,n2816);
nand (n3133,n3134,n3139);
or (n3134,n419,n3135);
not (n3135,n3136);
nand (n3136,n3137,n3138);
or (n3137,n645,n188);
or (n3138,n187,n646);
or (n3139,n2822,n420);
and (n3140,n3119,n3126);
and (n3141,n3095,n3115);
xor (n3142,n2877,n2886);
and (n3143,n3018,n3092);
and (n3144,n3013,n3014);
xor (n3145,n2702,n2705);
xor (n3146,n2793,n2912);
and (n3147,n3010,n3145);
and (n3148,n3005,n3006);
xor (n3149,n2784,n2787);
and (n3150,n3001,n3002);
nor (n3151,n3152,n3179);
xor (n3152,n3153,n3176);
xor (n3153,n3154,n3161);
xor (n3154,n3155,n3160);
xor (n3155,n3156,n3157);
xor (n3156,n1574,n1577);
or (n3157,n3158,n3159);
and (n3158,n2776,n2781);
and (n3159,n2777,n2778);
xor (n3160,n1749,n1796);
xor (n3161,n3162,n3173);
xor (n3162,n3163,n3166);
or (n3163,n3164,n3165);
and (n3164,n2739,n2746);
and (n3165,n2740,n2743);
xor (n3166,n3167,n3170);
xor (n3167,n3168,n3169);
xor (n3168,n684,n831);
xor (n3169,n1518,n1528);
or (n3170,n3171,n3172);
and (n3171,n2747,n2750);
and (n3172,n2748,n2749);
or (n3173,n3174,n3175);
and (n3174,n2762,n2775);
and (n3175,n2763,n2764);
or (n3176,n3177,n3178);
and (n3177,n2710,n2761);
and (n3178,n2711,n2738);
or (n3179,n3180,n3181);
and (n3180,n2024,n2782);
and (n3181,n2025,n2709);
nand (n3182,n3183,n4578,n4584);
nand (n3183,n3184,n3677);
nor (n3184,n3185,n3656);
nor (n3185,n3186,n3460);
xor (n3186,n3187,n3277);
xor (n3187,n3188,n3189);
xor (n3188,n3009,n3146);
xor (n3189,n3190,n3264);
xor (n3190,n3191,n3263);
or (n3191,n3192,n3262);
and (n3192,n3193,n3261);
xor (n3193,n3194,n3195);
xor (n3194,n2797,n2875);
or (n3195,n3196,n3260);
and (n3196,n3197,n3253);
xor (n3197,n3198,n3252);
or (n3198,n3199,n3251);
and (n3199,n3200,n3250);
xor (n3200,n3201,n3226);
or (n3201,n3202,n3225);
and (n3202,n3203,n3218);
xor (n3203,n3204,n3211);
nand (n3204,n3205,n3210);
or (n3205,n3206,n216);
not (n3206,n3207);
nor (n3207,n3208,n3209);
and (n3208,n159,n852);
and (n3209,n853,n160);
nand (n3210,n2892,n221);
nand (n3211,n3212,n3217);
or (n3212,n3213,n730);
not (n3213,n3214);
nor (n3214,n3215,n3216);
and (n3215,n495,n728);
and (n3216,n496,n266);
nand (n3217,n2899,n741);
nand (n3218,n3219,n3224);
or (n3219,n198,n3220);
not (n3220,n3221);
nor (n3221,n3222,n3223);
and (n3222,n119,n2194);
and (n3223,n1317,n120);
or (n3224,n2905,n184);
and (n3225,n3204,n3211);
or (n3226,n3227,n3249);
and (n3227,n3228,n3243);
xor (n3228,n3229,n3236);
nand (n3229,n3230,n3235);
or (n3230,n3231,n475);
not (n3231,n3232);
nand (n3232,n3233,n3234);
or (n3233,n85,n1262);
nand (n3234,n85,n1262);
nand (n3235,n2855,n488);
nand (n3236,n3237,n3242);
or (n3237,n3238,n588);
not (n3238,n3239);
nand (n3239,n3240,n3241);
or (n3240,n272,n455);
nand (n3241,n455,n272);
nand (n3242,n2862,n262);
not (n3243,n3244);
nor (n3244,n3245,n3246);
and (n3245,n253,n2869);
and (n3246,n3247,n3248);
not (n3247,n241);
xor (n3248,n286,n143);
and (n3249,n3229,n3236);
xor (n3250,n2851,n2866);
and (n3251,n3201,n3226);
xor (n3252,n2919,n2967);
or (n3253,n3254,n3259);
and (n3254,n3255,n3258);
xor (n3255,n3256,n3257);
xor (n3256,n2888,n2903);
xor (n3257,n2922,n2936);
xor (n3258,n2804,n2819);
and (n3259,n3256,n3257);
and (n3260,n3198,n3252);
xor (n3261,n2976,n2985);
and (n3262,n3194,n3195);
xor (n3263,n2973,n2994);
or (n3264,n3265,n3276);
and (n3265,n3266,n3275);
xor (n3266,n3267,n3274);
or (n3267,n3268,n3273);
and (n3268,n3269,n3272);
xor (n3269,n3270,n3271);
xor (n3270,n2801,n2849);
xor (n3271,n2979,n2982);
xor (n3272,n2987,n2990);
and (n3273,n3270,n3271);
xor (n3274,n2914,n2917);
xor (n3275,n3012,n3015);
and (n3276,n3267,n3274);
or (n3277,n3278,n3459);
and (n3278,n3279,n3411);
xor (n3279,n3280,n3410);
or (n3280,n3281,n3409);
and (n3281,n3282,n3327);
xor (n3282,n3283,n3326);
or (n3283,n3284,n3325);
and (n3284,n3285,n3288);
xor (n3285,n3286,n3287);
xor (n3286,n2946,n2960);
xor (n3287,n2828,n2842);
or (n3288,n3289,n3324);
and (n3289,n3290,n3299);
xor (n3290,n3291,n3298);
or (n3291,n3292,n3297);
and (n3292,n3293,n3296);
xor (n3293,n3294,n3295);
nor (n3294,n523,n1821);
and (n3295,n98,n1835);
nor (n3296,n342,n2051);
and (n3297,n3294,n3295);
xor (n3298,n3097,n3109);
or (n3299,n3300,n3323);
and (n3300,n3301,n3316);
xor (n3301,n3302,n3309);
nand (n3302,n3303,n3308);
or (n3303,n1552,n3304);
not (n3304,n3305);
nor (n3305,n3306,n3307);
and (n3306,n666,n513);
and (n3307,n106,n667);
nand (n3308,n3074,n1266);
nand (n3309,n3310,n3315);
or (n3310,n3311,n399);
not (n3311,n3312);
nor (n3312,n3313,n3314);
and (n3313,n535,n223);
and (n3314,n537,n225);
nand (n3315,n3034,n394);
nand (n3316,n3317,n3322);
or (n3317,n3318,n198);
not (n3318,n3319);
nor (n3319,n3320,n3321);
and (n3320,n1780,n120);
and (n3321,n1779,n119);
nand (n3322,n185,n3221);
and (n3323,n3302,n3309);
and (n3324,n3291,n3298);
and (n3325,n3286,n3287);
xor (n3326,n3017,n3142);
or (n3327,n3328,n3408);
and (n3328,n3329,n3407);
xor (n3329,n3330,n3331);
xor (n3330,n3094,n3116);
or (n3331,n3332,n3406);
and (n3332,n3333,n3382);
xor (n3333,n3334,n3358);
or (n3334,n3335,n3357);
and (n3335,n3336,n3351);
xor (n3336,n3337,n3344);
nand (n3337,n3338,n3343);
or (n3338,n3339,n137);
not (n3339,n3340);
nor (n3340,n3341,n3342);
and (n3341,n132,n655);
and (n3342,n653,n133);
nand (n3343,n3063,n139);
nand (n3344,n3345,n3350);
or (n3345,n3346,n156);
not (n3346,n3347);
nand (n3347,n3348,n3349);
or (n3348,n167,n2130);
nand (n3349,n167,n2130);
or (n3350,n3041,n157);
nand (n3351,n3352,n3356);
or (n3352,n3353,n1731);
nor (n3353,n3354,n3355);
and (n3354,n678,n77);
and (n3355,n679,n80);
or (n3356,n3128,n1733);
and (n3357,n3337,n3344);
or (n3358,n3359,n3381);
and (n3359,n3360,n3375);
xor (n3360,n3361,n3368);
nand (n3361,n3362,n3367);
or (n3362,n3363,n730);
not (n3363,n3364);
nand (n3364,n3365,n3366);
or (n3365,n463,n266);
or (n3366,n728,n461);
nand (n3367,n741,n3214);
nand (n3368,n3369,n3374);
or (n3369,n3370,n419);
not (n3370,n3371);
nor (n3371,n3372,n3373);
and (n3372,n187,n639);
and (n3373,n640,n188);
nand (n3374,n3136,n434);
nand (n3375,n3376,n3380);
or (n3376,n790,n3377);
nor (n3377,n3378,n3379);
and (n3378,n244,n303);
and (n3379,n245,n561);
or (n3380,n798,n3121);
and (n3381,n3361,n3368);
or (n3382,n3383,n3405);
and (n3383,n3384,n3399);
xor (n3384,n3385,n3392);
nand (n3385,n3386,n3391);
or (n3386,n3387,n588);
not (n3387,n3388);
nand (n3388,n3389,n3390);
or (n3389,n272,n965);
nand (n3390,n965,n272);
nand (n3391,n262,n3239);
nand (n3392,n3393,n3398);
or (n3393,n3394,n241);
not (n3394,n3395);
nor (n3395,n3396,n3397);
and (n3396,n615,n143);
and (n3397,n1033,n240);
nand (n3398,n3248,n253);
nand (n3399,n3400,n3404);
or (n3400,n216,n3401);
nor (n3401,n3402,n3403);
and (n3402,n159,n847);
and (n3403,n160,n846);
or (n3404,n3206,n232);
and (n3405,n3385,n3392);
and (n3406,n3334,n3358);
xor (n3407,n3200,n3250);
and (n3408,n3330,n3331);
and (n3409,n3283,n3326);
xor (n3410,n3193,n3261);
or (n3411,n3412,n3458);
and (n3412,n3413,n3457);
xor (n3413,n3414,n3456);
or (n3414,n3415,n3455);
and (n3415,n3416,n3448);
xor (n3416,n3417,n3447);
or (n3417,n3418,n3446);
and (n3418,n3419,n3445);
xor (n3419,n3420,n3444);
or (n3420,n3421,n3443);
and (n3421,n3422,n3437);
xor (n3422,n3423,n3430);
nand (n3423,n3424,n3429);
or (n3424,n3425,n475);
not (n3425,n3426);
nand (n3426,n3427,n3428);
or (n3427,n1559,n84);
nand (n3428,n1559,n84);
nand (n3429,n3232,n488);
nand (n3430,n3431,n3436);
or (n3431,n3432,n674);
not (n3432,n3433);
nor (n3433,n3434,n3435);
and (n3434,n34,n50);
and (n3435,n51,n35);
or (n3436,n3051,n37);
nand (n3437,n3438,n3442);
or (n3438,n3439,n1588);
nor (n3439,n3440,n3441);
and (n3440,n380,n42);
and (n3441,n379,n39);
or (n3442,n3056,n2067);
and (n3443,n3423,n3430);
xor (n3444,n3228,n3243);
xor (n3445,n3203,n3218);
and (n3446,n3420,n3444);
xor (n3447,n3020,n3068);
or (n3448,n3449,n3454);
and (n3449,n3450,n3453);
xor (n3450,n3451,n3452);
xor (n3451,n3023,n3038);
xor (n3452,n3118,n3133);
xor (n3453,n3070,n3084);
and (n3454,n3451,n3452);
and (n3455,n3417,n3447);
xor (n3456,n3197,n3253);
xor (n3457,n3269,n3272);
and (n3458,n3414,n3456);
and (n3459,n3280,n3410);
or (n3460,n3461,n3655);
and (n3461,n3462,n3654);
xor (n3462,n3463,n3464);
xor (n3463,n3266,n3275);
or (n3464,n3465,n3653);
and (n3465,n3466,n3604);
xor (n3466,n3467,n3603);
or (n3467,n3468,n3602);
and (n3468,n3469,n3601);
xor (n3469,n3470,n3471);
xor (n3470,n3255,n3258);
or (n3471,n3472,n3600);
and (n3472,n3473,n3548);
xor (n3473,n3474,n3475);
xor (n3474,n3047,n3060);
or (n3475,n3476,n3547);
and (n3476,n3477,n3524);
xor (n3477,n3478,n3501);
or (n3478,n3479,n3500);
and (n3479,n3480,n3494);
xor (n3480,n3481,n3488);
nand (n3481,n3482,n3487);
or (n3482,n3483,n137);
not (n3483,n3484);
nand (n3484,n3485,n3486);
or (n3485,n133,n1262);
nand (n3486,n1262,n133);
nand (n3487,n3340,n139);
nand (n3488,n3489,n3493);
or (n3489,n156,n3490);
nor (n3490,n3491,n3492);
and (n3491,n2051,n167);
and (n3492,n1829,n166);
nand (n3493,n358,n3347);
nand (n3494,n3495,n3499);
or (n3495,n3496,n1731);
nor (n3496,n3497,n3498);
and (n3497,n678,n565);
and (n3498,n679,n567);
or (n3499,n3353,n1733);
and (n3500,n3481,n3488);
or (n3501,n3502,n3523);
and (n3502,n3503,n3517);
xor (n3503,n3504,n3511);
nand (n3504,n3505,n3510);
or (n3505,n3506,n588);
not (n3506,n3507);
nand (n3507,n3508,n3509);
or (n3508,n646,n271);
nand (n3509,n646,n271);
nand (n3510,n3388,n262);
nand (n3511,n3512,n3513);
or (n3512,n242,n3394);
nand (n3513,n3247,n3514);
nand (n3514,n3515,n3516);
or (n3515,n143,n659);
nand (n3516,n143,n659);
nand (n3517,n3518,n3522);
or (n3518,n216,n3519);
nor (n3519,n3520,n3521);
and (n3520,n159,n1241);
and (n3521,n1240,n160);
or (n3522,n3401,n232);
and (n3523,n3504,n3511);
or (n3524,n3525,n3546);
and (n3525,n3526,n3540);
xor (n3526,n3527,n3533);
nand (n3527,n3528,n3532);
or (n3528,n3529,n1552);
nor (n3529,n3530,n3531);
and (n3530,n666,n496);
and (n3531,n667,n495);
or (n3532,n3304,n1272);
nand (n3533,n3534,n3535);
or (n3534,n403,n3311);
or (n3535,n399,n3536);
not (n3536,n3537);
nand (n3537,n3538,n3539);
or (n3538,n853,n225);
nand (n3539,n225,n853);
nand (n3540,n3541,n3545);
or (n3541,n198,n3542);
nor (n3542,n3543,n3544);
and (n3543,n1821,n120);
and (n3544,n1822,n119);
or (n3545,n3318,n184);
and (n3546,n3527,n3533);
and (n3547,n3478,n3501);
or (n3548,n3549,n3599);
and (n3549,n3550,n3575);
xor (n3550,n3551,n3574);
or (n3551,n3552,n3573);
and (n3552,n3553,n3566);
xor (n3553,n3554,n3561);
and (n3554,n3555,n120);
nand (n3555,n3556,n3559);
nand (n3556,n3557,n187);
not (n3557,n3558);
and (n3558,n1822,n189);
nand (n3559,n1821,n3560);
not (n3560,n189);
and (n3561,n3562,n85);
nand (n3562,n3563,n3564);
or (n3563,n1835,n478);
nand (n3564,n3565,n132);
nand (n3565,n1835,n478);
nor (n3566,n3567,n166);
and (n3567,n3568,n3571);
not (n3568,n3569);
nor (n3569,n3570,n160);
and (n3570,n1829,n161);
not (n3571,n3572);
nor (n3572,n1829,n161);
and (n3573,n3554,n3561);
xor (n3574,n3293,n3296);
or (n3575,n3576,n3598);
and (n3576,n3577,n3591);
xor (n3577,n3578,n3585);
nand (n3578,n3579,n3584);
or (n3579,n3580,n730);
not (n3580,n3581);
nand (n3581,n3582,n3583);
or (n3582,n455,n266);
or (n3583,n728,n456);
nand (n3584,n741,n3364);
nand (n3585,n3586,n3590);
or (n3586,n419,n3587);
nor (n3587,n3588,n3589);
and (n3588,n1317,n187);
and (n3589,n2194,n188);
or (n3590,n420,n3370);
nand (n3591,n3592,n3597);
or (n3592,n790,n3593);
not (n3593,n3594);
nor (n3594,n3595,n3596);
and (n3595,n286,n245);
and (n3596,n285,n244);
or (n3597,n3377,n798);
and (n3598,n3578,n3585);
and (n3599,n3551,n3574);
and (n3600,n3474,n3475);
xor (n3601,n3285,n3288);
and (n3602,n3470,n3471);
xor (n3603,n3282,n3327);
or (n3604,n3605,n3652);
and (n3605,n3606,n3651);
xor (n3606,n3607,n3650);
or (n3607,n3608,n3649);
and (n3608,n3609,n3618);
xor (n3609,n3610,n3611);
xor (n3610,n3290,n3299);
or (n3611,n3612,n3617);
and (n3612,n3613,n3616);
xor (n3613,n3614,n3615);
xor (n3614,n3301,n3316);
xor (n3615,n3384,n3399);
xor (n3616,n3360,n3375);
and (n3617,n3614,n3615);
or (n3618,n3619,n3648);
and (n3619,n3620,n3647);
xor (n3620,n3621,n3646);
or (n3621,n3622,n3645);
and (n3622,n3623,n3638);
xor (n3623,n3624,n3631);
nand (n3624,n3625,n3630);
or (n3625,n3626,n475);
not (n3626,n3627);
nand (n3627,n3628,n3629);
or (n3628,n84,n1835);
or (n3629,n1837,n85);
nand (n3630,n3426,n488);
nand (n3631,n3632,n3637);
or (n3632,n3633,n674);
not (n3633,n3634);
nand (n3634,n3635,n3636);
or (n3635,n325,n35);
or (n3636,n323,n34);
nand (n3637,n3433,n677);
nand (n3638,n3639,n3644);
or (n3639,n1588,n3640);
not (n3640,n3641);
nand (n3641,n3642,n3643);
or (n3642,n68,n39);
or (n3643,n69,n42);
or (n3644,n3439,n2067);
and (n3645,n3624,n3631);
xor (n3646,n3336,n3351);
xor (n3647,n3422,n3437);
and (n3648,n3621,n3646);
and (n3649,n3610,n3611);
xor (n3650,n3329,n3407);
xor (n3651,n3416,n3448);
and (n3652,n3607,n3650);
and (n3653,n3467,n3603);
xor (n3654,n3279,n3411);
and (n3655,n3463,n3464);
nor (n3656,n3657,n3658);
xor (n3657,n3462,n3654);
or (n3658,n3659,n3676);
and (n3659,n3660,n3675);
xor (n3660,n3661,n3662);
xor (n3661,n3413,n3457);
or (n3662,n3663,n3674);
and (n3663,n3664,n3673);
xor (n3664,n3665,n3672);
or (n3665,n3666,n3671);
and (n3666,n3667,n3670);
xor (n3667,n3668,n3669);
xor (n3668,n3333,n3382);
xor (n3669,n3450,n3453);
xor (n3670,n3419,n3445);
and (n3671,n3668,n3669);
xor (n3672,n3469,n3601);
xor (n3673,n3606,n3651);
and (n3674,n3665,n3672);
xor (n3675,n3466,n3604);
and (n3676,n3661,n3662);
nor (n3677,n3678,n4557);
and (n3678,n3679,n4325);
nor (n3679,n3680,n4321);
and (n3680,n3681,n4219);
nor (n3681,n3682,n4099);
nor (n3682,n3683,n3981);
xor (n3683,n3684,n3968);
xor (n3684,n3685,n3814);
xor (n3685,n3686,n3801);
xor (n3686,n3687,n3800);
or (n3687,n3688,n3799);
and (n3688,n3689,n3798);
xor (n3689,n3690,n3763);
or (n3690,n3691,n3762);
and (n3691,n3692,n3740);
xor (n3692,n3693,n3717);
or (n3693,n3694,n3716);
and (n3694,n3695,n3710);
xor (n3695,n3696,n3703);
nand (n3696,n3697,n3702);
or (n3697,n3698,n241);
not (n3698,n3699);
nand (n3699,n3700,n3701);
or (n3700,n143,n655);
nand (n3701,n143,n655);
nand (n3702,n3514,n253);
nand (n3703,n3704,n3709);
or (n3704,n3705,n588);
not (n3705,n3706);
nor (n3706,n3707,n3708);
and (n3707,n271,n639);
and (n3708,n640,n272);
nand (n3709,n3507,n262);
nand (n3710,n3711,n3712);
or (n3711,n2067,n3640);
or (n3712,n3713,n1588);
nor (n3713,n3714,n3715);
and (n3714,n51,n42);
and (n3715,n39,n50);
and (n3716,n3696,n3703);
or (n3717,n3718,n3739);
and (n3718,n3719,n3733);
xor (n3719,n3720,n3727);
nand (n3720,n3721,n3726);
or (n3721,n3722,n399);
not (n3722,n3723);
nor (n3723,n3724,n3725);
and (n3724,n225,n846);
and (n3725,n847,n223);
nand (n3726,n3537,n394);
nand (n3727,n3728,n3732);
or (n3728,n419,n3729);
nor (n3729,n3730,n3731);
and (n3730,n188,n1779);
and (n3731,n187,n1780);
or (n3732,n3587,n420);
nand (n3733,n3734,n3735);
or (n3734,n37,n3633);
or (n3735,n674,n3736);
nor (n3736,n3737,n3738);
and (n3737,n34,n535);
and (n3738,n35,n537);
and (n3739,n3720,n3727);
or (n3740,n3741,n3761);
and (n3741,n3742,n3755);
xor (n3742,n3743,n3749);
nand (n3743,n3744,n3748);
or (n3744,n216,n3745);
nor (n3745,n3746,n3747);
and (n3746,n1633,n159);
and (n3747,n2130,n160);
or (n3748,n3519,n232);
nand (n3749,n3750,n3754);
or (n3750,n3751,n1731);
nor (n3751,n3752,n3753);
and (n3752,n679,n561);
and (n3753,n678,n303);
or (n3754,n3496,n1733);
nand (n3755,n3756,n3760);
or (n3756,n3757,n1552);
nor (n3757,n3758,n3759);
and (n3758,n461,n666);
and (n3759,n463,n667);
or (n3760,n3529,n1272);
and (n3761,n3743,n3749);
and (n3762,n3693,n3717);
or (n3763,n3764,n3797);
and (n3764,n3765,n3774);
xor (n3765,n3766,n3773);
or (n3766,n3767,n3772);
and (n3767,n3768,n3771);
xor (n3768,n3769,n3770);
and (n3769,n185,n1822);
and (n3770,n358,n1829);
and (n3771,n488,n1835);
and (n3772,n3769,n3770);
xor (n3773,n3553,n3566);
or (n3774,n3775,n3796);
and (n3775,n3776,n3790);
xor (n3776,n3777,n3784);
nand (n3777,n3778,n3783);
or (n3778,n3779,n790);
not (n3779,n3780);
nor (n3780,n3781,n3782);
and (n3781,n615,n245);
and (n3782,n1033,n244);
nand (n3783,n3594,n802);
nand (n3784,n3785,n3786);
or (n3785,n737,n3580);
nand (n3786,n731,n3787);
nor (n3787,n3788,n3789);
and (n3788,n965,n728);
and (n3789,n761,n266);
nand (n3790,n3791,n3792);
or (n3791,n3483,n138);
or (n3792,n137,n3793);
nor (n3793,n3794,n3795);
and (n3794,n1559,n132);
and (n3795,n1558,n133);
and (n3796,n3777,n3784);
and (n3797,n3766,n3773);
xor (n3798,n3550,n3575);
and (n3799,n3690,n3763);
xor (n3800,n3473,n3548);
or (n3801,n3802,n3813);
and (n3802,n3803,n3812);
xor (n3803,n3804,n3811);
or (n3804,n3805,n3810);
and (n3805,n3806,n3809);
xor (n3806,n3807,n3808);
xor (n3807,n3623,n3638);
xor (n3808,n3480,n3494);
xor (n3809,n3503,n3517);
and (n3810,n3807,n3808);
xor (n3811,n3477,n3524);
xor (n3812,n3620,n3647);
and (n3813,n3804,n3811);
or (n3814,n3815,n3967);
and (n3815,n3816,n3874);
xor (n3816,n3817,n3873);
or (n3817,n3818,n3872);
and (n3818,n3819,n3871);
xor (n3819,n3820,n3821);
xor (n3820,n3765,n3774);
or (n3821,n3822,n3870);
and (n3822,n3823,n3847);
xor (n3823,n3824,n3846);
or (n3824,n3825,n3845);
and (n3825,n3826,n3838);
xor (n3826,n3827,n3833);
and (n3827,n3828,n188);
nand (n3828,n3829,n3832);
nand (n3829,n3830,n271);
not (n3830,n3831);
and (n3831,n1822,n423);
nand (n3832,n1821,n422);
and (n3833,n3834,n160);
nand (n3834,n3835,n3836);
or (n3835,n1829,n220);
nand (n3836,n3837,n225);
nand (n3837,n1829,n220);
nor (n3838,n3839,n132);
and (n3839,n3840,n3843);
not (n3840,n3841);
nor (n3841,n3842,n143);
and (n3842,n1835,n142);
not (n3843,n3844);
nor (n3844,n1835,n142);
and (n3845,n3827,n3833);
xor (n3846,n3768,n3771);
or (n3847,n3848,n3869);
and (n3848,n3849,n3863);
xor (n3849,n3850,n3857);
nand (n3850,n3851,n3856);
or (n3851,n3852,n399);
not (n3852,n3853);
nor (n3853,n3854,n3855);
and (n3854,n1241,n223);
and (n3855,n1240,n225);
nand (n3856,n3723,n394);
nand (n3857,n3858,n3862);
or (n3858,n137,n3859);
nor (n3859,n3860,n3861);
and (n3860,n1837,n133);
and (n3861,n132,n1835);
or (n3862,n138,n3793);
nand (n3863,n3864,n3868);
or (n3864,n3865,n1552);
nor (n3865,n3866,n3867);
and (n3866,n456,n666);
and (n3867,n455,n667);
or (n3868,n3757,n1272);
and (n3869,n3850,n3857);
and (n3870,n3824,n3846);
xor (n3871,n3692,n3740);
and (n3872,n3820,n3821);
xor (n3873,n3803,n3812);
or (n3874,n3875,n3966);
and (n3875,n3876,n3885);
xor (n3876,n3877,n3884);
or (n3877,n3878,n3883);
and (n3878,n3879,n3882);
xor (n3879,n3880,n3881);
xor (n3880,n3776,n3790);
xor (n3881,n3742,n3755);
xor (n3882,n3695,n3710);
and (n3883,n3880,n3881);
xor (n3884,n3806,n3809);
xor (n3885,n3886,n3889);
xor (n3886,n3887,n3888);
xor (n3887,n3526,n3540);
xor (n3888,n3577,n3591);
or (n3889,n3890,n3965);
and (n3890,n3891,n3943);
xor (n3891,n3892,n3917);
or (n3892,n3893,n3916);
and (n3893,n3894,n3909);
xor (n3894,n3895,n3902);
nand (n3895,n3896,n3901);
or (n3896,n3897,n241);
not (n3897,n3898);
nor (n3898,n3899,n3900);
and (n3899,n1260,n143);
and (n3900,n1262,n240);
nand (n3901,n253,n3699);
nand (n3902,n3903,n3908);
or (n3903,n588,n3904);
not (n3904,n3905);
nand (n3905,n3906,n3907);
or (n3906,n1317,n271);
nand (n3907,n1317,n271);
or (n3908,n261,n3705);
nand (n3909,n3910,n3915);
or (n3910,n3911,n1588);
not (n3911,n3912);
nor (n3912,n3913,n3914);
and (n3913,n42,n325);
and (n3914,n323,n39);
or (n3915,n3713,n2067);
and (n3916,n3895,n3902);
or (n3917,n3918,n3942);
and (n3918,n3919,n3934);
xor (n3919,n3920,n3927);
nand (n3920,n3921,n3926);
or (n3921,n3922,n790);
not (n3922,n3923);
nor (n3923,n3924,n3925);
and (n3924,n244,n659);
and (n3925,n660,n245);
nand (n3926,n3780,n802);
nand (n3927,n3928,n3933);
or (n3928,n3929,n419);
not (n3929,n3930);
nand (n3930,n3931,n3932);
or (n3931,n1822,n187);
or (n3932,n1821,n188);
or (n3933,n420,n3729);
nand (n3934,n3935,n3940);
or (n3935,n730,n3936);
not (n3936,n3937);
nor (n3937,n3938,n3939);
and (n3938,n645,n728);
and (n3939,n646,n266);
or (n3940,n3941,n737);
not (n3941,n3787);
and (n3942,n3920,n3927);
or (n3943,n3944,n3964);
and (n3944,n3945,n3958);
xor (n3945,n3946,n3952);
nand (n3946,n3947,n3951);
or (n3947,n216,n3948);
nor (n3948,n3949,n3950);
and (n3949,n2051,n160);
and (n3950,n159,n1829);
or (n3951,n3745,n232);
nand (n3952,n3953,n3957);
or (n3953,n3954,n1731);
nor (n3954,n3955,n3956);
and (n3955,n678,n286);
and (n3956,n679,n285);
or (n3957,n3751,n1733);
nand (n3958,n3959,n3963);
or (n3959,n674,n3960);
nor (n3960,n3961,n3962);
and (n3961,n34,n853);
and (n3962,n35,n852);
or (n3963,n3736,n37);
and (n3964,n3946,n3952);
and (n3965,n3892,n3917);
and (n3966,n3877,n3884);
and (n3967,n3817,n3873);
xor (n3968,n3969,n3972);
xor (n3969,n3970,n3971);
xor (n3970,n3609,n3618);
xor (n3971,n3667,n3670);
or (n3972,n3973,n3980);
and (n3973,n3974,n3979);
xor (n3974,n3975,n3976);
xor (n3975,n3613,n3616);
or (n3976,n3977,n3978);
and (n3977,n3886,n3889);
and (n3978,n3887,n3888);
xor (n3979,n3689,n3798);
and (n3980,n3975,n3976);
or (n3981,n3982,n4098);
and (n3982,n3983,n4097);
xor (n3983,n3984,n3985);
xor (n3984,n3974,n3979);
or (n3985,n3986,n4096);
and (n3986,n3987,n4095);
xor (n3987,n3988,n4030);
or (n3988,n3989,n4029);
and (n3989,n3990,n3993);
xor (n3990,n3991,n3992);
xor (n3991,n3719,n3733);
xor (n3992,n3823,n3847);
or (n3993,n3994,n4028);
and (n3994,n3995,n4004);
xor (n3995,n3996,n4003);
or (n3996,n3997,n4002);
and (n3997,n3998,n4001);
xor (n3998,n3999,n4000);
and (n3999,n434,n1822);
and (n4000,n221,n1829);
nor (n4001,n138,n1837);
and (n4002,n3999,n4000);
xor (n4003,n3826,n3838);
or (n4004,n4005,n4027);
and (n4005,n4006,n4021);
xor (n4006,n4007,n4014);
nand (n4007,n4008,n4013);
or (n4008,n1588,n4009);
not (n4009,n4010);
nand (n4010,n4011,n4012);
or (n4011,n535,n42);
nand (n4012,n535,n42);
nand (n4013,n3912,n1590);
nand (n4014,n4015,n4020);
or (n4015,n4016,n399);
not (n4016,n4017);
nor (n4017,n4018,n4019);
and (n4018,n1633,n223);
and (n4019,n2130,n225);
nand (n4020,n3853,n394);
nand (n4021,n4022,n4026);
or (n4022,n4023,n1731);
nor (n4023,n4024,n4025);
and (n4024,n678,n615);
and (n4025,n679,n1033);
or (n4026,n3954,n1733);
and (n4027,n4007,n4014);
and (n4028,n3996,n4003);
and (n4029,n3991,n3992);
or (n4030,n4031,n4094);
and (n4031,n4032,n4087);
xor (n4032,n4033,n4034);
xor (n4033,n3891,n3943);
or (n4034,n4035,n4086);
and (n4035,n4036,n4085);
xor (n4036,n4037,n4061);
or (n4037,n4038,n4060);
and (n4038,n4039,n4054);
xor (n4039,n4040,n4047);
nand (n4040,n4041,n4046);
or (n4041,n4042,n588);
not (n4042,n4043);
nand (n4043,n4044,n4045);
or (n4044,n1780,n271);
nand (n4045,n271,n1780);
nand (n4046,n262,n3905);
nand (n4047,n4048,n4053);
or (n4048,n4049,n730);
not (n4049,n4050);
nand (n4050,n4051,n4052);
or (n4051,n640,n728);
nand (n4052,n728,n640);
nand (n4053,n741,n3937);
nand (n4054,n4055,n4059);
or (n4055,n674,n4056);
nor (n4056,n4057,n4058);
and (n4057,n34,n847);
and (n4058,n846,n35);
or (n4059,n3960,n37);
and (n4060,n4040,n4047);
or (n4061,n4062,n4084);
and (n4062,n4063,n4078);
xor (n4063,n4064,n4071);
nand (n4064,n4065,n4070);
or (n4065,n4066,n790);
not (n4066,n4067);
nor (n4067,n4068,n4069);
and (n4068,n244,n655);
and (n4069,n653,n245);
nand (n4070,n802,n3923);
nand (n4071,n4072,n4077);
or (n4072,n4073,n1552);
not (n4073,n4074);
nand (n4074,n4075,n4076);
or (n4075,n666,n761);
nand (n4076,n761,n666);
or (n4077,n3865,n1272);
nand (n4078,n4079,n4083);
or (n4079,n241,n4080);
nor (n4080,n4081,n4082);
and (n4081,n240,n1559);
and (n4082,n143,n1558);
or (n4083,n242,n3897);
and (n4084,n4064,n4071);
xor (n4085,n3919,n3934);
and (n4086,n4037,n4061);
or (n4087,n4088,n4093);
and (n4088,n4089,n4092);
xor (n4089,n4090,n4091);
xor (n4090,n3894,n3909);
xor (n4091,n3945,n3958);
xor (n4092,n3849,n3863);
and (n4093,n4090,n4091);
and (n4094,n4033,n4034);
xor (n4095,n3819,n3871);
and (n4096,n3988,n4030);
xor (n4097,n3816,n3874);
and (n4098,n3984,n3985);
nor (n4099,n4100,n4101);
xor (n4100,n3983,n4097);
or (n4101,n4102,n4218);
and (n4102,n4103,n4217);
xor (n4103,n4104,n4105);
xor (n4104,n3876,n3885);
or (n4105,n4106,n4216);
and (n4106,n4107,n4215);
xor (n4107,n4108,n4109);
xor (n4108,n3879,n3882);
or (n4109,n4110,n4214);
and (n4110,n4111,n4163);
xor (n4111,n4112,n4162);
or (n4112,n4113,n4161);
and (n4113,n4114,n4137);
xor (n4114,n4115,n4136);
or (n4115,n4116,n4135);
and (n4116,n4117,n4130);
xor (n4117,n4118,n4123);
nor (n4118,n4119,n271);
nor (n4119,n4120,n4122);
and (n4120,n4121,n728);
nand (n4121,n1822,n265);
nor (n4122,n1822,n265);
nor (n4123,n4124,n225);
and (n4124,n4125,n4128);
not (n4125,n4126);
nor (n4126,n4127,n35);
and (n4127,n1829,n396);
not (n4128,n4129);
nor (n4129,n1829,n396);
nor (n4130,n4131,n240);
nor (n4131,n4132,n4134);
and (n4132,n4133,n244);
nand (n4133,n1835,n246);
and (n4134,n1837,n248);
and (n4135,n4118,n4123);
xor (n4136,n3998,n4001);
or (n4137,n4138,n4160);
and (n4138,n4139,n4154);
xor (n4139,n4140,n4147);
nand (n4140,n4141,n4146);
or (n4141,n4142,n790);
not (n4142,n4143);
nand (n4143,n4144,n4145);
or (n4144,n1260,n244);
nand (n4145,n1260,n244);
nand (n4146,n4067,n802);
nand (n4147,n4148,n4153);
or (n4148,n1552,n4149);
not (n4149,n4150);
nor (n4150,n4151,n4152);
and (n4151,n666,n645);
and (n4152,n646,n667);
nand (n4153,n4074,n1266);
nand (n4154,n4155,n4159);
or (n4155,n241,n4156);
nor (n4156,n4157,n4158);
and (n4157,n1837,n143);
and (n4158,n240,n1835);
or (n4159,n4080,n242);
and (n4160,n4140,n4147);
and (n4161,n4115,n4136);
xor (n4162,n3995,n4004);
or (n4163,n4164,n4213);
and (n4164,n4165,n4212);
xor (n4165,n4166,n4189);
or (n4166,n4167,n4188);
and (n4167,n4168,n4182);
xor (n4168,n4169,n4176);
nand (n4169,n4170,n4175);
or (n4170,n4171,n588);
not (n4171,n4172);
nand (n4172,n4173,n4174);
or (n4173,n271,n1822);
or (n4174,n1821,n272);
nand (n4175,n262,n4043);
nand (n4176,n4177,n4181);
or (n4177,n730,n4178);
nor (n4178,n4179,n4180);
and (n4179,n1317,n728);
and (n4180,n2194,n266);
nand (n4181,n741,n4050);
nand (n4182,n4183,n4187);
or (n4183,n674,n4184);
nor (n4184,n4185,n4186);
and (n4185,n34,n1241);
and (n4186,n35,n1240);
or (n4187,n4056,n37);
and (n4188,n4169,n4176);
or (n4189,n4190,n4211);
and (n4190,n4191,n4205);
xor (n4191,n4192,n4198);
nand (n4192,n4193,n4197);
or (n4193,n4194,n1588);
nor (n4194,n4195,n4196);
and (n4195,n42,n853);
and (n4196,n39,n852);
or (n4197,n4009,n2067);
nand (n4198,n4199,n4204);
or (n4199,n4200,n399);
not (n4200,n4201);
nand (n4201,n4202,n4203);
or (n4202,n225,n1829);
or (n4203,n2051,n223);
nand (n4204,n4017,n394);
nand (n4205,n4206,n4210);
or (n4206,n4207,n1731);
nor (n4207,n4208,n4209);
and (n4208,n660,n678);
and (n4209,n659,n679);
or (n4210,n4023,n1733);
and (n4211,n4192,n4198);
xor (n4212,n4063,n4078);
and (n4213,n4166,n4189);
and (n4214,n4112,n4162);
xor (n4215,n3990,n3993);
and (n4216,n4108,n4109);
xor (n4217,n3987,n4095);
and (n4218,n4104,n4105);
nand (n4219,n4220,n4320);
or (n4220,n4221,n4276);
nor (n4221,n4222,n4223);
xor (n4222,n4103,n4217);
or (n4223,n4224,n4275);
and (n4224,n4225,n4274);
xor (n4225,n4226,n4227);
xor (n4226,n4032,n4087);
or (n4227,n4228,n4273);
and (n4228,n4229,n4232);
xor (n4229,n4230,n4231);
xor (n4230,n4036,n4085);
xor (n4231,n4089,n4092);
or (n4232,n4233,n4272);
and (n4233,n4234,n4237);
xor (n4234,n4235,n4236);
xor (n4235,n4006,n4021);
xor (n4236,n4039,n4054);
or (n4237,n4238,n4271);
and (n4238,n4239,n4248);
xor (n4239,n4240,n4247);
or (n4240,n4241,n4246);
and (n4241,n4242,n4245);
xor (n4242,n4243,n4244);
and (n4243,n262,n1822);
and (n4244,n253,n1835);
nor (n4245,n403,n2051);
and (n4246,n4243,n4244);
xor (n4247,n4117,n4130);
or (n4248,n4249,n4270);
and (n4249,n4250,n4264);
xor (n4250,n4251,n4258);
nand (n4251,n4252,n4257);
or (n4252,n4253,n1731);
not (n4253,n4254);
nor (n4254,n4255,n4256);
and (n4255,n653,n679);
and (n4256,n678,n655);
or (n4257,n4207,n1733);
nand (n4258,n4259,n4263);
or (n4259,n674,n4260);
nor (n4260,n4261,n4262);
and (n4261,n34,n1633);
and (n4262,n2130,n35);
or (n4263,n4184,n37);
nand (n4264,n4265,n4269);
or (n4265,n730,n4266);
nor (n4266,n4267,n4268);
and (n4267,n728,n1780);
and (n4268,n266,n1779);
or (n4269,n737,n4178);
and (n4270,n4251,n4258);
and (n4271,n4240,n4247);
and (n4272,n4235,n4236);
and (n4273,n4230,n4231);
xor (n4274,n4107,n4215);
and (n4275,n4226,n4227);
nand (n4276,n4277,n4278);
xor (n4277,n4225,n4274);
or (n4278,n4279,n4319);
and (n4279,n4280,n4318);
xor (n4280,n4281,n4282);
xor (n4281,n4111,n4163);
or (n4282,n4283,n4317);
and (n4283,n4284,n4316);
xor (n4284,n4285,n4286);
xor (n4285,n4114,n4137);
or (n4286,n4287,n4315);
and (n4287,n4288,n4314);
xor (n4288,n4289,n4313);
or (n4289,n4290,n4312);
and (n4290,n4291,n4305);
xor (n4291,n4292,n4299);
nand (n4292,n4293,n4298);
or (n4293,n4294,n790);
not (n4294,n4295);
nor (n4295,n4296,n4297);
and (n4296,n1559,n245);
and (n4297,n1558,n244);
nand (n4298,n4143,n802);
nand (n4299,n4300,n4304);
or (n4300,n4301,n1588);
nor (n4301,n4302,n4303);
and (n4302,n42,n847);
and (n4303,n846,n39);
or (n4304,n4194,n2067);
nand (n4305,n4306,n4311);
or (n4306,n1552,n4307);
not (n4307,n4308);
nor (n4308,n4309,n4310);
and (n4309,n640,n667);
and (n4310,n639,n666);
or (n4311,n4149,n1272);
and (n4312,n4292,n4299);
xor (n4313,n4139,n4154);
xor (n4314,n4191,n4205);
and (n4315,n4289,n4313);
xor (n4316,n4165,n4212);
and (n4317,n4285,n4286);
xor (n4318,n4229,n4232);
and (n4319,n4281,n4282);
nand (n4320,n4222,n4223);
nor (n4321,n4322,n3682);
and (n4322,n4323,n4324);
nand (n4323,n3683,n3981);
nand (n4324,n4100,n4101);
nand (n4325,n3681,n4326);
nor (n4326,n4327,n4330);
nand (n4327,n4328,n4329);
or (n4328,n4278,n4277);
not (n4329,n4221);
nor (n4330,n4331,n4520,n4551);
and (n4331,n4332,n4436);
not (n4332,n4333);
nand (n4333,n4334,n4429);
or (n4334,n4335,n4422);
or (n4335,n4336,n4421);
and (n4336,n4337,n4369);
xor (n4337,n4338,n4368);
or (n4338,n4339,n4367);
and (n4339,n4340,n4366);
xor (n4340,n4341,n4365);
or (n4341,n4342,n4364);
and (n4342,n4343,n4357);
xor (n4343,n4344,n4351);
nand (n4344,n4345,n4350);
or (n4345,n1731,n4346);
not (n4346,n4347);
nor (n4347,n4348,n4349);
and (n4348,n1260,n679);
and (n4349,n1262,n678);
nand (n4350,n4254,n1734);
nand (n4351,n4352,n4353);
or (n4352,n1272,n4307);
nand (n4353,n4354,n1271);
nand (n4354,n4355,n4356);
or (n4355,n1317,n666);
nand (n4356,n666,n1317);
nand (n4357,n4358,n4363);
or (n4358,n4359,n674);
not (n4359,n4360);
nand (n4360,n4361,n4362);
or (n4361,n34,n1829);
or (n4362,n2051,n35);
or (n4363,n4260,n37);
and (n4364,n4344,n4351);
xor (n4365,n4291,n4305);
xor (n4366,n4250,n4264);
and (n4367,n4341,n4365);
xor (n4368,n4288,n4314);
xor (n4369,n4370,n4420);
xor (n4370,n4371,n4372);
xor (n4371,n4168,n4182);
or (n4372,n4373,n4419);
and (n4373,n4374,n4396);
xor (n4374,n4375,n4395);
or (n4375,n4376,n4394);
and (n4376,n4377,n4389);
xor (n4377,n4378,n4383);
nor (n4378,n4379,n728);
nor (n4379,n4380,n4381);
and (n4380,n1821,n734);
and (n4381,n4382,n666);
nand (n4382,n1822,n735);
and (n4383,n4384,n245);
nand (n4384,n4385,n4386);
or (n4385,n1835,n794);
nand (n4386,n4387,n678);
not (n4387,n4388);
and (n4388,n1835,n794);
nor (n4389,n4390,n34);
nor (n4390,n4391,n4393);
and (n4391,n4392,n42);
nand (n4392,n1829,n33);
and (n4393,n2051,n40);
and (n4394,n4378,n4383);
xor (n4395,n4242,n4245);
or (n4396,n4397,n4418);
and (n4397,n4398,n4412);
xor (n4398,n4399,n4405);
nand (n4399,n4400,n4404);
or (n4400,n790,n4401);
nor (n4401,n4402,n4403);
and (n4402,n1837,n245);
and (n4403,n1835,n244);
or (n4404,n798,n4294);
nand (n4405,n4406,n4411);
or (n4406,n1588,n4407);
not (n4407,n4408);
nor (n4408,n4409,n4410);
and (n4409,n42,n1240);
and (n4410,n1241,n39);
or (n4411,n4301,n2067);
nand (n4412,n4413,n4417);
or (n4413,n730,n4414);
nor (n4414,n4415,n4416);
and (n4415,n1821,n266);
and (n4416,n1822,n728);
or (n4417,n737,n4266);
and (n4418,n4399,n4405);
and (n4419,n4375,n4395);
xor (n4420,n4239,n4248);
and (n4421,n4338,n4368);
xor (n4422,n4423,n4428);
xor (n4423,n4424,n4427);
or (n4424,n4425,n4426);
and (n4425,n4370,n4420);
and (n4426,n4371,n4372);
xor (n4427,n4234,n4237);
xor (n4428,n4284,n4316);
nand (n4429,n4430,n4432);
not (n4430,n4431);
xor (n4431,n4280,n4318);
not (n4432,n4433);
or (n4433,n4434,n4435);
and (n4434,n4423,n4428);
and (n4435,n4424,n4427);
nand (n4436,n4437,n4517);
or (n4437,n4438,n4481);
nor (n4438,n4439,n4480);
or (n4439,n4440,n4479);
and (n4440,n4441,n4478);
xor (n4441,n4442,n4477);
or (n4442,n4443,n4476);
and (n4443,n4444,n4453);
xor (n4444,n4445,n4452);
or (n4445,n4446,n4451);
and (n4446,n4447,n4450);
xor (n4447,n4448,n4449);
and (n4448,n741,n1822);
and (n4449,n677,n1829);
nor (n4450,n798,n1837);
and (n4451,n4448,n4449);
xor (n4452,n4377,n4389);
or (n4453,n4454,n4475);
and (n4454,n4455,n4469);
xor (n4455,n4456,n4463);
nand (n4456,n4457,n4461);
or (n4457,n4458,n1552);
nor (n4458,n4459,n4460);
and (n4459,n666,n1780);
and (n4460,n667,n1779);
or (n4461,n4462,n1272);
not (n4462,n4354);
nand (n4463,n4464,n4465);
or (n4464,n1733,n4346);
or (n4465,n4466,n1731);
nor (n4466,n4467,n4468);
and (n4467,n678,n1559);
and (n4468,n1558,n679);
nand (n4469,n4470,n4471);
or (n4470,n2067,n4407);
or (n4471,n4472,n1588);
nor (n4472,n4473,n4474);
and (n4473,n39,n2130);
and (n4474,n42,n1633);
and (n4475,n4456,n4463);
and (n4476,n4445,n4452);
xor (n4477,n4374,n4396);
xor (n4478,n4340,n4366);
and (n4479,n4442,n4477);
xor (n4480,n4337,n4369);
nand (n4481,n4482,n4516);
or (n4482,n4483,n4515);
and (n4483,n4484,n4487);
xor (n4484,n4485,n4486);
xor (n4485,n4343,n4357);
xor (n4486,n4398,n4412);
or (n4487,n4488,n4514);
and (n4488,n4489,n4501);
xor (n4489,n4490,n4500);
or (n4490,n4491,n4499);
and (n4491,n4492,n4497);
xor (n4492,n4493,n4495);
and (n4493,n4494,n667);
nand (n4494,n1822,n1266);
nor (n4495,n4496,n42);
and (n4496,n1829,n1590);
nor (n4497,n4498,n678);
and (n4498,n1835,n1734);
and (n4499,n4493,n4495);
xor (n4500,n4447,n4450);
or (n4501,n4502,n4513);
and (n4502,n4503,n4510);
xor (n4503,n4504,n4507);
nand (n4504,n4505,n4506);
or (n4505,n4458,n1272);
or (n4506,n1552,n1822);
nand (n4507,n4508,n4509);
or (n4508,n4472,n2067);
or (n4509,n1588,n1829);
nand (n4510,n4511,n4512);
or (n4511,n1835,n1731);
or (n4512,n4466,n1733);
and (n4513,n4504,n4507);
and (n4514,n4490,n4500);
and (n4515,n4485,n4486);
xor (n4516,n4441,n4478);
or (n4517,n4518,n4519);
not (n4518,n4480);
not (n4519,n4439);
nor (n4520,n4333,n4521);
nand (n4521,n4522,n4523);
not (n4522,n4438);
nor (n4523,n4524,n4548);
and (n4524,n4525,n4533);
nor (n4525,n4526,n4532);
and (n4526,n4527,n4530,n4531);
or (n4527,n4528,n4529);
xor (n4528,n4484,n4487);
xor (n4529,n4444,n4453);
xor (n4530,n4489,n4501);
xor (n4531,n4455,n4469);
and (n4532,n4528,n4529);
nand (n4533,n4527,n4534);
nor (n4534,n4535,n4540,n4541);
and (n4535,n4536,n4538);
not (n4536,n4537);
xor (n4537,n4503,n4510);
not (n4538,n4539);
xor (n4539,n4492,n4497);
nor (n4540,n4530,n4531);
nor (n4541,n4542,n4543,n4544);
and (n4542,n4496,n4498);
nor (n4543,n4536,n4538);
nor (n4544,n4545,n4494);
and (n4545,n4546,n4547);
not (n4546,n4498);
not (n4547,n4496);
and (n4548,n4549,n4550);
not (n4549,n4516);
not (n4550,n4482);
nand (n4551,n4552,n4556);
or (n4552,n4553,n4554,n4555);
not (n4553,n4429);
not (n4554,n4422);
not (n4555,n4335);
nand (n4556,n4431,n4433);
nand (n4557,n4558,n4571);
or (n4558,n4559,n4562);
or (n4559,n4560,n4561);
and (n4560,n3684,n3968);
and (n4561,n3685,n3814);
xor (n4562,n4563,n4570);
xor (n4563,n4564,n4567);
or (n4564,n4565,n4566);
and (n4565,n3686,n3801);
and (n4566,n3687,n3800);
or (n4567,n4568,n4569);
and (n4568,n3969,n3972);
and (n4569,n3970,n3971);
xor (n4570,n3664,n3673);
nand (n4571,n4572,n4574);
not (n4572,n4573);
xor (n4573,n3660,n3675);
not (n4574,n4575);
or (n4575,n4576,n4577);
and (n4576,n4563,n4570);
and (n4577,n4564,n4567);
nand (n4578,n3184,n4579);
nand (n4579,n4580,n4581);
or (n4580,n4574,n4572);
or (n4581,n4582,n4583);
not (n4582,n4571);
nand (n4583,n4562,n4559);
nand (n4584,n4585,n4586);
not (n4585,n3185);
nand (n4586,n4587,n4590);
or (n4587,n4588,n4589);
not (n4588,n3460);
not (n4589,n3186);
nand (n4590,n3657,n3658);
nor (n4591,n4592,n4603);
nor (n4592,n4593,n4594);
xor (n4593,n3000,n3149);
or (n4594,n4595,n4602);
and (n4595,n4596,n4601);
xor (n4596,n4597,n4598);
xor (n4597,n2789,n2971);
or (n4598,n4599,n4600);
and (n4599,n3190,n3264);
and (n4600,n3191,n3263);
xor (n4601,n3004,n3007);
and (n4602,n4597,n4598);
nor (n4603,n4604,n4605);
xor (n4604,n4596,n4601);
or (n4605,n4606,n4607);
and (n4606,n3187,n3277);
and (n4607,n3188,n3189);
nand (n4608,n4609,n4616);
or (n4609,n4610,n4615);
not (n4610,n4611);
nand (n4611,n4612,n4614);
or (n4612,n4592,n4613);
nand (n4613,n4604,n4605);
nand (n4614,n4593,n4594);
not (n4615,n2021);
nand (n4616,n4617,n4622);
or (n4617,n4618,n4620);
not (n4618,n4619);
nand (n4619,n3152,n3179);
not (n4620,n4621);
nand (n4621,n2023,n2998);
not (n4622,n3151);
not (n4623,n4624);
nor (n4624,n4625,n4650);
nor (n4625,n4626,n4641);
xor (n4626,n4627,n4630);
xor (n4627,n4628,n4629);
xor (n4628,n19,n985);
xor (n4629,n1511,n1569);
or (n4630,n4631,n4640);
and (n4631,n4632,n4637);
xor (n4632,n4633,n4634);
xor (n4633,n1515,n1567);
or (n4634,n4635,n4636);
and (n4635,n3167,n3170);
and (n4636,n3168,n3169);
or (n4637,n4638,n4639);
and (n4638,n3155,n3160);
and (n4639,n3156,n3157);
and (n4640,n4633,n4634);
or (n4641,n4642,n4649);
and (n4642,n4643,n4646);
xor (n4643,n4644,n4645);
xor (n4644,n1571,n1844);
xor (n4645,n4632,n4637);
or (n4646,n4647,n4648);
and (n4647,n3162,n3173);
and (n4648,n3163,n3166);
and (n4649,n4644,n4645);
nor (n4650,n4651,n4652);
xor (n4651,n4643,n4646);
or (n4652,n4653,n4654);
and (n4653,n3153,n3176);
and (n4654,n3154,n3161);
nand (n4655,n4656,n4661);
or (n4656,n4657,n4659);
not (n4657,n4658);
nand (n4658,n4651,n4652);
not (n4659,n4660);
nand (n4660,n4626,n4641);
not (n4661,n4625);
not (n4662,n4663);
nor (n4663,n4664,n4667);
or (n4664,n4665,n4666);
and (n4665,n4627,n4630);
and (n4666,n4628,n4629);
xor (n4667,n16,n1509);
not (n4668,n4669);
nand (n4669,n4664,n4667);
nand (n4670,n2014,n11);
or (n4671,n4672,n1);
and (n4672,n4673,n3);
xor (n4673,n4674,n8699);
xor (n4674,n4675,n7379);
xor (n4675,n4676,n7247);
xor (n4676,n4677,n5965);
xor (n4677,n4678,n5845);
xor (n4678,n4679,n5963);
xor (n4679,n4680,n5840);
xor (n4680,n4681,n5956);
xor (n4681,n4682,n1242);
xor (n4682,n4683,n5944);
xor (n4683,n4684,n848);
xor (n4684,n4685,n5927);
xor (n4685,n4686,n854);
xor (n4686,n4687,n5905);
xor (n4687,n4688,n5819);
xor (n4688,n4689,n5878);
xor (n4689,n4690,n5813);
xor (n4690,n4691,n5846);
xor (n4691,n4692,n5807);
xor (n4692,n4693,n5804);
xor (n4693,n4694,n5803);
xor (n4694,n4695,n5753);
xor (n4695,n4696,n5752);
xor (n4696,n4697,n5699);
xor (n4697,n4698,n1480);
xor (n4698,n4699,n5636);
xor (n4699,n4700,n5635);
xor (n4700,n4701,n5568);
xor (n4701,n4702,n1458);
xor (n4702,n4703,n5493);
xor (n4703,n4704,n5492);
xor (n4704,n4705,n5415);
xor (n4705,n4706,n1464);
xor (n4706,n4707,n5329);
xor (n4707,n4708,n5328);
or (n4708,n4709,n5242);
and (n4709,n4710,n5241);
or (n4710,n4711,n5152);
and (n4711,n4712,n5151);
or (n4712,n4713,n5071);
and (n4713,n4714,n5070);
or (n4714,n4715,n4982);
and (n4715,n4716,n4981);
or (n4716,n4717,n4895);
and (n4717,n4718,n4894);
or (n4718,n4719,n4805);
and (n4719,n4720,n4804);
and (n4720,n1594,n4721);
or (n4721,n4722,n4724);
and (n4722,n4723,n2065);
and (n4723,n388,n1590);
and (n4724,n4725,n4726);
xor (n4725,n4723,n2065);
or (n4726,n4727,n4729);
and (n4727,n4728,n2108);
and (n4728,n229,n1590);
and (n4729,n4730,n4731);
xor (n4730,n4728,n2108);
or (n4731,n4732,n4735);
and (n4732,n4733,n4734);
and (n4733,n214,n1590);
and (n4734,n177,n39);
and (n4735,n4736,n4737);
xor (n4736,n4733,n4734);
or (n4737,n4738,n4741);
and (n4738,n4739,n4740);
and (n4739,n177,n1590);
and (n4740,n171,n39);
and (n4741,n4742,n4743);
xor (n4742,n4739,n4740);
or (n4743,n4744,n4747);
and (n4744,n4745,n4746);
and (n4745,n171,n1590);
and (n4746,n338,n39);
and (n4747,n4748,n4749);
xor (n4748,n4745,n4746);
or (n4749,n4750,n4753);
and (n4750,n4751,n4752);
and (n4751,n338,n1590);
and (n4752,n380,n39);
and (n4753,n4754,n4755);
xor (n4754,n4751,n4752);
or (n4755,n4756,n4759);
and (n4756,n4757,n4758);
and (n4757,n380,n1590);
and (n4758,n69,n39);
and (n4759,n4760,n4761);
xor (n4760,n4757,n4758);
or (n4761,n4762,n4765);
and (n4762,n4763,n4764);
and (n4763,n69,n1590);
and (n4764,n51,n39);
and (n4765,n4766,n4767);
xor (n4766,n4763,n4764);
or (n4767,n4768,n4770);
and (n4768,n4769,n3914);
and (n4769,n51,n1590);
and (n4770,n4771,n4772);
xor (n4771,n4769,n3914);
or (n4772,n4773,n4776);
and (n4773,n4774,n4775);
and (n4774,n323,n1590);
and (n4775,n535,n39);
and (n4776,n4777,n4778);
xor (n4777,n4774,n4775);
or (n4778,n4779,n4782);
and (n4779,n4780,n4781);
and (n4780,n535,n1590);
and (n4781,n853,n39);
and (n4782,n4783,n4784);
xor (n4783,n4780,n4781);
or (n4784,n4785,n4788);
and (n4785,n4786,n4787);
and (n4786,n853,n1590);
and (n4787,n847,n39);
and (n4788,n4789,n4790);
xor (n4789,n4786,n4787);
or (n4790,n4791,n4793);
and (n4791,n4792,n4410);
and (n4792,n847,n1590);
and (n4793,n4794,n4795);
xor (n4794,n4792,n4410);
or (n4795,n4796,n4799);
and (n4796,n4797,n4798);
and (n4797,n1241,n1590);
and (n4798,n1633,n39);
and (n4799,n4800,n4801);
xor (n4800,n4797,n4798);
and (n4801,n4802,n4803);
and (n4802,n1633,n1590);
and (n4803,n1829,n39);
and (n4804,n388,n33);
and (n4805,n4806,n4807);
xor (n4806,n4720,n4804);
or (n4807,n4808,n4811);
and (n4808,n4809,n4810);
xor (n4809,n1594,n4721);
and (n4810,n229,n33);
and (n4811,n4812,n4813);
xor (n4812,n4809,n4810);
or (n4813,n4814,n4817);
and (n4814,n4815,n4816);
xor (n4815,n4725,n4726);
and (n4816,n214,n33);
and (n4817,n4818,n4819);
xor (n4818,n4815,n4816);
or (n4819,n4820,n4823);
and (n4820,n4821,n4822);
xor (n4821,n4730,n4731);
and (n4822,n177,n33);
and (n4823,n4824,n4825);
xor (n4824,n4821,n4822);
or (n4825,n4826,n4829);
and (n4826,n4827,n4828);
xor (n4827,n4736,n4737);
and (n4828,n171,n33);
and (n4829,n4830,n4831);
xor (n4830,n4827,n4828);
or (n4831,n4832,n4835);
and (n4832,n4833,n4834);
xor (n4833,n4742,n4743);
and (n4834,n338,n33);
and (n4835,n4836,n4837);
xor (n4836,n4833,n4834);
or (n4837,n4838,n4841);
and (n4838,n4839,n4840);
xor (n4839,n4748,n4749);
and (n4840,n380,n33);
and (n4841,n4842,n4843);
xor (n4842,n4839,n4840);
or (n4843,n4844,n4847);
and (n4844,n4845,n4846);
xor (n4845,n4754,n4755);
and (n4846,n69,n33);
and (n4847,n4848,n4849);
xor (n4848,n4845,n4846);
or (n4849,n4850,n4853);
and (n4850,n4851,n4852);
xor (n4851,n4760,n4761);
and (n4852,n51,n33);
and (n4853,n4854,n4855);
xor (n4854,n4851,n4852);
or (n4855,n4856,n4859);
and (n4856,n4857,n4858);
xor (n4857,n4766,n4767);
and (n4858,n323,n33);
and (n4859,n4860,n4861);
xor (n4860,n4857,n4858);
or (n4861,n4862,n4865);
and (n4862,n4863,n4864);
xor (n4863,n4771,n4772);
and (n4864,n535,n33);
and (n4865,n4866,n4867);
xor (n4866,n4863,n4864);
or (n4867,n4868,n4871);
and (n4868,n4869,n4870);
xor (n4869,n4777,n4778);
and (n4870,n853,n33);
and (n4871,n4872,n4873);
xor (n4872,n4869,n4870);
or (n4873,n4874,n4877);
and (n4874,n4875,n4876);
xor (n4875,n4783,n4784);
and (n4876,n847,n33);
and (n4877,n4878,n4879);
xor (n4878,n4875,n4876);
or (n4879,n4880,n4883);
and (n4880,n4881,n4882);
xor (n4881,n4789,n4790);
and (n4882,n1241,n33);
and (n4883,n4884,n4885);
xor (n4884,n4881,n4882);
or (n4885,n4886,n4889);
and (n4886,n4887,n4888);
xor (n4887,n4794,n4795);
and (n4888,n1633,n33);
and (n4889,n4890,n4891);
xor (n4890,n4887,n4888);
and (n4891,n4892,n4893);
xor (n4892,n4800,n4801);
not (n4893,n4392);
and (n4894,n388,n35);
and (n4895,n4896,n4897);
xor (n4896,n4718,n4894);
or (n4897,n4898,n4901);
and (n4898,n4899,n4900);
xor (n4899,n4806,n4807);
and (n4900,n229,n35);
and (n4901,n4902,n4903);
xor (n4902,n4899,n4900);
or (n4903,n4904,n4907);
and (n4904,n4905,n4906);
xor (n4905,n4812,n4813);
and (n4906,n214,n35);
and (n4907,n4908,n4909);
xor (n4908,n4905,n4906);
or (n4909,n4910,n4912);
and (n4910,n4911,n2428);
xor (n4911,n4818,n4819);
and (n4912,n4913,n4914);
xor (n4913,n4911,n2428);
or (n4914,n4915,n4918);
and (n4915,n4916,n4917);
xor (n4916,n4824,n4825);
and (n4917,n171,n35);
and (n4918,n4919,n4920);
xor (n4919,n4916,n4917);
or (n4920,n4921,n4923);
and (n4921,n4922,n2205);
xor (n4922,n4830,n4831);
and (n4923,n4924,n4925);
xor (n4924,n4922,n2205);
or (n4925,n4926,n4929);
and (n4926,n4927,n4928);
xor (n4927,n4836,n4837);
and (n4928,n380,n35);
and (n4929,n4930,n4931);
xor (n4930,n4927,n4928);
or (n4931,n4932,n4935);
and (n4932,n4933,n4934);
xor (n4933,n4842,n4843);
and (n4934,n69,n35);
and (n4935,n4936,n4937);
xor (n4936,n4933,n4934);
or (n4937,n4938,n4940);
and (n4938,n4939,n3435);
xor (n4939,n4848,n4849);
and (n4940,n4941,n4942);
xor (n4941,n4939,n3435);
or (n4942,n4943,n4946);
and (n4943,n4944,n4945);
xor (n4944,n4854,n4855);
and (n4945,n323,n35);
and (n4946,n4947,n4948);
xor (n4947,n4944,n4945);
or (n4948,n4949,n4952);
and (n4949,n4950,n4951);
xor (n4950,n4860,n4861);
and (n4951,n535,n35);
and (n4952,n4953,n4954);
xor (n4953,n4950,n4951);
or (n4954,n4955,n4958);
and (n4955,n4956,n4957);
xor (n4956,n4866,n4867);
and (n4957,n853,n35);
and (n4958,n4959,n4960);
xor (n4959,n4956,n4957);
or (n4960,n4961,n4964);
and (n4961,n4962,n4963);
xor (n4962,n4872,n4873);
and (n4963,n847,n35);
and (n4964,n4965,n4966);
xor (n4965,n4962,n4963);
or (n4966,n4967,n4970);
and (n4967,n4968,n4969);
xor (n4968,n4878,n4879);
and (n4969,n1241,n35);
and (n4970,n4971,n4972);
xor (n4971,n4968,n4969);
or (n4972,n4973,n4976);
and (n4973,n4974,n4975);
xor (n4974,n4884,n4885);
and (n4975,n1633,n35);
and (n4976,n4977,n4978);
xor (n4977,n4974,n4975);
and (n4978,n4979,n4980);
xor (n4979,n4890,n4891);
and (n4980,n1829,n35);
and (n4981,n388,n396);
and (n4982,n4983,n4984);
xor (n4983,n4716,n4981);
or (n4984,n4985,n4988);
and (n4985,n4986,n4987);
xor (n4986,n4896,n4897);
and (n4987,n229,n396);
and (n4988,n4989,n4990);
xor (n4989,n4986,n4987);
or (n4990,n4991,n4994);
and (n4991,n4992,n4993);
xor (n4992,n4902,n4903);
and (n4993,n214,n396);
and (n4994,n4995,n4996);
xor (n4995,n4992,n4993);
or (n4996,n4997,n5000);
and (n4997,n4998,n4999);
xor (n4998,n4908,n4909);
and (n4999,n177,n396);
and (n5000,n5001,n5002);
xor (n5001,n4998,n4999);
or (n5002,n5003,n5006);
and (n5003,n5004,n5005);
xor (n5004,n4913,n4914);
and (n5005,n171,n396);
and (n5006,n5007,n5008);
xor (n5007,n5004,n5005);
or (n5008,n5009,n5012);
and (n5009,n5010,n5011);
xor (n5010,n4919,n4920);
and (n5011,n338,n396);
and (n5012,n5013,n5014);
xor (n5013,n5010,n5011);
or (n5014,n5015,n5018);
and (n5015,n5016,n5017);
xor (n5016,n4924,n4925);
and (n5017,n380,n396);
and (n5018,n5019,n5020);
xor (n5019,n5016,n5017);
or (n5020,n5021,n5024);
and (n5021,n5022,n5023);
xor (n5022,n4930,n4931);
and (n5023,n69,n396);
and (n5024,n5025,n5026);
xor (n5025,n5022,n5023);
or (n5026,n5027,n5030);
and (n5027,n5028,n5029);
xor (n5028,n4936,n4937);
and (n5029,n51,n396);
and (n5030,n5031,n5032);
xor (n5031,n5028,n5029);
or (n5032,n5033,n5036);
and (n5033,n5034,n5035);
xor (n5034,n4941,n4942);
and (n5035,n323,n396);
and (n5036,n5037,n5038);
xor (n5037,n5034,n5035);
or (n5038,n5039,n5042);
and (n5039,n5040,n5041);
xor (n5040,n4947,n4948);
and (n5041,n535,n396);
and (n5042,n5043,n5044);
xor (n5043,n5040,n5041);
or (n5044,n5045,n5048);
and (n5045,n5046,n5047);
xor (n5046,n4953,n4954);
and (n5047,n853,n396);
and (n5048,n5049,n5050);
xor (n5049,n5046,n5047);
or (n5050,n5051,n5054);
and (n5051,n5052,n5053);
xor (n5052,n4959,n4960);
and (n5053,n847,n396);
and (n5054,n5055,n5056);
xor (n5055,n5052,n5053);
or (n5056,n5057,n5060);
and (n5057,n5058,n5059);
xor (n5058,n4965,n4966);
and (n5059,n1241,n396);
and (n5060,n5061,n5062);
xor (n5061,n5058,n5059);
or (n5062,n5063,n5066);
and (n5063,n5064,n5065);
xor (n5064,n4971,n4972);
and (n5065,n1633,n396);
and (n5066,n5067,n5068);
xor (n5067,n5064,n5065);
and (n5068,n5069,n4127);
xor (n5069,n4977,n4978);
and (n5070,n388,n223);
and (n5071,n5072,n5073);
xor (n5072,n4714,n5070);
or (n5073,n5074,n5077);
and (n5074,n5075,n5076);
xor (n5075,n4983,n4984);
and (n5076,n229,n223);
and (n5077,n5078,n5079);
xor (n5078,n5075,n5076);
or (n5079,n5080,n5083);
and (n5080,n5081,n5082);
xor (n5081,n4989,n4990);
and (n5082,n214,n223);
and (n5083,n5084,n5085);
xor (n5084,n5081,n5082);
or (n5085,n5086,n5088);
and (n5086,n5087,n1343);
xor (n5087,n4995,n4996);
and (n5088,n5089,n5090);
xor (n5089,n5087,n1343);
or (n5090,n5091,n5093);
and (n5091,n5092,n1608);
xor (n5092,n5001,n5002);
and (n5093,n5094,n5095);
xor (n5094,n5092,n1608);
or (n5095,n5096,n5099);
and (n5096,n5097,n5098);
xor (n5097,n5007,n5008);
and (n5098,n338,n223);
and (n5099,n5100,n5101);
xor (n5100,n5097,n5098);
or (n5101,n5102,n5104);
and (n5102,n5103,n2271);
xor (n5103,n5013,n5014);
and (n5104,n5105,n5106);
xor (n5105,n5103,n2271);
or (n5106,n5107,n5109);
and (n5107,n5108,n2266);
xor (n5108,n5019,n5020);
and (n5109,n5110,n5111);
xor (n5110,n5108,n2266);
or (n5111,n5112,n5115);
and (n5112,n5113,n5114);
xor (n5113,n5025,n5026);
and (n5114,n51,n223);
and (n5115,n5116,n5117);
xor (n5116,n5113,n5114);
or (n5117,n5118,n5120);
and (n5118,n5119,n3036);
xor (n5119,n5031,n5032);
and (n5120,n5121,n5122);
xor (n5121,n5119,n3036);
or (n5122,n5123,n5125);
and (n5123,n5124,n3313);
xor (n5124,n5037,n5038);
and (n5125,n5126,n5127);
xor (n5126,n5124,n3313);
or (n5127,n5128,n5131);
and (n5128,n5129,n5130);
xor (n5129,n5043,n5044);
and (n5130,n853,n223);
and (n5131,n5132,n5133);
xor (n5132,n5129,n5130);
or (n5133,n5134,n5136);
and (n5134,n5135,n3725);
xor (n5135,n5049,n5050);
and (n5136,n5137,n5138);
xor (n5137,n5135,n3725);
or (n5138,n5139,n5141);
and (n5139,n5140,n3854);
xor (n5140,n5055,n5056);
and (n5141,n5142,n5143);
xor (n5142,n5140,n3854);
or (n5143,n5144,n5146);
and (n5144,n5145,n4018);
xor (n5145,n5061,n5062);
and (n5146,n5147,n5148);
xor (n5147,n5145,n4018);
and (n5148,n5149,n5150);
xor (n5149,n5067,n5068);
and (n5150,n1829,n223);
and (n5151,n388,n220);
and (n5152,n5153,n5154);
xor (n5153,n4712,n5151);
or (n5154,n5155,n5158);
and (n5155,n5156,n5157);
xor (n5156,n5072,n5073);
and (n5157,n229,n220);
and (n5158,n5159,n5160);
xor (n5159,n5156,n5157);
or (n5160,n5161,n5164);
and (n5161,n5162,n5163);
xor (n5162,n5078,n5079);
and (n5163,n214,n220);
and (n5164,n5165,n5166);
xor (n5165,n5162,n5163);
or (n5166,n5167,n5170);
and (n5167,n5168,n5169);
xor (n5168,n5084,n5085);
and (n5169,n177,n220);
and (n5170,n5171,n5172);
xor (n5171,n5168,n5169);
or (n5172,n5173,n5176);
and (n5173,n5174,n5175);
xor (n5174,n5089,n5090);
and (n5175,n171,n220);
and (n5176,n5177,n5178);
xor (n5177,n5174,n5175);
or (n5178,n5179,n5182);
and (n5179,n5180,n5181);
xor (n5180,n5094,n5095);
and (n5181,n338,n220);
and (n5182,n5183,n5184);
xor (n5183,n5180,n5181);
or (n5184,n5185,n5188);
and (n5185,n5186,n5187);
xor (n5186,n5100,n5101);
and (n5187,n380,n220);
and (n5188,n5189,n5190);
xor (n5189,n5186,n5187);
or (n5190,n5191,n5194);
and (n5191,n5192,n5193);
xor (n5192,n5105,n5106);
and (n5193,n69,n220);
and (n5194,n5195,n5196);
xor (n5195,n5192,n5193);
or (n5196,n5197,n5200);
and (n5197,n5198,n5199);
xor (n5198,n5110,n5111);
and (n5199,n51,n220);
and (n5200,n5201,n5202);
xor (n5201,n5198,n5199);
or (n5202,n5203,n5206);
and (n5203,n5204,n5205);
xor (n5204,n5116,n5117);
and (n5205,n323,n220);
and (n5206,n5207,n5208);
xor (n5207,n5204,n5205);
or (n5208,n5209,n5212);
and (n5209,n5210,n5211);
xor (n5210,n5121,n5122);
and (n5211,n535,n220);
and (n5212,n5213,n5214);
xor (n5213,n5210,n5211);
or (n5214,n5215,n5218);
and (n5215,n5216,n5217);
xor (n5216,n5126,n5127);
and (n5217,n853,n220);
and (n5218,n5219,n5220);
xor (n5219,n5216,n5217);
or (n5220,n5221,n5224);
and (n5221,n5222,n5223);
xor (n5222,n5132,n5133);
and (n5223,n847,n220);
and (n5224,n5225,n5226);
xor (n5225,n5222,n5223);
or (n5226,n5227,n5230);
and (n5227,n5228,n5229);
xor (n5228,n5137,n5138);
and (n5229,n1241,n220);
and (n5230,n5231,n5232);
xor (n5231,n5228,n5229);
or (n5232,n5233,n5236);
and (n5233,n5234,n5235);
xor (n5234,n5142,n5143);
and (n5235,n1633,n220);
and (n5236,n5237,n5238);
xor (n5237,n5234,n5235);
and (n5238,n5239,n5240);
xor (n5239,n5147,n5148);
not (n5240,n3837);
and (n5241,n388,n160);
and (n5242,n5243,n5244);
xor (n5243,n4710,n5241);
or (n5244,n5245,n5248);
and (n5245,n5246,n5247);
xor (n5246,n5153,n5154);
and (n5247,n229,n160);
and (n5248,n5249,n5250);
xor (n5249,n5246,n5247);
or (n5250,n5251,n5253);
and (n5251,n5252,n215);
xor (n5252,n5159,n5160);
and (n5253,n5254,n5255);
xor (n5254,n5252,n215);
or (n5255,n5256,n5259);
and (n5256,n5257,n5258);
xor (n5257,n5165,n5166);
and (n5258,n177,n160);
and (n5259,n5260,n5261);
xor (n5260,n5257,n5258);
or (n5261,n5262,n5265);
and (n5262,n5263,n5264);
xor (n5263,n5171,n5172);
and (n5264,n171,n160);
and (n5265,n5266,n5267);
xor (n5266,n5263,n5264);
or (n5267,n5268,n5271);
and (n5268,n5269,n5270);
xor (n5269,n5177,n5178);
and (n5270,n338,n160);
and (n5271,n5272,n5273);
xor (n5272,n5269,n5270);
or (n5273,n5274,n5277);
and (n5274,n5275,n5276);
xor (n5275,n5183,n5184);
and (n5276,n380,n160);
and (n5277,n5278,n5279);
xor (n5278,n5275,n5276);
or (n5279,n5280,n5283);
and (n5280,n5281,n5282);
xor (n5281,n5189,n5190);
and (n5282,n69,n160);
and (n5283,n5284,n5285);
xor (n5284,n5281,n5282);
or (n5285,n5286,n5289);
and (n5286,n5287,n5288);
xor (n5287,n5195,n5196);
and (n5288,n51,n160);
and (n5289,n5290,n5291);
xor (n5290,n5287,n5288);
or (n5291,n5292,n5295);
and (n5292,n5293,n5294);
xor (n5293,n5201,n5202);
and (n5294,n323,n160);
and (n5295,n5296,n5297);
xor (n5296,n5293,n5294);
or (n5297,n5298,n5300);
and (n5298,n5299,n2894);
xor (n5299,n5207,n5208);
and (n5300,n5301,n5302);
xor (n5301,n5299,n2894);
or (n5302,n5303,n5305);
and (n5303,n5304,n3209);
xor (n5304,n5213,n5214);
and (n5305,n5306,n5307);
xor (n5306,n5304,n3209);
or (n5307,n5308,n5311);
and (n5308,n5309,n5310);
xor (n5309,n5219,n5220);
and (n5310,n847,n160);
and (n5311,n5312,n5313);
xor (n5312,n5309,n5310);
or (n5313,n5314,n5317);
and (n5314,n5315,n5316);
xor (n5315,n5225,n5226);
and (n5316,n1241,n160);
and (n5317,n5318,n5319);
xor (n5318,n5315,n5316);
or (n5319,n5320,n5323);
and (n5320,n5321,n5322);
xor (n5321,n5231,n5232);
and (n5322,n1633,n160);
and (n5323,n5324,n5325);
xor (n5324,n5321,n5322);
and (n5325,n5326,n5327);
xor (n5326,n5237,n5238);
and (n5327,n1829,n160);
and (n5328,n388,n161);
or (n5329,n5330,n5333);
and (n5330,n5331,n5332);
xor (n5331,n5243,n5244);
and (n5332,n229,n161);
and (n5333,n5334,n5335);
xor (n5334,n5331,n5332);
or (n5335,n5336,n5339);
and (n5336,n5337,n5338);
xor (n5337,n5249,n5250);
and (n5338,n214,n161);
and (n5339,n5340,n5341);
xor (n5340,n5337,n5338);
or (n5341,n5342,n5345);
and (n5342,n5343,n5344);
xor (n5343,n5254,n5255);
and (n5344,n177,n161);
and (n5345,n5346,n5347);
xor (n5346,n5343,n5344);
or (n5347,n5348,n5351);
and (n5348,n5349,n5350);
xor (n5349,n5260,n5261);
and (n5350,n171,n161);
and (n5351,n5352,n5353);
xor (n5352,n5349,n5350);
or (n5353,n5354,n5357);
and (n5354,n5355,n5356);
xor (n5355,n5266,n5267);
and (n5356,n338,n161);
and (n5357,n5358,n5359);
xor (n5358,n5355,n5356);
or (n5359,n5360,n5363);
and (n5360,n5361,n5362);
xor (n5361,n5272,n5273);
and (n5362,n380,n161);
and (n5363,n5364,n5365);
xor (n5364,n5361,n5362);
or (n5365,n5366,n5369);
and (n5366,n5367,n5368);
xor (n5367,n5278,n5279);
and (n5368,n69,n161);
and (n5369,n5370,n5371);
xor (n5370,n5367,n5368);
or (n5371,n5372,n5375);
and (n5372,n5373,n5374);
xor (n5373,n5284,n5285);
and (n5374,n51,n161);
and (n5375,n5376,n5377);
xor (n5376,n5373,n5374);
or (n5377,n5378,n5381);
and (n5378,n5379,n5380);
xor (n5379,n5290,n5291);
and (n5380,n323,n161);
and (n5381,n5382,n5383);
xor (n5382,n5379,n5380);
or (n5383,n5384,n5387);
and (n5384,n5385,n5386);
xor (n5385,n5296,n5297);
and (n5386,n535,n161);
and (n5387,n5388,n5389);
xor (n5388,n5385,n5386);
or (n5389,n5390,n5393);
and (n5390,n5391,n5392);
xor (n5391,n5301,n5302);
and (n5392,n853,n161);
and (n5393,n5394,n5395);
xor (n5394,n5391,n5392);
or (n5395,n5396,n5399);
and (n5396,n5397,n5398);
xor (n5397,n5306,n5307);
and (n5398,n847,n161);
and (n5399,n5400,n5401);
xor (n5400,n5397,n5398);
or (n5401,n5402,n5405);
and (n5402,n5403,n5404);
xor (n5403,n5312,n5313);
and (n5404,n1241,n161);
and (n5405,n5406,n5407);
xor (n5406,n5403,n5404);
or (n5407,n5408,n5411);
and (n5408,n5409,n5410);
xor (n5409,n5318,n5319);
and (n5410,n1633,n161);
and (n5411,n5412,n5413);
xor (n5412,n5409,n5410);
and (n5413,n5414,n3570);
xor (n5414,n5324,n5325);
or (n5415,n5416,n5418);
and (n5416,n5417,n361);
xor (n5417,n5334,n5335);
and (n5418,n5419,n5420);
xor (n5419,n5417,n361);
or (n5420,n5421,n5424);
and (n5421,n5422,n5423);
xor (n5422,n5340,n5341);
and (n5423,n177,n167);
and (n5424,n5425,n5426);
xor (n5425,n5422,n5423);
or (n5426,n5427,n5430);
and (n5427,n5428,n5429);
xor (n5428,n5346,n5347);
and (n5429,n171,n167);
and (n5430,n5431,n5432);
xor (n5431,n5428,n5429);
or (n5432,n5433,n5436);
and (n5433,n5434,n5435);
xor (n5434,n5352,n5353);
and (n5435,n338,n167);
and (n5436,n5437,n5438);
xor (n5437,n5434,n5435);
or (n5438,n5439,n5442);
and (n5439,n5440,n5441);
xor (n5440,n5358,n5359);
and (n5441,n380,n167);
and (n5442,n5443,n5444);
xor (n5443,n5440,n5441);
or (n5444,n5445,n5447);
and (n5445,n5446,n1232);
xor (n5446,n5364,n5365);
and (n5447,n5448,n5449);
xor (n5448,n5446,n1232);
or (n5449,n5450,n5453);
and (n5450,n5451,n5452);
xor (n5451,n5370,n5371);
and (n5452,n51,n167);
and (n5453,n5454,n5455);
xor (n5454,n5451,n5452);
or (n5455,n5456,n5458);
and (n5456,n5457,n2511);
xor (n5457,n5376,n5377);
and (n5458,n5459,n5460);
xor (n5459,n5457,n2511);
or (n5460,n5461,n5464);
and (n5461,n5462,n5463);
xor (n5462,n5382,n5383);
and (n5463,n535,n167);
and (n5464,n5465,n5466);
xor (n5465,n5462,n5463);
or (n5466,n5467,n5469);
and (n5467,n5468,n2301);
xor (n5468,n5388,n5389);
and (n5469,n5470,n5471);
xor (n5470,n5468,n2301);
or (n5471,n5472,n5475);
and (n5472,n5473,n5474);
xor (n5473,n5394,n5395);
and (n5474,n847,n167);
and (n5475,n5476,n5477);
xor (n5476,n5473,n5474);
or (n5477,n5478,n5481);
and (n5478,n5479,n5480);
xor (n5479,n5400,n5401);
and (n5480,n1241,n167);
and (n5481,n5482,n5483);
xor (n5482,n5479,n5480);
or (n5483,n5484,n5487);
and (n5484,n5485,n5486);
xor (n5485,n5406,n5407);
and (n5486,n1633,n167);
and (n5487,n5488,n5489);
xor (n5488,n5485,n5486);
and (n5489,n5490,n5491);
xor (n5490,n5412,n5413);
and (n5491,n1829,n167);
and (n5492,n214,n344);
or (n5493,n5494,n5497);
and (n5494,n5495,n5496);
xor (n5495,n5419,n5420);
and (n5496,n177,n344);
and (n5497,n5498,n5499);
xor (n5498,n5495,n5496);
or (n5499,n5500,n5503);
and (n5500,n5501,n5502);
xor (n5501,n5425,n5426);
and (n5502,n171,n344);
and (n5503,n5504,n5505);
xor (n5504,n5501,n5502);
or (n5505,n5506,n5509);
and (n5506,n5507,n5508);
xor (n5507,n5431,n5432);
and (n5508,n338,n344);
and (n5509,n5510,n5511);
xor (n5510,n5507,n5508);
or (n5511,n5512,n5515);
and (n5512,n5513,n5514);
xor (n5513,n5437,n5438);
and (n5514,n380,n344);
and (n5515,n5516,n5517);
xor (n5516,n5513,n5514);
or (n5517,n5518,n5521);
and (n5518,n5519,n5520);
xor (n5519,n5443,n5444);
and (n5520,n69,n344);
and (n5521,n5522,n5523);
xor (n5522,n5519,n5520);
or (n5523,n5524,n5527);
and (n5524,n5525,n5526);
xor (n5525,n5448,n5449);
and (n5526,n51,n344);
and (n5527,n5528,n5529);
xor (n5528,n5525,n5526);
or (n5529,n5530,n5533);
and (n5530,n5531,n5532);
xor (n5531,n5454,n5455);
and (n5532,n323,n344);
and (n5533,n5534,n5535);
xor (n5534,n5531,n5532);
or (n5535,n5536,n5539);
and (n5536,n5537,n5538);
xor (n5537,n5459,n5460);
and (n5538,n535,n344);
and (n5539,n5540,n5541);
xor (n5540,n5537,n5538);
or (n5541,n5542,n5545);
and (n5542,n5543,n5544);
xor (n5543,n5465,n5466);
and (n5544,n853,n344);
and (n5545,n5546,n5547);
xor (n5546,n5543,n5544);
or (n5547,n5548,n5551);
and (n5548,n5549,n5550);
xor (n5549,n5470,n5471);
and (n5550,n847,n344);
and (n5551,n5552,n5553);
xor (n5552,n5549,n5550);
or (n5553,n5554,n5557);
and (n5554,n5555,n5556);
xor (n5555,n5476,n5477);
and (n5556,n1241,n344);
and (n5557,n5558,n5559);
xor (n5558,n5555,n5556);
or (n5559,n5560,n5563);
and (n5560,n5561,n5562);
xor (n5561,n5482,n5483);
and (n5562,n1633,n344);
and (n5563,n5564,n5565);
xor (n5564,n5561,n5562);
and (n5565,n5566,n5567);
xor (n5566,n5488,n5489);
not (n5567,n3112);
or (n5568,n5569,n5572);
and (n5569,n5570,n5571);
xor (n5570,n5498,n5499);
and (n5571,n171,n63);
and (n5572,n5573,n5574);
xor (n5573,n5570,n5571);
or (n5574,n5575,n5577);
and (n5575,n5576,n339);
xor (n5576,n5504,n5505);
and (n5577,n5578,n5579);
xor (n5578,n5576,n339);
or (n5579,n5580,n5582);
and (n5580,n5581,n543);
xor (n5581,n5510,n5511);
and (n5582,n5583,n5584);
xor (n5583,n5581,n543);
or (n5584,n5585,n5588);
and (n5585,n5586,n5587);
xor (n5586,n5516,n5517);
and (n5587,n69,n63);
and (n5588,n5589,n5590);
xor (n5589,n5586,n5587);
or (n5590,n5591,n5594);
and (n5591,n5592,n5593);
xor (n5592,n5522,n5523);
and (n5593,n51,n63);
and (n5594,n5595,n5596);
xor (n5595,n5592,n5593);
or (n5596,n5597,n5600);
and (n5597,n5598,n5599);
xor (n5598,n5528,n5529);
and (n5599,n323,n63);
and (n5600,n5601,n5602);
xor (n5601,n5598,n5599);
or (n5602,n5603,n5606);
and (n5603,n5604,n5605);
xor (n5604,n5534,n5535);
and (n5605,n535,n63);
and (n5606,n5607,n5608);
xor (n5607,n5604,n5605);
or (n5608,n5609,n5612);
and (n5609,n5610,n5611);
xor (n5610,n5540,n5541);
and (n5611,n853,n63);
and (n5612,n5613,n5614);
xor (n5613,n5610,n5611);
or (n5614,n5615,n5618);
and (n5615,n5616,n5617);
xor (n5616,n5546,n5547);
and (n5617,n847,n63);
and (n5618,n5619,n5620);
xor (n5619,n5616,n5617);
or (n5620,n5621,n5624);
and (n5621,n5622,n5623);
xor (n5622,n5552,n5553);
and (n5623,n1241,n63);
and (n5624,n5625,n5626);
xor (n5625,n5622,n5623);
or (n5626,n5627,n5630);
and (n5627,n5628,n5629);
xor (n5628,n5558,n5559);
and (n5629,n1633,n63);
and (n5630,n5631,n5632);
xor (n5631,n5628,n5629);
and (n5632,n5633,n5634);
xor (n5633,n5564,n5565);
and (n5634,n1829,n63);
and (n5635,n171,n58);
or (n5636,n5637,n5640);
and (n5637,n5638,n5639);
xor (n5638,n5573,n5574);
and (n5639,n338,n58);
and (n5640,n5641,n5642);
xor (n5641,n5638,n5639);
or (n5642,n5643,n5646);
and (n5643,n5644,n5645);
xor (n5644,n5578,n5579);
and (n5645,n380,n58);
and (n5646,n5647,n5648);
xor (n5647,n5644,n5645);
or (n5648,n5649,n5652);
and (n5649,n5650,n5651);
xor (n5650,n5583,n5584);
and (n5651,n69,n58);
and (n5652,n5653,n5654);
xor (n5653,n5650,n5651);
or (n5654,n5655,n5658);
and (n5655,n5656,n5657);
xor (n5656,n5589,n5590);
and (n5657,n51,n58);
and (n5658,n5659,n5660);
xor (n5659,n5656,n5657);
or (n5660,n5661,n5664);
and (n5661,n5662,n5663);
xor (n5662,n5595,n5596);
and (n5663,n323,n58);
and (n5664,n5665,n5666);
xor (n5665,n5662,n5663);
or (n5666,n5667,n5670);
and (n5667,n5668,n5669);
xor (n5668,n5601,n5602);
and (n5669,n535,n58);
and (n5670,n5671,n5672);
xor (n5671,n5668,n5669);
or (n5672,n5673,n5676);
and (n5673,n5674,n5675);
xor (n5674,n5607,n5608);
and (n5675,n853,n58);
and (n5676,n5677,n5678);
xor (n5677,n5674,n5675);
or (n5678,n5679,n5682);
and (n5679,n5680,n5681);
xor (n5680,n5613,n5614);
and (n5681,n847,n58);
and (n5682,n5683,n5684);
xor (n5683,n5680,n5681);
or (n5684,n5685,n5688);
and (n5685,n5686,n5687);
xor (n5686,n5619,n5620);
and (n5687,n1241,n58);
and (n5688,n5689,n5690);
xor (n5689,n5686,n5687);
or (n5690,n5691,n5694);
and (n5691,n5692,n5693);
xor (n5692,n5625,n5626);
and (n5693,n1633,n58);
and (n5694,n5695,n5696);
xor (n5695,n5692,n5693);
and (n5696,n5697,n5698);
xor (n5697,n5631,n5632);
not (n5698,n2360);
or (n5699,n5700,n5703);
and (n5700,n5701,n5702);
xor (n5701,n5641,n5642);
and (n5702,n380,n49);
and (n5703,n5704,n5705);
xor (n5704,n5701,n5702);
or (n5705,n5706,n5708);
and (n5706,n5707,n70);
xor (n5707,n5647,n5648);
and (n5708,n5709,n5710);
xor (n5709,n5707,n70);
or (n5710,n5711,n5713);
and (n5711,n5712,n52);
xor (n5712,n5653,n5654);
and (n5713,n5714,n5715);
xor (n5714,n5712,n52);
or (n5715,n5716,n5718);
and (n5716,n5717,n898);
xor (n5717,n5659,n5660);
and (n5718,n5719,n5720);
xor (n5719,n5717,n898);
or (n5720,n5721,n5724);
and (n5721,n5722,n5723);
xor (n5722,n5665,n5666);
and (n5723,n535,n49);
and (n5724,n5725,n5726);
xor (n5725,n5722,n5723);
or (n5726,n5727,n5730);
and (n5727,n5728,n5729);
xor (n5728,n5671,n5672);
and (n5729,n853,n49);
and (n5730,n5731,n5732);
xor (n5731,n5728,n5729);
or (n5732,n5733,n5735);
and (n5733,n5734,n1740);
xor (n5734,n5677,n5678);
and (n5735,n5736,n5737);
xor (n5736,n5734,n1740);
or (n5737,n5738,n5741);
and (n5738,n5739,n5740);
xor (n5739,n5683,n5684);
and (n5740,n1241,n49);
and (n5741,n5742,n5743);
xor (n5742,n5739,n5740);
or (n5743,n5744,n5747);
and (n5744,n5745,n5746);
xor (n5745,n5689,n5690);
and (n5746,n1633,n49);
and (n5747,n5748,n5749);
xor (n5748,n5745,n5746);
and (n5749,n5750,n5751);
xor (n5750,n5695,n5696);
and (n5751,n1829,n49);
and (n5752,n380,n312);
or (n5753,n5754,n5757);
and (n5754,n5755,n5756);
xor (n5755,n5704,n5705);
and (n5756,n69,n312);
and (n5757,n5758,n5759);
xor (n5758,n5755,n5756);
or (n5759,n5760,n5763);
and (n5760,n5761,n5762);
xor (n5761,n5709,n5710);
and (n5762,n51,n312);
and (n5763,n5764,n5765);
xor (n5764,n5761,n5762);
or (n5765,n5766,n5769);
and (n5766,n5767,n5768);
xor (n5767,n5714,n5715);
and (n5768,n323,n312);
and (n5769,n5770,n5771);
xor (n5770,n5767,n5768);
or (n5771,n5772,n5775);
and (n5772,n5773,n5774);
xor (n5773,n5719,n5720);
and (n5774,n535,n312);
and (n5775,n5776,n5777);
xor (n5776,n5773,n5774);
or (n5777,n5778,n5781);
and (n5778,n5779,n5780);
xor (n5779,n5725,n5726);
and (n5780,n853,n312);
and (n5781,n5782,n5783);
xor (n5782,n5779,n5780);
or (n5783,n5784,n5787);
and (n5784,n5785,n5786);
xor (n5785,n5731,n5732);
and (n5786,n847,n312);
and (n5787,n5788,n5789);
xor (n5788,n5785,n5786);
or (n5789,n5790,n5793);
and (n5790,n5791,n5792);
xor (n5791,n5736,n5737);
and (n5792,n1241,n312);
and (n5793,n5794,n5795);
xor (n5794,n5791,n5792);
or (n5795,n5796,n5799);
and (n5796,n5797,n5798);
xor (n5797,n5742,n5743);
and (n5798,n1633,n312);
and (n5799,n5800,n5801);
xor (n5800,n5797,n5798);
and (n5801,n5802,n1828);
xor (n5802,n5748,n5749);
and (n5803,n69,n313);
or (n5804,n5805,n5808);
and (n5805,n5806,n5807);
xor (n5806,n5758,n5759);
and (n5807,n51,n313);
and (n5808,n5809,n5810);
xor (n5809,n5806,n5807);
or (n5810,n5811,n5814);
and (n5811,n5812,n5813);
xor (n5812,n5764,n5765);
and (n5813,n323,n313);
and (n5814,n5815,n5816);
xor (n5815,n5812,n5813);
or (n5816,n5817,n5820);
and (n5817,n5818,n5819);
xor (n5818,n5770,n5771);
and (n5819,n535,n313);
and (n5820,n5821,n5822);
xor (n5821,n5818,n5819);
or (n5822,n5823,n5825);
and (n5823,n5824,n854);
xor (n5824,n5776,n5777);
and (n5825,n5826,n5827);
xor (n5826,n5824,n854);
or (n5827,n5828,n5830);
and (n5828,n5829,n848);
xor (n5829,n5782,n5783);
and (n5830,n5831,n5832);
xor (n5831,n5829,n848);
or (n5832,n5833,n5835);
and (n5833,n5834,n1242);
xor (n5834,n5788,n5789);
and (n5835,n5836,n5837);
xor (n5836,n5834,n1242);
or (n5837,n5838,n5841);
and (n5838,n5839,n5840);
xor (n5839,n5794,n5795);
and (n5840,n1633,n313);
and (n5841,n5842,n5843);
xor (n5842,n5839,n5840);
and (n5843,n5844,n5845);
xor (n5844,n5800,n5801);
and (n5845,n1829,n313);
or (n5846,n5847,n5849);
and (n5847,n5848,n5813);
xor (n5848,n5809,n5810);
and (n5849,n5850,n5851);
xor (n5850,n5848,n5813);
or (n5851,n5852,n5854);
and (n5852,n5853,n5819);
xor (n5853,n5815,n5816);
and (n5854,n5855,n5856);
xor (n5855,n5853,n5819);
or (n5856,n5857,n5859);
and (n5857,n5858,n854);
xor (n5858,n5821,n5822);
and (n5859,n5860,n5861);
xor (n5860,n5858,n854);
or (n5861,n5862,n5864);
and (n5862,n5863,n848);
xor (n5863,n5826,n5827);
and (n5864,n5865,n5866);
xor (n5865,n5863,n848);
or (n5866,n5867,n5869);
and (n5867,n5868,n1242);
xor (n5868,n5831,n5832);
and (n5869,n5870,n5871);
xor (n5870,n5868,n1242);
or (n5871,n5872,n5874);
and (n5872,n5873,n5840);
xor (n5873,n5836,n5837);
and (n5874,n5875,n5876);
xor (n5875,n5873,n5840);
and (n5876,n5877,n5845);
xor (n5877,n5842,n5843);
or (n5878,n5879,n5881);
and (n5879,n5880,n5819);
xor (n5880,n5850,n5851);
and (n5881,n5882,n5883);
xor (n5882,n5880,n5819);
or (n5883,n5884,n5886);
and (n5884,n5885,n854);
xor (n5885,n5855,n5856);
and (n5886,n5887,n5888);
xor (n5887,n5885,n854);
or (n5888,n5889,n5891);
and (n5889,n5890,n848);
xor (n5890,n5860,n5861);
and (n5891,n5892,n5893);
xor (n5892,n5890,n848);
or (n5893,n5894,n5896);
and (n5894,n5895,n1242);
xor (n5895,n5865,n5866);
and (n5896,n5897,n5898);
xor (n5897,n5895,n1242);
or (n5898,n5899,n5901);
and (n5899,n5900,n5840);
xor (n5900,n5870,n5871);
and (n5901,n5902,n5903);
xor (n5902,n5900,n5840);
and (n5903,n5904,n5845);
xor (n5904,n5875,n5876);
or (n5905,n5906,n5908);
and (n5906,n5907,n854);
xor (n5907,n5882,n5883);
and (n5908,n5909,n5910);
xor (n5909,n5907,n854);
or (n5910,n5911,n5913);
and (n5911,n5912,n848);
xor (n5912,n5887,n5888);
and (n5913,n5914,n5915);
xor (n5914,n5912,n848);
or (n5915,n5916,n5918);
and (n5916,n5917,n1242);
xor (n5917,n5892,n5893);
and (n5918,n5919,n5920);
xor (n5919,n5917,n1242);
or (n5920,n5921,n5923);
and (n5921,n5922,n5840);
xor (n5922,n5897,n5898);
and (n5923,n5924,n5925);
xor (n5924,n5922,n5840);
and (n5925,n5926,n5845);
xor (n5926,n5902,n5903);
or (n5927,n5928,n5930);
and (n5928,n5929,n848);
xor (n5929,n5909,n5910);
and (n5930,n5931,n5932);
xor (n5931,n5929,n848);
or (n5932,n5933,n5935);
and (n5933,n5934,n1242);
xor (n5934,n5914,n5915);
and (n5935,n5936,n5937);
xor (n5936,n5934,n1242);
or (n5937,n5938,n5940);
and (n5938,n5939,n5840);
xor (n5939,n5919,n5920);
and (n5940,n5941,n5942);
xor (n5941,n5939,n5840);
and (n5942,n5943,n5845);
xor (n5943,n5924,n5925);
or (n5944,n5945,n5947);
and (n5945,n5946,n1242);
xor (n5946,n5931,n5932);
and (n5947,n5948,n5949);
xor (n5948,n5946,n1242);
or (n5949,n5950,n5952);
and (n5950,n5951,n5840);
xor (n5951,n5936,n5937);
and (n5952,n5953,n5954);
xor (n5953,n5951,n5840);
and (n5954,n5955,n5845);
xor (n5955,n5941,n5942);
or (n5956,n5957,n5959);
and (n5957,n5958,n5840);
xor (n5958,n5948,n5949);
and (n5959,n5960,n5961);
xor (n5960,n5958,n5840);
and (n5961,n5962,n5845);
xor (n5962,n5953,n5954);
and (n5963,n5964,n5845);
xor (n5964,n5960,n5961);
xor (n5965,n5966,n2599);
xor (n5966,n5967,n7245);
xor (n5967,n5968,n1560);
xor (n5968,n5969,n7238);
xor (n5969,n5970,n7118);
xor (n5970,n5971,n7226);
xor (n5971,n5972,n652);
xor (n5972,n5973,n7209);
xor (n5973,n5974,n661);
xor (n5974,n5975,n7187);
xor (n5975,n5976,n1034);
xor (n5976,n5977,n7160);
xor (n5977,n5978,n287);
xor (n5978,n5979,n7128);
xor (n5979,n5980,n7092);
xor (n5980,n5981,n7089);
xor (n5981,n5982,n1425);
xor (n5982,n5983,n7038);
xor (n5983,n5984,n7037);
xor (n5984,n5985,n6982);
xor (n5985,n5986,n6981);
xor (n5986,n5987,n6918);
xor (n5987,n5988,n6917);
xor (n5988,n5989,n6854);
xor (n5989,n5990,n6853);
xor (n5990,n5991,n6779);
xor (n5991,n5992,n6778);
xor (n5992,n5993,n6702);
xor (n5993,n5994,n1400);
xor (n5994,n5995,n6615);
xor (n5995,n5996,n6614);
or (n5996,n5997,n6531);
and (n5997,n5998,n6530);
or (n5998,n5999,n6442);
and (n5999,n6000,n6441);
or (n6000,n6001,n6354);
and (n6001,n6002,n6353);
or (n6002,n6003,n6264);
and (n6003,n6004,n6263);
or (n6004,n6005,n6180);
and (n6005,n6006,n6179);
or (n6006,n6007,n6091);
and (n6007,n6008,n6090);
and (n6008,n1730,n6009);
or (n6009,n6010,n6012);
and (n6010,n6011,n2075);
and (n6011,n238,n1734);
and (n6012,n6013,n6014);
xor (n6013,n6011,n2075);
or (n6014,n6015,n6017);
and (n6015,n6016,n2229);
and (n6016,n152,n1734);
and (n6017,n6018,n6019);
xor (n6018,n6016,n2229);
or (n6019,n6020,n6022);
and (n6020,n6021,n2233);
and (n6021,n134,n1734);
and (n6022,n6023,n6024);
xor (n6023,n6021,n2233);
or (n6024,n6025,n6027);
and (n6025,n6026,n2818);
and (n6026,n473,n1734);
and (n6027,n6028,n6029);
xor (n6028,n6026,n2818);
or (n6029,n6030,n6033);
and (n6030,n6031,n6032);
and (n6031,n368,n1734);
and (n6032,n96,n679);
and (n6033,n6034,n6035);
xor (n6034,n6031,n6032);
or (n6035,n6036,n6039);
and (n6036,n6037,n6038);
and (n6037,n96,n1734);
and (n6038,n77,n679);
and (n6039,n6040,n6041);
xor (n6040,n6037,n6038);
or (n6041,n6042,n6045);
and (n6042,n6043,n6044);
and (n6043,n77,n1734);
and (n6044,n565,n679);
and (n6045,n6046,n6047);
xor (n6046,n6043,n6044);
or (n6047,n6048,n6051);
and (n6048,n6049,n6050);
and (n6049,n565,n1734);
and (n6050,n303,n679);
and (n6051,n6052,n6053);
xor (n6052,n6049,n6050);
or (n6053,n6054,n6057);
and (n6054,n6055,n6056);
and (n6055,n303,n1734);
and (n6056,n286,n679);
and (n6057,n6058,n6059);
xor (n6058,n6055,n6056);
or (n6059,n6060,n6063);
and (n6060,n6061,n6062);
and (n6061,n286,n1734);
and (n6062,n615,n679);
and (n6063,n6064,n6065);
xor (n6064,n6061,n6062);
or (n6065,n6066,n6069);
and (n6066,n6067,n6068);
and (n6067,n615,n1734);
and (n6068,n660,n679);
and (n6069,n6070,n6071);
xor (n6070,n6067,n6068);
or (n6071,n6072,n6074);
and (n6072,n6073,n4255);
and (n6073,n660,n1734);
and (n6074,n6075,n6076);
xor (n6075,n6073,n4255);
or (n6076,n6077,n6079);
and (n6077,n6078,n4348);
and (n6078,n653,n1734);
and (n6079,n6080,n6081);
xor (n6080,n6078,n4348);
or (n6081,n6082,n6085);
and (n6082,n6083,n6084);
and (n6083,n1260,n1734);
and (n6084,n1559,n679);
and (n6085,n6086,n6087);
xor (n6086,n6083,n6084);
and (n6087,n6088,n6089);
and (n6088,n1559,n1734);
and (n6089,n1835,n679);
and (n6090,n238,n794);
and (n6091,n6092,n6093);
xor (n6092,n6008,n6090);
or (n6093,n6094,n6097);
and (n6094,n6095,n6096);
xor (n6095,n1730,n6009);
and (n6096,n152,n794);
and (n6097,n6098,n6099);
xor (n6098,n6095,n6096);
or (n6099,n6100,n6103);
and (n6100,n6101,n6102);
xor (n6101,n6013,n6014);
and (n6102,n134,n794);
and (n6103,n6104,n6105);
xor (n6104,n6101,n6102);
or (n6105,n6106,n6109);
and (n6106,n6107,n6108);
xor (n6107,n6018,n6019);
and (n6108,n473,n794);
and (n6109,n6110,n6111);
xor (n6110,n6107,n6108);
or (n6111,n6112,n6115);
and (n6112,n6113,n6114);
xor (n6113,n6023,n6024);
and (n6114,n368,n794);
and (n6115,n6116,n6117);
xor (n6116,n6113,n6114);
or (n6117,n6118,n6121);
and (n6118,n6119,n6120);
xor (n6119,n6028,n6029);
and (n6120,n96,n794);
and (n6121,n6122,n6123);
xor (n6122,n6119,n6120);
or (n6123,n6124,n6127);
and (n6124,n6125,n6126);
xor (n6125,n6034,n6035);
and (n6126,n77,n794);
and (n6127,n6128,n6129);
xor (n6128,n6125,n6126);
or (n6129,n6130,n6133);
and (n6130,n6131,n6132);
xor (n6131,n6040,n6041);
and (n6132,n565,n794);
and (n6133,n6134,n6135);
xor (n6134,n6131,n6132);
or (n6135,n6136,n6139);
and (n6136,n6137,n6138);
xor (n6137,n6046,n6047);
and (n6138,n303,n794);
and (n6139,n6140,n6141);
xor (n6140,n6137,n6138);
or (n6141,n6142,n6145);
and (n6142,n6143,n6144);
xor (n6143,n6052,n6053);
and (n6144,n286,n794);
and (n6145,n6146,n6147);
xor (n6146,n6143,n6144);
or (n6147,n6148,n6151);
and (n6148,n6149,n6150);
xor (n6149,n6058,n6059);
and (n6150,n615,n794);
and (n6151,n6152,n6153);
xor (n6152,n6149,n6150);
or (n6153,n6154,n6157);
and (n6154,n6155,n6156);
xor (n6155,n6064,n6065);
and (n6156,n660,n794);
and (n6157,n6158,n6159);
xor (n6158,n6155,n6156);
or (n6159,n6160,n6163);
and (n6160,n6161,n6162);
xor (n6161,n6070,n6071);
and (n6162,n653,n794);
and (n6163,n6164,n6165);
xor (n6164,n6161,n6162);
or (n6165,n6166,n6169);
and (n6166,n6167,n6168);
xor (n6167,n6075,n6076);
and (n6168,n1260,n794);
and (n6169,n6170,n6171);
xor (n6170,n6167,n6168);
or (n6171,n6172,n6175);
and (n6172,n6173,n6174);
xor (n6173,n6080,n6081);
and (n6174,n1559,n794);
and (n6175,n6176,n6177);
xor (n6176,n6173,n6174);
and (n6177,n6178,n4388);
xor (n6178,n6086,n6087);
and (n6179,n238,n245);
and (n6180,n6181,n6182);
xor (n6181,n6006,n6179);
or (n6182,n6183,n6186);
and (n6183,n6184,n6185);
xor (n6184,n6092,n6093);
and (n6185,n152,n245);
and (n6186,n6187,n6188);
xor (n6187,n6184,n6185);
or (n6188,n6189,n6192);
and (n6189,n6190,n6191);
xor (n6190,n6098,n6099);
and (n6191,n134,n245);
and (n6192,n6193,n6194);
xor (n6193,n6190,n6191);
or (n6194,n6195,n6198);
and (n6195,n6196,n6197);
xor (n6196,n6104,n6105);
and (n6197,n473,n245);
and (n6198,n6199,n6200);
xor (n6199,n6196,n6197);
or (n6200,n6201,n6204);
and (n6201,n6202,n6203);
xor (n6202,n6110,n6111);
and (n6203,n368,n245);
and (n6204,n6205,n6206);
xor (n6205,n6202,n6203);
or (n6206,n6207,n6209);
and (n6207,n6208,n2387);
xor (n6208,n6116,n6117);
and (n6209,n6210,n6211);
xor (n6210,n6208,n2387);
or (n6211,n6212,n6215);
and (n6212,n6213,n6214);
xor (n6213,n6122,n6123);
and (n6214,n77,n245);
and (n6215,n6216,n6217);
xor (n6216,n6213,n6214);
or (n6217,n6218,n6221);
and (n6218,n6219,n6220);
xor (n6219,n6128,n6129);
and (n6220,n565,n245);
and (n6221,n6222,n6223);
xor (n6222,n6219,n6220);
or (n6223,n6224,n6227);
and (n6224,n6225,n6226);
xor (n6225,n6134,n6135);
and (n6226,n303,n245);
and (n6227,n6228,n6229);
xor (n6228,n6225,n6226);
or (n6229,n6230,n6232);
and (n6230,n6231,n3595);
xor (n6231,n6140,n6141);
and (n6232,n6233,n6234);
xor (n6233,n6231,n3595);
or (n6234,n6235,n6237);
and (n6235,n6236,n3781);
xor (n6236,n6146,n6147);
and (n6237,n6238,n6239);
xor (n6238,n6236,n3781);
or (n6239,n6240,n6242);
and (n6240,n6241,n3925);
xor (n6241,n6152,n6153);
and (n6242,n6243,n6244);
xor (n6243,n6241,n3925);
or (n6244,n6245,n6247);
and (n6245,n6246,n4069);
xor (n6246,n6158,n6159);
and (n6247,n6248,n6249);
xor (n6248,n6246,n4069);
or (n6249,n6250,n6253);
and (n6250,n6251,n6252);
xor (n6251,n6164,n6165);
and (n6252,n1260,n245);
and (n6253,n6254,n6255);
xor (n6254,n6251,n6252);
or (n6255,n6256,n6258);
and (n6256,n6257,n4296);
xor (n6257,n6170,n6171);
and (n6258,n6259,n6260);
xor (n6259,n6257,n4296);
and (n6260,n6261,n6262);
xor (n6261,n6176,n6177);
and (n6262,n1835,n245);
and (n6263,n238,n246);
and (n6264,n6265,n6266);
xor (n6265,n6004,n6263);
or (n6266,n6267,n6270);
and (n6267,n6268,n6269);
xor (n6268,n6181,n6182);
and (n6269,n152,n246);
and (n6270,n6271,n6272);
xor (n6271,n6268,n6269);
or (n6272,n6273,n6276);
and (n6273,n6274,n6275);
xor (n6274,n6187,n6188);
and (n6275,n134,n246);
and (n6276,n6277,n6278);
xor (n6277,n6274,n6275);
or (n6278,n6279,n6282);
and (n6279,n6280,n6281);
xor (n6280,n6193,n6194);
and (n6281,n473,n246);
and (n6282,n6283,n6284);
xor (n6283,n6280,n6281);
or (n6284,n6285,n6288);
and (n6285,n6286,n6287);
xor (n6286,n6199,n6200);
and (n6287,n368,n246);
and (n6288,n6289,n6290);
xor (n6289,n6286,n6287);
or (n6290,n6291,n6294);
and (n6291,n6292,n6293);
xor (n6292,n6205,n6206);
and (n6293,n96,n246);
and (n6294,n6295,n6296);
xor (n6295,n6292,n6293);
or (n6296,n6297,n6300);
and (n6297,n6298,n6299);
xor (n6298,n6210,n6211);
and (n6299,n77,n246);
and (n6300,n6301,n6302);
xor (n6301,n6298,n6299);
or (n6302,n6303,n6306);
and (n6303,n6304,n6305);
xor (n6304,n6216,n6217);
and (n6305,n565,n246);
and (n6306,n6307,n6308);
xor (n6307,n6304,n6305);
or (n6308,n6309,n6312);
and (n6309,n6310,n6311);
xor (n6310,n6222,n6223);
and (n6311,n303,n246);
and (n6312,n6313,n6314);
xor (n6313,n6310,n6311);
or (n6314,n6315,n6318);
and (n6315,n6316,n6317);
xor (n6316,n6228,n6229);
and (n6317,n286,n246);
and (n6318,n6319,n6320);
xor (n6319,n6316,n6317);
or (n6320,n6321,n6324);
and (n6321,n6322,n6323);
xor (n6322,n6233,n6234);
and (n6323,n615,n246);
and (n6324,n6325,n6326);
xor (n6325,n6322,n6323);
or (n6326,n6327,n6330);
and (n6327,n6328,n6329);
xor (n6328,n6238,n6239);
and (n6329,n660,n246);
and (n6330,n6331,n6332);
xor (n6331,n6328,n6329);
or (n6332,n6333,n6336);
and (n6333,n6334,n6335);
xor (n6334,n6243,n6244);
and (n6335,n653,n246);
and (n6336,n6337,n6338);
xor (n6337,n6334,n6335);
or (n6338,n6339,n6342);
and (n6339,n6340,n6341);
xor (n6340,n6248,n6249);
and (n6341,n1260,n246);
and (n6342,n6343,n6344);
xor (n6343,n6340,n6341);
or (n6344,n6345,n6348);
and (n6345,n6346,n6347);
xor (n6346,n6254,n6255);
and (n6347,n1559,n246);
and (n6348,n6349,n6350);
xor (n6349,n6346,n6347);
and (n6350,n6351,n6352);
xor (n6351,n6259,n6260);
not (n6352,n4133);
and (n6353,n238,n143);
and (n6354,n6355,n6356);
xor (n6355,n6002,n6353);
or (n6356,n6357,n6360);
and (n6357,n6358,n6359);
xor (n6358,n6265,n6266);
and (n6359,n152,n143);
and (n6360,n6361,n6362);
xor (n6361,n6358,n6359);
or (n6362,n6363,n6366);
and (n6363,n6364,n6365);
xor (n6364,n6271,n6272);
and (n6365,n134,n143);
and (n6366,n6367,n6368);
xor (n6367,n6364,n6365);
or (n6368,n6369,n6372);
and (n6369,n6370,n6371);
xor (n6370,n6277,n6278);
and (n6371,n473,n143);
and (n6372,n6373,n6374);
xor (n6373,n6370,n6371);
or (n6374,n6375,n6378);
and (n6375,n6376,n6377);
xor (n6376,n6283,n6284);
and (n6377,n368,n143);
and (n6378,n6379,n6380);
xor (n6379,n6376,n6377);
or (n6380,n6381,n6384);
and (n6381,n6382,n6383);
xor (n6382,n6289,n6290);
and (n6383,n96,n143);
and (n6384,n6385,n6386);
xor (n6385,n6382,n6383);
or (n6386,n6387,n6390);
and (n6387,n6388,n6389);
xor (n6388,n6295,n6296);
and (n6389,n77,n143);
and (n6390,n6391,n6392);
xor (n6391,n6388,n6389);
or (n6392,n6393,n6396);
and (n6393,n6394,n6395);
xor (n6394,n6301,n6302);
and (n6395,n565,n143);
and (n6396,n6397,n6398);
xor (n6397,n6394,n6395);
or (n6398,n6399,n6402);
and (n6399,n6400,n6401);
xor (n6400,n6307,n6308);
and (n6401,n303,n143);
and (n6402,n6403,n6404);
xor (n6403,n6400,n6401);
or (n6404,n6405,n6408);
and (n6405,n6406,n6407);
xor (n6406,n6313,n6314);
and (n6407,n286,n143);
and (n6408,n6409,n6410);
xor (n6409,n6406,n6407);
or (n6410,n6411,n6413);
and (n6411,n6412,n3396);
xor (n6412,n6319,n6320);
and (n6413,n6414,n6415);
xor (n6414,n6412,n3396);
or (n6415,n6416,n6419);
and (n6416,n6417,n6418);
xor (n6417,n6325,n6326);
and (n6418,n660,n143);
and (n6419,n6420,n6421);
xor (n6420,n6417,n6418);
or (n6421,n6422,n6425);
and (n6422,n6423,n6424);
xor (n6423,n6331,n6332);
and (n6424,n653,n143);
and (n6425,n6426,n6427);
xor (n6426,n6423,n6424);
or (n6427,n6428,n6430);
and (n6428,n6429,n3899);
xor (n6429,n6337,n6338);
and (n6430,n6431,n6432);
xor (n6431,n6429,n3899);
or (n6432,n6433,n6436);
and (n6433,n6434,n6435);
xor (n6434,n6343,n6344);
and (n6435,n1559,n143);
and (n6436,n6437,n6438);
xor (n6437,n6434,n6435);
and (n6438,n6439,n6440);
xor (n6439,n6349,n6350);
and (n6440,n1835,n143);
and (n6441,n238,n142);
and (n6442,n6443,n6444);
xor (n6443,n6000,n6441);
or (n6444,n6445,n6448);
and (n6445,n6446,n6447);
xor (n6446,n6355,n6356);
and (n6447,n152,n142);
and (n6448,n6449,n6450);
xor (n6449,n6446,n6447);
or (n6450,n6451,n6454);
and (n6451,n6452,n6453);
xor (n6452,n6361,n6362);
and (n6453,n134,n142);
and (n6454,n6455,n6456);
xor (n6455,n6452,n6453);
or (n6456,n6457,n6460);
and (n6457,n6458,n6459);
xor (n6458,n6367,n6368);
and (n6459,n473,n142);
and (n6460,n6461,n6462);
xor (n6461,n6458,n6459);
or (n6462,n6463,n6466);
and (n6463,n6464,n6465);
xor (n6464,n6373,n6374);
and (n6465,n368,n142);
and (n6466,n6467,n6468);
xor (n6467,n6464,n6465);
or (n6468,n6469,n6472);
and (n6469,n6470,n6471);
xor (n6470,n6379,n6380);
and (n6471,n96,n142);
and (n6472,n6473,n6474);
xor (n6473,n6470,n6471);
or (n6474,n6475,n6478);
and (n6475,n6476,n6477);
xor (n6476,n6385,n6386);
and (n6477,n77,n142);
and (n6478,n6479,n6480);
xor (n6479,n6476,n6477);
or (n6480,n6481,n6484);
and (n6481,n6482,n6483);
xor (n6482,n6391,n6392);
and (n6483,n565,n142);
and (n6484,n6485,n6486);
xor (n6485,n6482,n6483);
or (n6486,n6487,n6490);
and (n6487,n6488,n6489);
xor (n6488,n6397,n6398);
and (n6489,n303,n142);
and (n6490,n6491,n6492);
xor (n6491,n6488,n6489);
or (n6492,n6493,n6496);
and (n6493,n6494,n6495);
xor (n6494,n6403,n6404);
and (n6495,n286,n142);
and (n6496,n6497,n6498);
xor (n6497,n6494,n6495);
or (n6498,n6499,n6502);
and (n6499,n6500,n6501);
xor (n6500,n6409,n6410);
and (n6501,n615,n142);
and (n6502,n6503,n6504);
xor (n6503,n6500,n6501);
or (n6504,n6505,n6508);
and (n6505,n6506,n6507);
xor (n6506,n6414,n6415);
and (n6507,n660,n142);
and (n6508,n6509,n6510);
xor (n6509,n6506,n6507);
or (n6510,n6511,n6514);
and (n6511,n6512,n6513);
xor (n6512,n6420,n6421);
and (n6513,n653,n142);
and (n6514,n6515,n6516);
xor (n6515,n6512,n6513);
or (n6516,n6517,n6520);
and (n6517,n6518,n6519);
xor (n6518,n6426,n6427);
and (n6519,n1260,n142);
and (n6520,n6521,n6522);
xor (n6521,n6518,n6519);
or (n6522,n6523,n6526);
and (n6523,n6524,n6525);
xor (n6524,n6431,n6432);
and (n6525,n1559,n142);
and (n6526,n6527,n6528);
xor (n6527,n6524,n6525);
and (n6528,n6529,n3842);
xor (n6529,n6437,n6438);
and (n6530,n238,n133);
and (n6531,n6532,n6533);
xor (n6532,n5998,n6530);
or (n6533,n6534,n6536);
and (n6534,n6535,n153);
xor (n6535,n6443,n6444);
and (n6536,n6537,n6538);
xor (n6537,n6535,n153);
or (n6538,n6539,n6542);
and (n6539,n6540,n6541);
xor (n6540,n6449,n6450);
and (n6541,n134,n133);
and (n6542,n6543,n6544);
xor (n6543,n6540,n6541);
or (n6544,n6545,n6548);
and (n6545,n6546,n6547);
xor (n6546,n6455,n6456);
and (n6547,n473,n133);
and (n6548,n6549,n6550);
xor (n6549,n6546,n6547);
or (n6550,n6551,n6553);
and (n6551,n6552,n695);
xor (n6552,n6461,n6462);
and (n6553,n6554,n6555);
xor (n6554,n6552,n695);
or (n6555,n6556,n6558);
and (n6556,n6557,n1294);
xor (n6557,n6467,n6468);
and (n6558,n6559,n6560);
xor (n6559,n6557,n1294);
or (n6560,n6561,n6563);
and (n6561,n6562,n1688);
xor (n6562,n6473,n6474);
and (n6563,n6564,n6565);
xor (n6564,n6562,n1688);
or (n6565,n6566,n6569);
and (n6566,n6567,n6568);
xor (n6567,n6479,n6480);
and (n6568,n565,n133);
and (n6569,n6570,n6571);
xor (n6570,n6567,n6568);
or (n6571,n6572,n6575);
and (n6572,n6573,n6574);
xor (n6573,n6485,n6486);
and (n6574,n303,n133);
and (n6575,n6576,n6577);
xor (n6576,n6573,n6574);
or (n6577,n6578,n6581);
and (n6578,n6579,n6580);
xor (n6579,n6491,n6492);
and (n6580,n286,n133);
and (n6581,n6582,n6583);
xor (n6582,n6579,n6580);
or (n6583,n6584,n6587);
and (n6584,n6585,n6586);
xor (n6585,n6497,n6498);
and (n6586,n615,n133);
and (n6587,n6588,n6589);
xor (n6588,n6585,n6586);
or (n6589,n6590,n6592);
and (n6590,n6591,n3065);
xor (n6591,n6503,n6504);
and (n6592,n6593,n6594);
xor (n6593,n6591,n3065);
or (n6594,n6595,n6597);
and (n6595,n6596,n3342);
xor (n6596,n6509,n6510);
and (n6597,n6598,n6599);
xor (n6598,n6596,n3342);
or (n6599,n6600,n6603);
and (n6600,n6601,n6602);
xor (n6601,n6515,n6516);
and (n6602,n1260,n133);
and (n6603,n6604,n6605);
xor (n6604,n6601,n6602);
or (n6605,n6606,n6609);
and (n6606,n6607,n6608);
xor (n6607,n6521,n6522);
and (n6608,n1559,n133);
and (n6609,n6610,n6611);
xor (n6610,n6607,n6608);
and (n6611,n6612,n6613);
xor (n6612,n6527,n6528);
and (n6613,n1835,n133);
and (n6614,n238,n478);
or (n6615,n6616,n6619);
and (n6616,n6617,n6618);
xor (n6617,n6532,n6533);
and (n6618,n152,n478);
and (n6619,n6620,n6621);
xor (n6620,n6617,n6618);
or (n6621,n6622,n6625);
and (n6622,n6623,n6624);
xor (n6623,n6537,n6538);
and (n6624,n134,n478);
and (n6625,n6626,n6627);
xor (n6626,n6623,n6624);
or (n6627,n6628,n6631);
and (n6628,n6629,n6630);
xor (n6629,n6543,n6544);
and (n6630,n473,n478);
and (n6631,n6632,n6633);
xor (n6632,n6629,n6630);
or (n6633,n6634,n6637);
and (n6634,n6635,n6636);
xor (n6635,n6549,n6550);
and (n6636,n368,n478);
and (n6637,n6638,n6639);
xor (n6638,n6635,n6636);
or (n6639,n6640,n6643);
and (n6640,n6641,n6642);
xor (n6641,n6554,n6555);
and (n6642,n96,n478);
and (n6643,n6644,n6645);
xor (n6644,n6641,n6642);
or (n6645,n6646,n6649);
and (n6646,n6647,n6648);
xor (n6647,n6559,n6560);
and (n6648,n77,n478);
and (n6649,n6650,n6651);
xor (n6650,n6647,n6648);
or (n6651,n6652,n6655);
and (n6652,n6653,n6654);
xor (n6653,n6564,n6565);
and (n6654,n565,n478);
and (n6655,n6656,n6657);
xor (n6656,n6653,n6654);
or (n6657,n6658,n6661);
and (n6658,n6659,n6660);
xor (n6659,n6570,n6571);
and (n6660,n303,n478);
and (n6661,n6662,n6663);
xor (n6662,n6659,n6660);
or (n6663,n6664,n6667);
and (n6664,n6665,n6666);
xor (n6665,n6576,n6577);
and (n6666,n286,n478);
and (n6667,n6668,n6669);
xor (n6668,n6665,n6666);
or (n6669,n6670,n6673);
and (n6670,n6671,n6672);
xor (n6671,n6582,n6583);
and (n6672,n615,n478);
and (n6673,n6674,n6675);
xor (n6674,n6671,n6672);
or (n6675,n6676,n6679);
and (n6676,n6677,n6678);
xor (n6677,n6588,n6589);
and (n6678,n660,n478);
and (n6679,n6680,n6681);
xor (n6680,n6677,n6678);
or (n6681,n6682,n6685);
and (n6682,n6683,n6684);
xor (n6683,n6593,n6594);
and (n6684,n653,n478);
and (n6685,n6686,n6687);
xor (n6686,n6683,n6684);
or (n6687,n6688,n6691);
and (n6688,n6689,n6690);
xor (n6689,n6598,n6599);
and (n6690,n1260,n478);
and (n6691,n6692,n6693);
xor (n6692,n6689,n6690);
or (n6693,n6694,n6697);
and (n6694,n6695,n6696);
xor (n6695,n6604,n6605);
and (n6696,n1559,n478);
and (n6697,n6698,n6699);
xor (n6698,n6695,n6696);
and (n6699,n6700,n6701);
xor (n6700,n6610,n6611);
not (n6701,n3565);
or (n6702,n6703,n6705);
and (n6703,n6704,n487);
xor (n6704,n6620,n6621);
and (n6705,n6706,n6707);
xor (n6706,n6704,n487);
or (n6707,n6708,n6710);
and (n6708,n6709,n474);
xor (n6709,n6626,n6627);
and (n6710,n6711,n6712);
xor (n6711,n6709,n474);
or (n6712,n6713,n6715);
and (n6713,n6714,n973);
xor (n6714,n6632,n6633);
and (n6715,n6716,n6717);
xor (n6716,n6714,n973);
or (n6717,n6718,n6721);
and (n6718,n6719,n6720);
xor (n6719,n6638,n6639);
and (n6720,n96,n85);
and (n6721,n6722,n6723);
xor (n6722,n6719,n6720);
or (n6723,n6724,n6727);
and (n6724,n6725,n6726);
xor (n6725,n6644,n6645);
and (n6726,n77,n85);
and (n6727,n6728,n6729);
xor (n6728,n6725,n6726);
or (n6729,n6730,n6733);
and (n6730,n6731,n6732);
xor (n6731,n6650,n6651);
and (n6732,n565,n85);
and (n6733,n6734,n6735);
xor (n6734,n6731,n6732);
or (n6735,n6736,n6739);
and (n6736,n6737,n6738);
xor (n6737,n6656,n6657);
and (n6738,n303,n85);
and (n6739,n6740,n6741);
xor (n6740,n6737,n6738);
or (n6741,n6742,n6745);
and (n6742,n6743,n6744);
xor (n6743,n6662,n6663);
and (n6744,n286,n85);
and (n6745,n6746,n6747);
xor (n6746,n6743,n6744);
or (n6747,n6748,n6750);
and (n6748,n6749,n2315);
xor (n6749,n6668,n6669);
and (n6750,n6751,n6752);
xor (n6751,n6749,n2315);
or (n6752,n6753,n6755);
and (n6753,n6754,n2311);
xor (n6754,n6674,n6675);
and (n6755,n6756,n6757);
xor (n6756,n6754,n2311);
or (n6757,n6758,n6761);
and (n6758,n6759,n6760);
xor (n6759,n6680,n6681);
and (n6760,n653,n85);
and (n6761,n6762,n6763);
xor (n6762,n6759,n6760);
or (n6763,n6764,n6767);
and (n6764,n6765,n6766);
xor (n6765,n6686,n6687);
and (n6766,n1260,n85);
and (n6767,n6768,n6769);
xor (n6768,n6765,n6766);
or (n6769,n6770,n6773);
and (n6770,n6771,n6772);
xor (n6771,n6692,n6693);
and (n6772,n1559,n85);
and (n6773,n6774,n6775);
xor (n6774,n6771,n6772);
and (n6775,n6776,n6777);
xor (n6776,n6698,n6699);
and (n6777,n1835,n85);
and (n6778,n134,n86);
or (n6779,n6780,n6783);
and (n6780,n6781,n6782);
xor (n6781,n6706,n6707);
and (n6782,n473,n86);
and (n6783,n6784,n6785);
xor (n6784,n6781,n6782);
or (n6785,n6786,n6789);
and (n6786,n6787,n6788);
xor (n6787,n6711,n6712);
and (n6788,n368,n86);
and (n6789,n6790,n6791);
xor (n6790,n6787,n6788);
or (n6791,n6792,n6795);
and (n6792,n6793,n6794);
xor (n6793,n6716,n6717);
and (n6794,n96,n86);
and (n6795,n6796,n6797);
xor (n6796,n6793,n6794);
or (n6797,n6798,n6801);
and (n6798,n6799,n6800);
xor (n6799,n6722,n6723);
and (n6800,n77,n86);
and (n6801,n6802,n6803);
xor (n6802,n6799,n6800);
or (n6803,n6804,n6807);
and (n6804,n6805,n6806);
xor (n6805,n6728,n6729);
and (n6806,n565,n86);
and (n6807,n6808,n6809);
xor (n6808,n6805,n6806);
or (n6809,n6810,n6813);
and (n6810,n6811,n6812);
xor (n6811,n6734,n6735);
and (n6812,n303,n86);
and (n6813,n6814,n6815);
xor (n6814,n6811,n6812);
or (n6815,n6816,n6819);
and (n6816,n6817,n6818);
xor (n6817,n6740,n6741);
and (n6818,n286,n86);
and (n6819,n6820,n6821);
xor (n6820,n6817,n6818);
or (n6821,n6822,n6825);
and (n6822,n6823,n6824);
xor (n6823,n6746,n6747);
and (n6824,n615,n86);
and (n6825,n6826,n6827);
xor (n6826,n6823,n6824);
or (n6827,n6828,n6831);
and (n6828,n6829,n6830);
xor (n6829,n6751,n6752);
and (n6830,n660,n86);
and (n6831,n6832,n6833);
xor (n6832,n6829,n6830);
or (n6833,n6834,n6837);
and (n6834,n6835,n6836);
xor (n6835,n6756,n6757);
and (n6836,n653,n86);
and (n6837,n6838,n6839);
xor (n6838,n6835,n6836);
or (n6839,n6840,n6843);
and (n6840,n6841,n6842);
xor (n6841,n6762,n6763);
and (n6842,n1260,n86);
and (n6843,n6844,n6845);
xor (n6844,n6841,n6842);
or (n6845,n6846,n6849);
and (n6846,n6847,n6848);
xor (n6847,n6768,n6769);
and (n6848,n1559,n86);
and (n6849,n6850,n6851);
xor (n6850,n6847,n6848);
and (n6851,n6852,n3108);
xor (n6852,n6774,n6775);
and (n6853,n473,n76);
or (n6854,n6855,n6858);
and (n6855,n6856,n6857);
xor (n6856,n6784,n6785);
and (n6857,n368,n76);
and (n6858,n6859,n6860);
xor (n6859,n6856,n6857);
or (n6860,n6861,n6864);
and (n6861,n6862,n6863);
xor (n6862,n6790,n6791);
and (n6863,n96,n76);
and (n6864,n6865,n6866);
xor (n6865,n6862,n6863);
or (n6866,n6867,n6869);
and (n6867,n6868,n75);
xor (n6868,n6796,n6797);
and (n6869,n6870,n6871);
xor (n6870,n6868,n75);
or (n6871,n6872,n6874);
and (n6872,n6873,n888);
xor (n6873,n6802,n6803);
and (n6874,n6875,n6876);
xor (n6875,n6873,n888);
or (n6876,n6877,n6879);
and (n6877,n6878,n884);
xor (n6878,n6808,n6809);
and (n6879,n6880,n6881);
xor (n6880,n6878,n884);
or (n6881,n6882,n6884);
and (n6882,n6883,n1190);
xor (n6883,n6814,n6815);
and (n6884,n6885,n6886);
xor (n6885,n6883,n1190);
or (n6886,n6887,n6889);
and (n6887,n6888,n1659);
xor (n6888,n6820,n6821);
and (n6889,n6890,n6891);
xor (n6890,n6888,n1659);
or (n6891,n6892,n6895);
and (n6892,n6893,n6894);
xor (n6893,n6826,n6827);
and (n6894,n660,n76);
and (n6895,n6896,n6897);
xor (n6896,n6893,n6894);
or (n6897,n6898,n6900);
and (n6898,n6899,n2223);
xor (n6899,n6832,n6833);
and (n6900,n6901,n6902);
xor (n6901,n6899,n2223);
or (n6902,n6903,n6906);
and (n6903,n6904,n6905);
xor (n6904,n6838,n6839);
and (n6905,n1260,n76);
and (n6906,n6907,n6908);
xor (n6907,n6904,n6905);
or (n6908,n6909,n6912);
and (n6909,n6910,n6911);
xor (n6910,n6844,n6845);
and (n6911,n1559,n76);
and (n6912,n6913,n6914);
xor (n6913,n6910,n6911);
and (n6914,n6915,n6916);
xor (n6915,n6850,n6851);
and (n6916,n1835,n76);
and (n6917,n368,n553);
or (n6918,n6919,n6922);
and (n6919,n6920,n6921);
xor (n6920,n6859,n6860);
and (n6921,n96,n553);
and (n6922,n6923,n6924);
xor (n6923,n6920,n6921);
or (n6924,n6925,n6928);
and (n6925,n6926,n6927);
xor (n6926,n6865,n6866);
and (n6927,n77,n553);
and (n6928,n6929,n6930);
xor (n6929,n6926,n6927);
or (n6930,n6931,n6934);
and (n6931,n6932,n6933);
xor (n6932,n6870,n6871);
and (n6933,n565,n553);
and (n6934,n6935,n6936);
xor (n6935,n6932,n6933);
or (n6936,n6937,n6940);
and (n6937,n6938,n6939);
xor (n6938,n6875,n6876);
and (n6939,n303,n553);
and (n6940,n6941,n6942);
xor (n6941,n6938,n6939);
or (n6942,n6943,n6946);
and (n6943,n6944,n6945);
xor (n6944,n6880,n6881);
and (n6945,n286,n553);
and (n6946,n6947,n6948);
xor (n6947,n6944,n6945);
or (n6948,n6949,n6952);
and (n6949,n6950,n6951);
xor (n6950,n6885,n6886);
and (n6951,n615,n553);
and (n6952,n6953,n6954);
xor (n6953,n6950,n6951);
or (n6954,n6955,n6958);
and (n6955,n6956,n6957);
xor (n6956,n6890,n6891);
and (n6957,n660,n553);
and (n6958,n6959,n6960);
xor (n6959,n6956,n6957);
or (n6960,n6961,n6964);
and (n6961,n6962,n6963);
xor (n6962,n6896,n6897);
and (n6963,n653,n553);
and (n6964,n6965,n6966);
xor (n6965,n6962,n6963);
or (n6966,n6967,n6970);
and (n6967,n6968,n6969);
xor (n6968,n6901,n6902);
and (n6969,n1260,n553);
and (n6970,n6971,n6972);
xor (n6971,n6968,n6969);
or (n6972,n6973,n6976);
and (n6973,n6974,n6975);
xor (n6974,n6907,n6908);
and (n6975,n1559,n553);
and (n6976,n6977,n6978);
xor (n6977,n6974,n6975);
and (n6978,n6979,n6980);
xor (n6979,n6913,n6914);
not (n6980,n2364);
and (n6981,n96,n298);
or (n6982,n6983,n6986);
and (n6983,n6984,n6985);
xor (n6984,n6923,n6924);
and (n6985,n77,n298);
and (n6986,n6987,n6988);
xor (n6987,n6984,n6985);
or (n6988,n6989,n6992);
and (n6989,n6990,n6991);
xor (n6990,n6929,n6930);
and (n6991,n565,n298);
and (n6992,n6993,n6994);
xor (n6993,n6990,n6991);
or (n6994,n6995,n6998);
and (n6995,n6996,n6997);
xor (n6996,n6935,n6936);
and (n6997,n303,n298);
and (n6998,n6999,n7000);
xor (n6999,n6996,n6997);
or (n7000,n7001,n7004);
and (n7001,n7002,n7003);
xor (n7002,n6941,n6942);
and (n7003,n286,n298);
and (n7004,n7005,n7006);
xor (n7005,n7002,n7003);
or (n7006,n7007,n7010);
and (n7007,n7008,n7009);
xor (n7008,n6947,n6948);
and (n7009,n615,n298);
and (n7010,n7011,n7012);
xor (n7011,n7008,n7009);
or (n7012,n7013,n7016);
and (n7013,n7014,n7015);
xor (n7014,n6953,n6954);
and (n7015,n660,n298);
and (n7016,n7017,n7018);
xor (n7017,n7014,n7015);
or (n7018,n7019,n7022);
and (n7019,n7020,n7021);
xor (n7020,n6959,n6960);
and (n7021,n653,n298);
and (n7022,n7023,n7024);
xor (n7023,n7020,n7021);
or (n7024,n7025,n7028);
and (n7025,n7026,n7027);
xor (n7026,n6965,n6966);
and (n7027,n1260,n298);
and (n7028,n7029,n7030);
xor (n7029,n7026,n7027);
or (n7030,n7031,n7033);
and (n7031,n7032,n2155);
xor (n7032,n6971,n6972);
and (n7033,n7034,n7035);
xor (n7034,n7032,n2155);
and (n7035,n7036,n2151);
xor (n7036,n6977,n6978);
and (n7037,n77,n292);
or (n7038,n7039,n7042);
and (n7039,n7040,n7041);
xor (n7040,n6987,n6988);
and (n7041,n565,n292);
and (n7042,n7043,n7044);
xor (n7043,n7040,n7041);
or (n7044,n7045,n7048);
and (n7045,n7046,n7047);
xor (n7046,n6993,n6994);
and (n7047,n303,n292);
and (n7048,n7049,n7050);
xor (n7049,n7046,n7047);
or (n7050,n7051,n7054);
and (n7051,n7052,n7053);
xor (n7052,n6999,n7000);
and (n7053,n286,n292);
and (n7054,n7055,n7056);
xor (n7055,n7052,n7053);
or (n7056,n7057,n7060);
and (n7057,n7058,n7059);
xor (n7058,n7005,n7006);
and (n7059,n615,n292);
and (n7060,n7061,n7062);
xor (n7061,n7058,n7059);
or (n7062,n7063,n7066);
and (n7063,n7064,n7065);
xor (n7064,n7011,n7012);
and (n7065,n660,n292);
and (n7066,n7067,n7068);
xor (n7067,n7064,n7065);
or (n7068,n7069,n7072);
and (n7069,n7070,n7071);
xor (n7070,n7017,n7018);
and (n7071,n653,n292);
and (n7072,n7073,n7074);
xor (n7073,n7070,n7071);
or (n7074,n7075,n7078);
and (n7075,n7076,n7077);
xor (n7076,n7023,n7024);
and (n7077,n1260,n292);
and (n7078,n7079,n7080);
xor (n7079,n7076,n7077);
or (n7080,n7081,n7084);
and (n7081,n7082,n7083);
xor (n7082,n7029,n7030);
and (n7083,n1559,n292);
and (n7084,n7085,n7086);
xor (n7085,n7082,n7083);
and (n7086,n7087,n7088);
xor (n7087,n7034,n7035);
not (n7088,n1834);
or (n7089,n7090,n7093);
and (n7090,n7091,n7092);
xor (n7091,n7043,n7044);
and (n7092,n303,n284);
and (n7093,n7094,n7095);
xor (n7094,n7091,n7092);
or (n7095,n7096,n7098);
and (n7096,n7097,n287);
xor (n7097,n7049,n7050);
and (n7098,n7099,n7100);
xor (n7099,n7097,n287);
or (n7100,n7101,n7103);
and (n7101,n7102,n1034);
xor (n7102,n7055,n7056);
and (n7103,n7104,n7105);
xor (n7104,n7102,n1034);
or (n7105,n7106,n7108);
and (n7106,n7107,n661);
xor (n7107,n7061,n7062);
and (n7108,n7109,n7110);
xor (n7109,n7107,n661);
or (n7110,n7111,n7113);
and (n7111,n7112,n652);
xor (n7112,n7067,n7068);
and (n7113,n7114,n7115);
xor (n7114,n7112,n652);
or (n7115,n7116,n7119);
and (n7116,n7117,n7118);
xor (n7117,n7073,n7074);
and (n7118,n1260,n284);
and (n7119,n7120,n7121);
xor (n7120,n7117,n7118);
or (n7121,n7122,n7124);
and (n7122,n7123,n1560);
xor (n7123,n7079,n7080);
and (n7124,n7125,n7126);
xor (n7125,n7123,n1560);
and (n7126,n7127,n2599);
xor (n7127,n7085,n7086);
or (n7128,n7129,n7131);
and (n7129,n7130,n287);
xor (n7130,n7094,n7095);
and (n7131,n7132,n7133);
xor (n7132,n7130,n287);
or (n7133,n7134,n7136);
and (n7134,n7135,n1034);
xor (n7135,n7099,n7100);
and (n7136,n7137,n7138);
xor (n7137,n7135,n1034);
or (n7138,n7139,n7141);
and (n7139,n7140,n661);
xor (n7140,n7104,n7105);
and (n7141,n7142,n7143);
xor (n7142,n7140,n661);
or (n7143,n7144,n7146);
and (n7144,n7145,n652);
xor (n7145,n7109,n7110);
and (n7146,n7147,n7148);
xor (n7147,n7145,n652);
or (n7148,n7149,n7151);
and (n7149,n7150,n7118);
xor (n7150,n7114,n7115);
and (n7151,n7152,n7153);
xor (n7152,n7150,n7118);
or (n7153,n7154,n7156);
and (n7154,n7155,n1560);
xor (n7155,n7120,n7121);
and (n7156,n7157,n7158);
xor (n7157,n7155,n1560);
and (n7158,n7159,n2599);
xor (n7159,n7125,n7126);
or (n7160,n7161,n7163);
and (n7161,n7162,n1034);
xor (n7162,n7132,n7133);
and (n7163,n7164,n7165);
xor (n7164,n7162,n1034);
or (n7165,n7166,n7168);
and (n7166,n7167,n661);
xor (n7167,n7137,n7138);
and (n7168,n7169,n7170);
xor (n7169,n7167,n661);
or (n7170,n7171,n7173);
and (n7171,n7172,n652);
xor (n7172,n7142,n7143);
and (n7173,n7174,n7175);
xor (n7174,n7172,n652);
or (n7175,n7176,n7178);
and (n7176,n7177,n7118);
xor (n7177,n7147,n7148);
and (n7178,n7179,n7180);
xor (n7179,n7177,n7118);
or (n7180,n7181,n7183);
and (n7181,n7182,n1560);
xor (n7182,n7152,n7153);
and (n7183,n7184,n7185);
xor (n7184,n7182,n1560);
and (n7185,n7186,n2599);
xor (n7186,n7157,n7158);
or (n7187,n7188,n7190);
and (n7188,n7189,n661);
xor (n7189,n7164,n7165);
and (n7190,n7191,n7192);
xor (n7191,n7189,n661);
or (n7192,n7193,n7195);
and (n7193,n7194,n652);
xor (n7194,n7169,n7170);
and (n7195,n7196,n7197);
xor (n7196,n7194,n652);
or (n7197,n7198,n7200);
and (n7198,n7199,n7118);
xor (n7199,n7174,n7175);
and (n7200,n7201,n7202);
xor (n7201,n7199,n7118);
or (n7202,n7203,n7205);
and (n7203,n7204,n1560);
xor (n7204,n7179,n7180);
and (n7205,n7206,n7207);
xor (n7206,n7204,n1560);
and (n7207,n7208,n2599);
xor (n7208,n7184,n7185);
or (n7209,n7210,n7212);
and (n7210,n7211,n652);
xor (n7211,n7191,n7192);
and (n7212,n7213,n7214);
xor (n7213,n7211,n652);
or (n7214,n7215,n7217);
and (n7215,n7216,n7118);
xor (n7216,n7196,n7197);
and (n7217,n7218,n7219);
xor (n7218,n7216,n7118);
or (n7219,n7220,n7222);
and (n7220,n7221,n1560);
xor (n7221,n7201,n7202);
and (n7222,n7223,n7224);
xor (n7223,n7221,n1560);
and (n7224,n7225,n2599);
xor (n7225,n7206,n7207);
or (n7226,n7227,n7229);
and (n7227,n7228,n7118);
xor (n7228,n7213,n7214);
and (n7229,n7230,n7231);
xor (n7230,n7228,n7118);
or (n7231,n7232,n7234);
and (n7232,n7233,n1560);
xor (n7233,n7218,n7219);
and (n7234,n7235,n7236);
xor (n7235,n7233,n1560);
and (n7236,n7237,n2599);
xor (n7237,n7223,n7224);
or (n7238,n7239,n7241);
and (n7239,n7240,n1560);
xor (n7240,n7230,n7231);
and (n7241,n7242,n7243);
xor (n7242,n7240,n1560);
and (n7243,n7244,n2599);
xor (n7244,n7235,n7236);
and (n7245,n7246,n2599);
xor (n7246,n7242,n7243);
or (n7247,n7248,n7251,n7378);
and (n7248,n7249,n7250);
xor (n7249,n5964,n5845);
xor (n7250,n7246,n2599);
and (n7251,n7250,n7252);
or (n7252,n7253,n7256,n7377);
and (n7253,n7254,n7255);
xor (n7254,n5962,n5845);
xor (n7255,n7244,n2599);
and (n7256,n7255,n7257);
or (n7257,n7258,n7261,n7376);
and (n7258,n7259,n7260);
xor (n7259,n5955,n5845);
xor (n7260,n7237,n2599);
and (n7261,n7260,n7262);
or (n7262,n7263,n7266,n7375);
and (n7263,n7264,n7265);
xor (n7264,n5943,n5845);
xor (n7265,n7225,n2599);
and (n7266,n7265,n7267);
or (n7267,n7268,n7271,n7374);
and (n7268,n7269,n7270);
xor (n7269,n5926,n5845);
xor (n7270,n7208,n2599);
and (n7271,n7270,n7272);
or (n7272,n7273,n7276,n7373);
and (n7273,n7274,n7275);
xor (n7274,n5904,n5845);
xor (n7275,n7186,n2599);
and (n7276,n7275,n7277);
or (n7277,n7278,n7281,n7372);
and (n7278,n7279,n7280);
xor (n7279,n5877,n5845);
xor (n7280,n7159,n2599);
and (n7281,n7280,n7282);
or (n7282,n7283,n7286,n7371);
and (n7283,n7284,n7285);
xor (n7284,n5844,n5845);
xor (n7285,n7127,n2599);
and (n7286,n7285,n7287);
or (n7287,n7288,n7291,n7370);
and (n7288,n7289,n7290);
xor (n7289,n5802,n1828);
xor (n7290,n7087,n7088);
and (n7291,n7290,n7292);
or (n7292,n7293,n7296,n7369);
and (n7293,n7294,n7295);
xor (n7294,n5750,n5751);
xor (n7295,n7036,n2151);
and (n7296,n7295,n7297);
or (n7297,n7298,n7301,n7368);
and (n7298,n7299,n7300);
xor (n7299,n5697,n5698);
xor (n7300,n6979,n6980);
and (n7301,n7300,n7302);
or (n7302,n7303,n7306,n7367);
and (n7303,n7304,n7305);
xor (n7304,n5633,n5634);
xor (n7305,n6915,n6916);
and (n7306,n7305,n7307);
or (n7307,n7308,n7311,n7366);
and (n7308,n7309,n7310);
xor (n7309,n5566,n5567);
xor (n7310,n6852,n3108);
and (n7311,n7310,n7312);
or (n7312,n7313,n7316,n7365);
and (n7313,n7314,n7315);
xor (n7314,n5490,n5491);
xor (n7315,n6776,n6777);
and (n7316,n7315,n7317);
or (n7317,n7318,n7321,n7364);
and (n7318,n7319,n7320);
xor (n7319,n5414,n3570);
xor (n7320,n6700,n6701);
and (n7321,n7320,n7322);
or (n7322,n7323,n7326,n7363);
and (n7323,n7324,n7325);
xor (n7324,n5326,n5327);
xor (n7325,n6612,n6613);
and (n7326,n7325,n7327);
or (n7327,n7328,n7331,n7362);
and (n7328,n7329,n7330);
xor (n7329,n5239,n5240);
xor (n7330,n6529,n3842);
and (n7331,n7330,n7332);
or (n7332,n7333,n7336,n7361);
and (n7333,n7334,n7335);
xor (n7334,n5149,n5150);
xor (n7335,n6439,n6440);
and (n7336,n7335,n7337);
or (n7337,n7338,n7341,n7360);
and (n7338,n7339,n7340);
xor (n7339,n5069,n4127);
xor (n7340,n6351,n6352);
and (n7341,n7340,n7342);
or (n7342,n7343,n7346,n7359);
and (n7343,n7344,n7345);
xor (n7344,n4979,n4980);
xor (n7345,n6261,n6262);
and (n7346,n7345,n7347);
or (n7347,n7348,n7351,n7358);
and (n7348,n7349,n7350);
xor (n7349,n4892,n4893);
xor (n7350,n6178,n4388);
and (n7351,n7350,n7352);
or (n7352,n7353,n7356,n7357);
and (n7353,n7354,n7355);
xor (n7354,n4802,n4803);
xor (n7355,n6088,n6089);
and (n7356,n7355,n4542);
and (n7357,n7354,n4542);
and (n7358,n7349,n7352);
and (n7359,n7344,n7347);
and (n7360,n7339,n7342);
and (n7361,n7334,n7337);
and (n7362,n7329,n7332);
and (n7363,n7324,n7327);
and (n7364,n7319,n7322);
and (n7365,n7314,n7317);
and (n7366,n7309,n7312);
and (n7367,n7304,n7307);
and (n7368,n7299,n7302);
and (n7369,n7294,n7297);
and (n7370,n7289,n7292);
and (n7371,n7284,n7287);
and (n7372,n7279,n7282);
and (n7373,n7274,n7277);
and (n7374,n7269,n7272);
and (n7375,n7264,n7267);
and (n7376,n7259,n7262);
and (n7377,n7254,n7257);
and (n7378,n7249,n7252);
xor (n7379,n7380,n2576);
xor (n7380,n7381,n8697);
xor (n7381,n7382,n8575);
xor (n7382,n7383,n8690);
xor (n7383,n7384,n8569);
xor (n7384,n7385,n8678);
xor (n7385,n7386,n8563);
xor (n7386,n7387,n8661);
xor (n7387,n7388,n647);
xor (n7388,n7389,n8639);
xor (n7389,n7390,n966);
xor (n7390,n7391,n8612);
xor (n7391,n7392,n457);
xor (n7392,n7393,n8580);
xor (n7393,n7394,n8542);
xor (n7394,n7395,n8539);
xor (n7395,n7396,n8538);
xor (n7396,n7397,n8488);
xor (n7397,n7398,n8487);
xor (n7398,n7399,n8432);
xor (n7399,n7400,n1407);
xor (n7400,n7401,n8370);
xor (n7401,n7402,n8369);
xor (n7402,n7403,n8304);
xor (n7403,n7404,n1413);
xor (n7404,n7405,n8230);
xor (n7405,n7406,n8229);
xor (n7406,n7407,n8154);
xor (n7407,n7408,n1491);
xor (n7408,n7409,n8068);
xor (n7409,n7410,n8067);
xor (n7410,n7411,n7980);
xor (n7411,n7412,n7979);
or (n7412,n7413,n7885);
and (n7413,n7414,n7884);
or (n7414,n7415,n7793);
and (n7415,n7416,n7792);
or (n7416,n7417,n7697);
and (n7417,n7418,n7696);
or (n7418,n7419,n7606);
and (n7419,n7420,n745);
or (n7420,n7421,n7511);
and (n7421,n7422,n7510);
and (n7422,n1270,n7423);
or (n7423,n7424,n7426);
and (n7424,n7425,n1551);
and (n7425,n270,n1266);
and (n7426,n7427,n7428);
xor (n7427,n7425,n1551);
or (n7428,n7429,n7431);
and (n7429,n7430,n2448);
and (n7430,n432,n1266);
and (n7431,n7432,n7433);
xor (n7432,n7430,n2448);
or (n7433,n7434,n7437);
and (n7434,n7435,n7436);
and (n7435,n417,n1266);
and (n7436,n583,n667);
and (n7437,n7438,n7439);
xor (n7438,n7435,n7436);
or (n7439,n7440,n7442);
and (n7440,n7441,n2239);
and (n7441,n583,n1266);
and (n7442,n7443,n7444);
xor (n7443,n7441,n2239);
or (n7444,n7445,n7448);
and (n7445,n7446,n7447);
and (n7446,n195,n1266);
and (n7447,n206,n667);
and (n7448,n7449,n7450);
xor (n7449,n7446,n7447);
or (n7450,n7451,n7454);
and (n7451,n7452,n7453);
and (n7452,n206,n1266);
and (n7453,n126,n667);
and (n7454,n7455,n7456);
xor (n7455,n7452,n7453);
or (n7456,n7457,n7459);
and (n7457,n7458,n3307);
and (n7458,n126,n1266);
and (n7459,n7460,n7461);
xor (n7460,n7458,n3307);
or (n7461,n7462,n7465);
and (n7462,n7463,n7464);
and (n7463,n106,n1266);
and (n7464,n496,n667);
and (n7465,n7466,n7467);
xor (n7466,n7463,n7464);
or (n7467,n7468,n7471);
and (n7468,n7469,n7470);
and (n7469,n496,n1266);
and (n7470,n461,n667);
and (n7471,n7472,n7473);
xor (n7472,n7469,n7470);
or (n7473,n7474,n7477);
and (n7474,n7475,n7476);
and (n7475,n461,n1266);
and (n7476,n456,n667);
and (n7477,n7478,n7479);
xor (n7478,n7475,n7476);
or (n7479,n7480,n7483);
and (n7480,n7481,n7482);
and (n7481,n456,n1266);
and (n7482,n761,n667);
and (n7483,n7484,n7485);
xor (n7484,n7481,n7482);
or (n7485,n7486,n7488);
and (n7486,n7487,n4152);
and (n7487,n761,n1266);
and (n7488,n7489,n7490);
xor (n7489,n7487,n4152);
or (n7490,n7491,n7493);
and (n7491,n7492,n4309);
and (n7492,n646,n1266);
and (n7493,n7494,n7495);
xor (n7494,n7492,n4309);
or (n7495,n7496,n7499);
and (n7496,n7497,n7498);
and (n7497,n640,n1266);
and (n7498,n1317,n667);
and (n7499,n7500,n7501);
xor (n7500,n7497,n7498);
or (n7501,n7502,n7505);
and (n7502,n7503,n7504);
and (n7503,n1317,n1266);
and (n7504,n1780,n667);
and (n7505,n7506,n7507);
xor (n7506,n7503,n7504);
and (n7507,n7508,n7509);
and (n7508,n1780,n1266);
and (n7509,n1822,n667);
and (n7510,n270,n735);
and (n7511,n7512,n7513);
xor (n7512,n7422,n7510);
or (n7513,n7514,n7517);
and (n7514,n7515,n7516);
xor (n7515,n1270,n7423);
and (n7516,n432,n735);
and (n7517,n7518,n7519);
xor (n7518,n7515,n7516);
or (n7519,n7520,n7523);
and (n7520,n7521,n7522);
xor (n7521,n7427,n7428);
and (n7522,n417,n735);
and (n7523,n7524,n7525);
xor (n7524,n7521,n7522);
or (n7525,n7526,n7529);
and (n7526,n7527,n7528);
xor (n7527,n7432,n7433);
and (n7528,n583,n735);
and (n7529,n7530,n7531);
xor (n7530,n7527,n7528);
or (n7531,n7532,n7535);
and (n7532,n7533,n7534);
xor (n7533,n7438,n7439);
and (n7534,n195,n735);
and (n7535,n7536,n7537);
xor (n7536,n7533,n7534);
or (n7537,n7538,n7541);
and (n7538,n7539,n7540);
xor (n7539,n7443,n7444);
and (n7540,n206,n735);
and (n7541,n7542,n7543);
xor (n7542,n7539,n7540);
or (n7543,n7544,n7547);
and (n7544,n7545,n7546);
xor (n7545,n7449,n7450);
and (n7546,n126,n735);
and (n7547,n7548,n7549);
xor (n7548,n7545,n7546);
or (n7549,n7550,n7553);
and (n7550,n7551,n7552);
xor (n7551,n7455,n7456);
and (n7552,n106,n735);
and (n7553,n7554,n7555);
xor (n7554,n7551,n7552);
or (n7555,n7556,n7559);
and (n7556,n7557,n7558);
xor (n7557,n7460,n7461);
and (n7558,n496,n735);
and (n7559,n7560,n7561);
xor (n7560,n7557,n7558);
or (n7561,n7562,n7565);
and (n7562,n7563,n7564);
xor (n7563,n7466,n7467);
and (n7564,n461,n735);
and (n7565,n7566,n7567);
xor (n7566,n7563,n7564);
or (n7567,n7568,n7571);
and (n7568,n7569,n7570);
xor (n7569,n7472,n7473);
and (n7570,n456,n735);
and (n7571,n7572,n7573);
xor (n7572,n7569,n7570);
or (n7573,n7574,n7577);
and (n7574,n7575,n7576);
xor (n7575,n7478,n7479);
and (n7576,n761,n735);
and (n7577,n7578,n7579);
xor (n7578,n7575,n7576);
or (n7579,n7580,n7583);
and (n7580,n7581,n7582);
xor (n7581,n7484,n7485);
and (n7582,n646,n735);
and (n7583,n7584,n7585);
xor (n7584,n7581,n7582);
or (n7585,n7586,n7589);
and (n7586,n7587,n7588);
xor (n7587,n7489,n7490);
and (n7588,n640,n735);
and (n7589,n7590,n7591);
xor (n7590,n7587,n7588);
or (n7591,n7592,n7595);
and (n7592,n7593,n7594);
xor (n7593,n7494,n7495);
and (n7594,n1317,n735);
and (n7595,n7596,n7597);
xor (n7596,n7593,n7594);
or (n7597,n7598,n7601);
and (n7598,n7599,n7600);
xor (n7599,n7500,n7501);
and (n7600,n1780,n735);
and (n7601,n7602,n7603);
xor (n7602,n7599,n7600);
and (n7603,n7604,n7605);
xor (n7604,n7506,n7507);
not (n7605,n4382);
and (n7606,n7607,n7608);
xor (n7607,n7420,n745);
or (n7608,n7609,n7612);
and (n7609,n7610,n7611);
xor (n7610,n7512,n7513);
and (n7611,n432,n266);
and (n7612,n7613,n7614);
xor (n7613,n7610,n7611);
or (n7614,n7615,n7618);
and (n7615,n7616,n7617);
xor (n7616,n7518,n7519);
and (n7617,n417,n266);
and (n7618,n7619,n7620);
xor (n7619,n7616,n7617);
or (n7620,n7621,n7624);
and (n7621,n7622,n7623);
xor (n7622,n7524,n7525);
and (n7623,n583,n266);
and (n7624,n7625,n7626);
xor (n7625,n7622,n7623);
or (n7626,n7627,n7630);
and (n7627,n7628,n7629);
xor (n7628,n7530,n7531);
and (n7629,n195,n266);
and (n7630,n7631,n7632);
xor (n7631,n7628,n7629);
or (n7632,n7633,n7635);
and (n7633,n7634,n2165);
xor (n7634,n7536,n7537);
and (n7635,n7636,n7637);
xor (n7636,n7634,n2165);
or (n7637,n7638,n7640);
and (n7638,n7639,n2161);
xor (n7639,n7542,n7543);
and (n7640,n7641,n7642);
xor (n7641,n7639,n2161);
or (n7642,n7643,n7646);
and (n7643,n7644,n7645);
xor (n7644,n7548,n7549);
and (n7645,n106,n266);
and (n7646,n7647,n7648);
xor (n7647,n7644,n7645);
or (n7648,n7649,n7651);
and (n7649,n7650,n3216);
xor (n7650,n7554,n7555);
and (n7651,n7652,n7653);
xor (n7652,n7650,n3216);
or (n7653,n7654,n7657);
and (n7654,n7655,n7656);
xor (n7655,n7560,n7561);
and (n7656,n461,n266);
and (n7657,n7658,n7659);
xor (n7658,n7655,n7656);
or (n7659,n7660,n7663);
and (n7660,n7661,n7662);
xor (n7661,n7566,n7567);
and (n7662,n456,n266);
and (n7663,n7664,n7665);
xor (n7664,n7661,n7662);
or (n7665,n7666,n7668);
and (n7666,n7667,n3789);
xor (n7667,n7572,n7573);
and (n7668,n7669,n7670);
xor (n7669,n7667,n3789);
or (n7670,n7671,n7673);
and (n7671,n7672,n3939);
xor (n7672,n7578,n7579);
and (n7673,n7674,n7675);
xor (n7674,n7672,n3939);
or (n7675,n7676,n7679);
and (n7676,n7677,n7678);
xor (n7677,n7584,n7585);
and (n7678,n640,n266);
and (n7679,n7680,n7681);
xor (n7680,n7677,n7678);
or (n7681,n7682,n7685);
and (n7682,n7683,n7684);
xor (n7683,n7590,n7591);
and (n7684,n1317,n266);
and (n7685,n7686,n7687);
xor (n7686,n7683,n7684);
or (n7687,n7688,n7691);
and (n7688,n7689,n7690);
xor (n7689,n7596,n7597);
and (n7690,n1780,n266);
and (n7691,n7692,n7693);
xor (n7692,n7689,n7690);
and (n7693,n7694,n7695);
xor (n7694,n7602,n7603);
and (n7695,n1822,n266);
and (n7696,n270,n265);
and (n7697,n7698,n7699);
xor (n7698,n7418,n7696);
or (n7699,n7700,n7703);
and (n7700,n7701,n7702);
xor (n7701,n7607,n7608);
and (n7702,n432,n265);
and (n7703,n7704,n7705);
xor (n7704,n7701,n7702);
or (n7705,n7706,n7709);
and (n7706,n7707,n7708);
xor (n7707,n7613,n7614);
and (n7708,n417,n265);
and (n7709,n7710,n7711);
xor (n7710,n7707,n7708);
or (n7711,n7712,n7715);
and (n7712,n7713,n7714);
xor (n7713,n7619,n7620);
and (n7714,n583,n265);
and (n7715,n7716,n7717);
xor (n7716,n7713,n7714);
or (n7717,n7718,n7721);
and (n7718,n7719,n7720);
xor (n7719,n7625,n7626);
and (n7720,n195,n265);
and (n7721,n7722,n7723);
xor (n7722,n7719,n7720);
or (n7723,n7724,n7727);
and (n7724,n7725,n7726);
xor (n7725,n7631,n7632);
and (n7726,n206,n265);
and (n7727,n7728,n7729);
xor (n7728,n7725,n7726);
or (n7729,n7730,n7733);
and (n7730,n7731,n7732);
xor (n7731,n7636,n7637);
and (n7732,n126,n265);
and (n7733,n7734,n7735);
xor (n7734,n7731,n7732);
or (n7735,n7736,n7739);
and (n7736,n7737,n7738);
xor (n7737,n7641,n7642);
and (n7738,n106,n265);
and (n7739,n7740,n7741);
xor (n7740,n7737,n7738);
or (n7741,n7742,n7745);
and (n7742,n7743,n7744);
xor (n7743,n7647,n7648);
and (n7744,n496,n265);
and (n7745,n7746,n7747);
xor (n7746,n7743,n7744);
or (n7747,n7748,n7751);
and (n7748,n7749,n7750);
xor (n7749,n7652,n7653);
and (n7750,n461,n265);
and (n7751,n7752,n7753);
xor (n7752,n7749,n7750);
or (n7753,n7754,n7757);
and (n7754,n7755,n7756);
xor (n7755,n7658,n7659);
and (n7756,n456,n265);
and (n7757,n7758,n7759);
xor (n7758,n7755,n7756);
or (n7759,n7760,n7763);
and (n7760,n7761,n7762);
xor (n7761,n7664,n7665);
and (n7762,n761,n265);
and (n7763,n7764,n7765);
xor (n7764,n7761,n7762);
or (n7765,n7766,n7769);
and (n7766,n7767,n7768);
xor (n7767,n7669,n7670);
and (n7768,n646,n265);
and (n7769,n7770,n7771);
xor (n7770,n7767,n7768);
or (n7771,n7772,n7775);
and (n7772,n7773,n7774);
xor (n7773,n7674,n7675);
and (n7774,n640,n265);
and (n7775,n7776,n7777);
xor (n7776,n7773,n7774);
or (n7777,n7778,n7781);
and (n7778,n7779,n7780);
xor (n7779,n7680,n7681);
and (n7780,n1317,n265);
and (n7781,n7782,n7783);
xor (n7782,n7779,n7780);
or (n7783,n7784,n7787);
and (n7784,n7785,n7786);
xor (n7785,n7686,n7687);
and (n7786,n1780,n265);
and (n7787,n7788,n7789);
xor (n7788,n7785,n7786);
and (n7789,n7790,n7791);
xor (n7790,n7692,n7693);
not (n7791,n4121);
and (n7792,n270,n272);
and (n7793,n7794,n7795);
xor (n7794,n7416,n7792);
or (n7795,n7796,n7799);
and (n7796,n7797,n7798);
xor (n7797,n7698,n7699);
and (n7798,n432,n272);
and (n7799,n7800,n7801);
xor (n7800,n7797,n7798);
or (n7801,n7802,n7805);
and (n7802,n7803,n7804);
xor (n7803,n7704,n7705);
and (n7804,n417,n272);
and (n7805,n7806,n7807);
xor (n7806,n7803,n7804);
or (n7807,n7808,n7811);
and (n7808,n7809,n7810);
xor (n7809,n7710,n7711);
and (n7810,n583,n272);
and (n7811,n7812,n7813);
xor (n7812,n7809,n7810);
or (n7813,n7814,n7817);
and (n7814,n7815,n7816);
xor (n7815,n7716,n7717);
and (n7816,n195,n272);
and (n7817,n7818,n7819);
xor (n7818,n7815,n7816);
or (n7819,n7820,n7823);
and (n7820,n7821,n7822);
xor (n7821,n7722,n7723);
and (n7822,n206,n272);
and (n7823,n7824,n7825);
xor (n7824,n7821,n7822);
or (n7825,n7826,n7828);
and (n7826,n7827,n2496);
xor (n7827,n7728,n7729);
and (n7828,n7829,n7830);
xor (n7829,n7827,n2496);
or (n7830,n7831,n7834);
and (n7831,n7832,n7833);
xor (n7832,n7734,n7735);
and (n7833,n106,n272);
and (n7834,n7835,n7836);
xor (n7835,n7832,n7833);
or (n7836,n7837,n7839);
and (n7837,n7838,n2276);
xor (n7838,n7740,n7741);
and (n7839,n7840,n7841);
xor (n7840,n7838,n2276);
or (n7841,n7842,n7844);
and (n7842,n7843,n2864);
xor (n7843,n7746,n7747);
and (n7844,n7845,n7846);
xor (n7845,n7843,n2864);
or (n7846,n7847,n7850);
and (n7847,n7848,n7849);
xor (n7848,n7752,n7753);
and (n7849,n456,n272);
and (n7850,n7851,n7852);
xor (n7851,n7848,n7849);
or (n7852,n7853,n7856);
and (n7853,n7854,n7855);
xor (n7854,n7758,n7759);
and (n7855,n761,n272);
and (n7856,n7857,n7858);
xor (n7857,n7854,n7855);
or (n7858,n7859,n7862);
and (n7859,n7860,n7861);
xor (n7860,n7764,n7765);
and (n7861,n646,n272);
and (n7862,n7863,n7864);
xor (n7863,n7860,n7861);
or (n7864,n7865,n7867);
and (n7865,n7866,n3708);
xor (n7866,n7770,n7771);
and (n7867,n7868,n7869);
xor (n7868,n7866,n3708);
or (n7869,n7870,n7873);
and (n7870,n7871,n7872);
xor (n7871,n7776,n7777);
and (n7872,n1317,n272);
and (n7873,n7874,n7875);
xor (n7874,n7871,n7872);
or (n7875,n7876,n7879);
and (n7876,n7877,n7878);
xor (n7877,n7782,n7783);
and (n7878,n1780,n272);
and (n7879,n7880,n7881);
xor (n7880,n7877,n7878);
and (n7881,n7882,n7883);
xor (n7882,n7788,n7789);
and (n7883,n1822,n272);
and (n7884,n270,n423);
and (n7885,n7886,n7887);
xor (n7886,n7414,n7884);
or (n7887,n7888,n7891);
and (n7888,n7889,n7890);
xor (n7889,n7794,n7795);
and (n7890,n432,n423);
and (n7891,n7892,n7893);
xor (n7892,n7889,n7890);
or (n7893,n7894,n7897);
and (n7894,n7895,n7896);
xor (n7895,n7800,n7801);
and (n7896,n417,n423);
and (n7897,n7898,n7899);
xor (n7898,n7895,n7896);
or (n7899,n7900,n7903);
and (n7900,n7901,n7902);
xor (n7901,n7806,n7807);
and (n7902,n583,n423);
and (n7903,n7904,n7905);
xor (n7904,n7901,n7902);
or (n7905,n7906,n7909);
and (n7906,n7907,n7908);
xor (n7907,n7812,n7813);
and (n7908,n195,n423);
and (n7909,n7910,n7911);
xor (n7910,n7907,n7908);
or (n7911,n7912,n7915);
and (n7912,n7913,n7914);
xor (n7913,n7818,n7819);
and (n7914,n206,n423);
and (n7915,n7916,n7917);
xor (n7916,n7913,n7914);
or (n7917,n7918,n7921);
and (n7918,n7919,n7920);
xor (n7919,n7824,n7825);
and (n7920,n126,n423);
and (n7921,n7922,n7923);
xor (n7922,n7919,n7920);
or (n7923,n7924,n7927);
and (n7924,n7925,n7926);
xor (n7925,n7829,n7830);
and (n7926,n106,n423);
and (n7927,n7928,n7929);
xor (n7928,n7925,n7926);
or (n7929,n7930,n7933);
and (n7930,n7931,n7932);
xor (n7931,n7835,n7836);
and (n7932,n496,n423);
and (n7933,n7934,n7935);
xor (n7934,n7931,n7932);
or (n7935,n7936,n7939);
and (n7936,n7937,n7938);
xor (n7937,n7840,n7841);
and (n7938,n461,n423);
and (n7939,n7940,n7941);
xor (n7940,n7937,n7938);
or (n7941,n7942,n7945);
and (n7942,n7943,n7944);
xor (n7943,n7845,n7846);
and (n7944,n456,n423);
and (n7945,n7946,n7947);
xor (n7946,n7943,n7944);
or (n7947,n7948,n7951);
and (n7948,n7949,n7950);
xor (n7949,n7851,n7852);
and (n7950,n761,n423);
and (n7951,n7952,n7953);
xor (n7952,n7949,n7950);
or (n7953,n7954,n7957);
and (n7954,n7955,n7956);
xor (n7955,n7857,n7858);
and (n7956,n646,n423);
and (n7957,n7958,n7959);
xor (n7958,n7955,n7956);
or (n7959,n7960,n7963);
and (n7960,n7961,n7962);
xor (n7961,n7863,n7864);
and (n7962,n640,n423);
and (n7963,n7964,n7965);
xor (n7964,n7961,n7962);
or (n7965,n7966,n7969);
and (n7966,n7967,n7968);
xor (n7967,n7868,n7869);
and (n7968,n1317,n423);
and (n7969,n7970,n7971);
xor (n7970,n7967,n7968);
or (n7971,n7972,n7975);
and (n7972,n7973,n7974);
xor (n7973,n7874,n7875);
and (n7974,n1780,n423);
and (n7975,n7976,n7977);
xor (n7976,n7973,n7974);
and (n7977,n7978,n3831);
xor (n7978,n7880,n7881);
and (n7979,n270,n188);
or (n7980,n7981,n7984);
and (n7981,n7982,n7983);
xor (n7982,n7886,n7887);
and (n7983,n432,n188);
and (n7984,n7985,n7986);
xor (n7985,n7982,n7983);
or (n7986,n7987,n7989);
and (n7987,n7988,n418);
xor (n7988,n7892,n7893);
and (n7989,n7990,n7991);
xor (n7990,n7988,n418);
or (n7991,n7992,n7994);
and (n7992,n7993,n584);
xor (n7993,n7898,n7899);
and (n7994,n7995,n7996);
xor (n7995,n7993,n584);
or (n7996,n7997,n7999);
and (n7997,n7998,n917);
xor (n7998,n7904,n7905);
and (n7999,n8000,n8001);
xor (n8000,n7998,n917);
or (n8001,n8002,n8005);
and (n8002,n8003,n8004);
xor (n8003,n7910,n7911);
and (n8004,n206,n188);
and (n8005,n8006,n8007);
xor (n8006,n8003,n8004);
or (n8007,n8008,n8011);
and (n8008,n8009,n8010);
xor (n8009,n7916,n7917);
and (n8010,n126,n188);
and (n8011,n8012,n8013);
xor (n8012,n8009,n8010);
or (n8013,n8014,n8017);
and (n8014,n8015,n8016);
xor (n8015,n7922,n7923);
and (n8016,n106,n188);
and (n8017,n8018,n8019);
xor (n8018,n8015,n8016);
or (n8019,n8020,n8023);
and (n8020,n8021,n8022);
xor (n8021,n7928,n7929);
and (n8022,n496,n188);
and (n8023,n8024,n8025);
xor (n8024,n8021,n8022);
or (n8025,n8026,n8028);
and (n8026,n8027,n2261);
xor (n8027,n7934,n7935);
and (n8028,n8029,n8030);
xor (n8029,n8027,n2261);
or (n8030,n8031,n8033);
and (n8031,n8032,n2257);
xor (n8032,n7940,n7941);
and (n8033,n8034,n8035);
xor (n8034,n8032,n2257);
or (n8035,n8036,n8039);
and (n8036,n8037,n8038);
xor (n8037,n7946,n7947);
and (n8038,n761,n188);
and (n8039,n8040,n8041);
xor (n8040,n8037,n8038);
or (n8041,n8042,n8045);
and (n8042,n8043,n8044);
xor (n8043,n7952,n7953);
and (n8044,n646,n188);
and (n8045,n8046,n8047);
xor (n8046,n8043,n8044);
or (n8047,n8048,n8050);
and (n8048,n8049,n3373);
xor (n8049,n7958,n7959);
and (n8050,n8051,n8052);
xor (n8051,n8049,n3373);
or (n8052,n8053,n8056);
and (n8053,n8054,n8055);
xor (n8054,n7964,n7965);
and (n8055,n1317,n188);
and (n8056,n8057,n8058);
xor (n8057,n8054,n8055);
or (n8058,n8059,n8062);
and (n8059,n8060,n8061);
xor (n8060,n7970,n7971);
and (n8061,n1780,n188);
and (n8062,n8063,n8064);
xor (n8063,n8060,n8061);
and (n8064,n8065,n8066);
xor (n8065,n7976,n7977);
and (n8066,n1822,n188);
and (n8067,n432,n189);
or (n8068,n8069,n8072);
and (n8069,n8070,n8071);
xor (n8070,n7985,n7986);
and (n8071,n417,n189);
and (n8072,n8073,n8074);
xor (n8073,n8070,n8071);
or (n8074,n8075,n8078);
and (n8075,n8076,n8077);
xor (n8076,n7990,n7991);
and (n8077,n583,n189);
and (n8078,n8079,n8080);
xor (n8079,n8076,n8077);
or (n8080,n8081,n8084);
and (n8081,n8082,n8083);
xor (n8082,n7995,n7996);
and (n8083,n195,n189);
and (n8084,n8085,n8086);
xor (n8085,n8082,n8083);
or (n8086,n8087,n8090);
and (n8087,n8088,n8089);
xor (n8088,n8000,n8001);
and (n8089,n206,n189);
and (n8090,n8091,n8092);
xor (n8091,n8088,n8089);
or (n8092,n8093,n8096);
and (n8093,n8094,n8095);
xor (n8094,n8006,n8007);
and (n8095,n126,n189);
and (n8096,n8097,n8098);
xor (n8097,n8094,n8095);
or (n8098,n8099,n8102);
and (n8099,n8100,n8101);
xor (n8100,n8012,n8013);
and (n8101,n106,n189);
and (n8102,n8103,n8104);
xor (n8103,n8100,n8101);
or (n8104,n8105,n8108);
and (n8105,n8106,n8107);
xor (n8106,n8018,n8019);
and (n8107,n496,n189);
and (n8108,n8109,n8110);
xor (n8109,n8106,n8107);
or (n8110,n8111,n8114);
and (n8111,n8112,n8113);
xor (n8112,n8024,n8025);
and (n8113,n461,n189);
and (n8114,n8115,n8116);
xor (n8115,n8112,n8113);
or (n8116,n8117,n8120);
and (n8117,n8118,n8119);
xor (n8118,n8029,n8030);
and (n8119,n456,n189);
and (n8120,n8121,n8122);
xor (n8121,n8118,n8119);
or (n8122,n8123,n8126);
and (n8123,n8124,n8125);
xor (n8124,n8034,n8035);
and (n8125,n761,n189);
and (n8126,n8127,n8128);
xor (n8127,n8124,n8125);
or (n8128,n8129,n8132);
and (n8129,n8130,n8131);
xor (n8130,n8040,n8041);
and (n8131,n646,n189);
and (n8132,n8133,n8134);
xor (n8133,n8130,n8131);
or (n8134,n8135,n8138);
and (n8135,n8136,n8137);
xor (n8136,n8046,n8047);
and (n8137,n640,n189);
and (n8138,n8139,n8140);
xor (n8139,n8136,n8137);
or (n8140,n8141,n8144);
and (n8141,n8142,n8143);
xor (n8142,n8051,n8052);
and (n8143,n1317,n189);
and (n8144,n8145,n8146);
xor (n8145,n8142,n8143);
or (n8146,n8147,n8150);
and (n8147,n8148,n8149);
xor (n8148,n8057,n8058);
and (n8149,n1780,n189);
and (n8150,n8151,n8152);
xor (n8151,n8148,n8149);
and (n8152,n8153,n3558);
xor (n8153,n8063,n8064);
or (n8154,n8155,n8157);
and (n8155,n8156,n1003);
xor (n8156,n8073,n8074);
and (n8157,n8158,n8159);
xor (n8158,n8156,n1003);
or (n8159,n8160,n8162);
and (n8160,n8161,n196);
xor (n8161,n8079,n8080);
and (n8162,n8163,n8164);
xor (n8163,n8161,n196);
or (n8164,n8165,n8168);
and (n8165,n8166,n8167);
xor (n8166,n8085,n8086);
and (n8167,n206,n120);
and (n8168,n8169,n8170);
xor (n8169,n8166,n8167);
or (n8170,n8171,n8174);
and (n8171,n8172,n8173);
xor (n8172,n8091,n8092);
and (n8173,n126,n120);
and (n8174,n8175,n8176);
xor (n8175,n8172,n8173);
or (n8176,n8177,n8180);
and (n8177,n8178,n8179);
xor (n8178,n8097,n8098);
and (n8179,n106,n120);
and (n8180,n8181,n8182);
xor (n8181,n8178,n8179);
or (n8182,n8183,n8186);
and (n8183,n8184,n8185);
xor (n8184,n8103,n8104);
and (n8185,n496,n120);
and (n8186,n8187,n8188);
xor (n8187,n8184,n8185);
or (n8188,n8189,n8191);
and (n8189,n8190,n1724);
xor (n8190,n8109,n8110);
and (n8191,n8192,n8193);
xor (n8192,n8190,n1724);
or (n8193,n8194,n8197);
and (n8194,n8195,n8196);
xor (n8195,n8115,n8116);
and (n8196,n456,n120);
and (n8197,n8198,n8199);
xor (n8198,n8195,n8196);
or (n8199,n8200,n8202);
and (n8200,n8201,n2114);
xor (n8201,n8121,n8122);
and (n8202,n8203,n8204);
xor (n8203,n8201,n2114);
or (n8204,n8205,n8208);
and (n8205,n8206,n8207);
xor (n8206,n8127,n8128);
and (n8207,n646,n120);
and (n8208,n8209,n8210);
xor (n8209,n8206,n8207);
or (n8210,n8211,n8214);
and (n8211,n8212,n8213);
xor (n8212,n8133,n8134);
and (n8213,n640,n120);
and (n8214,n8215,n8216);
xor (n8215,n8212,n8213);
or (n8216,n8217,n8219);
and (n8217,n8218,n3223);
xor (n8218,n8139,n8140);
and (n8219,n8220,n8221);
xor (n8220,n8218,n3223);
or (n8221,n8222,n8224);
and (n8222,n8223,n3320);
xor (n8223,n8145,n8146);
and (n8224,n8225,n8226);
xor (n8225,n8223,n3320);
and (n8226,n8227,n8228);
xor (n8227,n8151,n8152);
and (n8228,n1822,n120);
and (n8229,n583,n115);
or (n8230,n8231,n8234);
and (n8231,n8232,n8233);
xor (n8232,n8158,n8159);
and (n8233,n195,n115);
and (n8234,n8235,n8236);
xor (n8235,n8232,n8233);
or (n8236,n8237,n8240);
and (n8237,n8238,n8239);
xor (n8238,n8163,n8164);
and (n8239,n206,n115);
and (n8240,n8241,n8242);
xor (n8241,n8238,n8239);
or (n8242,n8243,n8246);
and (n8243,n8244,n8245);
xor (n8244,n8169,n8170);
and (n8245,n126,n115);
and (n8246,n8247,n8248);
xor (n8247,n8244,n8245);
or (n8248,n8249,n8252);
and (n8249,n8250,n8251);
xor (n8250,n8175,n8176);
and (n8251,n106,n115);
and (n8252,n8253,n8254);
xor (n8253,n8250,n8251);
or (n8254,n8255,n8258);
and (n8255,n8256,n8257);
xor (n8256,n8181,n8182);
and (n8257,n496,n115);
and (n8258,n8259,n8260);
xor (n8259,n8256,n8257);
or (n8260,n8261,n8264);
and (n8261,n8262,n8263);
xor (n8262,n8187,n8188);
and (n8263,n461,n115);
and (n8264,n8265,n8266);
xor (n8265,n8262,n8263);
or (n8266,n8267,n8270);
and (n8267,n8268,n8269);
xor (n8268,n8192,n8193);
and (n8269,n456,n115);
and (n8270,n8271,n8272);
xor (n8271,n8268,n8269);
or (n8272,n8273,n8276);
and (n8273,n8274,n8275);
xor (n8274,n8198,n8199);
and (n8275,n761,n115);
and (n8276,n8277,n8278);
xor (n8277,n8274,n8275);
or (n8278,n8279,n8282);
and (n8279,n8280,n8281);
xor (n8280,n8203,n8204);
and (n8281,n646,n115);
and (n8282,n8283,n8284);
xor (n8283,n8280,n8281);
or (n8284,n8285,n8288);
and (n8285,n8286,n8287);
xor (n8286,n8209,n8210);
and (n8287,n640,n115);
and (n8288,n8289,n8290);
xor (n8289,n8286,n8287);
or (n8290,n8291,n8294);
and (n8291,n8292,n8293);
xor (n8292,n8215,n8216);
and (n8293,n1317,n115);
and (n8294,n8295,n8296);
xor (n8295,n8292,n8293);
or (n8296,n8297,n8300);
and (n8297,n8298,n8299);
xor (n8298,n8220,n8221);
and (n8299,n1780,n115);
and (n8300,n8301,n8302);
xor (n8301,n8298,n8299);
and (n8302,n8303,n3101);
xor (n8303,n8225,n8226);
or (n8304,n8305,n8307);
and (n8305,n8306,n522);
xor (n8306,n8235,n8236);
and (n8307,n8308,n8309);
xor (n8308,n8306,n522);
or (n8309,n8310,n8312);
and (n8310,n8311,n127);
xor (n8311,n8241,n8242);
and (n8312,n8313,n8314);
xor (n8313,n8311,n127);
or (n8314,n8315,n8318);
and (n8315,n8316,n8317);
xor (n8316,n8247,n8248);
and (n8317,n106,n108);
and (n8318,n8319,n8320);
xor (n8319,n8316,n8317);
or (n8320,n8321,n8324);
and (n8321,n8322,n8323);
xor (n8322,n8253,n8254);
and (n8323,n496,n108);
and (n8324,n8325,n8326);
xor (n8325,n8322,n8323);
or (n8326,n8327,n8330);
and (n8327,n8328,n8329);
xor (n8328,n8259,n8260);
and (n8329,n461,n108);
and (n8330,n8331,n8332);
xor (n8331,n8328,n8329);
or (n8332,n8333,n8336);
and (n8333,n8334,n8335);
xor (n8334,n8265,n8266);
and (n8335,n456,n108);
and (n8336,n8337,n8338);
xor (n8337,n8334,n8335);
or (n8338,n8339,n8342);
and (n8339,n8340,n8341);
xor (n8340,n8271,n8272);
and (n8341,n761,n108);
and (n8342,n8343,n8344);
xor (n8343,n8340,n8341);
or (n8344,n8345,n8348);
and (n8345,n8346,n8347);
xor (n8346,n8277,n8278);
and (n8347,n646,n108);
and (n8348,n8349,n8350);
xor (n8349,n8346,n8347);
or (n8350,n8351,n8353);
and (n8351,n8352,n2199);
xor (n8352,n8283,n8284);
and (n8353,n8354,n8355);
xor (n8354,n8352,n2199);
or (n8355,n8356,n8358);
and (n8356,n8357,n2195);
xor (n8357,n8289,n8290);
and (n8358,n8359,n8360);
xor (n8359,n8357,n2195);
or (n8360,n8361,n8364);
and (n8361,n8362,n8363);
xor (n8362,n8295,n8296);
and (n8363,n1780,n108);
and (n8364,n8365,n8366);
xor (n8365,n8362,n8363);
and (n8366,n8367,n8368);
xor (n8367,n8301,n8302);
and (n8368,n1822,n108);
and (n8369,n206,n502);
or (n8370,n8371,n8374);
and (n8371,n8372,n8373);
xor (n8372,n8308,n8309);
and (n8373,n126,n502);
and (n8374,n8375,n8376);
xor (n8375,n8372,n8373);
or (n8376,n8377,n8380);
and (n8377,n8378,n8379);
xor (n8378,n8313,n8314);
and (n8379,n106,n502);
and (n8380,n8381,n8382);
xor (n8381,n8378,n8379);
or (n8382,n8383,n8386);
and (n8383,n8384,n8385);
xor (n8384,n8319,n8320);
and (n8385,n496,n502);
and (n8386,n8387,n8388);
xor (n8387,n8384,n8385);
or (n8388,n8389,n8392);
and (n8389,n8390,n8391);
xor (n8390,n8325,n8326);
and (n8391,n461,n502);
and (n8392,n8393,n8394);
xor (n8393,n8390,n8391);
or (n8394,n8395,n8398);
and (n8395,n8396,n8397);
xor (n8396,n8331,n8332);
and (n8397,n456,n502);
and (n8398,n8399,n8400);
xor (n8399,n8396,n8397);
or (n8400,n8401,n8404);
and (n8401,n8402,n8403);
xor (n8402,n8337,n8338);
and (n8403,n761,n502);
and (n8404,n8405,n8406);
xor (n8405,n8402,n8403);
or (n8406,n8407,n8410);
and (n8407,n8408,n8409);
xor (n8408,n8343,n8344);
and (n8409,n646,n502);
and (n8410,n8411,n8412);
xor (n8411,n8408,n8409);
or (n8412,n8413,n8416);
and (n8413,n8414,n8415);
xor (n8414,n8349,n8350);
and (n8415,n640,n502);
and (n8416,n8417,n8418);
xor (n8417,n8414,n8415);
or (n8418,n8419,n8422);
and (n8419,n8420,n8421);
xor (n8420,n8354,n8355);
and (n8421,n1317,n502);
and (n8422,n8423,n8424);
xor (n8423,n8420,n8421);
or (n8424,n8425,n8428);
and (n8425,n8426,n8427);
xor (n8426,n8359,n8360);
and (n8427,n1780,n502);
and (n8428,n8429,n8430);
xor (n8429,n8426,n8427);
and (n8430,n8431,n2354);
xor (n8431,n8365,n8366);
or (n8432,n8433,n8435);
and (n8433,n8434,n514);
xor (n8434,n8375,n8376);
and (n8435,n8436,n8437);
xor (n8436,n8434,n514);
or (n8437,n8438,n8440);
and (n8438,n8439,n497);
xor (n8439,n8381,n8382);
and (n8440,n8441,n8442);
xor (n8441,n8439,n497);
or (n8442,n8443,n8446);
and (n8443,n8444,n8445);
xor (n8444,n8387,n8388);
and (n8445,n461,n450);
and (n8446,n8447,n8448);
xor (n8447,n8444,n8445);
or (n8448,n8449,n8452);
and (n8449,n8450,n8451);
xor (n8450,n8393,n8394);
and (n8451,n456,n450);
and (n8452,n8453,n8454);
xor (n8453,n8450,n8451);
or (n8454,n8455,n8458);
and (n8455,n8456,n8457);
xor (n8456,n8399,n8400);
and (n8457,n761,n450);
and (n8458,n8459,n8460);
xor (n8459,n8456,n8457);
or (n8460,n8461,n8464);
and (n8461,n8462,n8463);
xor (n8462,n8405,n8406);
and (n8463,n646,n450);
and (n8464,n8465,n8466);
xor (n8465,n8462,n8463);
or (n8466,n8467,n8470);
and (n8467,n8468,n8469);
xor (n8468,n8411,n8412);
and (n8469,n640,n450);
and (n8470,n8471,n8472);
xor (n8471,n8468,n8469);
or (n8472,n8473,n8476);
and (n8473,n8474,n8475);
xor (n8474,n8417,n8418);
and (n8475,n1317,n450);
and (n8476,n8477,n8478);
xor (n8477,n8474,n8475);
or (n8478,n8479,n8482);
and (n8479,n8480,n8481);
xor (n8480,n8423,n8424);
and (n8481,n1780,n450);
and (n8482,n8483,n8484);
xor (n8483,n8480,n8481);
and (n8484,n8485,n8486);
xor (n8485,n8429,n8430);
and (n8486,n1822,n450);
and (n8487,n106,n445);
or (n8488,n8489,n8492);
and (n8489,n8490,n8491);
xor (n8490,n8436,n8437);
and (n8491,n496,n445);
and (n8492,n8493,n8494);
xor (n8493,n8490,n8491);
or (n8494,n8495,n8498);
and (n8495,n8496,n8497);
xor (n8496,n8441,n8442);
and (n8497,n461,n445);
and (n8498,n8499,n8500);
xor (n8499,n8496,n8497);
or (n8500,n8501,n8504);
and (n8501,n8502,n8503);
xor (n8502,n8447,n8448);
and (n8503,n456,n445);
and (n8504,n8505,n8506);
xor (n8505,n8502,n8503);
or (n8506,n8507,n8510);
and (n8507,n8508,n8509);
xor (n8508,n8453,n8454);
and (n8509,n761,n445);
and (n8510,n8511,n8512);
xor (n8511,n8508,n8509);
or (n8512,n8513,n8516);
and (n8513,n8514,n8515);
xor (n8514,n8459,n8460);
and (n8515,n646,n445);
and (n8516,n8517,n8518);
xor (n8517,n8514,n8515);
or (n8518,n8519,n8522);
and (n8519,n8520,n8521);
xor (n8520,n8465,n8466);
and (n8521,n640,n445);
and (n8522,n8523,n8524);
xor (n8523,n8520,n8521);
or (n8524,n8525,n8528);
and (n8525,n8526,n8527);
xor (n8526,n8471,n8472);
and (n8527,n1317,n445);
and (n8528,n8529,n8530);
xor (n8529,n8526,n8527);
or (n8530,n8531,n8534);
and (n8531,n8532,n8533);
xor (n8532,n8477,n8478);
and (n8533,n1780,n445);
and (n8534,n8535,n8536);
xor (n8535,n8532,n8533);
and (n8536,n8537,n1824);
xor (n8537,n8483,n8484);
and (n8538,n496,n444);
or (n8539,n8540,n8543);
and (n8540,n8541,n8542);
xor (n8541,n8493,n8494);
and (n8542,n461,n444);
and (n8543,n8544,n8545);
xor (n8544,n8541,n8542);
or (n8545,n8546,n8548);
and (n8546,n8547,n457);
xor (n8547,n8499,n8500);
and (n8548,n8549,n8550);
xor (n8549,n8547,n457);
or (n8550,n8551,n8553);
and (n8551,n8552,n966);
xor (n8552,n8505,n8506);
and (n8553,n8554,n8555);
xor (n8554,n8552,n966);
or (n8555,n8556,n8558);
and (n8556,n8557,n647);
xor (n8557,n8511,n8512);
and (n8558,n8559,n8560);
xor (n8559,n8557,n647);
or (n8560,n8561,n8564);
and (n8561,n8562,n8563);
xor (n8562,n8517,n8518);
and (n8563,n640,n444);
and (n8564,n8565,n8566);
xor (n8565,n8562,n8563);
or (n8566,n8567,n8570);
and (n8567,n8568,n8569);
xor (n8568,n8523,n8524);
and (n8569,n1317,n444);
and (n8570,n8571,n8572);
xor (n8571,n8568,n8569);
or (n8572,n8573,n8576);
and (n8573,n8574,n8575);
xor (n8574,n8529,n8530);
and (n8575,n1780,n444);
and (n8576,n8577,n8578);
xor (n8577,n8574,n8575);
and (n8578,n8579,n2576);
xor (n8579,n8535,n8536);
or (n8580,n8581,n8583);
and (n8581,n8582,n457);
xor (n8582,n8544,n8545);
and (n8583,n8584,n8585);
xor (n8584,n8582,n457);
or (n8585,n8586,n8588);
and (n8586,n8587,n966);
xor (n8587,n8549,n8550);
and (n8588,n8589,n8590);
xor (n8589,n8587,n966);
or (n8590,n8591,n8593);
and (n8591,n8592,n647);
xor (n8592,n8554,n8555);
and (n8593,n8594,n8595);
xor (n8594,n8592,n647);
or (n8595,n8596,n8598);
and (n8596,n8597,n8563);
xor (n8597,n8559,n8560);
and (n8598,n8599,n8600);
xor (n8599,n8597,n8563);
or (n8600,n8601,n8603);
and (n8601,n8602,n8569);
xor (n8602,n8565,n8566);
and (n8603,n8604,n8605);
xor (n8604,n8602,n8569);
or (n8605,n8606,n8608);
and (n8606,n8607,n8575);
xor (n8607,n8571,n8572);
and (n8608,n8609,n8610);
xor (n8609,n8607,n8575);
and (n8610,n8611,n2576);
xor (n8611,n8577,n8578);
or (n8612,n8613,n8615);
and (n8613,n8614,n966);
xor (n8614,n8584,n8585);
and (n8615,n8616,n8617);
xor (n8616,n8614,n966);
or (n8617,n8618,n8620);
and (n8618,n8619,n647);
xor (n8619,n8589,n8590);
and (n8620,n8621,n8622);
xor (n8621,n8619,n647);
or (n8622,n8623,n8625);
and (n8623,n8624,n8563);
xor (n8624,n8594,n8595);
and (n8625,n8626,n8627);
xor (n8626,n8624,n8563);
or (n8627,n8628,n8630);
and (n8628,n8629,n8569);
xor (n8629,n8599,n8600);
and (n8630,n8631,n8632);
xor (n8631,n8629,n8569);
or (n8632,n8633,n8635);
and (n8633,n8634,n8575);
xor (n8634,n8604,n8605);
and (n8635,n8636,n8637);
xor (n8636,n8634,n8575);
and (n8637,n8638,n2576);
xor (n8638,n8609,n8610);
or (n8639,n8640,n8642);
and (n8640,n8641,n647);
xor (n8641,n8616,n8617);
and (n8642,n8643,n8644);
xor (n8643,n8641,n647);
or (n8644,n8645,n8647);
and (n8645,n8646,n8563);
xor (n8646,n8621,n8622);
and (n8647,n8648,n8649);
xor (n8648,n8646,n8563);
or (n8649,n8650,n8652);
and (n8650,n8651,n8569);
xor (n8651,n8626,n8627);
and (n8652,n8653,n8654);
xor (n8653,n8651,n8569);
or (n8654,n8655,n8657);
and (n8655,n8656,n8575);
xor (n8656,n8631,n8632);
and (n8657,n8658,n8659);
xor (n8658,n8656,n8575);
and (n8659,n8660,n2576);
xor (n8660,n8636,n8637);
or (n8661,n8662,n8664);
and (n8662,n8663,n8563);
xor (n8663,n8643,n8644);
and (n8664,n8665,n8666);
xor (n8665,n8663,n8563);
or (n8666,n8667,n8669);
and (n8667,n8668,n8569);
xor (n8668,n8648,n8649);
and (n8669,n8670,n8671);
xor (n8670,n8668,n8569);
or (n8671,n8672,n8674);
and (n8672,n8673,n8575);
xor (n8673,n8653,n8654);
and (n8674,n8675,n8676);
xor (n8675,n8673,n8575);
and (n8676,n8677,n2576);
xor (n8677,n8658,n8659);
or (n8678,n8679,n8681);
and (n8679,n8680,n8569);
xor (n8680,n8665,n8666);
and (n8681,n8682,n8683);
xor (n8682,n8680,n8569);
or (n8683,n8684,n8686);
and (n8684,n8685,n8575);
xor (n8685,n8670,n8671);
and (n8686,n8687,n8688);
xor (n8687,n8685,n8575);
and (n8688,n8689,n2576);
xor (n8689,n8675,n8676);
or (n8690,n8691,n8693);
and (n8691,n8692,n8575);
xor (n8692,n8682,n8683);
and (n8693,n8694,n8695);
xor (n8694,n8692,n8575);
and (n8695,n8696,n2576);
xor (n8696,n8687,n8688);
and (n8697,n8698,n2576);
xor (n8698,n8694,n8695);
or (n8699,n8700,n8704,n8855);
and (n8700,n8701,n8703);
xor (n8701,n8702,n7252);
xor (n8702,n7249,n7250);
xor (n8703,n8698,n2576);
and (n8704,n8703,n8705);
or (n8705,n8706,n8710,n8854);
and (n8706,n8707,n8709);
xor (n8707,n8708,n7257);
xor (n8708,n7254,n7255);
xor (n8709,n8696,n2576);
and (n8710,n8709,n8711);
or (n8711,n8712,n8716,n8853);
and (n8712,n8713,n8715);
xor (n8713,n8714,n7262);
xor (n8714,n7259,n7260);
xor (n8715,n8689,n2576);
and (n8716,n8715,n8717);
or (n8717,n8718,n8722,n8852);
and (n8718,n8719,n8721);
xor (n8719,n8720,n7267);
xor (n8720,n7264,n7265);
xor (n8721,n8677,n2576);
and (n8722,n8721,n8723);
or (n8723,n8724,n8728,n8851);
and (n8724,n8725,n8727);
xor (n8725,n8726,n7272);
xor (n8726,n7269,n7270);
xor (n8727,n8660,n2576);
and (n8728,n8727,n8729);
or (n8729,n8730,n8734,n8850);
and (n8730,n8731,n8733);
xor (n8731,n8732,n7277);
xor (n8732,n7274,n7275);
xor (n8733,n8638,n2576);
and (n8734,n8733,n8735);
or (n8735,n8736,n8740,n8849);
and (n8736,n8737,n8739);
xor (n8737,n8738,n7282);
xor (n8738,n7279,n7280);
xor (n8739,n8611,n2576);
and (n8740,n8739,n8741);
or (n8741,n8742,n8746,n8848);
and (n8742,n8743,n8745);
xor (n8743,n8744,n7287);
xor (n8744,n7284,n7285);
xor (n8745,n8579,n2576);
and (n8746,n8745,n8747);
or (n8747,n8748,n8752,n8847);
and (n8748,n8749,n8751);
xor (n8749,n8750,n7292);
xor (n8750,n7289,n7290);
xor (n8751,n8537,n1824);
and (n8752,n8751,n8753);
or (n8753,n8754,n8758,n8846);
and (n8754,n8755,n8757);
xor (n8755,n8756,n7297);
xor (n8756,n7294,n7295);
xor (n8757,n8485,n8486);
and (n8758,n8757,n8759);
or (n8759,n8760,n8764,n8845);
and (n8760,n8761,n8763);
xor (n8761,n8762,n7302);
xor (n8762,n7299,n7300);
xor (n8763,n8431,n2354);
and (n8764,n8763,n8765);
or (n8765,n8766,n8770,n8844);
and (n8766,n8767,n8769);
xor (n8767,n8768,n7307);
xor (n8768,n7304,n7305);
xor (n8769,n8367,n8368);
and (n8770,n8769,n8771);
or (n8771,n8772,n8776,n8843);
and (n8772,n8773,n8775);
xor (n8773,n8774,n7312);
xor (n8774,n7309,n7310);
xor (n8775,n8303,n3101);
and (n8776,n8775,n8777);
or (n8777,n8778,n8782,n8842);
and (n8778,n8779,n8781);
xor (n8779,n8780,n7317);
xor (n8780,n7314,n7315);
xor (n8781,n8227,n8228);
and (n8782,n8781,n8783);
or (n8783,n8784,n8788,n8841);
and (n8784,n8785,n8787);
xor (n8785,n8786,n7322);
xor (n8786,n7319,n7320);
xor (n8787,n8153,n3558);
and (n8788,n8787,n8789);
or (n8789,n8790,n8794,n8840);
and (n8790,n8791,n8793);
xor (n8791,n8792,n7327);
xor (n8792,n7324,n7325);
xor (n8793,n8065,n8066);
and (n8794,n8793,n8795);
or (n8795,n8796,n8800,n8839);
and (n8796,n8797,n8799);
xor (n8797,n8798,n7332);
xor (n8798,n7329,n7330);
xor (n8799,n7978,n3831);
and (n8800,n8799,n8801);
or (n8801,n8802,n8806,n8838);
and (n8802,n8803,n8805);
xor (n8803,n8804,n7337);
xor (n8804,n7334,n7335);
xor (n8805,n7882,n7883);
and (n8806,n8805,n8807);
or (n8807,n8808,n8812,n8837);
and (n8808,n8809,n8811);
xor (n8809,n8810,n7342);
xor (n8810,n7339,n7340);
xor (n8811,n7790,n7791);
and (n8812,n8811,n8813);
or (n8813,n8814,n8818,n8836);
and (n8814,n8815,n8817);
xor (n8815,n8816,n7347);
xor (n8816,n7344,n7345);
xor (n8817,n7694,n7695);
and (n8818,n8817,n8819);
or (n8819,n8820,n8824,n8835);
and (n8820,n8821,n8823);
xor (n8821,n8822,n7352);
xor (n8822,n7349,n7350);
xor (n8823,n7604,n7605);
and (n8824,n8823,n8825);
or (n8825,n8826,n8830,n8834);
and (n8826,n8827,n8829);
xor (n8827,n8828,n4542);
xor (n8828,n7354,n7355);
xor (n8829,n7508,n7509);
and (n8830,n8829,n8831);
and (n8831,n8832,n8833);
xor (n8832,n4496,n4498);
not (n8833,n4494);
and (n8834,n8827,n8831);
and (n8835,n8821,n8825);
and (n8836,n8815,n8819);
and (n8837,n8809,n8813);
and (n8838,n8803,n8807);
and (n8839,n8797,n8801);
and (n8840,n8791,n8795);
and (n8841,n8785,n8789);
and (n8842,n8779,n8783);
and (n8843,n8773,n8777);
and (n8844,n8767,n8771);
and (n8845,n8761,n8765);
and (n8846,n8755,n8759);
and (n8847,n8749,n8753);
and (n8848,n8743,n8747);
and (n8849,n8737,n8741);
and (n8850,n8731,n8735);
and (n8851,n8725,n8729);
and (n8852,n8719,n8723);
and (n8853,n8713,n8717);
and (n8854,n8707,n8711);
and (n8855,n8701,n8705);
endmodule
