module top (out,n20,n25,n26,n27,n29,n30,n41,n44,n47
        ,n50,n53,n56,n59,n62,n65,n67,n70,n81,n91
        ,n96,n99,n102,n105,n108,n111,n114,n116,n118,n126
        ,n140,n145,n178,n183,n186,n189,n192,n205,n258,n263
        ,n266,n269,n272,n275,n278,n294,n404,n415);
output out;
input n20;
input n25;
input n26;
input n27;
input n29;
input n30;
input n41;
input n44;
input n47;
input n50;
input n53;
input n56;
input n59;
input n62;
input n65;
input n67;
input n70;
input n81;
input n91;
input n96;
input n99;
input n102;
input n105;
input n108;
input n111;
input n114;
input n116;
input n118;
input n126;
input n140;
input n145;
input n178;
input n183;
input n186;
input n189;
input n192;
input n205;
input n258;
input n263;
input n266;
input n269;
input n272;
input n275;
input n278;
input n294;
input n404;
input n415;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n21;
wire n22;
wire n23;
wire n24;
wire n28;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n42;
wire n43;
wire n45;
wire n46;
wire n48;
wire n49;
wire n51;
wire n52;
wire n54;
wire n55;
wire n57;
wire n58;
wire n60;
wire n61;
wire n63;
wire n64;
wire n66;
wire n68;
wire n69;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n92;
wire n93;
wire n94;
wire n95;
wire n97;
wire n98;
wire n100;
wire n101;
wire n103;
wire n104;
wire n106;
wire n107;
wire n109;
wire n110;
wire n112;
wire n113;
wire n115;
wire n117;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n141;
wire n142;
wire n143;
wire n144;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n179;
wire n180;
wire n181;
wire n182;
wire n184;
wire n185;
wire n187;
wire n188;
wire n190;
wire n191;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n259;
wire n260;
wire n261;
wire n262;
wire n264;
wire n265;
wire n267;
wire n268;
wire n270;
wire n271;
wire n273;
wire n274;
wire n276;
wire n277;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
xor (out,n0,n1505);
nand (n0,n1,n1504);
or (n1,n2,n800);
not (n2,n3);
nand (n3,n4,n799);
not (n4,n5);
nor (n5,n6,n720);
xor (n6,n7,n661);
xor (n7,n8,n487);
xor (n8,n9,n389);
xor (n9,n10,n224);
xor (n10,n11,n171);
xor (n11,n12,n132);
nand (n12,n13,n121);
or (n13,n14,n87);
nand (n14,n15,n77);
or (n15,n16,n74);
and (n16,n17,n71);
wire s0n17,s1n17,notn17;
or (n17,s0n17,s1n17);
not(notn17,n68);
and (s0n17,notn17,n18);
and (s1n17,n68,n37);
wire s0n18,s1n18,notn18;
or (n18,s0n18,s1n18);
not(notn18,n21);
and (s0n18,notn18,1'b0);
and (s1n18,n21,n20);
or (n21,n22,n33);
or (n22,n23,n31);
nor (n23,n24,n26,n27,n28,n30);
not (n24,n25);
not (n28,n29);
nor (n31,n25,n32,n27,n28,n30);
not (n32,n26);
or (n33,n34,n36);
and (n34,n24,n26,n27,n28,n35);
not (n35,n30);
nor (n36,n24,n32,n27,n28,n30);
xor (n37,n38,n39);
not (n38,n20);
and (n39,n40,n42);
not (n40,n41);
and (n42,n43,n45);
not (n43,n44);
and (n45,n46,n48);
not (n46,n47);
and (n48,n49,n51);
not (n49,n50);
and (n51,n52,n54);
not (n52,n53);
and (n54,n55,n57);
not (n55,n56);
and (n57,n58,n60);
not (n58,n59);
and (n60,n61,n63);
not (n61,n62);
and (n63,n64,n66);
not (n64,n65);
not (n66,n67);
and (n68,n69,n70);
or (n69,n23,n34);
wire s0n71,s1n71,notn71;
or (n71,s0n71,s1n71);
not(notn71,n68);
and (s0n71,notn71,n72);
and (s1n71,n68,n73);
wire s0n72,s1n72,notn72;
or (n72,s0n72,s1n72);
not(notn72,n21);
and (s0n72,notn72,1'b0);
and (s1n72,n21,n41);
xor (n73,n40,n42);
and (n74,n75,n76);
not (n75,n17);
not (n76,n71);
nand (n77,n78,n85);
or (n78,n75,n79);
wire s0n79,s1n79,notn79;
or (n79,s0n79,s1n79);
not(notn79,n68);
and (s0n79,notn79,n80);
and (s1n79,n68,n82);
wire s0n80,s1n80,notn80;
or (n80,s0n80,s1n80);
not(notn80,n21);
and (s0n80,notn80,1'b0);
and (s1n80,n21,n81);
xor (n82,n83,n84);
not (n83,n81);
and (n84,n38,n39);
or (n85,n86,n17);
not (n86,n79);
nor (n87,n88,n119);
and (n88,n86,n89);
wire s0n89,s1n89,notn89;
or (n89,s0n89,s1n89);
not(notn89,n117);
and (s0n89,notn89,n90);
and (s1n89,n117,n92);
wire s0n90,s1n90,notn90;
or (n90,s0n90,s1n90);
not(notn90,n21);
and (s0n90,notn90,1'b0);
and (s1n90,n21,n91);
xor (n92,n93,n94);
not (n93,n91);
and (n94,n95,n97);
not (n95,n96);
and (n97,n98,n100);
not (n98,n99);
and (n100,n101,n103);
not (n101,n102);
and (n103,n104,n106);
not (n104,n105);
and (n106,n107,n109);
not (n107,n108);
and (n109,n110,n112);
not (n110,n111);
and (n112,n113,n115);
not (n113,n114);
not (n115,n116);
and (n117,n69,n118);
and (n119,n79,n120);
not (n120,n89);
or (n121,n15,n122);
nor (n122,n123,n130);
and (n123,n86,n124);
wire s0n124,s1n124,notn124;
or (n124,s0n124,s1n124);
not(notn124,n117);
and (s0n124,notn124,n125);
and (s1n124,n117,n127);
wire s0n125,s1n125,notn125;
or (n125,s0n125,s1n125);
not(notn125,n21);
and (s0n125,notn125,1'b0);
and (s1n125,n21,n126);
xor (n127,n128,n129);
not (n128,n126);
and (n129,n93,n94);
and (n130,n79,n131);
not (n131,n124);
nand (n132,n133,n162);
or (n133,n134,n155);
or (n134,n135,n152);
nor (n135,n136,n150);
and (n136,n137,n147);
not (n137,n138);
wire s0n138,s1n138,notn138;
or (n138,s0n138,s1n138);
not(notn138,n68);
and (s0n138,notn138,n139);
and (s1n138,n68,n141);
wire s0n139,s1n139,notn139;
or (n139,s0n139,s1n139);
not(notn139,n21);
and (s0n139,notn139,1'b0);
and (s1n139,n21,n140);
xor (n141,n142,n143);
not (n142,n140);
and (n143,n144,n146);
not (n144,n145);
and (n146,n83,n84);
wire s0n147,s1n147,notn147;
or (n147,s0n147,s1n147);
not(notn147,n68);
and (s0n147,notn147,n148);
and (s1n147,n68,n149);
wire s0n148,s1n148,notn148;
or (n148,s0n148,s1n148);
not(notn148,n21);
and (s0n148,notn148,1'b0);
and (s1n148,n21,n145);
xor (n149,n144,n146);
and (n150,n151,n138);
not (n151,n147);
nor (n152,n153,n154);
and (n153,n147,n79);
and (n154,n151,n86);
nor (n155,n156,n160);
and (n156,n137,n157);
wire s0n157,s1n157,notn157;
or (n157,s0n157,s1n157);
not(notn157,n117);
and (s0n157,notn157,n158);
and (s1n157,n117,n159);
wire s0n158,s1n158,notn158;
or (n158,s0n158,s1n158);
not(notn158,n21);
and (s0n158,notn158,1'b0);
and (s1n158,n21,n99);
xor (n159,n98,n100);
and (n160,n138,n161);
not (n161,n157);
or (n162,n163,n170);
nor (n163,n164,n168);
and (n164,n137,n165);
wire s0n165,s1n165,notn165;
or (n165,s0n165,s1n165);
not(notn165,n117);
and (s0n165,notn165,n166);
and (s1n165,n117,n167);
wire s0n166,s1n166,notn166;
or (n166,s0n166,s1n166);
not(notn166,n21);
and (s0n166,notn166,1'b0);
and (s1n166,n21,n96);
xor (n167,n95,n97);
and (n168,n138,n169);
not (n169,n165);
not (n170,n152);
nand (n171,n172,n215);
or (n172,n173,n210);
or (n173,n174,n200);
nor (n174,n175,n197);
and (n175,n176,n194);
wire s0n176,s1n176,notn176;
or (n176,s0n176,s1n176);
not(notn176,n68);
and (s0n176,notn176,n177);
and (s1n176,n68,n179);
wire s0n177,s1n177,notn177;
or (n177,s0n177,s1n177);
not(notn177,n21);
and (s0n177,notn177,1'b0);
and (s1n177,n21,n178);
xor (n179,n180,n181);
not (n180,n178);
and (n181,n182,n184);
not (n182,n183);
and (n184,n185,n187);
not (n185,n186);
and (n187,n188,n190);
not (n188,n189);
and (n190,n191,n193);
not (n191,n192);
and (n193,n142,n143);
wire s0n194,s1n194,notn194;
or (n194,s0n194,s1n194);
not(notn194,n68);
and (s0n194,notn194,n195);
and (s1n194,n68,n196);
wire s0n195,s1n195,notn195;
or (n195,s0n195,s1n195);
not(notn195,n21);
and (s0n195,notn195,1'b0);
and (s1n195,n21,n183);
xor (n196,n182,n184);
and (n197,n198,n199);
not (n198,n176);
not (n199,n194);
nor (n200,n201,n209);
and (n201,n176,n202);
not (n202,n203);
wire s0n203,s1n203,notn203;
or (n203,s0n203,s1n203);
not(notn203,n68);
and (s0n203,notn203,n204);
and (s1n203,n68,n206);
wire s0n204,s1n204,notn204;
or (n204,s0n204,s1n204);
not(notn204,n21);
and (s0n204,notn204,1'b0);
and (s1n204,n21,n205);
xor (n206,n207,n208);
not (n207,n205);
and (n208,n180,n181);
and (n209,n198,n203);
nor (n210,n211,n214);
and (n211,n203,n212);
not (n212,n213);
wire s0n213,s1n213,notn213;
or (n213,s0n213,s1n213);
not(notn213,n21);
and (s0n213,notn213,1'b0);
and (s1n213,n21,n116);
and (n214,n202,n213);
or (n215,n216,n217);
not (n216,n174);
nor (n217,n218,n222);
and (n218,n219,n202);
wire s0n219,s1n219,notn219;
or (n219,s0n219,s1n219);
not(notn219,n117);
and (s0n219,notn219,n220);
and (s1n219,n117,n221);
wire s0n220,s1n220,notn220;
or (n220,s0n220,s1n220);
not(notn220,n21);
and (s0n220,notn220,1'b0);
and (s1n220,n21,n114);
xor (n221,n113,n115);
and (n222,n223,n203);
not (n223,n219);
or (n224,n225,n388);
and (n225,n226,n300);
xor (n226,n227,n237);
nand (n227,n228,n236);
or (n228,n134,n229);
nor (n229,n230,n234);
and (n230,n137,n231);
wire s0n231,s1n231,notn231;
or (n231,s0n231,s1n231);
not(notn231,n117);
and (s0n231,notn231,n232);
and (s1n231,n117,n233);
wire s0n232,s1n232,notn232;
or (n232,s0n232,s1n232);
not(notn232,n21);
and (s0n232,notn232,1'b0);
and (s1n232,n21,n102);
xor (n233,n101,n103);
and (n234,n138,n235);
not (n235,n231);
or (n236,n155,n170);
and (n237,n238,n252);
nor (n238,n239,n199);
nor (n239,n240,n250);
and (n240,n241,n245);
not (n241,n242);
wire s0n242,s1n242,notn242;
or (n242,s0n242,s1n242);
not(notn242,n68);
and (s0n242,notn242,n243);
and (s1n242,n68,n244);
wire s0n243,s1n243,notn243;
or (n243,s0n243,s1n243);
not(notn243,n21);
and (s0n243,notn243,1'b0);
and (s1n243,n21,n189);
xor (n244,n188,n190);
not (n245,n246);
and (n246,n213,n247);
wire s0n247,s1n247,notn247;
or (n247,s0n247,s1n247);
not(notn247,n68);
and (s0n247,notn247,n248);
and (s1n247,n68,n249);
wire s0n248,s1n248,notn248;
or (n248,s0n248,s1n248);
not(notn248,n21);
and (s0n248,notn248,1'b0);
and (s1n248,n21,n186);
xor (n249,n185,n187);
and (n250,n251,n212);
not (n251,n247);
nand (n252,n253,n289);
or (n253,n254,n286);
nor (n254,n255,n284);
and (n255,n256,n280);
wire s0n256,s1n256,notn256;
or (n256,s0n256,s1n256);
not(notn256,n117);
and (s0n256,notn256,n257);
and (s1n256,n117,n259);
wire s0n257,s1n257,notn257;
or (n257,s0n257,s1n257);
not(notn257,n21);
and (s0n257,notn257,1'b0);
and (s1n257,n21,n258);
xor (n259,n260,n261);
not (n260,n258);
and (n261,n262,n264);
not (n262,n263);
and (n264,n265,n267);
not (n265,n266);
and (n267,n268,n270);
not (n268,n269);
and (n270,n271,n273);
not (n271,n272);
and (n273,n274,n276);
not (n274,n275);
and (n276,n277,n279);
not (n277,n278);
and (n279,n128,n129);
not (n280,n281);
wire s0n281,s1n281,notn281;
or (n281,s0n281,s1n281);
not(notn281,n68);
and (s0n281,notn281,n282);
and (s1n281,n68,n283);
wire s0n282,s1n282,notn282;
or (n282,s0n282,s1n282);
not(notn282,n21);
and (s0n282,notn282,1'b0);
and (s1n282,n21,n65);
xor (n283,n64,n66);
and (n284,n285,n281);
not (n285,n256);
nand (n286,n281,n287);
not (n287,n288);
wire s0n288,s1n288,notn288;
or (n288,s0n288,s1n288);
not(notn288,n21);
and (s0n288,notn288,1'b0);
and (s1n288,n21,n67);
or (n289,n290,n287);
nor (n290,n291,n298);
and (n291,n292,n280);
wire s0n292,s1n292,notn292;
or (n292,s0n292,s1n292);
not(notn292,n117);
and (s0n292,notn292,n293);
and (s1n292,n117,n295);
wire s0n293,s1n293,notn293;
or (n293,s0n293,s1n293);
not(notn293,n21);
and (s0n293,notn293,1'b0);
and (s1n293,n21,n294);
xor (n295,n296,n297);
not (n296,n294);
and (n297,n260,n261);
and (n298,n299,n281);
not (n299,n292);
or (n300,n301,n387);
and (n301,n302,n369);
xor (n302,n303,n339);
nand (n303,n304,n331);
or (n304,n305,n324);
nand (n305,n306,n317);
or (n306,n307,n314);
and (n307,n308,n311);
wire s0n308,s1n308,notn308;
or (n308,s0n308,s1n308);
not(notn308,n68);
and (s0n308,notn308,n309);
and (s1n308,n68,n310);
wire s0n309,s1n309,notn309;
or (n309,s0n309,s1n309);
not(notn309,n21);
and (s0n309,notn309,1'b0);
and (s1n309,n21,n53);
xor (n310,n52,n54);
wire s0n311,s1n311,notn311;
or (n311,s0n311,s1n311);
not(notn311,n68);
and (s0n311,notn311,n312);
and (s1n311,n68,n313);
wire s0n312,s1n312,notn312;
or (n312,s0n312,s1n312);
not(notn312,n21);
and (s0n312,notn312,1'b0);
and (s1n312,n21,n50);
xor (n313,n49,n51);
and (n314,n315,n316);
not (n315,n308);
not (n316,n311);
nor (n317,n318,n322);
and (n318,n319,n311);
wire s0n319,s1n319,notn319;
or (n319,s0n319,s1n319);
not(notn319,n68);
and (s0n319,notn319,n320);
and (s1n319,n68,n321);
wire s0n320,s1n320,notn320;
or (n320,s0n320,s1n320);
not(notn320,n21);
and (s0n320,notn320,1'b0);
and (s1n320,n21,n47);
xor (n321,n46,n48);
and (n322,n323,n316);
not (n323,n319);
nor (n324,n325,n329);
and (n325,n326,n323);
wire s0n326,s1n326,notn326;
or (n326,s0n326,s1n326);
not(notn326,n117);
and (s0n326,notn326,n327);
and (s1n326,n117,n328);
wire s0n327,s1n327,notn327;
or (n327,s0n327,s1n327);
not(notn327,n21);
and (s0n327,notn327,1'b0);
and (s1n327,n21,n278);
xor (n328,n277,n279);
and (n329,n330,n319);
not (n330,n326);
or (n331,n332,n306);
nor (n332,n333,n337);
and (n333,n334,n323);
wire s0n334,s1n334,notn334;
or (n334,s0n334,s1n334);
not(notn334,n117);
and (s0n334,notn334,n335);
and (s1n334,n117,n336);
wire s0n335,s1n335,notn335;
or (n335,s0n335,s1n335);
not(notn335,n21);
and (s0n335,notn335,1'b0);
and (s1n335,n21,n275);
xor (n336,n274,n276);
and (n337,n338,n319);
not (n338,n334);
nand (n339,n340,n360);
or (n340,n341,n353);
not (n341,n342);
nor (n342,n343,n349);
nand (n343,n344,n348);
or (n344,n137,n345);
wire s0n345,s1n345,notn345;
or (n345,s0n345,s1n345);
not(notn345,n68);
and (s0n345,notn345,n346);
and (s1n345,n68,n347);
wire s0n346,s1n346,notn346;
or (n346,s0n346,s1n346);
not(notn346,n21);
and (s0n346,notn346,1'b0);
and (s1n346,n21,n192);
xor (n347,n191,n193);
nand (n348,n137,n345);
nor (n349,n350,n351);
and (n350,n241,n345);
and (n351,n352,n242);
not (n352,n345);
nor (n353,n354,n358);
and (n354,n355,n241);
wire s0n355,s1n355,notn355;
or (n355,s0n355,s1n355);
not(notn355,n117);
and (s0n355,notn355,n356);
and (s1n355,n117,n357);
wire s0n356,s1n356,notn356;
or (n356,s0n356,s1n356);
not(notn356,n21);
and (s0n356,notn356,1'b0);
and (s1n356,n21,n111);
xor (n357,n110,n112);
and (n358,n359,n242);
not (n359,n355);
or (n360,n361,n362);
not (n361,n343);
nor (n362,n363,n367);
and (n363,n364,n241);
wire s0n364,s1n364,notn364;
or (n364,s0n364,s1n364);
not(notn364,n117);
and (s0n364,notn364,n365);
and (s1n364,n117,n366);
wire s0n365,s1n365,notn365;
or (n365,s0n365,s1n365);
not(notn365,n21);
and (s0n365,notn365,1'b0);
and (s1n365,n21,n108);
xor (n366,n107,n109);
and (n367,n368,n242);
not (n368,n364);
nand (n369,n370,n383);
or (n370,n371,n375);
not (n371,n372);
nand (n372,n373,n374);
or (n373,n199,n213);
or (n374,n194,n212);
not (n375,n376);
and (n376,n377,n380);
nor (n377,n378,n379);
and (n378,n242,n251);
and (n379,n241,n247);
nand (n380,n381,n382);
or (n381,n251,n194);
or (n382,n199,n247);
or (n383,n384,n377);
nor (n384,n385,n386);
and (n385,n219,n199);
and (n386,n223,n194);
and (n387,n303,n339);
and (n388,n227,n237);
xor (n389,n390,n439);
xor (n390,n391,n421);
xor (n391,n392,n398);
nor (n392,n393,n202);
nor (n393,n394,n397);
and (n394,n395,n199);
not (n395,n396);
and (n396,n213,n176);
and (n397,n198,n212);
nand (n398,n399,n410);
or (n399,n400,n286);
nor (n400,n401,n408);
and (n401,n402,n280);
wire s0n402,s1n402,notn402;
or (n402,s0n402,s1n402);
not(notn402,n117);
and (s0n402,notn402,n403);
and (s1n402,n117,n405);
wire s0n403,s1n403,notn403;
or (n403,s0n403,s1n403);
not(notn403,n21);
and (s0n403,notn403,1'b0);
and (s1n403,n21,n404);
xor (n405,n406,n407);
not (n406,n404);
and (n407,n296,n297);
and (n408,n409,n281);
not (n409,n402);
or (n410,n411,n287);
nor (n411,n412,n419);
and (n412,n413,n280);
wire s0n413,s1n413,notn413;
or (n413,s0n413,s1n413);
not(notn413,n117);
and (s0n413,notn413,n414);
and (s1n413,n117,n416);
wire s0n414,s1n414,notn414;
or (n414,s0n414,s1n414);
not(notn414,n21);
and (s0n414,notn414,1'b0);
and (s1n414,n21,n415);
xor (n416,n417,n418);
not (n417,n415);
and (n418,n406,n407);
and (n419,n420,n281);
not (n420,n413);
or (n421,n422,n438);
and (n422,n423,n428);
xor (n423,n424,n425);
nor (n424,n216,n212);
nand (n425,n426,n427);
or (n426,n290,n286);
or (n427,n400,n287);
nand (n428,n429,n437);
or (n429,n430,n306);
nor (n430,n431,n435);
and (n431,n432,n323);
wire s0n432,s1n432,notn432;
or (n432,s0n432,s1n432);
not(notn432,n117);
and (s0n432,notn432,n433);
and (s1n432,n117,n434);
wire s0n433,s1n433,notn433;
or (n433,s0n433,s1n433);
not(notn433,n21);
and (s0n433,notn433,1'b0);
and (s1n433,n21,n272);
xor (n434,n271,n273);
and (n435,n436,n319);
not (n436,n432);
or (n437,n305,n332);
and (n438,n424,n425);
or (n439,n440,n486);
and (n440,n441,n458);
xor (n441,n442,n452);
nand (n442,n443,n444);
or (n443,n341,n362);
or (n444,n445,n361);
nor (n445,n446,n450);
and (n446,n241,n447);
wire s0n447,s1n447,notn447;
or (n447,s0n447,s1n447);
not(notn447,n117);
and (s0n447,notn447,n448);
and (s1n447,n117,n449);
wire s0n448,s1n448,notn448;
or (n448,s0n448,s1n448);
not(notn448,n21);
and (s0n448,notn448,1'b0);
and (s1n448,n21,n105);
xor (n449,n104,n106);
and (n450,n451,n242);
not (n451,n447);
nand (n452,n453,n454);
or (n453,n375,n384);
or (n454,n455,n377);
nor (n455,n456,n457);
and (n456,n355,n199);
and (n457,n359,n194);
nand (n458,n459,n482);
or (n459,n460,n475);
nand (n460,n461,n468);
nor (n461,n462,n466);
and (n462,n280,n463);
wire s0n463,s1n463,notn463;
or (n463,s0n463,s1n463);
not(notn463,n68);
and (s0n463,notn463,n464);
and (s1n463,n68,n465);
wire s0n464,s1n464,notn464;
or (n464,s0n464,s1n464);
not(notn464,n21);
and (s0n464,notn464,1'b0);
and (s1n464,n21,n62);
xor (n465,n61,n63);
and (n466,n281,n467);
not (n467,n463);
nand (n468,n469,n474);
or (n469,n470,n463);
not (n470,n471);
wire s0n471,s1n471,notn471;
or (n471,s0n471,s1n471);
not(notn471,n68);
and (s0n471,notn471,n472);
and (s1n471,n68,n473);
wire s0n472,s1n472,notn472;
or (n472,s0n472,s1n472);
not(notn472,n21);
and (s0n472,notn472,1'b0);
and (s1n472,n21,n59);
xor (n473,n58,n60);
nand (n474,n470,n463);
nor (n475,n476,n480);
and (n476,n470,n477);
wire s0n477,s1n477,notn477;
or (n477,s0n477,s1n477);
not(notn477,n117);
and (s0n477,notn477,n478);
and (s1n477,n117,n479);
wire s0n478,s1n478,notn478;
or (n478,s0n478,s1n478);
not(notn478,n21);
and (s0n478,notn478,1'b0);
and (s1n478,n21,n263);
xor (n479,n262,n264);
and (n480,n481,n471);
not (n481,n477);
or (n482,n461,n483);
nor (n483,n484,n485);
and (n484,n470,n256);
and (n485,n285,n471);
and (n486,n442,n452);
or (n487,n488,n660);
and (n488,n489,n637);
xor (n489,n490,n603);
or (n490,n491,n602);
and (n491,n492,n565);
xor (n492,n493,n521);
or (n493,n494,n520);
and (n494,n495,n503);
xor (n495,n496,n497);
nor (n496,n377,n212);
nand (n497,n498,n502);
or (n498,n499,n286);
nor (n499,n500,n501);
and (n500,n477,n280);
and (n501,n481,n281);
or (n502,n254,n287);
nand (n503,n504,n512);
or (n504,n460,n505);
nor (n505,n506,n510);
and (n506,n470,n507);
wire s0n507,s1n507,notn507;
or (n507,s0n507,s1n507);
not(notn507,n117);
and (s0n507,notn507,n508);
and (s1n507,n117,n509);
wire s0n508,s1n508,notn508;
or (n508,s0n508,s1n508);
not(notn508,n21);
and (s0n508,notn508,1'b0);
and (s1n508,n21,n269);
xor (n509,n268,n270);
and (n510,n511,n471);
not (n511,n507);
or (n512,n461,n513);
nor (n513,n514,n518);
and (n514,n470,n515);
wire s0n515,s1n515,notn515;
or (n515,s0n515,s1n515);
not(notn515,n117);
and (s0n515,notn515,n516);
and (s1n515,n117,n517);
wire s0n516,s1n516,notn516;
or (n516,s0n516,s1n516);
not(notn516,n21);
and (s0n516,notn516,1'b0);
and (s1n516,n21,n266);
xor (n517,n265,n267);
and (n518,n519,n471);
not (n519,n515);
and (n520,n496,n497);
or (n521,n522,n564);
and (n522,n523,n555);
xor (n523,n524,n545);
nand (n524,n525,n541);
or (n525,n526,n538);
nand (n526,n527,n534);
not (n527,n528);
nand (n528,n529,n533);
or (n529,n470,n530);
wire s0n530,s1n530,notn530;
or (n530,s0n530,s1n530);
not(notn530,n68);
and (s0n530,notn530,n531);
and (s1n530,n68,n532);
wire s0n531,s1n531,notn531;
or (n531,s0n531,s1n531);
not(notn531,n21);
and (s0n531,notn531,1'b0);
and (s1n531,n21,n56);
xor (n532,n55,n57);
nand (n533,n530,n470);
nor (n534,n535,n537);
and (n535,n315,n536);
not (n536,n530);
and (n537,n308,n530);
nor (n538,n539,n540);
and (n539,n334,n315);
and (n540,n338,n308);
or (n541,n527,n542);
nor (n542,n543,n544);
and (n543,n432,n315);
and (n544,n436,n308);
nand (n545,n546,n551);
or (n546,n547,n14);
not (n547,n548);
nand (n548,n549,n550);
or (n549,n235,n79);
or (n550,n86,n231);
or (n551,n552,n15);
nor (n552,n553,n554);
and (n553,n86,n157);
and (n554,n79,n161);
nand (n555,n556,n560);
or (n556,n134,n557);
nor (n557,n558,n559);
and (n558,n364,n137);
and (n559,n368,n138);
or (n560,n561,n170);
nor (n561,n562,n563);
and (n562,n137,n447);
and (n563,n451,n138);
and (n564,n524,n545);
or (n565,n566,n601);
and (n566,n567,n580);
xor (n567,n568,n574);
nand (n568,n569,n573);
or (n569,n341,n570);
nor (n570,n571,n572);
and (n571,n219,n241);
and (n572,n223,n242);
or (n573,n353,n361);
nand (n574,n575,n579);
or (n575,n305,n576);
nor (n576,n577,n578);
and (n577,n124,n323);
and (n578,n131,n319);
or (n579,n324,n306);
nand (n580,n581,n597);
or (n581,n582,n594);
nand (n582,n583,n590);
nor (n583,n584,n588);
and (n584,n585,n71);
wire s0n585,s1n585,notn585;
or (n585,s0n585,s1n585);
not(notn585,n68);
and (s0n585,notn585,n586);
and (s1n585,n68,n587);
wire s0n586,s1n586,notn586;
or (n586,s0n586,s1n586);
not(notn586,n21);
and (s0n586,notn586,1'b0);
and (s1n586,n21,n44);
xor (n587,n43,n45);
and (n588,n589,n76);
not (n589,n585);
not (n590,n591);
nor (n591,n592,n593);
and (n592,n319,n585);
and (n593,n323,n589);
nor (n594,n595,n596);
and (n595,n76,n165);
and (n596,n71,n169);
or (n597,n598,n590);
nor (n598,n599,n600);
and (n599,n76,n89);
and (n600,n71,n120);
and (n601,n568,n574);
and (n602,n493,n521);
or (n603,n604,n636);
and (n604,n605,n624);
xor (n605,n606,n607);
xor (n606,n302,n369);
xor (n607,n608,n618);
xor (n608,n609,n612);
nand (n609,n610,n611);
or (n610,n460,n513);
or (n611,n461,n475);
nand (n612,n613,n614);
or (n613,n582,n598);
or (n614,n615,n590);
nor (n615,n616,n617);
and (n616,n76,n124);
and (n617,n71,n131);
nand (n618,n619,n620);
or (n619,n542,n526);
or (n620,n527,n621);
nor (n621,n622,n623);
and (n622,n507,n315);
and (n623,n511,n308);
xor (n624,n625,n635);
xor (n625,n626,n632);
nand (n626,n627,n628);
or (n627,n14,n552);
or (n628,n629,n15);
nor (n629,n630,n631);
and (n630,n86,n165);
and (n631,n79,n169);
nand (n632,n633,n634);
or (n633,n134,n561);
or (n634,n170,n229);
xor (n635,n238,n252);
and (n636,n606,n607);
xor (n637,n638,n659);
xor (n638,n639,n642);
or (n639,n640,n641);
and (n640,n608,n618);
and (n641,n609,n612);
xor (n642,n643,n656);
xor (n643,n644,n650);
nand (n644,n645,n646);
or (n645,n582,n615);
or (n646,n647,n590);
nor (n647,n648,n649);
and (n648,n76,n326);
and (n649,n71,n330);
nand (n650,n651,n652);
or (n651,n526,n621);
or (n652,n527,n653);
nor (n653,n654,n655);
and (n654,n515,n315);
and (n655,n519,n308);
nand (n656,n657,n658);
or (n657,n14,n629);
or (n658,n15,n87);
xor (n659,n423,n428);
and (n660,n490,n603);
xor (n661,n662,n711);
xor (n662,n663,n666);
or (n663,n664,n665);
and (n664,n638,n659);
and (n665,n639,n642);
xor (n666,n667,n691);
xor (n667,n668,n671);
or (n668,n669,n670);
and (n669,n643,n656);
and (n670,n644,n650);
xor (n671,n672,n685);
xor (n672,n673,n679);
nand (n673,n674,n675);
or (n674,n460,n483);
or (n675,n676,n461);
nor (n676,n677,n678);
and (n677,n292,n470);
and (n678,n299,n471);
nand (n679,n680,n681);
or (n680,n582,n647);
or (n681,n682,n590);
nor (n682,n683,n684);
and (n683,n76,n334);
and (n684,n71,n338);
nand (n685,n686,n687);
or (n686,n526,n653);
or (n687,n527,n688);
nor (n688,n689,n690);
and (n689,n477,n315);
and (n690,n481,n308);
xor (n691,n692,n705);
xor (n692,n693,n699);
nand (n693,n694,n695);
or (n694,n305,n430);
or (n695,n306,n696);
nor (n696,n697,n698);
and (n697,n507,n323);
and (n698,n511,n319);
nand (n699,n700,n701);
or (n700,n341,n445);
or (n701,n361,n702);
nor (n702,n703,n704);
and (n703,n231,n241);
and (n704,n235,n242);
nand (n705,n706,n707);
or (n706,n375,n455);
or (n707,n708,n377);
nor (n708,n709,n710);
and (n709,n364,n199);
and (n710,n368,n194);
or (n711,n712,n719);
and (n712,n713,n718);
xor (n713,n714,n715);
xor (n714,n441,n458);
or (n715,n716,n717);
and (n716,n625,n635);
and (n717,n626,n632);
xor (n718,n226,n300);
and (n719,n714,n715);
or (n720,n721,n798);
and (n721,n722,n797);
xor (n722,n723,n724);
xor (n723,n713,n718);
or (n724,n725,n796);
and (n725,n726,n768);
xor (n726,n727,n767);
or (n727,n728,n766);
and (n728,n729,n744);
xor (n729,n730,n743);
and (n730,n731,n737);
nand (n731,n732,n736);
or (n732,n733,n286);
nor (n733,n734,n735);
and (n734,n515,n280);
and (n735,n519,n281);
or (n736,n499,n287);
nor (n737,n738,n241);
nor (n738,n739,n742);
and (n739,n137,n740);
not (n740,n741);
and (n741,n213,n345);
and (n742,n352,n212);
xor (n743,n495,n503);
or (n744,n745,n765);
and (n745,n746,n759);
xor (n746,n747,n753);
nand (n747,n748,n752);
or (n748,n460,n749);
nor (n749,n750,n751);
and (n750,n432,n470);
and (n751,n436,n471);
or (n752,n461,n505);
nand (n753,n754,n758);
or (n754,n341,n755);
nor (n755,n756,n757);
and (n756,n242,n212);
and (n757,n241,n213);
or (n758,n570,n361);
nand (n759,n760,n761);
or (n760,n576,n306);
or (n761,n305,n762);
nor (n762,n763,n764);
and (n763,n89,n323);
and (n764,n120,n319);
and (n765,n747,n753);
and (n766,n730,n743);
xor (n767,n492,n565);
or (n768,n769,n795);
and (n769,n770,n794);
xor (n770,n771,n793);
or (n771,n772,n792);
and (n772,n773,n786);
xor (n773,n774,n780);
nand (n774,n775,n779);
or (n775,n582,n776);
nor (n776,n777,n778);
and (n777,n76,n157);
and (n778,n71,n161);
or (n779,n594,n590);
nand (n780,n781,n785);
or (n781,n526,n782);
nor (n782,n783,n784);
and (n783,n326,n315);
and (n784,n330,n308);
or (n785,n527,n538);
nand (n786,n787,n788);
or (n787,n15,n547);
or (n788,n14,n789);
nor (n789,n790,n791);
and (n790,n86,n447);
and (n791,n79,n451);
and (n792,n774,n780);
xor (n793,n523,n555);
xor (n794,n567,n580);
and (n795,n771,n793);
and (n796,n727,n767);
xor (n797,n489,n637);
and (n798,n723,n724);
nand (n799,n6,n720);
not (n800,n801);
nand (n801,n802,n1502);
or (n802,n803,n1497);
nor (n803,n804,n1493);
not (n804,n805);
nand (n805,n806,n1462);
or (n806,n807,n1461);
and (n807,n808,n1051);
xor (n808,n809,n1022);
or (n809,n810,n1021);
and (n810,n811,n970);
xor (n811,n812,n889);
xor (n812,n813,n858);
xor (n813,n814,n829);
xor (n814,n815,n823);
xor (n815,n816,n817);
nor (n816,n361,n212);
nand (n817,n818,n822);
or (n818,n819,n286);
nor (n819,n820,n821);
and (n820,n280,n507);
and (n821,n511,n281);
or (n822,n733,n287);
nand (n823,n824,n828);
or (n824,n460,n825);
nor (n825,n826,n827);
and (n826,n470,n334);
and (n827,n338,n471);
or (n828,n461,n749);
or (n829,n830,n857);
and (n830,n831,n847);
xor (n831,n832,n838);
nand (n832,n833,n837);
or (n833,n460,n834);
nor (n834,n835,n836);
and (n835,n470,n326);
and (n836,n330,n471);
or (n837,n461,n825);
nand (n838,n839,n843);
or (n839,n305,n840);
nor (n840,n841,n842);
and (n841,n157,n323);
and (n842,n161,n319);
or (n843,n306,n844);
nor (n844,n845,n846);
and (n845,n165,n323);
and (n846,n169,n319);
nand (n847,n848,n853);
or (n848,n849,n582);
not (n849,n850);
nand (n850,n851,n852);
or (n851,n71,n451);
or (n852,n76,n447);
or (n853,n854,n590);
nor (n854,n855,n856);
and (n855,n76,n231);
and (n856,n71,n235);
and (n857,n832,n838);
or (n858,n859,n888);
and (n859,n860,n879);
xor (n860,n861,n870);
nand (n861,n862,n866);
or (n862,n526,n863);
nor (n863,n864,n865);
and (n864,n89,n315);
and (n865,n120,n308);
or (n866,n867,n527);
nor (n867,n868,n869);
and (n868,n124,n315);
and (n869,n131,n308);
nand (n870,n871,n875);
or (n871,n14,n872);
nor (n872,n873,n874);
and (n873,n355,n86);
and (n874,n359,n79);
or (n875,n876,n15);
nor (n876,n877,n878);
and (n877,n364,n86);
and (n878,n368,n79);
nand (n879,n880,n884);
or (n880,n170,n881);
nor (n881,n882,n883);
and (n882,n219,n137);
and (n883,n223,n138);
or (n884,n134,n885);
nor (n885,n886,n887);
and (n886,n138,n212);
and (n887,n137,n213);
and (n888,n861,n870);
xor (n889,n890,n926);
xor (n890,n891,n915);
xor (n891,n892,n902);
xor (n892,n893,n896);
nand (n893,n894,n895);
or (n894,n14,n876);
or (n895,n789,n15);
nand (n896,n897,n898);
or (n897,n134,n881);
or (n898,n899,n170);
nor (n899,n900,n901);
and (n900,n355,n137);
and (n901,n359,n138);
and (n902,n903,n909);
nand (n903,n904,n908);
or (n904,n905,n286);
nor (n905,n906,n907);
and (n906,n280,n432);
and (n907,n436,n281);
or (n908,n819,n287);
nor (n909,n910,n137);
nor (n910,n911,n914);
and (n911,n86,n912);
not (n912,n913);
and (n913,n213,n147);
and (n914,n151,n212);
xor (n915,n916,n923);
xor (n916,n917,n920);
nand (n917,n918,n919);
or (n918,n305,n844);
or (n919,n762,n306);
nand (n920,n921,n922);
or (n921,n582,n854);
or (n922,n776,n590);
nand (n923,n924,n925);
or (n924,n527,n782);
or (n925,n526,n867);
or (n926,n927,n969);
and (n927,n928,n947);
xor (n928,n929,n930);
xor (n929,n903,n909);
or (n930,n931,n946);
and (n931,n932,n940);
xor (n932,n933,n934);
nor (n933,n170,n212);
nand (n934,n935,n939);
or (n935,n936,n286);
nor (n936,n937,n938);
and (n937,n280,n334);
and (n938,n338,n281);
or (n939,n905,n287);
nand (n940,n941,n942);
or (n941,n461,n834);
or (n942,n460,n943);
nor (n943,n944,n945);
and (n944,n124,n470);
and (n945,n131,n471);
and (n946,n933,n934);
or (n947,n948,n968);
and (n948,n949,n962);
xor (n949,n950,n956);
nand (n950,n951,n955);
or (n951,n305,n952);
nor (n952,n953,n954);
and (n953,n231,n323);
and (n954,n235,n319);
or (n955,n840,n306);
nand (n956,n957,n958);
or (n957,n590,n849);
or (n958,n582,n959);
nor (n959,n960,n961);
and (n960,n76,n364);
and (n961,n71,n368);
nand (n962,n963,n964);
or (n963,n15,n872);
or (n964,n14,n965);
nor (n965,n966,n967);
and (n966,n219,n86);
and (n967,n223,n79);
and (n968,n950,n956);
and (n969,n929,n930);
or (n970,n971,n1020);
and (n971,n972,n975);
xor (n972,n973,n974);
xor (n973,n860,n879);
xor (n974,n831,n847);
or (n975,n976,n1019);
and (n976,n977,n997);
xor (n977,n978,n984);
nand (n978,n979,n983);
or (n979,n526,n980);
nor (n980,n981,n982);
and (n981,n165,n315);
and (n982,n169,n308);
or (n983,n527,n863);
and (n984,n985,n991);
nand (n985,n986,n990);
or (n986,n987,n286);
nor (n987,n988,n989);
and (n988,n326,n280);
and (n989,n330,n281);
or (n990,n936,n287);
nor (n991,n992,n86);
nor (n992,n993,n996);
and (n993,n76,n994);
not (n994,n995);
and (n995,n213,n17);
and (n996,n75,n212);
or (n997,n998,n1018);
and (n998,n999,n1012);
xor (n999,n1000,n1006);
nand (n1000,n1001,n1005);
or (n1001,n460,n1002);
nor (n1002,n1003,n1004);
and (n1003,n89,n470);
and (n1004,n120,n471);
or (n1005,n461,n943);
nand (n1006,n1007,n1011);
or (n1007,n305,n1008);
nor (n1008,n1009,n1010);
and (n1009,n447,n323);
and (n1010,n451,n319);
or (n1011,n952,n306);
nand (n1012,n1013,n1017);
or (n1013,n582,n1014);
nor (n1014,n1015,n1016);
and (n1015,n355,n76);
and (n1016,n359,n71);
or (n1017,n959,n590);
and (n1018,n1000,n1006);
and (n1019,n978,n984);
and (n1020,n973,n974);
and (n1021,n812,n889);
xor (n1022,n1023,n1036);
xor (n1023,n1024,n1033);
xor (n1024,n1025,n1032);
xor (n1025,n1026,n1029);
or (n1026,n1027,n1028);
and (n1027,n916,n923);
and (n1028,n917,n920);
or (n1029,n1030,n1031);
and (n1030,n892,n902);
and (n1031,n893,n896);
xor (n1032,n773,n786);
or (n1033,n1034,n1035);
and (n1034,n890,n926);
and (n1035,n891,n915);
xor (n1036,n1037,n1042);
xor (n1037,n1038,n1039);
xor (n1038,n746,n759);
or (n1039,n1040,n1041);
and (n1040,n813,n858);
and (n1041,n814,n829);
xor (n1042,n1043,n1048);
xor (n1043,n1044,n1047);
nand (n1044,n1045,n1046);
or (n1045,n134,n899);
or (n1046,n557,n170);
xor (n1047,n731,n737);
or (n1048,n1049,n1050);
and (n1049,n815,n823);
and (n1050,n816,n817);
or (n1051,n1052,n1460);
and (n1052,n1053,n1084);
xor (n1053,n1054,n1083);
or (n1054,n1055,n1082);
and (n1055,n1056,n1081);
xor (n1056,n1057,n1080);
or (n1057,n1058,n1079);
and (n1058,n1059,n1062);
xor (n1059,n1060,n1061);
xor (n1060,n932,n940);
xor (n1061,n949,n962);
or (n1062,n1063,n1078);
and (n1063,n1064,n1077);
xor (n1064,n1065,n1071);
nand (n1065,n1066,n1070);
or (n1066,n14,n1067);
nor (n1067,n1068,n1069);
and (n1068,n79,n212);
and (n1069,n86,n213);
or (n1070,n965,n15);
nand (n1071,n1072,n1076);
or (n1072,n526,n1073);
nor (n1073,n1074,n1075);
and (n1074,n157,n315);
and (n1075,n161,n308);
or (n1076,n980,n527);
xor (n1077,n985,n991);
and (n1078,n1065,n1071);
and (n1079,n1060,n1061);
xor (n1080,n928,n947);
xor (n1081,n972,n975);
and (n1082,n1057,n1080);
xor (n1083,n811,n970);
nand (n1084,n1085,n1457,n1459);
or (n1085,n1086,n1452);
nand (n1086,n1087,n1441);
or (n1087,n1088,n1440);
and (n1088,n1089,n1210);
xor (n1089,n1090,n1195);
or (n1090,n1091,n1194);
and (n1091,n1092,n1160);
xor (n1092,n1093,n1115);
xor (n1093,n1094,n1109);
xor (n1094,n1095,n1102);
nand (n1095,n1096,n1101);
or (n1096,n305,n1097);
not (n1097,n1098);
nor (n1098,n1099,n1100);
and (n1099,n323,n368);
and (n1100,n364,n319);
or (n1101,n1008,n306);
nand (n1102,n1103,n1108);
or (n1103,n1104,n582);
not (n1104,n1105);
nand (n1105,n1106,n1107);
or (n1106,n223,n71);
or (n1107,n219,n76);
or (n1108,n1014,n590);
nand (n1109,n1110,n1114);
or (n1110,n526,n1111);
nor (n1111,n1112,n1113);
and (n1112,n231,n315);
and (n1113,n235,n308);
or (n1114,n527,n1073);
or (n1115,n1116,n1159);
and (n1116,n1117,n1139);
xor (n1117,n1118,n1124);
nand (n1118,n1119,n1123);
or (n1119,n526,n1120);
nor (n1120,n1121,n1122);
and (n1121,n447,n315);
and (n1122,n451,n308);
or (n1123,n1111,n527);
xor (n1124,n1125,n1131);
nor (n1125,n1126,n76);
nor (n1126,n1127,n1130);
and (n1127,n1128,n323);
not (n1128,n1129);
and (n1129,n213,n585);
and (n1130,n589,n212);
nand (n1131,n1132,n1135);
or (n1132,n286,n1133);
not (n1133,n1134);
xnor (n1134,n89,n280);
or (n1135,n1136,n287);
nor (n1136,n1137,n1138);
and (n1137,n280,n124);
and (n1138,n131,n281);
or (n1139,n1140,n1158);
and (n1140,n1141,n1149);
xor (n1141,n1142,n1143);
nor (n1142,n590,n212);
nand (n1143,n1144,n1145);
or (n1144,n287,n1133);
or (n1145,n1146,n286);
nor (n1146,n1147,n1148);
and (n1147,n280,n165);
and (n1148,n169,n281);
nand (n1149,n1150,n1154);
or (n1150,n305,n1151);
nor (n1151,n1152,n1153);
and (n1152,n219,n323);
and (n1153,n223,n319);
or (n1154,n1155,n306);
nor (n1155,n1156,n1157);
and (n1156,n355,n323);
and (n1157,n359,n319);
and (n1158,n1142,n1143);
and (n1159,n1118,n1124);
xor (n1160,n1161,n1175);
xor (n1161,n1162,n1163);
and (n1162,n1125,n1131);
xor (n1163,n1164,n1169);
xor (n1164,n1165,n1166);
nor (n1165,n15,n212);
nand (n1166,n1167,n1168);
or (n1167,n1136,n286);
or (n1168,n987,n287);
nand (n1169,n1170,n1174);
or (n1170,n460,n1171);
nor (n1171,n1172,n1173);
and (n1172,n165,n470);
and (n1173,n169,n471);
or (n1174,n461,n1002);
or (n1175,n1176,n1193);
and (n1176,n1177,n1187);
xor (n1177,n1178,n1184);
nand (n1178,n1179,n1183);
or (n1179,n460,n1180);
nor (n1180,n1181,n1182);
and (n1181,n470,n157);
and (n1182,n161,n471);
or (n1183,n1171,n461);
nand (n1184,n1185,n1186);
or (n1185,n306,n1097);
or (n1186,n1155,n305);
nand (n1187,n1188,n1189);
or (n1188,n590,n1104);
or (n1189,n582,n1190);
nor (n1190,n1191,n1192);
and (n1191,n71,n212);
and (n1192,n76,n213);
and (n1193,n1178,n1184);
and (n1194,n1093,n1115);
xor (n1195,n1196,n1201);
xor (n1196,n1197,n1198);
xor (n1197,n999,n1012);
or (n1198,n1199,n1200);
and (n1199,n1161,n1175);
and (n1200,n1162,n1163);
xor (n1201,n1202,n1209);
xor (n1202,n1203,n1206);
or (n1203,n1204,n1205);
and (n1204,n1164,n1169);
and (n1205,n1165,n1166);
or (n1206,n1207,n1208);
and (n1207,n1094,n1109);
and (n1208,n1095,n1102);
xor (n1209,n1064,n1077);
or (n1210,n1211,n1439);
and (n1211,n1212,n1249);
xor (n1212,n1213,n1248);
or (n1213,n1214,n1247);
and (n1214,n1215,n1246);
xor (n1215,n1216,n1245);
or (n1216,n1217,n1244);
and (n1217,n1218,n1231);
xor (n1218,n1219,n1225);
nand (n1219,n1220,n1224);
or (n1220,n460,n1221);
nor (n1221,n1222,n1223);
and (n1222,n231,n470);
and (n1223,n471,n235);
or (n1224,n1180,n461);
nand (n1225,n1226,n1230);
or (n1226,n526,n1227);
nor (n1227,n1228,n1229);
and (n1228,n364,n315);
and (n1229,n368,n308);
or (n1230,n1120,n527);
and (n1231,n1232,n1238);
nor (n1232,n1233,n323);
nor (n1233,n1234,n1237);
and (n1234,n1235,n315);
not (n1235,n1236);
and (n1236,n213,n311);
and (n1237,n316,n212);
nand (n1238,n1239,n1243);
or (n1239,n1240,n286);
nor (n1240,n1241,n1242);
and (n1241,n280,n157);
and (n1242,n161,n281);
or (n1243,n1146,n287);
and (n1244,n1219,n1225);
xor (n1245,n1177,n1187);
xor (n1246,n1117,n1139);
and (n1247,n1216,n1245);
xor (n1248,n1092,n1160);
nand (n1249,n1250,n1436,n1438);
or (n1250,n1251,n1309);
nand (n1251,n1252,n1304);
not (n1252,n1253);
nor (n1253,n1254,n1280);
xor (n1254,n1255,n1279);
xor (n1255,n1256,n1278);
or (n1256,n1257,n1277);
and (n1257,n1258,n1271);
xor (n1258,n1259,n1265);
nand (n1259,n1260,n1264);
or (n1260,n305,n1261);
nor (n1261,n1262,n1263);
and (n1262,n319,n212);
and (n1263,n323,n213);
or (n1264,n1151,n306);
nand (n1265,n1266,n1270);
or (n1266,n1267,n460);
nor (n1267,n1268,n1269);
and (n1268,n471,n451);
and (n1269,n470,n447);
or (n1270,n1221,n461);
nand (n1271,n1272,n1276);
or (n1272,n526,n1273);
nor (n1273,n1274,n1275);
and (n1274,n355,n315);
and (n1275,n359,n308);
or (n1276,n1227,n527);
and (n1277,n1259,n1265);
xor (n1278,n1141,n1149);
xor (n1279,n1218,n1231);
or (n1280,n1281,n1303);
and (n1281,n1282,n1302);
xor (n1282,n1283,n1284);
xor (n1283,n1232,n1238);
or (n1284,n1285,n1301);
and (n1285,n1286,n1295);
xor (n1286,n1287,n1288);
nor (n1287,n306,n212);
nand (n1288,n1289,n1294);
or (n1289,n1290,n286);
not (n1290,n1291);
nand (n1291,n1292,n1293);
or (n1292,n281,n235);
nand (n1293,n235,n281);
or (n1294,n1240,n287);
nand (n1295,n1296,n1300);
or (n1296,n460,n1297);
nor (n1297,n1298,n1299);
and (n1298,n470,n364);
and (n1299,n471,n368);
or (n1300,n1267,n461);
and (n1301,n1287,n1288);
xor (n1302,n1258,n1271);
and (n1303,n1283,n1284);
or (n1304,n1305,n1306);
xor (n1305,n1215,n1246);
or (n1306,n1307,n1308);
and (n1307,n1255,n1279);
and (n1308,n1256,n1278);
nor (n1309,n1310,n1435);
and (n1310,n1311,n1430);
or (n1311,n1312,n1429);
and (n1312,n1313,n1354);
xor (n1313,n1314,n1347);
or (n1314,n1315,n1346);
and (n1315,n1316,n1332);
xor (n1316,n1317,n1323);
nand (n1317,n1318,n1322);
or (n1318,n460,n1319);
nor (n1319,n1320,n1321);
and (n1320,n471,n359);
and (n1321,n470,n355);
or (n1322,n1297,n461);
or (n1323,n1324,n1328);
nor (n1324,n1325,n527);
nor (n1325,n1326,n1327);
and (n1326,n315,n219);
and (n1327,n308,n223);
nor (n1328,n526,n1329);
nor (n1329,n1330,n1331);
and (n1330,n308,n212);
and (n1331,n315,n213);
xor (n1332,n1333,n1339);
nor (n1333,n1334,n315);
nor (n1334,n1335,n1338);
and (n1335,n1336,n470);
not (n1336,n1337);
and (n1337,n213,n530);
and (n1338,n536,n212);
nand (n1339,n1340,n1345);
or (n1340,n286,n1341);
not (n1341,n1342);
nand (n1342,n1343,n1344);
or (n1343,n280,n447);
nand (n1344,n447,n280);
nand (n1345,n1291,n288);
and (n1346,n1317,n1323);
xor (n1347,n1348,n1353);
xor (n1348,n1349,n1352);
nand (n1349,n1350,n1351);
or (n1350,n526,n1325);
or (n1351,n1273,n527);
and (n1352,n1333,n1339);
xor (n1353,n1286,n1295);
or (n1354,n1355,n1428);
and (n1355,n1356,n1376);
xor (n1356,n1357,n1375);
or (n1357,n1358,n1374);
and (n1358,n1359,n1368);
xor (n1359,n1360,n1361);
and (n1360,n528,n213);
nand (n1361,n1362,n1367);
or (n1362,n286,n1363);
not (n1363,n1364);
nand (n1364,n1365,n1366);
or (n1365,n281,n368);
nand (n1366,n368,n281);
nand (n1367,n1342,n288);
nand (n1368,n1369,n1373);
or (n1369,n460,n1370);
nor (n1370,n1371,n1372);
and (n1371,n470,n219);
and (n1372,n471,n223);
or (n1373,n1319,n461);
and (n1374,n1360,n1361);
xor (n1375,n1316,n1332);
or (n1376,n1377,n1427);
and (n1377,n1378,n1395);
xor (n1378,n1379,n1394);
and (n1379,n1380,n1386);
and (n1380,n1381,n471);
nand (n1381,n1382,n1385);
nand (n1382,n1383,n280);
not (n1383,n1384);
and (n1384,n213,n463);
nand (n1385,n467,n212);
nand (n1386,n1387,n1388);
or (n1387,n287,n1363);
nand (n1388,n1389,n1393);
not (n1389,n1390);
nor (n1390,n1391,n1392);
and (n1391,n359,n281);
and (n1392,n355,n280);
not (n1393,n286);
xor (n1394,n1359,n1368);
or (n1395,n1396,n1426);
and (n1396,n1397,n1405);
xor (n1397,n1398,n1404);
nand (n1398,n1399,n1403);
or (n1399,n460,n1400);
nor (n1400,n1401,n1402);
and (n1401,n471,n212);
and (n1402,n470,n213);
or (n1403,n1370,n461);
xor (n1404,n1380,n1386);
or (n1405,n1406,n1425);
and (n1406,n1407,n1415);
xor (n1407,n1408,n1409);
nor (n1408,n461,n212);
nand (n1409,n1410,n1414);
or (n1410,n1411,n286);
or (n1411,n1412,n1413);
and (n1412,n280,n223);
and (n1413,n219,n281);
or (n1414,n1390,n287);
nor (n1415,n1416,n1423);
nor (n1416,n1417,n1419);
and (n1417,n1418,n288);
not (n1418,n1411);
and (n1419,n1420,n1393);
nand (n1420,n1421,n1422);
or (n1421,n280,n213);
or (n1422,n281,n212);
or (n1423,n280,n1424);
and (n1424,n213,n288);
and (n1425,n1408,n1409);
and (n1426,n1398,n1404);
and (n1427,n1379,n1394);
and (n1428,n1357,n1375);
and (n1429,n1314,n1347);
or (n1430,n1431,n1432);
xor (n1431,n1282,n1302);
or (n1432,n1433,n1434);
and (n1433,n1348,n1353);
and (n1434,n1349,n1352);
and (n1435,n1431,n1432);
nand (n1436,n1304,n1437);
and (n1437,n1254,n1280);
nand (n1438,n1305,n1306);
and (n1439,n1213,n1248);
and (n1440,n1090,n1195);
or (n1441,n1442,n1449);
xor (n1442,n1443,n1448);
xor (n1443,n1444,n1445);
xor (n1444,n977,n997);
or (n1445,n1446,n1447);
and (n1446,n1202,n1209);
and (n1447,n1203,n1206);
xor (n1448,n1059,n1062);
or (n1449,n1450,n1451);
and (n1450,n1196,n1201);
and (n1451,n1197,n1198);
nor (n1452,n1453,n1454);
xor (n1453,n1056,n1081);
or (n1454,n1455,n1456);
and (n1455,n1443,n1448);
and (n1456,n1444,n1445);
or (n1457,n1452,n1458);
nand (n1458,n1442,n1449);
nand (n1459,n1453,n1454);
and (n1460,n1054,n1083);
and (n1461,n809,n1022);
nor (n1462,n1463,n1488);
nor (n1463,n1464,n1479);
xor (n1464,n1465,n1478);
xor (n1465,n1466,n1467);
xor (n1466,n605,n624);
or (n1467,n1468,n1477);
and (n1468,n1469,n1476);
xor (n1469,n1470,n1473);
or (n1470,n1471,n1472);
and (n1471,n1043,n1048);
and (n1472,n1044,n1047);
or (n1473,n1474,n1475);
and (n1474,n1025,n1032);
and (n1475,n1026,n1029);
xor (n1476,n729,n744);
and (n1477,n1470,n1473);
xor (n1478,n726,n768);
or (n1479,n1480,n1487);
and (n1480,n1481,n1486);
xor (n1481,n1482,n1483);
xor (n1482,n770,n794);
or (n1483,n1484,n1485);
and (n1484,n1037,n1042);
and (n1485,n1038,n1039);
xor (n1486,n1469,n1476);
and (n1487,n1482,n1483);
nor (n1488,n1489,n1490);
xor (n1489,n1481,n1486);
or (n1490,n1491,n1492);
and (n1491,n1023,n1036);
and (n1492,n1024,n1033);
nand (n1493,n1494,n1496);
or (n1494,n1463,n1495);
nand (n1495,n1489,n1490);
nand (n1496,n1464,n1479);
nor (n1497,n1498,n1501);
or (n1498,n1499,n1500);
and (n1499,n1465,n1478);
and (n1500,n1466,n1467);
xor (n1501,n722,n797);
not (n1502,n1503);
and (n1503,n1498,n1501);
or (n1504,n801,n3);
xor (n1505,n1506,n2522);
xor (n1506,n1507,n2520);
xor (n1507,n1508,n2519);
xor (n1508,n1509,n2510);
xor (n1509,n1510,n2509);
xor (n1510,n1511,n2495);
xor (n1511,n1512,n2494);
xor (n1512,n1513,n2473);
xor (n1513,n1514,n2472);
xor (n1514,n1515,n2446);
xor (n1515,n1516,n2445);
xor (n1516,n1517,n2412);
xor (n1517,n1518,n2411);
xor (n1518,n1519,n2373);
xor (n1519,n1520,n2372);
xor (n1520,n1521,n2327);
xor (n1521,n1522,n2326);
xor (n1522,n1523,n2276);
xor (n1523,n1524,n2275);
xor (n1524,n1525,n2218);
xor (n1525,n1526,n2217);
xor (n1526,n1527,n2155);
xor (n1527,n1528,n2154);
xor (n1528,n1529,n2086);
xor (n1529,n1530,n2085);
xor (n1530,n1531,n2011);
xor (n1531,n1532,n2010);
xor (n1532,n1533,n1929);
xor (n1533,n1534,n1928);
xor (n1534,n1535,n1842);
xor (n1535,n1536,n1841);
xor (n1536,n1537,n1748);
xor (n1537,n1538,n1747);
xor (n1538,n1539,n1649);
xor (n1539,n1540,n1648);
xor (n1540,n1541,n1544);
xor (n1541,n1542,n1543);
and (n1542,n413,n288);
and (n1543,n402,n281);
or (n1544,n1545,n1548);
and (n1545,n1546,n1547);
and (n1546,n402,n288);
and (n1547,n292,n281);
and (n1548,n1549,n1550);
xor (n1549,n1546,n1547);
or (n1550,n1551,n1554);
and (n1551,n1552,n1553);
and (n1552,n292,n288);
and (n1553,n256,n281);
and (n1554,n1555,n1556);
xor (n1555,n1552,n1553);
or (n1556,n1557,n1560);
and (n1557,n1558,n1559);
and (n1558,n256,n288);
and (n1559,n477,n281);
and (n1560,n1561,n1562);
xor (n1561,n1558,n1559);
or (n1562,n1563,n1566);
and (n1563,n1564,n1565);
and (n1564,n477,n288);
and (n1565,n515,n281);
and (n1566,n1567,n1568);
xor (n1567,n1564,n1565);
or (n1568,n1569,n1572);
and (n1569,n1570,n1571);
and (n1570,n515,n288);
and (n1571,n507,n281);
and (n1572,n1573,n1574);
xor (n1573,n1570,n1571);
or (n1574,n1575,n1578);
and (n1575,n1576,n1577);
and (n1576,n507,n288);
and (n1577,n432,n281);
and (n1578,n1579,n1580);
xor (n1579,n1576,n1577);
or (n1580,n1581,n1584);
and (n1581,n1582,n1583);
and (n1582,n432,n288);
and (n1583,n334,n281);
and (n1584,n1585,n1586);
xor (n1585,n1582,n1583);
or (n1586,n1587,n1590);
and (n1587,n1588,n1589);
and (n1588,n334,n288);
and (n1589,n326,n281);
and (n1590,n1591,n1592);
xor (n1591,n1588,n1589);
or (n1592,n1593,n1596);
and (n1593,n1594,n1595);
and (n1594,n326,n288);
and (n1595,n124,n281);
and (n1596,n1597,n1598);
xor (n1597,n1594,n1595);
or (n1598,n1599,n1602);
and (n1599,n1600,n1601);
and (n1600,n124,n288);
and (n1601,n89,n281);
and (n1602,n1603,n1604);
xor (n1603,n1600,n1601);
or (n1604,n1605,n1608);
and (n1605,n1606,n1607);
and (n1606,n89,n288);
and (n1607,n165,n281);
and (n1608,n1609,n1610);
xor (n1609,n1606,n1607);
or (n1610,n1611,n1614);
and (n1611,n1612,n1613);
and (n1612,n165,n288);
and (n1613,n157,n281);
and (n1614,n1615,n1616);
xor (n1615,n1612,n1613);
or (n1616,n1617,n1620);
and (n1617,n1618,n1619);
and (n1618,n157,n288);
and (n1619,n231,n281);
and (n1620,n1621,n1622);
xor (n1621,n1618,n1619);
or (n1622,n1623,n1626);
and (n1623,n1624,n1625);
and (n1624,n231,n288);
and (n1625,n447,n281);
and (n1626,n1627,n1628);
xor (n1627,n1624,n1625);
or (n1628,n1629,n1632);
and (n1629,n1630,n1631);
and (n1630,n447,n288);
and (n1631,n364,n281);
and (n1632,n1633,n1634);
xor (n1633,n1630,n1631);
or (n1634,n1635,n1638);
and (n1635,n1636,n1637);
and (n1636,n364,n288);
and (n1637,n355,n281);
and (n1638,n1639,n1640);
xor (n1639,n1636,n1637);
or (n1640,n1641,n1643);
and (n1641,n1642,n1413);
and (n1642,n355,n288);
and (n1643,n1644,n1645);
xor (n1644,n1642,n1413);
and (n1645,n1646,n1647);
and (n1646,n219,n288);
and (n1647,n213,n281);
and (n1648,n292,n463);
or (n1649,n1650,n1653);
and (n1650,n1651,n1652);
xor (n1651,n1549,n1550);
and (n1652,n256,n463);
and (n1653,n1654,n1655);
xor (n1654,n1651,n1652);
or (n1655,n1656,n1659);
and (n1656,n1657,n1658);
xor (n1657,n1555,n1556);
and (n1658,n477,n463);
and (n1659,n1660,n1661);
xor (n1660,n1657,n1658);
or (n1661,n1662,n1665);
and (n1662,n1663,n1664);
xor (n1663,n1561,n1562);
and (n1664,n515,n463);
and (n1665,n1666,n1667);
xor (n1666,n1663,n1664);
or (n1667,n1668,n1671);
and (n1668,n1669,n1670);
xor (n1669,n1567,n1568);
and (n1670,n507,n463);
and (n1671,n1672,n1673);
xor (n1672,n1669,n1670);
or (n1673,n1674,n1677);
and (n1674,n1675,n1676);
xor (n1675,n1573,n1574);
and (n1676,n432,n463);
and (n1677,n1678,n1679);
xor (n1678,n1675,n1676);
or (n1679,n1680,n1683);
and (n1680,n1681,n1682);
xor (n1681,n1579,n1580);
and (n1682,n334,n463);
and (n1683,n1684,n1685);
xor (n1684,n1681,n1682);
or (n1685,n1686,n1689);
and (n1686,n1687,n1688);
xor (n1687,n1585,n1586);
and (n1688,n326,n463);
and (n1689,n1690,n1691);
xor (n1690,n1687,n1688);
or (n1691,n1692,n1695);
and (n1692,n1693,n1694);
xor (n1693,n1591,n1592);
and (n1694,n124,n463);
and (n1695,n1696,n1697);
xor (n1696,n1693,n1694);
or (n1697,n1698,n1701);
and (n1698,n1699,n1700);
xor (n1699,n1597,n1598);
and (n1700,n89,n463);
and (n1701,n1702,n1703);
xor (n1702,n1699,n1700);
or (n1703,n1704,n1707);
and (n1704,n1705,n1706);
xor (n1705,n1603,n1604);
and (n1706,n165,n463);
and (n1707,n1708,n1709);
xor (n1708,n1705,n1706);
or (n1709,n1710,n1713);
and (n1710,n1711,n1712);
xor (n1711,n1609,n1610);
and (n1712,n157,n463);
and (n1713,n1714,n1715);
xor (n1714,n1711,n1712);
or (n1715,n1716,n1719);
and (n1716,n1717,n1718);
xor (n1717,n1615,n1616);
and (n1718,n231,n463);
and (n1719,n1720,n1721);
xor (n1720,n1717,n1718);
or (n1721,n1722,n1725);
and (n1722,n1723,n1724);
xor (n1723,n1621,n1622);
and (n1724,n447,n463);
and (n1725,n1726,n1727);
xor (n1726,n1723,n1724);
or (n1727,n1728,n1731);
and (n1728,n1729,n1730);
xor (n1729,n1627,n1628);
and (n1730,n364,n463);
and (n1731,n1732,n1733);
xor (n1732,n1729,n1730);
or (n1733,n1734,n1737);
and (n1734,n1735,n1736);
xor (n1735,n1633,n1634);
and (n1736,n355,n463);
and (n1737,n1738,n1739);
xor (n1738,n1735,n1736);
or (n1739,n1740,n1743);
and (n1740,n1741,n1742);
xor (n1741,n1639,n1640);
and (n1742,n219,n463);
and (n1743,n1744,n1745);
xor (n1744,n1741,n1742);
and (n1745,n1746,n1384);
xor (n1746,n1644,n1645);
and (n1747,n256,n471);
or (n1748,n1749,n1752);
and (n1749,n1750,n1751);
xor (n1750,n1654,n1655);
and (n1751,n477,n471);
and (n1752,n1753,n1754);
xor (n1753,n1750,n1751);
or (n1754,n1755,n1758);
and (n1755,n1756,n1757);
xor (n1756,n1660,n1661);
and (n1757,n515,n471);
and (n1758,n1759,n1760);
xor (n1759,n1756,n1757);
or (n1760,n1761,n1764);
and (n1761,n1762,n1763);
xor (n1762,n1666,n1667);
and (n1763,n507,n471);
and (n1764,n1765,n1766);
xor (n1765,n1762,n1763);
or (n1766,n1767,n1770);
and (n1767,n1768,n1769);
xor (n1768,n1672,n1673);
and (n1769,n432,n471);
and (n1770,n1771,n1772);
xor (n1771,n1768,n1769);
or (n1772,n1773,n1776);
and (n1773,n1774,n1775);
xor (n1774,n1678,n1679);
and (n1775,n334,n471);
and (n1776,n1777,n1778);
xor (n1777,n1774,n1775);
or (n1778,n1779,n1782);
and (n1779,n1780,n1781);
xor (n1780,n1684,n1685);
and (n1781,n326,n471);
and (n1782,n1783,n1784);
xor (n1783,n1780,n1781);
or (n1784,n1785,n1788);
and (n1785,n1786,n1787);
xor (n1786,n1690,n1691);
and (n1787,n124,n471);
and (n1788,n1789,n1790);
xor (n1789,n1786,n1787);
or (n1790,n1791,n1794);
and (n1791,n1792,n1793);
xor (n1792,n1696,n1697);
and (n1793,n89,n471);
and (n1794,n1795,n1796);
xor (n1795,n1792,n1793);
or (n1796,n1797,n1800);
and (n1797,n1798,n1799);
xor (n1798,n1702,n1703);
and (n1799,n165,n471);
and (n1800,n1801,n1802);
xor (n1801,n1798,n1799);
or (n1802,n1803,n1806);
and (n1803,n1804,n1805);
xor (n1804,n1708,n1709);
and (n1805,n157,n471);
and (n1806,n1807,n1808);
xor (n1807,n1804,n1805);
or (n1808,n1809,n1812);
and (n1809,n1810,n1811);
xor (n1810,n1714,n1715);
and (n1811,n231,n471);
and (n1812,n1813,n1814);
xor (n1813,n1810,n1811);
or (n1814,n1815,n1818);
and (n1815,n1816,n1817);
xor (n1816,n1720,n1721);
and (n1817,n447,n471);
and (n1818,n1819,n1820);
xor (n1819,n1816,n1817);
or (n1820,n1821,n1824);
and (n1821,n1822,n1823);
xor (n1822,n1726,n1727);
and (n1823,n364,n471);
and (n1824,n1825,n1826);
xor (n1825,n1822,n1823);
or (n1826,n1827,n1830);
and (n1827,n1828,n1829);
xor (n1828,n1732,n1733);
and (n1829,n355,n471);
and (n1830,n1831,n1832);
xor (n1831,n1828,n1829);
or (n1832,n1833,n1836);
and (n1833,n1834,n1835);
xor (n1834,n1738,n1739);
and (n1835,n219,n471);
and (n1836,n1837,n1838);
xor (n1837,n1834,n1835);
and (n1838,n1839,n1840);
xor (n1839,n1744,n1745);
and (n1840,n213,n471);
and (n1841,n477,n530);
or (n1842,n1843,n1846);
and (n1843,n1844,n1845);
xor (n1844,n1753,n1754);
and (n1845,n515,n530);
and (n1846,n1847,n1848);
xor (n1847,n1844,n1845);
or (n1848,n1849,n1852);
and (n1849,n1850,n1851);
xor (n1850,n1759,n1760);
and (n1851,n507,n530);
and (n1852,n1853,n1854);
xor (n1853,n1850,n1851);
or (n1854,n1855,n1858);
and (n1855,n1856,n1857);
xor (n1856,n1765,n1766);
and (n1857,n432,n530);
and (n1858,n1859,n1860);
xor (n1859,n1856,n1857);
or (n1860,n1861,n1864);
and (n1861,n1862,n1863);
xor (n1862,n1771,n1772);
and (n1863,n334,n530);
and (n1864,n1865,n1866);
xor (n1865,n1862,n1863);
or (n1866,n1867,n1870);
and (n1867,n1868,n1869);
xor (n1868,n1777,n1778);
and (n1869,n326,n530);
and (n1870,n1871,n1872);
xor (n1871,n1868,n1869);
or (n1872,n1873,n1876);
and (n1873,n1874,n1875);
xor (n1874,n1783,n1784);
and (n1875,n124,n530);
and (n1876,n1877,n1878);
xor (n1877,n1874,n1875);
or (n1878,n1879,n1882);
and (n1879,n1880,n1881);
xor (n1880,n1789,n1790);
and (n1881,n89,n530);
and (n1882,n1883,n1884);
xor (n1883,n1880,n1881);
or (n1884,n1885,n1888);
and (n1885,n1886,n1887);
xor (n1886,n1795,n1796);
and (n1887,n165,n530);
and (n1888,n1889,n1890);
xor (n1889,n1886,n1887);
or (n1890,n1891,n1894);
and (n1891,n1892,n1893);
xor (n1892,n1801,n1802);
and (n1893,n157,n530);
and (n1894,n1895,n1896);
xor (n1895,n1892,n1893);
or (n1896,n1897,n1900);
and (n1897,n1898,n1899);
xor (n1898,n1807,n1808);
and (n1899,n231,n530);
and (n1900,n1901,n1902);
xor (n1901,n1898,n1899);
or (n1902,n1903,n1906);
and (n1903,n1904,n1905);
xor (n1904,n1813,n1814);
and (n1905,n447,n530);
and (n1906,n1907,n1908);
xor (n1907,n1904,n1905);
or (n1908,n1909,n1912);
and (n1909,n1910,n1911);
xor (n1910,n1819,n1820);
and (n1911,n364,n530);
and (n1912,n1913,n1914);
xor (n1913,n1910,n1911);
or (n1914,n1915,n1918);
and (n1915,n1916,n1917);
xor (n1916,n1825,n1826);
and (n1917,n355,n530);
and (n1918,n1919,n1920);
xor (n1919,n1916,n1917);
or (n1920,n1921,n1924);
and (n1921,n1922,n1923);
xor (n1922,n1831,n1832);
and (n1923,n219,n530);
and (n1924,n1925,n1926);
xor (n1925,n1922,n1923);
and (n1926,n1927,n1337);
xor (n1927,n1837,n1838);
and (n1928,n515,n308);
or (n1929,n1930,n1933);
and (n1930,n1931,n1932);
xor (n1931,n1847,n1848);
and (n1932,n507,n308);
and (n1933,n1934,n1935);
xor (n1934,n1931,n1932);
or (n1935,n1936,n1939);
and (n1936,n1937,n1938);
xor (n1937,n1853,n1854);
and (n1938,n432,n308);
and (n1939,n1940,n1941);
xor (n1940,n1937,n1938);
or (n1941,n1942,n1945);
and (n1942,n1943,n1944);
xor (n1943,n1859,n1860);
and (n1944,n334,n308);
and (n1945,n1946,n1947);
xor (n1946,n1943,n1944);
or (n1947,n1948,n1951);
and (n1948,n1949,n1950);
xor (n1949,n1865,n1866);
and (n1950,n326,n308);
and (n1951,n1952,n1953);
xor (n1952,n1949,n1950);
or (n1953,n1954,n1957);
and (n1954,n1955,n1956);
xor (n1955,n1871,n1872);
and (n1956,n124,n308);
and (n1957,n1958,n1959);
xor (n1958,n1955,n1956);
or (n1959,n1960,n1963);
and (n1960,n1961,n1962);
xor (n1961,n1877,n1878);
and (n1962,n89,n308);
and (n1963,n1964,n1965);
xor (n1964,n1961,n1962);
or (n1965,n1966,n1969);
and (n1966,n1967,n1968);
xor (n1967,n1883,n1884);
and (n1968,n165,n308);
and (n1969,n1970,n1971);
xor (n1970,n1967,n1968);
or (n1971,n1972,n1975);
and (n1972,n1973,n1974);
xor (n1973,n1889,n1890);
and (n1974,n157,n308);
and (n1975,n1976,n1977);
xor (n1976,n1973,n1974);
or (n1977,n1978,n1981);
and (n1978,n1979,n1980);
xor (n1979,n1895,n1896);
and (n1980,n231,n308);
and (n1981,n1982,n1983);
xor (n1982,n1979,n1980);
or (n1983,n1984,n1987);
and (n1984,n1985,n1986);
xor (n1985,n1901,n1902);
and (n1986,n447,n308);
and (n1987,n1988,n1989);
xor (n1988,n1985,n1986);
or (n1989,n1990,n1993);
and (n1990,n1991,n1992);
xor (n1991,n1907,n1908);
and (n1992,n364,n308);
and (n1993,n1994,n1995);
xor (n1994,n1991,n1992);
or (n1995,n1996,n1999);
and (n1996,n1997,n1998);
xor (n1997,n1913,n1914);
and (n1998,n355,n308);
and (n1999,n2000,n2001);
xor (n2000,n1997,n1998);
or (n2001,n2002,n2005);
and (n2002,n2003,n2004);
xor (n2003,n1919,n1920);
and (n2004,n219,n308);
and (n2005,n2006,n2007);
xor (n2006,n2003,n2004);
and (n2007,n2008,n2009);
xor (n2008,n1925,n1926);
and (n2009,n213,n308);
and (n2010,n507,n311);
or (n2011,n2012,n2015);
and (n2012,n2013,n2014);
xor (n2013,n1934,n1935);
and (n2014,n432,n311);
and (n2015,n2016,n2017);
xor (n2016,n2013,n2014);
or (n2017,n2018,n2021);
and (n2018,n2019,n2020);
xor (n2019,n1940,n1941);
and (n2020,n334,n311);
and (n2021,n2022,n2023);
xor (n2022,n2019,n2020);
or (n2023,n2024,n2027);
and (n2024,n2025,n2026);
xor (n2025,n1946,n1947);
and (n2026,n326,n311);
and (n2027,n2028,n2029);
xor (n2028,n2025,n2026);
or (n2029,n2030,n2033);
and (n2030,n2031,n2032);
xor (n2031,n1952,n1953);
and (n2032,n124,n311);
and (n2033,n2034,n2035);
xor (n2034,n2031,n2032);
or (n2035,n2036,n2039);
and (n2036,n2037,n2038);
xor (n2037,n1958,n1959);
and (n2038,n89,n311);
and (n2039,n2040,n2041);
xor (n2040,n2037,n2038);
or (n2041,n2042,n2045);
and (n2042,n2043,n2044);
xor (n2043,n1964,n1965);
and (n2044,n165,n311);
and (n2045,n2046,n2047);
xor (n2046,n2043,n2044);
or (n2047,n2048,n2051);
and (n2048,n2049,n2050);
xor (n2049,n1970,n1971);
and (n2050,n157,n311);
and (n2051,n2052,n2053);
xor (n2052,n2049,n2050);
or (n2053,n2054,n2057);
and (n2054,n2055,n2056);
xor (n2055,n1976,n1977);
and (n2056,n231,n311);
and (n2057,n2058,n2059);
xor (n2058,n2055,n2056);
or (n2059,n2060,n2063);
and (n2060,n2061,n2062);
xor (n2061,n1982,n1983);
and (n2062,n447,n311);
and (n2063,n2064,n2065);
xor (n2064,n2061,n2062);
or (n2065,n2066,n2069);
and (n2066,n2067,n2068);
xor (n2067,n1988,n1989);
and (n2068,n364,n311);
and (n2069,n2070,n2071);
xor (n2070,n2067,n2068);
or (n2071,n2072,n2075);
and (n2072,n2073,n2074);
xor (n2073,n1994,n1995);
and (n2074,n355,n311);
and (n2075,n2076,n2077);
xor (n2076,n2073,n2074);
or (n2077,n2078,n2081);
and (n2078,n2079,n2080);
xor (n2079,n2000,n2001);
and (n2080,n219,n311);
and (n2081,n2082,n2083);
xor (n2082,n2079,n2080);
and (n2083,n2084,n1236);
xor (n2084,n2006,n2007);
and (n2085,n432,n319);
or (n2086,n2087,n2090);
and (n2087,n2088,n2089);
xor (n2088,n2016,n2017);
and (n2089,n334,n319);
and (n2090,n2091,n2092);
xor (n2091,n2088,n2089);
or (n2092,n2093,n2096);
and (n2093,n2094,n2095);
xor (n2094,n2022,n2023);
and (n2095,n326,n319);
and (n2096,n2097,n2098);
xor (n2097,n2094,n2095);
or (n2098,n2099,n2102);
and (n2099,n2100,n2101);
xor (n2100,n2028,n2029);
and (n2101,n124,n319);
and (n2102,n2103,n2104);
xor (n2103,n2100,n2101);
or (n2104,n2105,n2108);
and (n2105,n2106,n2107);
xor (n2106,n2034,n2035);
and (n2107,n89,n319);
and (n2108,n2109,n2110);
xor (n2109,n2106,n2107);
or (n2110,n2111,n2114);
and (n2111,n2112,n2113);
xor (n2112,n2040,n2041);
and (n2113,n165,n319);
and (n2114,n2115,n2116);
xor (n2115,n2112,n2113);
or (n2116,n2117,n2120);
and (n2117,n2118,n2119);
xor (n2118,n2046,n2047);
and (n2119,n157,n319);
and (n2120,n2121,n2122);
xor (n2121,n2118,n2119);
or (n2122,n2123,n2126);
and (n2123,n2124,n2125);
xor (n2124,n2052,n2053);
and (n2125,n231,n319);
and (n2126,n2127,n2128);
xor (n2127,n2124,n2125);
or (n2128,n2129,n2132);
and (n2129,n2130,n2131);
xor (n2130,n2058,n2059);
and (n2131,n447,n319);
and (n2132,n2133,n2134);
xor (n2133,n2130,n2131);
or (n2134,n2135,n2137);
and (n2135,n2136,n1100);
xor (n2136,n2064,n2065);
and (n2137,n2138,n2139);
xor (n2138,n2136,n1100);
or (n2139,n2140,n2143);
and (n2140,n2141,n2142);
xor (n2141,n2070,n2071);
and (n2142,n355,n319);
and (n2143,n2144,n2145);
xor (n2144,n2141,n2142);
or (n2145,n2146,n2149);
and (n2146,n2147,n2148);
xor (n2147,n2076,n2077);
and (n2148,n219,n319);
and (n2149,n2150,n2151);
xor (n2150,n2147,n2148);
and (n2151,n2152,n2153);
xor (n2152,n2082,n2083);
and (n2153,n213,n319);
and (n2154,n334,n585);
or (n2155,n2156,n2159);
and (n2156,n2157,n2158);
xor (n2157,n2091,n2092);
and (n2158,n326,n585);
and (n2159,n2160,n2161);
xor (n2160,n2157,n2158);
or (n2161,n2162,n2165);
and (n2162,n2163,n2164);
xor (n2163,n2097,n2098);
and (n2164,n124,n585);
and (n2165,n2166,n2167);
xor (n2166,n2163,n2164);
or (n2167,n2168,n2171);
and (n2168,n2169,n2170);
xor (n2169,n2103,n2104);
and (n2170,n89,n585);
and (n2171,n2172,n2173);
xor (n2172,n2169,n2170);
or (n2173,n2174,n2177);
and (n2174,n2175,n2176);
xor (n2175,n2109,n2110);
and (n2176,n165,n585);
and (n2177,n2178,n2179);
xor (n2178,n2175,n2176);
or (n2179,n2180,n2183);
and (n2180,n2181,n2182);
xor (n2181,n2115,n2116);
and (n2182,n157,n585);
and (n2183,n2184,n2185);
xor (n2184,n2181,n2182);
or (n2185,n2186,n2189);
and (n2186,n2187,n2188);
xor (n2187,n2121,n2122);
and (n2188,n231,n585);
and (n2189,n2190,n2191);
xor (n2190,n2187,n2188);
or (n2191,n2192,n2195);
and (n2192,n2193,n2194);
xor (n2193,n2127,n2128);
and (n2194,n447,n585);
and (n2195,n2196,n2197);
xor (n2196,n2193,n2194);
or (n2197,n2198,n2201);
and (n2198,n2199,n2200);
xor (n2199,n2133,n2134);
and (n2200,n364,n585);
and (n2201,n2202,n2203);
xor (n2202,n2199,n2200);
or (n2203,n2204,n2207);
and (n2204,n2205,n2206);
xor (n2205,n2138,n2139);
and (n2206,n355,n585);
and (n2207,n2208,n2209);
xor (n2208,n2205,n2206);
or (n2209,n2210,n2213);
and (n2210,n2211,n2212);
xor (n2211,n2144,n2145);
and (n2212,n219,n585);
and (n2213,n2214,n2215);
xor (n2214,n2211,n2212);
and (n2215,n2216,n1129);
xor (n2216,n2150,n2151);
and (n2217,n326,n71);
or (n2218,n2219,n2222);
and (n2219,n2220,n2221);
xor (n2220,n2160,n2161);
and (n2221,n124,n71);
and (n2222,n2223,n2224);
xor (n2223,n2220,n2221);
or (n2224,n2225,n2228);
and (n2225,n2226,n2227);
xor (n2226,n2166,n2167);
and (n2227,n89,n71);
and (n2228,n2229,n2230);
xor (n2229,n2226,n2227);
or (n2230,n2231,n2234);
and (n2231,n2232,n2233);
xor (n2232,n2172,n2173);
and (n2233,n165,n71);
and (n2234,n2235,n2236);
xor (n2235,n2232,n2233);
or (n2236,n2237,n2240);
and (n2237,n2238,n2239);
xor (n2238,n2178,n2179);
and (n2239,n157,n71);
and (n2240,n2241,n2242);
xor (n2241,n2238,n2239);
or (n2242,n2243,n2246);
and (n2243,n2244,n2245);
xor (n2244,n2184,n2185);
and (n2245,n231,n71);
and (n2246,n2247,n2248);
xor (n2247,n2244,n2245);
or (n2248,n2249,n2252);
and (n2249,n2250,n2251);
xor (n2250,n2190,n2191);
and (n2251,n447,n71);
and (n2252,n2253,n2254);
xor (n2253,n2250,n2251);
or (n2254,n2255,n2258);
and (n2255,n2256,n2257);
xor (n2256,n2196,n2197);
and (n2257,n364,n71);
and (n2258,n2259,n2260);
xor (n2259,n2256,n2257);
or (n2260,n2261,n2264);
and (n2261,n2262,n2263);
xor (n2262,n2202,n2203);
and (n2263,n355,n71);
and (n2264,n2265,n2266);
xor (n2265,n2262,n2263);
or (n2266,n2267,n2270);
and (n2267,n2268,n2269);
xor (n2268,n2208,n2209);
and (n2269,n219,n71);
and (n2270,n2271,n2272);
xor (n2271,n2268,n2269);
and (n2272,n2273,n2274);
xor (n2273,n2214,n2215);
and (n2274,n213,n71);
and (n2275,n124,n17);
or (n2276,n2277,n2280);
and (n2277,n2278,n2279);
xor (n2278,n2223,n2224);
and (n2279,n89,n17);
and (n2280,n2281,n2282);
xor (n2281,n2278,n2279);
or (n2282,n2283,n2286);
and (n2283,n2284,n2285);
xor (n2284,n2229,n2230);
and (n2285,n165,n17);
and (n2286,n2287,n2288);
xor (n2287,n2284,n2285);
or (n2288,n2289,n2292);
and (n2289,n2290,n2291);
xor (n2290,n2235,n2236);
and (n2291,n157,n17);
and (n2292,n2293,n2294);
xor (n2293,n2290,n2291);
or (n2294,n2295,n2298);
and (n2295,n2296,n2297);
xor (n2296,n2241,n2242);
and (n2297,n231,n17);
and (n2298,n2299,n2300);
xor (n2299,n2296,n2297);
or (n2300,n2301,n2304);
and (n2301,n2302,n2303);
xor (n2302,n2247,n2248);
and (n2303,n447,n17);
and (n2304,n2305,n2306);
xor (n2305,n2302,n2303);
or (n2306,n2307,n2310);
and (n2307,n2308,n2309);
xor (n2308,n2253,n2254);
and (n2309,n364,n17);
and (n2310,n2311,n2312);
xor (n2311,n2308,n2309);
or (n2312,n2313,n2316);
and (n2313,n2314,n2315);
xor (n2314,n2259,n2260);
and (n2315,n355,n17);
and (n2316,n2317,n2318);
xor (n2317,n2314,n2315);
or (n2318,n2319,n2322);
and (n2319,n2320,n2321);
xor (n2320,n2265,n2266);
and (n2321,n219,n17);
and (n2322,n2323,n2324);
xor (n2323,n2320,n2321);
and (n2324,n2325,n995);
xor (n2325,n2271,n2272);
and (n2326,n89,n79);
or (n2327,n2328,n2331);
and (n2328,n2329,n2330);
xor (n2329,n2281,n2282);
and (n2330,n165,n79);
and (n2331,n2332,n2333);
xor (n2332,n2329,n2330);
or (n2333,n2334,n2337);
and (n2334,n2335,n2336);
xor (n2335,n2287,n2288);
and (n2336,n157,n79);
and (n2337,n2338,n2339);
xor (n2338,n2335,n2336);
or (n2339,n2340,n2343);
and (n2340,n2341,n2342);
xor (n2341,n2293,n2294);
and (n2342,n231,n79);
and (n2343,n2344,n2345);
xor (n2344,n2341,n2342);
or (n2345,n2346,n2349);
and (n2346,n2347,n2348);
xor (n2347,n2299,n2300);
and (n2348,n447,n79);
and (n2349,n2350,n2351);
xor (n2350,n2347,n2348);
or (n2351,n2352,n2355);
and (n2352,n2353,n2354);
xor (n2353,n2305,n2306);
and (n2354,n364,n79);
and (n2355,n2356,n2357);
xor (n2356,n2353,n2354);
or (n2357,n2358,n2361);
and (n2358,n2359,n2360);
xor (n2359,n2311,n2312);
and (n2360,n355,n79);
and (n2361,n2362,n2363);
xor (n2362,n2359,n2360);
or (n2363,n2364,n2367);
and (n2364,n2365,n2366);
xor (n2365,n2317,n2318);
and (n2366,n219,n79);
and (n2367,n2368,n2369);
xor (n2368,n2365,n2366);
and (n2369,n2370,n2371);
xor (n2370,n2323,n2324);
and (n2371,n213,n79);
and (n2372,n165,n147);
or (n2373,n2374,n2377);
and (n2374,n2375,n2376);
xor (n2375,n2332,n2333);
and (n2376,n157,n147);
and (n2377,n2378,n2379);
xor (n2378,n2375,n2376);
or (n2379,n2380,n2383);
and (n2380,n2381,n2382);
xor (n2381,n2338,n2339);
and (n2382,n231,n147);
and (n2383,n2384,n2385);
xor (n2384,n2381,n2382);
or (n2385,n2386,n2389);
and (n2386,n2387,n2388);
xor (n2387,n2344,n2345);
and (n2388,n447,n147);
and (n2389,n2390,n2391);
xor (n2390,n2387,n2388);
or (n2391,n2392,n2395);
and (n2392,n2393,n2394);
xor (n2393,n2350,n2351);
and (n2394,n364,n147);
and (n2395,n2396,n2397);
xor (n2396,n2393,n2394);
or (n2397,n2398,n2401);
and (n2398,n2399,n2400);
xor (n2399,n2356,n2357);
and (n2400,n355,n147);
and (n2401,n2402,n2403);
xor (n2402,n2399,n2400);
or (n2403,n2404,n2407);
and (n2404,n2405,n2406);
xor (n2405,n2362,n2363);
and (n2406,n219,n147);
and (n2407,n2408,n2409);
xor (n2408,n2405,n2406);
and (n2409,n2410,n913);
xor (n2410,n2368,n2369);
and (n2411,n157,n138);
or (n2412,n2413,n2416);
and (n2413,n2414,n2415);
xor (n2414,n2378,n2379);
and (n2415,n231,n138);
and (n2416,n2417,n2418);
xor (n2417,n2414,n2415);
or (n2418,n2419,n2422);
and (n2419,n2420,n2421);
xor (n2420,n2384,n2385);
and (n2421,n447,n138);
and (n2422,n2423,n2424);
xor (n2423,n2420,n2421);
or (n2424,n2425,n2428);
and (n2425,n2426,n2427);
xor (n2426,n2390,n2391);
and (n2427,n364,n138);
and (n2428,n2429,n2430);
xor (n2429,n2426,n2427);
or (n2430,n2431,n2434);
and (n2431,n2432,n2433);
xor (n2432,n2396,n2397);
and (n2433,n355,n138);
and (n2434,n2435,n2436);
xor (n2435,n2432,n2433);
or (n2436,n2437,n2440);
and (n2437,n2438,n2439);
xor (n2438,n2402,n2403);
and (n2439,n219,n138);
and (n2440,n2441,n2442);
xor (n2441,n2438,n2439);
and (n2442,n2443,n2444);
xor (n2443,n2408,n2409);
and (n2444,n213,n138);
and (n2445,n231,n345);
or (n2446,n2447,n2450);
and (n2447,n2448,n2449);
xor (n2448,n2417,n2418);
and (n2449,n447,n345);
and (n2450,n2451,n2452);
xor (n2451,n2448,n2449);
or (n2452,n2453,n2456);
and (n2453,n2454,n2455);
xor (n2454,n2423,n2424);
and (n2455,n364,n345);
and (n2456,n2457,n2458);
xor (n2457,n2454,n2455);
or (n2458,n2459,n2462);
and (n2459,n2460,n2461);
xor (n2460,n2429,n2430);
and (n2461,n355,n345);
and (n2462,n2463,n2464);
xor (n2463,n2460,n2461);
or (n2464,n2465,n2468);
and (n2465,n2466,n2467);
xor (n2466,n2435,n2436);
and (n2467,n219,n345);
and (n2468,n2469,n2470);
xor (n2469,n2466,n2467);
and (n2470,n2471,n741);
xor (n2471,n2441,n2442);
and (n2472,n447,n242);
or (n2473,n2474,n2477);
and (n2474,n2475,n2476);
xor (n2475,n2451,n2452);
and (n2476,n364,n242);
and (n2477,n2478,n2479);
xor (n2478,n2475,n2476);
or (n2479,n2480,n2483);
and (n2480,n2481,n2482);
xor (n2481,n2457,n2458);
and (n2482,n355,n242);
and (n2483,n2484,n2485);
xor (n2484,n2481,n2482);
or (n2485,n2486,n2489);
and (n2486,n2487,n2488);
xor (n2487,n2463,n2464);
and (n2488,n219,n242);
and (n2489,n2490,n2491);
xor (n2490,n2487,n2488);
and (n2491,n2492,n2493);
xor (n2492,n2469,n2470);
and (n2493,n213,n242);
and (n2494,n364,n247);
or (n2495,n2496,n2499);
and (n2496,n2497,n2498);
xor (n2497,n2478,n2479);
and (n2498,n355,n247);
and (n2499,n2500,n2501);
xor (n2500,n2497,n2498);
or (n2501,n2502,n2505);
and (n2502,n2503,n2504);
xor (n2503,n2484,n2485);
and (n2504,n219,n247);
and (n2505,n2506,n2507);
xor (n2506,n2503,n2504);
and (n2507,n2508,n246);
xor (n2508,n2490,n2491);
and (n2509,n355,n194);
or (n2510,n2511,n2514);
and (n2511,n2512,n2513);
xor (n2512,n2500,n2501);
and (n2513,n219,n194);
and (n2514,n2515,n2516);
xor (n2515,n2512,n2513);
and (n2516,n2517,n2518);
xor (n2517,n2506,n2507);
and (n2518,n213,n194);
and (n2519,n219,n176);
and (n2520,n2521,n396);
xor (n2521,n2515,n2516);
and (n2522,n213,n203);
endmodule
