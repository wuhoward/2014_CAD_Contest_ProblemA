module top (out,n3,n22,n25,n26,n34,n35,n41,n42,n47
        ,n55,n57,n58,n67,n68,n78,n93,n94,n97,n103
        ,n125,n126,n133,n241,n242,n250,n307,n313,n362,n373
        ,n379,n389,n395,n402,n407);
output out;
input n3;
input n22;
input n25;
input n26;
input n34;
input n35;
input n41;
input n42;
input n47;
input n55;
input n57;
input n58;
input n67;
input n68;
input n78;
input n93;
input n94;
input n97;
input n103;
input n125;
input n126;
input n133;
input n241;
input n242;
input n250;
input n307;
input n313;
input n362;
input n373;
input n379;
input n389;
input n395;
input n402;
input n407;
wire n0;
wire n1;
wire n2;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n23;
wire n24;
wire n27;
wire n28;
wire n29;
wire n30;
wire n31;
wire n32;
wire n33;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n43;
wire n44;
wire n45;
wire n46;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n56;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n95;
wire n96;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n306;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n403;
wire n404;
wire n405;
wire n406;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
xor (out,n0,n771);
nand (n0,n1,n343);
or (n1,n2,n4);
not (n2,n3);
not (n4,n5);
nand (n5,n6,n342);
or (n6,n7,n289);
not (n7,n8);
nor (n8,n9,n287);
and (n9,n10,n230);
or (n10,n11,n229);
and (n11,n12,n145);
xor (n12,n13,n108);
or (n13,n14,n107);
and (n14,n15,n81);
xor (n15,n16,n50);
nand (n16,n17,n44);
or (n17,n18,n28);
not (n18,n19);
nor (n19,n20,n27);
and (n20,n21,n23);
not (n21,n22);
not (n23,n24);
wire s0n24,s1n24,notn24;
or (n24,s0n24,s1n24);
not(notn24,n3);
and (s0n24,notn24,n25);
and (s1n24,n3,n26);
and (n27,n22,n24);
not (n28,n29);
and (n29,n30,n37);
nand (n30,n31,n36);
or (n31,n32,n24);
not (n32,n33);
wire s0n33,s1n33,notn33;
or (n33,s0n33,s1n33);
not(notn33,n3);
and (s0n33,notn33,n34);
and (s1n33,n3,n35);
nand (n36,n24,n32);
not (n37,n38);
nand (n38,n39,n43);
or (n39,n32,n40);
wire s0n40,s1n40,notn40;
or (n40,s0n40,s1n40);
not(notn40,n3);
and (s0n40,notn40,n41);
and (s1n40,n3,n42);
nand (n43,n40,n32);
nand (n44,n38,n45);
nor (n45,n46,n48);
and (n46,n47,n24);
and (n48,n23,n49);
not (n49,n47);
nand (n50,n51,n70);
or (n51,n52,n62);
not (n52,n53);
nor (n53,n54,n59);
and (n54,n55,n56);
wire s0n56,s1n56,notn56;
or (n56,s0n56,s1n56);
not(notn56,n3);
and (s0n56,notn56,n57);
and (s1n56,n3,n58);
and (n59,n60,n61);
not (n60,n55);
not (n61,n56);
not (n62,n63);
nand (n63,n64,n69);
or (n64,n65,n24);
not (n65,n66);
wire s0n66,s1n66,notn66;
or (n66,s0n66,s1n66);
not(notn66,n3);
and (s0n66,notn66,n67);
and (s1n66,n3,n68);
nand (n69,n24,n65);
nand (n70,n71,n76);
not (n71,n72);
nand (n72,n62,n73);
nand (n73,n74,n75);
or (n74,n65,n56);
nand (n75,n56,n65);
nand (n76,n77,n79);
or (n77,n61,n78);
or (n79,n56,n80);
not (n80,n78);
xor (n81,n82,n87);
and (n82,n83,n56);
nand (n83,n84,n86);
or (n84,n24,n85);
and (n85,n78,n66);
or (n86,n66,n78);
nand (n87,n88,n100);
or (n88,n89,n95);
not (n89,n90);
nor (n90,n91,n92);
not (n91,n40);
wire s0n92,s1n92,notn92;
or (n92,s0n92,s1n92);
not(notn92,n3);
and (s0n92,notn92,n93);
and (s1n92,n3,n94);
nor (n95,n96,n98);
and (n96,n91,n97);
and (n98,n40,n99);
not (n99,n97);
or (n100,n101,n106);
nor (n101,n102,n104);
and (n102,n103,n91);
and (n104,n105,n40);
not (n105,n103);
not (n106,n92);
and (n107,n16,n50);
xor (n108,n109,n117);
xor (n109,n110,n116);
nand (n110,n111,n112);
or (n111,n52,n72);
or (n112,n62,n113);
nor (n113,n114,n115);
and (n114,n61,n22);
and (n115,n56,n21);
and (n116,n82,n87);
xor (n117,n118,n138);
xor (n118,n119,n128);
and (n119,n120,n78);
not (n120,n121);
nor (n121,n122,n127);
and (n122,n123,n56);
not (n123,n124);
wire s0n124,s1n124,notn124;
or (n124,s0n124,s1n124);
not(notn124,n3);
and (s0n124,notn124,n125);
and (s1n124,n3,n126);
and (n127,n124,n61);
nand (n128,n129,n136);
or (n129,n106,n130);
not (n130,n131);
nor (n131,n132,n134);
and (n132,n133,n40);
and (n134,n135,n91);
not (n135,n133);
nand (n136,n137,n90);
not (n137,n101);
nand (n138,n139,n141);
or (n139,n140,n28);
not (n140,n45);
nand (n141,n38,n142);
nand (n142,n143,n144);
or (n143,n24,n99);
or (n144,n23,n97);
or (n145,n146,n228);
and (n146,n147,n168);
xor (n147,n148,n167);
or (n148,n149,n166);
and (n149,n150,n159);
xor (n150,n151,n152);
and (n151,n63,n78);
nand (n152,n153,n158);
or (n153,n154,n28);
not (n154,n155);
nor (n155,n156,n157);
and (n156,n55,n24);
and (n157,n60,n23);
nand (n158,n19,n38);
nand (n159,n160,n165);
or (n160,n89,n161);
not (n161,n162);
nor (n162,n163,n164);
and (n163,n49,n91);
and (n164,n47,n40);
or (n165,n95,n106);
and (n166,n151,n152);
xor (n167,n15,n81);
or (n168,n169,n227);
and (n169,n170,n226);
xor (n170,n171,n185);
nor (n171,n172,n180);
not (n172,n173);
nand (n173,n174,n179);
or (n174,n175,n89);
not (n175,n176);
nand (n176,n177,n178);
or (n177,n21,n40);
nand (n178,n40,n21);
nand (n179,n162,n92);
nand (n180,n181,n24);
nand (n181,n182,n184);
or (n182,n40,n183);
and (n183,n78,n33);
or (n184,n33,n78);
nand (n185,n186,n224);
or (n186,n187,n210);
not (n187,n188);
nand (n188,n189,n209);
or (n189,n190,n199);
nor (n190,n191,n198);
nand (n191,n192,n197);
or (n192,n193,n89);
not (n193,n194);
nand (n194,n195,n196);
or (n195,n60,n40);
nand (n196,n40,n60);
nand (n197,n176,n92);
nor (n198,n37,n80);
nand (n199,n200,n207);
nand (n200,n201,n206);
or (n201,n202,n89);
not (n202,n203);
nand (n203,n204,n205);
or (n204,n91,n78);
or (n205,n40,n80);
nand (n206,n194,n92);
nor (n207,n208,n91);
and (n208,n78,n92);
nand (n209,n191,n198);
not (n210,n211);
nand (n211,n212,n220);
not (n212,n213);
nand (n213,n214,n219);
or (n214,n215,n28);
not (n215,n216);
nand (n216,n217,n218);
or (n217,n23,n78);
or (n218,n24,n80);
nand (n219,n38,n155);
nor (n220,n221,n223);
and (n221,n172,n222);
not (n222,n180);
and (n223,n173,n180);
nand (n224,n225,n213);
not (n225,n220);
xor (n226,n150,n159);
and (n227,n171,n185);
and (n228,n148,n167);
and (n229,n13,n108);
or (n230,n231,n284);
xor (n231,n232,n255);
xor (n232,n233,n252);
xor (n233,n234,n243);
nor (n234,n235,n239);
nor (n235,n236,n238);
and (n236,n61,n237);
nand (n237,n124,n78);
and (n238,n123,n80);
not (n239,n240);
wire s0n240,s1n240,notn240;
or (n240,s0n240,s1n240);
not(notn240,n3);
and (s0n240,notn240,n241);
and (s1n240,n3,n242);
nand (n243,n244,n245);
or (n244,n130,n89);
nand (n245,n246,n92);
not (n246,n247);
nor (n247,n248,n251);
and (n248,n249,n40);
not (n249,n250);
and (n251,n250,n91);
or (n252,n253,n254);
and (n253,n118,n138);
and (n254,n119,n128);
xor (n255,n256,n278);
xor (n256,n257,n271);
nand (n257,n258,n267);
or (n258,n259,n263);
not (n259,n260);
nand (n260,n261,n262);
or (n261,n239,n78);
or (n262,n240,n80);
nand (n263,n121,n264);
nand (n264,n265,n266);
or (n265,n123,n240);
nand (n266,n240,n123);
or (n267,n121,n268);
nor (n268,n269,n270);
and (n269,n55,n239);
and (n270,n60,n240);
nand (n271,n272,n274);
or (n272,n273,n28);
not (n273,n142);
nand (n274,n38,n275);
nor (n275,n276,n277);
and (n276,n103,n24);
and (n277,n105,n23);
nand (n278,n279,n280);
or (n279,n72,n113);
or (n280,n62,n281);
nor (n281,n282,n283);
and (n282,n61,n47);
and (n283,n56,n49);
or (n284,n285,n286);
and (n285,n109,n117);
and (n286,n110,n116);
not (n287,n288);
nand (n288,n231,n284);
not (n289,n290);
nor (n290,n291,n341);
not (n291,n292);
nand (n292,n293,n338);
xor (n293,n294,n322);
xor (n294,n295,n298);
or (n295,n296,n297);
and (n296,n256,n278);
and (n297,n257,n271);
xor (n298,n299,n316);
xor (n299,n300,n308);
and (n300,n301,n78);
not (n301,n302);
nand (n302,n240,n303);
not (n303,n304);
wire s0n304,s1n304,notn304;
or (n304,s0n304,s1n304);
not(notn304,n3);
and (s0n304,notn304,1'b0);
and (s1n304,n3,n306);
and (n306,n307,n242);
nand (n308,n309,n310);
or (n309,n89,n247);
or (n310,n311,n106);
nor (n311,n312,n314);
and (n312,n91,n313);
and (n314,n40,n315);
not (n315,n313);
nand (n316,n317,n318);
or (n317,n263,n268);
or (n318,n121,n319);
nor (n319,n320,n321);
and (n320,n22,n239);
and (n321,n21,n240);
xor (n322,n323,n337);
xor (n323,n324,n331);
nand (n324,n325,n327);
or (n325,n28,n326);
not (n326,n275);
or (n327,n37,n328);
nor (n328,n329,n330);
and (n329,n23,n133);
and (n330,n24,n135);
nand (n331,n332,n333);
or (n332,n72,n281);
or (n333,n62,n334);
nor (n334,n335,n336);
and (n335,n61,n97);
and (n336,n56,n99);
and (n337,n234,n243);
or (n338,n339,n340);
and (n339,n232,n255);
and (n340,n233,n252);
nor (n341,n293,n338);
or (n342,n290,n8);
nand (n343,n344,n2);
xor (n344,n345,n528);
and (n345,n346,n526);
not (n346,n347);
nor (n347,n348,n481);
or (n348,n349,n480);
and (n349,n350,n442);
xor (n350,n351,n382);
xor (n351,n352,n369);
xor (n352,n353,n365);
nand (n353,n354,n359);
or (n354,n355,n263);
not (n355,n356);
nor (n356,n357,n358);
and (n357,n313,n240);
and (n358,n315,n239);
nand (n359,n120,n360);
nor (n360,n361,n363);
and (n361,n362,n240);
and (n363,n364,n239);
not (n364,n362);
nor (n365,n302,n366);
nor (n366,n367,n368);
and (n367,n304,n249);
and (n368,n303,n250);
nand (n369,n370,n376);
or (n370,n72,n371);
nor (n371,n372,n374);
and (n372,n61,n373);
and (n374,n56,n375);
not (n375,n373);
or (n376,n62,n377);
nor (n377,n378,n380);
and (n378,n61,n379);
and (n380,n56,n381);
not (n381,n379);
xor (n382,n383,n422);
xor (n383,n384,n408);
xor (n384,n385,n398);
nand (n385,n386,n392);
or (n386,n89,n387);
nor (n387,n388,n390);
and (n388,n91,n389);
and (n390,n40,n391);
not (n391,n389);
or (n392,n393,n106);
nor (n393,n394,n396);
and (n394,n91,n395);
and (n396,n40,n397);
not (n397,n395);
nand (n398,n399,n405);
or (n399,n28,n400);
nor (n400,n401,n403);
and (n401,n23,n402);
and (n403,n24,n404);
not (n404,n402);
or (n405,n406,n37);
xor (n406,n407,n23);
and (n408,n409,n416);
nand (n409,n410,n415);
or (n410,n89,n411);
nor (n411,n412,n413);
and (n412,n91,n407);
and (n413,n40,n414);
not (n414,n407);
or (n415,n387,n106);
nand (n416,n417,n421);
or (n417,n28,n418);
nor (n418,n419,n420);
and (n419,n23,n379);
and (n420,n24,n381);
or (n421,n37,n400);
or (n422,n423,n441);
and (n423,n424,n435);
xor (n424,n425,n431);
nand (n425,n426,n430);
or (n426,n427,n263);
nor (n427,n428,n429);
and (n428,n250,n239);
and (n429,n249,n240);
nand (n430,n120,n356);
nor (n431,n302,n432);
nor (n432,n433,n434);
and (n433,n304,n135);
and (n434,n303,n133);
nand (n435,n436,n440);
or (n436,n72,n437);
nor (n437,n438,n439);
and (n438,n61,n362);
and (n439,n56,n364);
or (n440,n62,n371);
and (n441,n425,n431);
or (n442,n443,n479);
and (n443,n444,n459);
xor (n444,n445,n446);
xor (n445,n409,n416);
and (n446,n447,n453);
nand (n447,n448,n452);
or (n448,n89,n449);
nor (n449,n450,n451);
and (n450,n91,n402);
and (n451,n40,n404);
or (n452,n411,n106);
nand (n453,n454,n458);
or (n454,n28,n455);
nor (n455,n456,n457);
and (n456,n23,n373);
and (n457,n24,n375);
or (n458,n418,n37);
or (n459,n460,n478);
and (n460,n461,n472);
xor (n461,n462,n468);
nand (n462,n463,n467);
or (n463,n263,n464);
nor (n464,n465,n466);
and (n465,n239,n133);
and (n466,n240,n135);
or (n467,n121,n427);
nor (n468,n302,n469);
nor (n469,n470,n471);
and (n470,n304,n105);
and (n471,n303,n103);
nand (n472,n473,n474);
or (n473,n437,n62);
or (n474,n72,n475);
nor (n475,n476,n477);
and (n476,n61,n313);
and (n477,n56,n315);
and (n478,n462,n468);
and (n479,n445,n446);
and (n480,n351,n382);
xor (n481,n482,n523);
xor (n482,n483,n502);
xor (n483,n484,n496);
xor (n484,n485,n492);
nand (n485,n486,n488);
or (n486,n487,n263);
not (n487,n360);
or (n488,n121,n489);
nor (n489,n490,n491);
and (n490,n239,n373);
and (n491,n240,n375);
nor (n492,n302,n493);
nor (n493,n494,n495);
and (n494,n304,n315);
and (n495,n303,n313);
nand (n496,n497,n498);
or (n497,n72,n377);
or (n498,n62,n499);
nor (n499,n500,n501);
and (n500,n61,n402);
and (n501,n56,n404);
xor (n502,n503,n520);
xor (n503,n504,n519);
xor (n504,n505,n513);
nand (n505,n506,n507);
or (n506,n89,n393);
or (n507,n508,n106);
nor (n508,n509,n511);
and (n509,n91,n510);
and (n510,n307,n395);
and (n511,n40,n512);
not (n512,n510);
nand (n513,n514,n515);
or (n514,n406,n28);
nand (n515,n38,n516);
nand (n516,n517,n518);
or (n517,n24,n391);
or (n518,n23,n389);
and (n519,n385,n398);
or (n520,n521,n522);
and (n521,n352,n369);
and (n522,n353,n365);
or (n523,n524,n525);
and (n524,n383,n422);
and (n525,n384,n408);
not (n526,n527);
and (n527,n348,n481);
nand (n528,n529,n760,n770);
nand (n529,n530,n681);
nand (n530,n531,n675,n680);
nand (n531,n532,n628);
nand (n532,n533,n627);
or (n533,n534,n582);
nor (n534,n535,n581);
and (n535,n536,n291);
not (n536,n537);
nor (n537,n538,n541);
or (n538,n539,n540);
and (n539,n294,n322);
and (n540,n295,n298);
xor (n541,n542,n564);
xor (n542,n543,n561);
xor (n543,n544,n555);
xor (n544,n545,n551);
nand (n545,n546,n547);
or (n546,n319,n263);
nand (n547,n548,n120);
nor (n548,n549,n550);
and (n549,n47,n240);
and (n550,n49,n239);
nor (n551,n302,n552);
nor (n552,n553,n554);
and (n553,n304,n60);
and (n554,n303,n55);
nand (n555,n556,n557);
or (n556,n89,n311);
or (n557,n558,n106);
nor (n558,n559,n560);
and (n559,n91,n362);
and (n560,n40,n364);
or (n561,n562,n563);
and (n562,n323,n337);
and (n563,n324,n331);
xor (n564,n565,n578);
xor (n565,n566,n572);
nand (n566,n567,n568);
or (n567,n72,n334);
or (n568,n62,n569);
nor (n569,n570,n571);
and (n570,n61,n103);
and (n571,n56,n105);
nand (n572,n573,n574);
or (n573,n28,n328);
or (n574,n575,n37);
nor (n575,n576,n577);
and (n576,n23,n250);
and (n577,n24,n249);
or (n578,n579,n580);
and (n579,n299,n316);
and (n580,n300,n308);
and (n581,n538,n541);
nor (n582,n583,n624);
xor (n583,n584,n621);
xor (n584,n585,n604);
xor (n585,n586,n598);
xor (n586,n587,n594);
nand (n587,n588,n590);
or (n588,n589,n263);
not (n589,n548);
nand (n590,n120,n591);
nor (n591,n592,n593);
and (n592,n97,n240);
and (n593,n99,n239);
nor (n594,n302,n595);
nor (n595,n596,n597);
and (n596,n304,n21);
and (n597,n303,n22);
nand (n598,n599,n600);
or (n599,n72,n569);
or (n600,n62,n601);
nor (n601,n602,n603);
and (n602,n61,n133);
and (n603,n56,n135);
xor (n604,n605,n618);
xor (n605,n606,n612);
nand (n606,n607,n608);
or (n607,n89,n558);
or (n608,n609,n106);
nor (n609,n610,n611);
and (n610,n91,n373);
and (n611,n40,n375);
nand (n612,n613,n614);
or (n613,n28,n575);
or (n614,n615,n37);
nor (n615,n616,n617);
and (n616,n23,n313);
and (n617,n24,n315);
or (n618,n619,n620);
and (n619,n544,n555);
and (n620,n545,n551);
or (n621,n622,n623);
and (n622,n565,n578);
and (n623,n566,n572);
or (n624,n625,n626);
and (n625,n542,n564);
and (n626,n543,n561);
nand (n627,n583,n624);
nand (n628,n629,n671);
not (n629,n630);
xor (n630,n631,n670);
xor (n631,n632,n651);
xor (n632,n633,n645);
xor (n633,n634,n641);
nand (n634,n635,n637);
or (n635,n636,n263);
not (n636,n591);
nand (n637,n120,n638);
nor (n638,n639,n640);
and (n639,n103,n240);
and (n640,n105,n239);
nor (n641,n302,n642);
nor (n642,n643,n644);
and (n643,n304,n49);
and (n644,n303,n47);
nand (n645,n646,n647);
or (n646,n72,n601);
or (n647,n62,n648);
nor (n648,n649,n650);
and (n649,n61,n250);
and (n650,n56,n249);
xor (n651,n652,n667);
xor (n652,n653,n666);
xor (n653,n654,n660);
nand (n654,n655,n656);
or (n655,n89,n609);
or (n656,n657,n106);
nor (n657,n658,n659);
and (n658,n91,n379);
and (n659,n40,n381);
nand (n660,n661,n662);
or (n661,n28,n615);
or (n662,n37,n663);
nor (n663,n664,n665);
and (n664,n23,n362);
and (n665,n24,n364);
and (n666,n606,n612);
or (n667,n668,n669);
and (n668,n586,n598);
and (n669,n587,n594);
and (n670,n605,n618);
not (n671,n672);
or (n672,n673,n674);
and (n673,n584,n621);
and (n674,n585,n604);
nand (n675,n628,n676,n679);
nor (n676,n8,n677);
nand (n677,n678,n536);
not (n678,n341);
not (n679,n582);
nand (n680,n630,n672);
nor (n681,n682,n739);
nand (n682,n683,n732);
not (n683,n684);
nor (n684,n685,n723);
xor (n685,n686,n714);
xor (n686,n687,n688);
xor (n687,n461,n472);
xor (n688,n689,n698);
xor (n689,n690,n691);
xor (n690,n447,n453);
and (n691,n692,n695);
nand (n692,n693,n694);
or (n693,n89,n657);
or (n694,n449,n106);
nand (n695,n696,n697);
or (n696,n28,n663);
or (n697,n455,n37);
or (n698,n699,n713);
and (n699,n700,n710);
xor (n700,n701,n706);
nand (n701,n702,n704);
or (n702,n703,n263);
not (n703,n638);
nand (n704,n705,n120);
not (n705,n464);
nor (n706,n302,n707);
nor (n707,n708,n709);
and (n708,n304,n99);
and (n709,n303,n97);
nand (n710,n711,n712);
or (n711,n72,n648);
or (n712,n62,n475);
and (n713,n701,n706);
or (n714,n715,n722);
and (n715,n716,n719);
xor (n716,n717,n718);
xor (n717,n692,n695);
and (n718,n654,n660);
or (n719,n720,n721);
and (n720,n633,n645);
and (n721,n634,n641);
and (n722,n717,n718);
or (n723,n724,n731);
and (n724,n725,n728);
xor (n725,n726,n727);
xor (n726,n700,n710);
xor (n727,n716,n719);
or (n728,n729,n730);
and (n729,n652,n667);
and (n730,n653,n666);
and (n731,n726,n727);
nand (n732,n733,n735);
not (n733,n734);
xor (n734,n725,n728);
not (n735,n736);
or (n736,n737,n738);
and (n737,n631,n670);
and (n738,n632,n651);
nand (n739,n740,n753);
nand (n740,n741,n749);
not (n741,n742);
xor (n742,n743,n746);
xor (n743,n744,n745);
xor (n744,n424,n435);
xor (n745,n444,n459);
or (n746,n747,n748);
and (n747,n689,n698);
and (n748,n690,n691);
not (n749,n750);
or (n750,n751,n752);
and (n751,n686,n714);
and (n752,n687,n688);
nand (n753,n754,n756);
not (n754,n755);
xor (n755,n350,n442);
not (n756,n757);
or (n757,n758,n759);
and (n758,n743,n746);
and (n759,n744,n745);
nand (n760,n761,n753);
nand (n761,n762,n769);
or (n762,n763,n764);
not (n763,n740);
not (n764,n765);
nand (n765,n766,n768);
or (n766,n684,n767);
nand (n767,n734,n736);
nand (n768,n685,n723);
nand (n769,n742,n750);
nand (n770,n757,n755);
wire s0n771,s1n771,notn771;
or (n771,s0n771,s1n771);
not(notn771,n3);
and (s0n771,notn771,n772);
and (s1n771,n3,n1445);
xor (n772,n773,n1325);
xor (n773,n774,n1443);
xor (n774,n775,n1320);
xor (n775,n776,n1436);
xor (n776,n777,n1314);
xor (n777,n778,n1424);
xor (n778,n779,n1308);
xor (n779,n780,n1407);
xor (n780,n781,n1302);
xor (n781,n782,n1385);
xor (n782,n783,n1296);
xor (n783,n784,n1358);
xor (n784,n785,n1290);
xor (n785,n786,n1326);
xor (n786,n787,n1284);
xor (n787,n788,n1281);
xor (n788,n789,n1280);
xor (n789,n790,n1233);
xor (n790,n791,n361);
xor (n791,n792,n1176);
xor (n792,n793,n1175);
xor (n793,n794,n1113);
xor (n794,n795,n1112);
xor (n795,n796,n1044);
xor (n796,n797,n1043);
xor (n797,n798,n972);
xor (n798,n799,n971);
xor (n799,n800,n891);
xor (n800,n801,n890);
xor (n801,n802,n805);
xor (n802,n803,n804);
and (n803,n510,n92);
and (n804,n395,n40);
or (n805,n806,n809);
and (n806,n807,n808);
and (n807,n395,n92);
and (n808,n389,n40);
and (n809,n810,n811);
xor (n810,n807,n808);
or (n811,n812,n815);
and (n812,n813,n814);
and (n813,n389,n92);
and (n814,n407,n40);
and (n815,n816,n817);
xor (n816,n813,n814);
or (n817,n818,n821);
and (n818,n819,n820);
and (n819,n407,n92);
and (n820,n402,n40);
and (n821,n822,n823);
xor (n822,n819,n820);
or (n823,n824,n827);
and (n824,n825,n826);
and (n825,n402,n92);
and (n826,n379,n40);
and (n827,n828,n829);
xor (n828,n825,n826);
or (n829,n830,n833);
and (n830,n831,n832);
and (n831,n379,n92);
and (n832,n373,n40);
and (n833,n834,n835);
xor (n834,n831,n832);
or (n835,n836,n839);
and (n836,n837,n838);
and (n837,n373,n92);
and (n838,n362,n40);
and (n839,n840,n841);
xor (n840,n837,n838);
or (n841,n842,n845);
and (n842,n843,n844);
and (n843,n362,n92);
and (n844,n313,n40);
and (n845,n846,n847);
xor (n846,n843,n844);
or (n847,n848,n851);
and (n848,n849,n850);
and (n849,n313,n92);
and (n850,n250,n40);
and (n851,n852,n853);
xor (n852,n849,n850);
or (n853,n854,n856);
and (n854,n855,n132);
and (n855,n250,n92);
and (n856,n857,n858);
xor (n857,n855,n132);
or (n858,n859,n862);
and (n859,n860,n861);
and (n860,n133,n92);
and (n861,n103,n40);
and (n862,n863,n864);
xor (n863,n860,n861);
or (n864,n865,n868);
and (n865,n866,n867);
and (n866,n103,n92);
and (n867,n97,n40);
and (n868,n869,n870);
xor (n869,n866,n867);
or (n870,n871,n873);
and (n871,n872,n164);
and (n872,n97,n92);
and (n873,n874,n875);
xor (n874,n872,n164);
or (n875,n876,n879);
and (n876,n877,n878);
and (n877,n47,n92);
and (n878,n22,n40);
and (n879,n880,n881);
xor (n880,n877,n878);
or (n881,n882,n885);
and (n882,n883,n884);
and (n883,n22,n92);
and (n884,n55,n40);
and (n885,n886,n887);
xor (n886,n883,n884);
and (n887,n888,n889);
and (n888,n55,n92);
and (n889,n78,n40);
and (n890,n389,n33);
or (n891,n892,n895);
and (n892,n893,n894);
xor (n893,n810,n811);
and (n894,n407,n33);
and (n895,n896,n897);
xor (n896,n893,n894);
or (n897,n898,n901);
and (n898,n899,n900);
xor (n899,n816,n817);
and (n900,n402,n33);
and (n901,n902,n903);
xor (n902,n899,n900);
or (n903,n904,n907);
and (n904,n905,n906);
xor (n905,n822,n823);
and (n906,n379,n33);
and (n907,n908,n909);
xor (n908,n905,n906);
or (n909,n910,n913);
and (n910,n911,n912);
xor (n911,n828,n829);
and (n912,n373,n33);
and (n913,n914,n915);
xor (n914,n911,n912);
or (n915,n916,n919);
and (n916,n917,n918);
xor (n917,n834,n835);
and (n918,n362,n33);
and (n919,n920,n921);
xor (n920,n917,n918);
or (n921,n922,n925);
and (n922,n923,n924);
xor (n923,n840,n841);
and (n924,n313,n33);
and (n925,n926,n927);
xor (n926,n923,n924);
or (n927,n928,n931);
and (n928,n929,n930);
xor (n929,n846,n847);
and (n930,n250,n33);
and (n931,n932,n933);
xor (n932,n929,n930);
or (n933,n934,n937);
and (n934,n935,n936);
xor (n935,n852,n853);
and (n936,n133,n33);
and (n937,n938,n939);
xor (n938,n935,n936);
or (n939,n940,n943);
and (n940,n941,n942);
xor (n941,n857,n858);
and (n942,n103,n33);
and (n943,n944,n945);
xor (n944,n941,n942);
or (n945,n946,n949);
and (n946,n947,n948);
xor (n947,n863,n864);
and (n948,n97,n33);
and (n949,n950,n951);
xor (n950,n947,n948);
or (n951,n952,n955);
and (n952,n953,n954);
xor (n953,n869,n870);
and (n954,n47,n33);
and (n955,n956,n957);
xor (n956,n953,n954);
or (n957,n958,n961);
and (n958,n959,n960);
xor (n959,n874,n875);
and (n960,n22,n33);
and (n961,n962,n963);
xor (n962,n959,n960);
or (n963,n964,n967);
and (n964,n965,n966);
xor (n965,n880,n881);
and (n966,n55,n33);
and (n967,n968,n969);
xor (n968,n965,n966);
and (n969,n970,n183);
xor (n970,n886,n887);
and (n971,n407,n24);
or (n972,n973,n976);
and (n973,n974,n975);
xor (n974,n896,n897);
and (n975,n402,n24);
and (n976,n977,n978);
xor (n977,n974,n975);
or (n978,n979,n982);
and (n979,n980,n981);
xor (n980,n902,n903);
and (n981,n379,n24);
and (n982,n983,n984);
xor (n983,n980,n981);
or (n984,n985,n988);
and (n985,n986,n987);
xor (n986,n908,n909);
and (n987,n373,n24);
and (n988,n989,n990);
xor (n989,n986,n987);
or (n990,n991,n994);
and (n991,n992,n993);
xor (n992,n914,n915);
and (n993,n362,n24);
and (n994,n995,n996);
xor (n995,n992,n993);
or (n996,n997,n1000);
and (n997,n998,n999);
xor (n998,n920,n921);
and (n999,n313,n24);
and (n1000,n1001,n1002);
xor (n1001,n998,n999);
or (n1002,n1003,n1006);
and (n1003,n1004,n1005);
xor (n1004,n926,n927);
and (n1005,n250,n24);
and (n1006,n1007,n1008);
xor (n1007,n1004,n1005);
or (n1008,n1009,n1012);
and (n1009,n1010,n1011);
xor (n1010,n932,n933);
and (n1011,n133,n24);
and (n1012,n1013,n1014);
xor (n1013,n1010,n1011);
or (n1014,n1015,n1017);
and (n1015,n1016,n276);
xor (n1016,n938,n939);
and (n1017,n1018,n1019);
xor (n1018,n1016,n276);
or (n1019,n1020,n1023);
and (n1020,n1021,n1022);
xor (n1021,n944,n945);
and (n1022,n97,n24);
and (n1023,n1024,n1025);
xor (n1024,n1021,n1022);
or (n1025,n1026,n1028);
and (n1026,n1027,n46);
xor (n1027,n950,n951);
and (n1028,n1029,n1030);
xor (n1029,n1027,n46);
or (n1030,n1031,n1033);
and (n1031,n1032,n27);
xor (n1032,n956,n957);
and (n1033,n1034,n1035);
xor (n1034,n1032,n27);
or (n1035,n1036,n1038);
and (n1036,n1037,n156);
xor (n1037,n962,n963);
and (n1038,n1039,n1040);
xor (n1039,n1037,n156);
and (n1040,n1041,n1042);
xor (n1041,n968,n969);
and (n1042,n78,n24);
and (n1043,n402,n66);
or (n1044,n1045,n1048);
and (n1045,n1046,n1047);
xor (n1046,n977,n978);
and (n1047,n379,n66);
and (n1048,n1049,n1050);
xor (n1049,n1046,n1047);
or (n1050,n1051,n1054);
and (n1051,n1052,n1053);
xor (n1052,n983,n984);
and (n1053,n373,n66);
and (n1054,n1055,n1056);
xor (n1055,n1052,n1053);
or (n1056,n1057,n1060);
and (n1057,n1058,n1059);
xor (n1058,n989,n990);
and (n1059,n362,n66);
and (n1060,n1061,n1062);
xor (n1061,n1058,n1059);
or (n1062,n1063,n1066);
and (n1063,n1064,n1065);
xor (n1064,n995,n996);
and (n1065,n313,n66);
and (n1066,n1067,n1068);
xor (n1067,n1064,n1065);
or (n1068,n1069,n1072);
and (n1069,n1070,n1071);
xor (n1070,n1001,n1002);
and (n1071,n250,n66);
and (n1072,n1073,n1074);
xor (n1073,n1070,n1071);
or (n1074,n1075,n1078);
and (n1075,n1076,n1077);
xor (n1076,n1007,n1008);
and (n1077,n133,n66);
and (n1078,n1079,n1080);
xor (n1079,n1076,n1077);
or (n1080,n1081,n1084);
and (n1081,n1082,n1083);
xor (n1082,n1013,n1014);
and (n1083,n103,n66);
and (n1084,n1085,n1086);
xor (n1085,n1082,n1083);
or (n1086,n1087,n1090);
and (n1087,n1088,n1089);
xor (n1088,n1018,n1019);
and (n1089,n97,n66);
and (n1090,n1091,n1092);
xor (n1091,n1088,n1089);
or (n1092,n1093,n1096);
and (n1093,n1094,n1095);
xor (n1094,n1024,n1025);
and (n1095,n47,n66);
and (n1096,n1097,n1098);
xor (n1097,n1094,n1095);
or (n1098,n1099,n1102);
and (n1099,n1100,n1101);
xor (n1100,n1029,n1030);
and (n1101,n22,n66);
and (n1102,n1103,n1104);
xor (n1103,n1100,n1101);
or (n1104,n1105,n1108);
and (n1105,n1106,n1107);
xor (n1106,n1034,n1035);
and (n1107,n55,n66);
and (n1108,n1109,n1110);
xor (n1109,n1106,n1107);
and (n1110,n1111,n85);
xor (n1111,n1039,n1040);
and (n1112,n379,n56);
or (n1113,n1114,n1117);
and (n1114,n1115,n1116);
xor (n1115,n1049,n1050);
and (n1116,n373,n56);
and (n1117,n1118,n1119);
xor (n1118,n1115,n1116);
or (n1119,n1120,n1123);
and (n1120,n1121,n1122);
xor (n1121,n1055,n1056);
and (n1122,n362,n56);
and (n1123,n1124,n1125);
xor (n1124,n1121,n1122);
or (n1125,n1126,n1129);
and (n1126,n1127,n1128);
xor (n1127,n1061,n1062);
and (n1128,n313,n56);
and (n1129,n1130,n1131);
xor (n1130,n1127,n1128);
or (n1131,n1132,n1135);
and (n1132,n1133,n1134);
xor (n1133,n1067,n1068);
and (n1134,n250,n56);
and (n1135,n1136,n1137);
xor (n1136,n1133,n1134);
or (n1137,n1138,n1141);
and (n1138,n1139,n1140);
xor (n1139,n1073,n1074);
and (n1140,n133,n56);
and (n1141,n1142,n1143);
xor (n1142,n1139,n1140);
or (n1143,n1144,n1147);
and (n1144,n1145,n1146);
xor (n1145,n1079,n1080);
and (n1146,n103,n56);
and (n1147,n1148,n1149);
xor (n1148,n1145,n1146);
or (n1149,n1150,n1153);
and (n1150,n1151,n1152);
xor (n1151,n1085,n1086);
and (n1152,n97,n56);
and (n1153,n1154,n1155);
xor (n1154,n1151,n1152);
or (n1155,n1156,n1159);
and (n1156,n1157,n1158);
xor (n1157,n1091,n1092);
and (n1158,n47,n56);
and (n1159,n1160,n1161);
xor (n1160,n1157,n1158);
or (n1161,n1162,n1165);
and (n1162,n1163,n1164);
xor (n1163,n1097,n1098);
and (n1164,n22,n56);
and (n1165,n1166,n1167);
xor (n1166,n1163,n1164);
or (n1167,n1168,n1170);
and (n1168,n1169,n54);
xor (n1169,n1103,n1104);
and (n1170,n1171,n1172);
xor (n1171,n1169,n54);
and (n1172,n1173,n1174);
xor (n1173,n1109,n1110);
and (n1174,n78,n56);
and (n1175,n373,n124);
or (n1176,n1177,n1180);
and (n1177,n1178,n1179);
xor (n1178,n1118,n1119);
and (n1179,n362,n124);
and (n1180,n1181,n1182);
xor (n1181,n1178,n1179);
or (n1182,n1183,n1186);
and (n1183,n1184,n1185);
xor (n1184,n1124,n1125);
and (n1185,n313,n124);
and (n1186,n1187,n1188);
xor (n1187,n1184,n1185);
or (n1188,n1189,n1192);
and (n1189,n1190,n1191);
xor (n1190,n1130,n1131);
and (n1191,n250,n124);
and (n1192,n1193,n1194);
xor (n1193,n1190,n1191);
or (n1194,n1195,n1198);
and (n1195,n1196,n1197);
xor (n1196,n1136,n1137);
and (n1197,n133,n124);
and (n1198,n1199,n1200);
xor (n1199,n1196,n1197);
or (n1200,n1201,n1204);
and (n1201,n1202,n1203);
xor (n1202,n1142,n1143);
and (n1203,n103,n124);
and (n1204,n1205,n1206);
xor (n1205,n1202,n1203);
or (n1206,n1207,n1210);
and (n1207,n1208,n1209);
xor (n1208,n1148,n1149);
and (n1209,n97,n124);
and (n1210,n1211,n1212);
xor (n1211,n1208,n1209);
or (n1212,n1213,n1216);
and (n1213,n1214,n1215);
xor (n1214,n1154,n1155);
and (n1215,n47,n124);
and (n1216,n1217,n1218);
xor (n1217,n1214,n1215);
or (n1218,n1219,n1222);
and (n1219,n1220,n1221);
xor (n1220,n1160,n1161);
and (n1221,n22,n124);
and (n1222,n1223,n1224);
xor (n1223,n1220,n1221);
or (n1224,n1225,n1228);
and (n1225,n1226,n1227);
xor (n1226,n1166,n1167);
and (n1227,n55,n124);
and (n1228,n1229,n1230);
xor (n1229,n1226,n1227);
and (n1230,n1231,n1232);
xor (n1231,n1171,n1172);
not (n1232,n237);
or (n1233,n1234,n1236);
and (n1234,n1235,n357);
xor (n1235,n1181,n1182);
and (n1236,n1237,n1238);
xor (n1237,n1235,n357);
or (n1238,n1239,n1242);
and (n1239,n1240,n1241);
xor (n1240,n1187,n1188);
and (n1241,n250,n240);
and (n1242,n1243,n1244);
xor (n1243,n1240,n1241);
or (n1244,n1245,n1248);
and (n1245,n1246,n1247);
xor (n1246,n1193,n1194);
and (n1247,n133,n240);
and (n1248,n1249,n1250);
xor (n1249,n1246,n1247);
or (n1250,n1251,n1253);
and (n1251,n1252,n639);
xor (n1252,n1199,n1200);
and (n1253,n1254,n1255);
xor (n1254,n1252,n639);
or (n1255,n1256,n1258);
and (n1256,n1257,n592);
xor (n1257,n1205,n1206);
and (n1258,n1259,n1260);
xor (n1259,n1257,n592);
or (n1260,n1261,n1263);
and (n1261,n1262,n549);
xor (n1262,n1211,n1212);
and (n1263,n1264,n1265);
xor (n1264,n1262,n549);
or (n1265,n1266,n1269);
and (n1266,n1267,n1268);
xor (n1267,n1217,n1218);
and (n1268,n22,n240);
and (n1269,n1270,n1271);
xor (n1270,n1267,n1268);
or (n1271,n1272,n1275);
and (n1272,n1273,n1274);
xor (n1273,n1223,n1224);
and (n1274,n55,n240);
and (n1275,n1276,n1277);
xor (n1276,n1273,n1274);
and (n1277,n1278,n1279);
xor (n1278,n1229,n1230);
and (n1279,n78,n240);
and (n1280,n313,n304);
or (n1281,n1282,n1285);
and (n1282,n1283,n1284);
xor (n1283,n1237,n1238);
and (n1284,n250,n304);
and (n1285,n1286,n1287);
xor (n1286,n1283,n1284);
or (n1287,n1288,n1291);
and (n1288,n1289,n1290);
xor (n1289,n1243,n1244);
and (n1290,n133,n304);
and (n1291,n1292,n1293);
xor (n1292,n1289,n1290);
or (n1293,n1294,n1297);
and (n1294,n1295,n1296);
xor (n1295,n1249,n1250);
and (n1296,n103,n304);
and (n1297,n1298,n1299);
xor (n1298,n1295,n1296);
or (n1299,n1300,n1303);
and (n1300,n1301,n1302);
xor (n1301,n1254,n1255);
and (n1302,n97,n304);
and (n1303,n1304,n1305);
xor (n1304,n1301,n1302);
or (n1305,n1306,n1309);
and (n1306,n1307,n1308);
xor (n1307,n1259,n1260);
and (n1308,n47,n304);
and (n1309,n1310,n1311);
xor (n1310,n1307,n1308);
or (n1311,n1312,n1315);
and (n1312,n1313,n1314);
xor (n1313,n1264,n1265);
and (n1314,n22,n304);
and (n1315,n1316,n1317);
xor (n1316,n1313,n1314);
or (n1317,n1318,n1321);
and (n1318,n1319,n1320);
xor (n1319,n1270,n1271);
and (n1320,n55,n304);
and (n1321,n1322,n1323);
xor (n1322,n1319,n1320);
and (n1323,n1324,n1325);
xor (n1324,n1276,n1277);
and (n1325,n78,n304);
or (n1326,n1327,n1329);
and (n1327,n1328,n1290);
xor (n1328,n1286,n1287);
and (n1329,n1330,n1331);
xor (n1330,n1328,n1290);
or (n1331,n1332,n1334);
and (n1332,n1333,n1296);
xor (n1333,n1292,n1293);
and (n1334,n1335,n1336);
xor (n1335,n1333,n1296);
or (n1336,n1337,n1339);
and (n1337,n1338,n1302);
xor (n1338,n1298,n1299);
and (n1339,n1340,n1341);
xor (n1340,n1338,n1302);
or (n1341,n1342,n1344);
and (n1342,n1343,n1308);
xor (n1343,n1304,n1305);
and (n1344,n1345,n1346);
xor (n1345,n1343,n1308);
or (n1346,n1347,n1349);
and (n1347,n1348,n1314);
xor (n1348,n1310,n1311);
and (n1349,n1350,n1351);
xor (n1350,n1348,n1314);
or (n1351,n1352,n1354);
and (n1352,n1353,n1320);
xor (n1353,n1316,n1317);
and (n1354,n1355,n1356);
xor (n1355,n1353,n1320);
and (n1356,n1357,n1325);
xor (n1357,n1322,n1323);
or (n1358,n1359,n1361);
and (n1359,n1360,n1296);
xor (n1360,n1330,n1331);
and (n1361,n1362,n1363);
xor (n1362,n1360,n1296);
or (n1363,n1364,n1366);
and (n1364,n1365,n1302);
xor (n1365,n1335,n1336);
and (n1366,n1367,n1368);
xor (n1367,n1365,n1302);
or (n1368,n1369,n1371);
and (n1369,n1370,n1308);
xor (n1370,n1340,n1341);
and (n1371,n1372,n1373);
xor (n1372,n1370,n1308);
or (n1373,n1374,n1376);
and (n1374,n1375,n1314);
xor (n1375,n1345,n1346);
and (n1376,n1377,n1378);
xor (n1377,n1375,n1314);
or (n1378,n1379,n1381);
and (n1379,n1380,n1320);
xor (n1380,n1350,n1351);
and (n1381,n1382,n1383);
xor (n1382,n1380,n1320);
and (n1383,n1384,n1325);
xor (n1384,n1355,n1356);
or (n1385,n1386,n1388);
and (n1386,n1387,n1302);
xor (n1387,n1362,n1363);
and (n1388,n1389,n1390);
xor (n1389,n1387,n1302);
or (n1390,n1391,n1393);
and (n1391,n1392,n1308);
xor (n1392,n1367,n1368);
and (n1393,n1394,n1395);
xor (n1394,n1392,n1308);
or (n1395,n1396,n1398);
and (n1396,n1397,n1314);
xor (n1397,n1372,n1373);
and (n1398,n1399,n1400);
xor (n1399,n1397,n1314);
or (n1400,n1401,n1403);
and (n1401,n1402,n1320);
xor (n1402,n1377,n1378);
and (n1403,n1404,n1405);
xor (n1404,n1402,n1320);
and (n1405,n1406,n1325);
xor (n1406,n1382,n1383);
or (n1407,n1408,n1410);
and (n1408,n1409,n1308);
xor (n1409,n1389,n1390);
and (n1410,n1411,n1412);
xor (n1411,n1409,n1308);
or (n1412,n1413,n1415);
and (n1413,n1414,n1314);
xor (n1414,n1394,n1395);
and (n1415,n1416,n1417);
xor (n1416,n1414,n1314);
or (n1417,n1418,n1420);
and (n1418,n1419,n1320);
xor (n1419,n1399,n1400);
and (n1420,n1421,n1422);
xor (n1421,n1419,n1320);
and (n1422,n1423,n1325);
xor (n1423,n1404,n1405);
or (n1424,n1425,n1427);
and (n1425,n1426,n1314);
xor (n1426,n1411,n1412);
and (n1427,n1428,n1429);
xor (n1428,n1426,n1314);
or (n1429,n1430,n1432);
and (n1430,n1431,n1320);
xor (n1431,n1416,n1417);
and (n1432,n1433,n1434);
xor (n1433,n1431,n1320);
and (n1434,n1435,n1325);
xor (n1435,n1421,n1422);
or (n1436,n1437,n1439);
and (n1437,n1438,n1320);
xor (n1438,n1428,n1429);
and (n1439,n1440,n1441);
xor (n1440,n1438,n1320);
and (n1441,n1442,n1325);
xor (n1442,n1433,n1434);
and (n1443,n1444,n1325);
xor (n1444,n1440,n1441);
xor (n1445,n1324,n1325);
endmodule
