module top (out,n7,n9,n10,n14,n22,n23,n30,n44,n63
        ,n65,n74,n75,n99,n100,n112,n165,n166,n170,n175
        ,n195,n197,n213,n267,n299,n428,n442,n443,n515,n524
        ,n525,n561,n633,n663,n664,n854,n858,n860,n886,n887
        ,n994,n1011,n1012,n1198,n1202,n1204,n1215,n1227,n1241);
output out;
input n7;
input n9;
input n10;
input n14;
input n22;
input n23;
input n30;
input n44;
input n63;
input n65;
input n74;
input n75;
input n99;
input n100;
input n112;
input n165;
input n166;
input n170;
input n175;
input n195;
input n197;
input n213;
input n267;
input n299;
input n428;
input n442;
input n443;
input n515;
input n524;
input n525;
input n561;
input n633;
input n663;
input n664;
input n854;
input n858;
input n860;
input n886;
input n887;
input n994;
input n1011;
input n1012;
input n1198;
input n1202;
input n1204;
input n1215;
input n1227;
input n1241;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n8;
wire n11;
wire n12;
wire n13;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n24;
wire n25;
wire n26;
wire n27;
wire n28;
wire n29;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n64;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n167;
wire n168;
wire n169;
wire n171;
wire n172;
wire n173;
wire n174;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n196;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n855;
wire n856;
wire n857;
wire n859;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1199;
wire n1200;
wire n1201;
wire n1203;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2988;
wire n2989;
wire n2990;
wire n2991;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2996;
wire n2997;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3003;
wire n3004;
wire n3005;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3010;
wire n3011;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3038;
wire n3039;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
wire n3056;
wire n3057;
wire n3058;
wire n3059;
wire n3060;
wire n3061;
wire n3062;
wire n3063;
wire n3064;
wire n3065;
wire n3066;
wire n3067;
wire n3068;
wire n3069;
wire n3070;
wire n3071;
wire n3072;
wire n3073;
wire n3074;
wire n3075;
wire n3076;
wire n3077;
wire n3078;
wire n3079;
wire n3080;
wire n3081;
wire n3082;
wire n3083;
wire n3084;
wire n3085;
wire n3086;
wire n3087;
wire n3088;
wire n3089;
wire n3090;
wire n3091;
wire n3092;
wire n3093;
wire n3094;
wire n3095;
wire n3096;
wire n3097;
wire n3098;
wire n3099;
wire n3100;
wire n3101;
wire n3102;
wire n3103;
wire n3104;
wire n3105;
wire n3106;
wire n3107;
wire n3108;
wire n3109;
wire n3110;
wire n3111;
wire n3112;
wire n3113;
wire n3114;
wire n3115;
wire n3116;
wire n3117;
wire n3118;
wire n3119;
wire n3120;
wire n3121;
wire n3122;
wire n3123;
wire n3124;
wire n3125;
wire n3126;
wire n3127;
wire n3128;
wire n3129;
wire n3130;
wire n3131;
wire n3132;
wire n3133;
wire n3134;
wire n3135;
wire n3136;
wire n3137;
wire n3138;
wire n3139;
wire n3140;
wire n3141;
wire n3142;
wire n3143;
wire n3144;
wire n3145;
wire n3146;
wire n3147;
wire n3148;
wire n3149;
wire n3150;
wire n3151;
wire n3152;
wire n3153;
wire n3154;
wire n3155;
wire n3156;
wire n3157;
wire n3158;
wire n3159;
wire n3160;
wire n3161;
wire n3162;
wire n3163;
wire n3164;
wire n3165;
wire n3166;
wire n3167;
wire n3168;
wire n3169;
wire n3170;
wire n3171;
wire n3172;
wire n3173;
wire n3174;
wire n3175;
wire n3176;
wire n3177;
wire n3178;
wire n3179;
wire n3180;
wire n3181;
wire n3182;
wire n3183;
wire n3184;
wire n3185;
wire n3186;
wire n3187;
wire n3188;
wire n3189;
wire n3190;
wire n3191;
wire n3192;
wire n3193;
wire n3194;
wire n3195;
wire n3196;
wire n3197;
wire n3198;
wire n3199;
wire n3200;
wire n3201;
wire n3202;
wire n3203;
wire n3204;
wire n3205;
wire n3206;
wire n3207;
wire n3208;
wire n3209;
wire n3210;
wire n3211;
wire n3212;
wire n3213;
wire n3214;
wire n3215;
wire n3216;
wire n3217;
wire n3218;
wire n3219;
wire n3220;
wire n3221;
wire n3222;
wire n3223;
wire n3224;
wire n3225;
wire n3226;
wire n3227;
wire n3228;
wire n3229;
wire n3230;
wire n3231;
wire n3232;
wire n3233;
wire n3234;
wire n3235;
wire n3236;
wire n3237;
wire n3238;
wire n3239;
wire n3240;
wire n3241;
wire n3242;
wire n3243;
wire n3244;
wire n3245;
wire n3246;
wire n3247;
wire n3248;
wire n3249;
wire n3250;
wire n3251;
wire n3252;
wire n3253;
wire n3254;
wire n3255;
wire n3256;
wire n3257;
wire n3258;
wire n3259;
wire n3260;
wire n3261;
wire n3262;
wire n3263;
wire n3264;
wire n3265;
wire n3266;
wire n3267;
wire n3268;
wire n3269;
wire n3270;
wire n3271;
wire n3272;
wire n3273;
wire n3274;
wire n3275;
wire n3276;
wire n3277;
wire n3278;
wire n3279;
wire n3280;
wire n3281;
wire n3282;
wire n3283;
wire n3284;
wire n3285;
wire n3286;
wire n3287;
wire n3288;
wire n3289;
wire n3290;
wire n3291;
wire n3292;
wire n3293;
wire n3294;
wire n3295;
wire n3296;
wire n3297;
wire n3298;
wire n3299;
wire n3300;
wire n3301;
wire n3302;
wire n3303;
wire n3304;
wire n3305;
wire n3306;
wire n3307;
wire n3308;
wire n3309;
wire n3310;
wire n3311;
wire n3312;
wire n3313;
wire n3314;
wire n3315;
wire n3316;
wire n3317;
wire n3318;
wire n3319;
wire n3320;
wire n3321;
wire n3322;
wire n3323;
wire n3324;
wire n3325;
wire n3326;
wire n3327;
wire n3328;
wire n3329;
wire n3330;
wire n3331;
wire n3332;
wire n3333;
wire n3334;
wire n3335;
wire n3336;
wire n3337;
wire n3338;
wire n3339;
wire n3340;
wire n3341;
wire n3342;
wire n3343;
wire n3344;
wire n3345;
wire n3346;
wire n3347;
wire n3348;
wire n3349;
wire n3350;
wire n3351;
wire n3352;
wire n3353;
wire n3354;
wire n3355;
wire n3356;
wire n3357;
wire n3358;
wire n3359;
wire n3360;
wire n3361;
wire n3362;
wire n3363;
wire n3364;
wire n3365;
wire n3366;
wire n3367;
wire n3368;
wire n3369;
wire n3370;
wire n3371;
wire n3372;
wire n3373;
wire n3374;
wire n3375;
wire n3376;
wire n3377;
wire n3378;
wire n3379;
wire n3380;
wire n3381;
wire n3382;
wire n3383;
wire n3384;
wire n3385;
wire n3386;
wire n3387;
wire n3388;
wire n3389;
wire n3390;
wire n3391;
wire n3392;
wire n3393;
wire n3394;
wire n3395;
wire n3396;
wire n3397;
wire n3398;
wire n3399;
wire n3400;
wire n3401;
wire n3402;
wire n3403;
wire n3404;
wire n3405;
wire n3406;
wire n3407;
wire n3408;
wire n3409;
wire n3410;
wire n3411;
wire n3412;
wire n3413;
wire n3414;
wire n3415;
wire n3416;
wire n3417;
wire n3418;
wire n3419;
wire n3420;
wire n3421;
wire n3422;
wire n3423;
wire n3424;
wire n3425;
wire n3426;
wire n3427;
wire n3428;
wire n3429;
wire n3430;
wire n3431;
wire n3432;
wire n3433;
wire n3434;
wire n3435;
wire n3436;
wire n3437;
wire n3438;
wire n3439;
wire n3440;
wire n3441;
wire n3442;
wire n3443;
wire n3444;
wire n3445;
wire n3446;
wire n3447;
wire n3448;
wire n3449;
wire n3450;
wire n3451;
wire n3452;
wire n3453;
wire n3454;
wire n3455;
wire n3456;
wire n3457;
wire n3458;
wire n3459;
wire n3460;
wire n3461;
wire n3462;
wire n3463;
wire n3464;
wire n3465;
wire n3466;
wire n3467;
wire n3468;
wire n3469;
wire n3470;
wire n3471;
wire n3472;
wire n3473;
wire n3474;
wire n3475;
wire n3476;
wire n3477;
wire n3478;
wire n3479;
wire n3480;
wire n3481;
wire n3482;
wire n3483;
wire n3484;
wire n3485;
wire n3486;
wire n3487;
wire n3488;
wire n3489;
wire n3490;
wire n3491;
wire n3492;
wire n3493;
wire n3494;
wire n3495;
wire n3496;
wire n3497;
wire n3498;
wire n3499;
wire n3500;
wire n3501;
wire n3502;
wire n3503;
wire n3504;
wire n3505;
wire n3506;
wire n3507;
wire n3508;
wire n3509;
wire n3510;
wire n3511;
wire n3512;
wire n3513;
wire n3514;
wire n3515;
wire n3516;
wire n3517;
wire n3518;
wire n3519;
wire n3520;
wire n3521;
wire n3522;
wire n3523;
wire n3524;
wire n3525;
wire n3526;
wire n3527;
wire n3528;
wire n3529;
wire n3530;
wire n3531;
wire n3532;
wire n3533;
wire n3534;
wire n3535;
wire n3536;
wire n3537;
wire n3538;
wire n3539;
wire n3540;
wire n3541;
wire n3542;
wire n3543;
wire n3544;
wire n3545;
wire n3546;
wire n3547;
wire n3548;
wire n3549;
wire n3550;
wire n3551;
wire n3552;
wire n3553;
wire n3554;
wire n3555;
wire n3556;
wire n3557;
wire n3558;
wire n3559;
wire n3560;
wire n3561;
wire n3562;
wire n3563;
wire n3564;
wire n3565;
wire n3566;
wire n3567;
wire n3568;
wire n3569;
wire n3570;
wire n3571;
wire n3572;
wire n3573;
wire n3574;
wire n3575;
wire n3576;
wire n3577;
wire n3578;
wire n3579;
wire n3580;
wire n3581;
wire n3582;
wire n3583;
wire n3584;
wire n3585;
wire n3586;
wire n3587;
wire n3588;
wire n3589;
wire n3590;
wire n3591;
wire n3592;
wire n3593;
wire n3594;
wire n3595;
wire n3596;
wire n3597;
wire n3598;
wire n3599;
wire n3600;
wire n3601;
wire n3602;
wire n3603;
wire n3604;
wire n3605;
wire n3606;
wire n3607;
wire n3608;
wire n3609;
wire n3610;
wire n3611;
wire n3612;
wire n3613;
wire n3614;
wire n3615;
wire n3616;
wire n3617;
wire n3618;
wire n3619;
wire n3620;
wire n3621;
wire n3622;
wire n3623;
wire n3624;
wire n3625;
wire n3626;
wire n3627;
wire n3628;
wire n3629;
wire n3630;
wire n3631;
wire n3632;
wire n3633;
wire n3634;
wire n3635;
wire n3636;
wire n3637;
wire n3638;
wire n3639;
wire n3640;
wire n3641;
wire n3642;
wire n3643;
wire n3644;
wire n3645;
wire n3646;
wire n3647;
wire n3648;
wire n3649;
wire n3650;
wire n3651;
wire n3652;
wire n3653;
wire n3654;
wire n3655;
wire n3656;
wire n3657;
wire n3658;
wire n3659;
wire n3660;
wire n3661;
wire n3662;
wire n3663;
wire n3664;
wire n3665;
wire n3666;
wire n3667;
wire n3668;
wire n3669;
wire n3670;
wire n3671;
wire n3672;
wire n3673;
wire n3674;
wire n3675;
wire n3676;
wire n3677;
wire n3678;
wire n3679;
wire n3680;
wire n3681;
wire n3682;
wire n3683;
wire n3684;
wire n3685;
wire n3686;
wire n3687;
wire n3688;
wire n3689;
wire n3690;
wire n3691;
wire n3692;
wire n3693;
wire n3694;
wire n3695;
wire n3696;
wire n3697;
wire n3698;
wire n3699;
wire n3700;
wire n3701;
wire n3702;
wire n3703;
wire n3704;
wire n3705;
wire n3706;
wire n3707;
wire n3708;
wire n3709;
wire n3710;
wire n3711;
wire n3712;
wire n3713;
wire n3714;
wire n3715;
wire n3716;
wire n3717;
wire n3718;
wire n3719;
wire n3720;
wire n3721;
wire n3722;
wire n3723;
wire n3724;
wire n3725;
wire n3726;
wire n3727;
wire n3728;
wire n3729;
wire n3730;
wire n3731;
wire n3732;
wire n3733;
wire n3734;
wire n3735;
wire n3736;
wire n3737;
wire n3738;
wire n3739;
wire n3740;
wire n3741;
wire n3742;
wire n3743;
wire n3744;
wire n3745;
wire n3746;
wire n3747;
wire n3748;
wire n3749;
wire n3750;
wire n3751;
wire n3752;
wire n3753;
wire n3754;
wire n3755;
wire n3756;
wire n3757;
wire n3758;
wire n3759;
wire n3760;
wire n3761;
wire n3762;
wire n3763;
wire n3764;
wire n3765;
wire n3766;
wire n3767;
wire n3768;
wire n3769;
wire n3770;
wire n3771;
wire n3772;
wire n3773;
wire n3774;
wire n3775;
wire n3776;
wire n3777;
wire n3778;
wire n3779;
wire n3780;
wire n3781;
wire n3782;
wire n3783;
wire n3784;
wire n3785;
wire n3786;
wire n3787;
wire n3788;
wire n3789;
wire n3790;
wire n3791;
wire n3792;
wire n3793;
wire n3794;
wire n3795;
wire n3796;
wire n3797;
wire n3798;
wire n3799;
wire n3800;
wire n3801;
wire n3802;
wire n3803;
wire n3804;
wire n3805;
wire n3806;
wire n3807;
wire n3808;
wire n3809;
wire n3810;
wire n3811;
wire n3812;
wire n3813;
wire n3814;
wire n3815;
wire n3816;
wire n3817;
wire n3818;
wire n3819;
wire n3820;
wire n3821;
wire n3822;
wire n3823;
wire n3824;
wire n3825;
wire n3826;
wire n3827;
wire n3828;
wire n3829;
wire n3830;
wire n3831;
wire n3832;
wire n3833;
wire n3834;
wire n3835;
wire n3836;
wire n3837;
wire n3838;
wire n3839;
wire n3840;
wire n3841;
wire n3842;
wire n3843;
wire n3844;
wire n3845;
wire n3846;
wire n3847;
wire n3848;
wire n3849;
wire n3850;
wire n3851;
wire n3852;
wire n3853;
wire n3854;
wire n3855;
wire n3856;
wire n3857;
wire n3858;
wire n3859;
wire n3860;
wire n3861;
wire n3862;
wire n3863;
wire n3864;
wire n3865;
wire n3866;
wire n3867;
wire n3868;
wire n3869;
wire n3870;
wire n3871;
wire n3872;
wire n3873;
wire n3874;
wire n3875;
wire n3876;
wire n3877;
wire n3878;
wire n3879;
wire n3880;
wire n3881;
wire n3882;
wire n3883;
wire n3884;
wire n3885;
wire n3886;
wire n3887;
wire n3888;
wire n3889;
wire n3890;
wire n3891;
wire n3892;
wire n3893;
wire n3894;
wire n3895;
xor (out,n0,n3143);
not (n0,n1);
nand (n1,n2,n47);
nand (n2,n3,n33);
xor (n3,n4,n15);
not (n4,n5);
or (n5,n6,n11);
and (n6,n7,n8);
xor (n8,n9,n10);
and (n11,n7,n12);
nor (n12,n8,n13);
xnor (n13,n14,n9);
nand (n15,n16,n31,n32);
nand (n16,n17,n27);
not (n17,n18);
xor (n18,n19,n10);
or (n19,n20,n24);
and (n20,n7,n21);
xor (n21,n22,n23);
and (n24,n7,n25);
nor (n25,n21,n26);
xnor (n26,n10,n22);
xor (n27,n28,n14);
or (n28,n6,n29);
and (n29,n30,n12);
nand (n31,n14,n27);
nand (n32,n17,n14);
nand (n33,n34,n37,n46);
nand (n34,n18,n35);
xor (n35,n36,n14);
xor (n36,n17,n27);
nand (n37,n38,n35);
nand (n38,n39,n32,n45);
nand (n39,n40,n14);
xor (n40,n41,n14);
or (n41,n42,n43);
and (n42,n30,n8);
and (n43,n44,n12);
nand (n45,n40,n17);
nand (n46,n18,n38);
nand (n47,n48,n3141);
nand (n48,n49,n145);
nor (n49,n50,n143);
nor (n50,n51,n136);
nand (n51,n52,n125);
nand (n52,n53,n89,n124);
nand (n53,n54,n68);
nand (n54,n55,n66,n67);
nand (n55,n56,n60);
xor (n56,n57,n10);
or (n57,n58,n59);
and (n58,n30,n21);
and (n59,n44,n25);
xor (n60,n61,n14);
or (n61,n62,n64);
and (n62,n63,n8);
and (n64,n65,n12);
nand (n66,n14,n60);
nand (n67,n56,n14);
xor (n68,n69,n79);
xor (n69,n14,n70);
xor (n70,n71,n23);
or (n71,n72,n76);
and (n72,n7,n73);
xor (n73,n74,n75);
and (n76,n7,n77);
nor (n77,n73,n78);
xnor (n78,n23,n74);
xor (n79,n80,n85);
xor (n80,n81,n82);
not (n81,n70);
xor (n82,n83,n10);
or (n83,n20,n84);
and (n84,n30,n25);
xor (n85,n86,n14);
or (n86,n87,n88);
and (n87,n44,n8);
and (n88,n63,n12);
nand (n89,n90,n68);
nand (n90,n91,n114,n123);
nand (n91,n81,n92);
nand (n92,n93,n107,n113);
nand (n93,n94,n104);
not (n94,n95);
xor (n95,n96,n75);
or (n96,n97,n101);
and (n97,n7,n98);
xor (n98,n99,n100);
and (n101,n7,n102);
nor (n102,n98,n103);
xnor (n103,n75,n99);
xor (n104,n105,n23);
or (n105,n72,n106);
and (n106,n30,n77);
nand (n107,n108,n104);
xor (n108,n109,n14);
or (n109,n110,n111);
and (n110,n65,n8);
and (n111,n112,n12);
nand (n113,n94,n108);
nand (n114,n115,n92);
nand (n115,n116,n121,n122);
nand (n116,n117,n14);
xor (n117,n118,n10);
or (n118,n119,n120);
and (n119,n44,n21);
and (n120,n63,n25);
nand (n121,n95,n14);
nand (n122,n117,n95);
nand (n123,n81,n115);
nand (n124,n54,n90);
xor (n125,n126,n132);
xor (n126,n127,n131);
nand (n127,n128,n129,n130);
nand (n128,n81,n82);
nand (n129,n85,n82);
nand (n130,n81,n85);
xor (n131,n41,n17);
nand (n132,n133,n134,n135);
nand (n133,n14,n70);
nand (n134,n79,n70);
nand (n135,n14,n79);
nor (n136,n137,n139);
xor (n137,n138,n38);
not (n138,n28);
nand (n139,n140,n141,n142);
nand (n140,n127,n131);
nand (n141,n132,n131);
nand (n142,n127,n132);
not (n143,n144);
nand (n144,n137,n139);
nand (n145,n146,n148);
nor (n146,n147,n136);
nor (n147,n52,n125);
nand (n148,n149,n403);
nor (n149,n150,n397);
nor (n150,n151,n373);
nor (n151,n152,n371);
nor (n152,n153,n346);
nand (n153,n154,n310);
nand (n154,n155,n256,n309);
nand (n155,n156,n215);
nand (n156,n157,n199,n214);
nand (n157,n158,n185);
nand (n158,n159,n179,n184);
nand (n159,n160,n171);
not (n160,n161);
xor (n161,n162,n170);
or (n162,n163,n167);
and (n163,n7,n164);
xor (n164,n165,n166);
and (n167,n7,n168);
nor (n168,n164,n169);
xnor (n169,n170,n165);
xor (n171,n172,n100);
or (n172,n173,n176);
and (n173,n7,n174);
xor (n174,n175,n170);
and (n176,n30,n177);
nor (n177,n174,n178);
xnor (n178,n100,n175);
nand (n179,n180,n171);
xor (n180,n181,n75);
or (n181,n182,n183);
and (n182,n44,n98);
and (n183,n63,n102);
nand (n184,n160,n180);
nand (n185,n186,n191,n198);
nand (n186,n187,n161);
xor (n187,n188,n23);
or (n188,n189,n190);
and (n189,n65,n73);
and (n190,n112,n77);
nand (n191,n192,n161);
xor (n192,n193,n10);
or (n193,n194,n196);
and (n194,n195,n21);
and (n196,n197,n25);
nand (n198,n187,n192);
nand (n199,n200,n185);
xor (n200,n201,n209);
xor (n201,n202,n205);
xor (n202,n203,n100);
or (n203,n173,n204);
and (n204,n7,n177);
xor (n205,n206,n10);
or (n206,n207,n208);
and (n207,n112,n21);
and (n208,n195,n25);
xor (n209,n210,n14);
or (n210,n211,n212);
and (n211,n197,n8);
and (n212,n213,n12);
nand (n214,n158,n200);
xor (n215,n216,n240);
xor (n216,n217,n230);
nand (n217,n218,n228,n229);
nand (n218,n219,n223);
xor (n219,n220,n23);
or (n220,n221,n222);
and (n221,n63,n73);
and (n222,n65,n77);
not (n223,n224);
xor (n224,n225,n75);
or (n225,n226,n227);
and (n226,n30,n98);
and (n227,n44,n102);
nand (n228,n14,n223);
nand (n229,n219,n14);
xor (n230,n231,n14);
xor (n231,n232,n236);
xor (n232,n233,n14);
or (n233,n234,n235);
and (n234,n195,n8);
and (n235,n197,n12);
xor (n236,n237,n23);
or (n237,n238,n239);
and (n238,n44,n73);
and (n239,n63,n77);
xor (n240,n241,n246);
xor (n241,n224,n242);
nand (n242,n243,n244,n245);
nand (n243,n202,n205);
nand (n244,n209,n205);
nand (n245,n202,n209);
xor (n246,n247,n252);
xor (n247,n248,n249);
not (n248,n202);
xor (n249,n250,n75);
or (n250,n97,n251);
and (n251,n30,n102);
xor (n252,n253,n10);
or (n253,n254,n255);
and (n254,n65,n21);
and (n255,n112,n25);
nand (n256,n257,n215);
nand (n257,n258,n286,n308);
nand (n258,n259,n261);
xor (n259,n260,n14);
xor (n260,n219,n223);
nand (n261,n262,n268,n285);
nand (n262,n263,n14);
xor (n263,n264,n14);
or (n264,n265,n266);
and (n265,n213,n8);
and (n266,n267,n12);
nand (n268,n269,n14);
nand (n269,n270,n279,n284);
nand (n270,n271,n275);
xor (n271,n272,n100);
or (n272,n273,n274);
and (n273,n30,n174);
and (n274,n44,n177);
xor (n275,n276,n75);
or (n276,n277,n278);
and (n277,n63,n98);
and (n278,n65,n102);
nand (n279,n280,n275);
xor (n280,n281,n23);
or (n281,n282,n283);
and (n282,n112,n73);
and (n283,n195,n77);
nand (n284,n271,n280);
nand (n285,n263,n269);
nand (n286,n287,n261);
nand (n287,n288,n304,n307);
nand (n288,n289,n302);
nand (n289,n290,n300,n301);
nand (n290,n291,n295);
xor (n291,n292,n10);
or (n292,n293,n294);
and (n293,n197,n21);
and (n294,n213,n25);
xor (n295,n296,n14);
or (n296,n297,n298);
and (n297,n267,n8);
and (n298,n299,n12);
nand (n300,n160,n295);
nand (n301,n291,n160);
xor (n302,n303,n180);
xor (n303,n160,n171);
nand (n304,n305,n302);
xor (n305,n306,n192);
xor (n306,n187,n161);
nand (n307,n289,n305);
nand (n308,n259,n287);
nand (n309,n156,n257);
xor (n310,n311,n342);
xor (n311,n312,n316);
nand (n312,n313,n314,n315);
nand (n313,n224,n242);
nand (n314,n246,n242);
nand (n315,n224,n246);
xor (n316,n317,n336);
xor (n317,n318,n332);
xor (n318,n319,n328);
xor (n319,n320,n324);
xor (n320,n321,n23);
or (n321,n322,n323);
and (n322,n30,n73);
and (n323,n44,n77);
xor (n324,n325,n14);
or (n325,n326,n327);
and (n326,n112,n8);
and (n327,n195,n12);
xor (n328,n329,n10);
or (n329,n330,n331);
and (n330,n63,n21);
and (n331,n65,n25);
nand (n332,n333,n334,n335);
nand (n333,n232,n236);
nand (n334,n14,n236);
nand (n335,n232,n14);
xor (n336,n337,n338);
xor (n337,n94,n14);
nand (n338,n339,n340,n341);
nand (n339,n248,n249);
nand (n340,n252,n249);
nand (n341,n248,n252);
nand (n342,n343,n344,n345);
nand (n343,n217,n230);
nand (n344,n240,n230);
nand (n345,n217,n240);
nor (n346,n347,n367);
xor (n347,n348,n363);
xor (n348,n349,n353);
nand (n349,n350,n351,n352);
nand (n350,n94,n14);
nand (n351,n338,n14);
nand (n352,n94,n338);
xor (n353,n354,n361);
xor (n354,n355,n359);
nand (n355,n356,n357,n358);
nand (n356,n320,n324);
nand (n357,n328,n324);
nand (n358,n320,n328);
xor (n359,n360,n108);
xor (n360,n94,n104);
xor (n361,n362,n95);
xor (n362,n117,n14);
nand (n363,n364,n365,n366);
nand (n364,n318,n332);
nand (n365,n336,n332);
nand (n366,n318,n336);
nand (n367,n368,n369,n370);
nand (n368,n312,n316);
nand (n369,n342,n316);
nand (n370,n312,n342);
not (n371,n372);
nand (n372,n347,n367);
not (n373,n374);
nor (n374,n375,n390);
nor (n375,n376,n386);
xor (n376,n377,n382);
xor (n377,n378,n380);
xor (n378,n379,n14);
xor (n379,n56,n60);
xor (n380,n381,n115);
xor (n381,n81,n92);
nand (n382,n383,n384,n385);
nand (n383,n355,n359);
nand (n384,n361,n359);
nand (n385,n355,n361);
nand (n386,n387,n388,n389);
nand (n387,n349,n353);
nand (n388,n363,n353);
nand (n389,n349,n363);
nor (n390,n391,n395);
nand (n391,n392,n393,n394);
nand (n392,n378,n380);
nand (n393,n382,n380);
nand (n394,n378,n382);
xor (n395,n396,n90);
xor (n396,n54,n68);
not (n397,n398);
nor (n398,n399,n401);
nor (n399,n400,n390);
nand (n400,n376,n386);
not (n401,n402);
nand (n402,n391,n395);
nand (n403,n404,n3137);
nand (n404,n405,n1175);
nor (n405,n406,n1160);
nor (n406,n407,n753);
nand (n407,n408,n730);
nor (n408,n409,n706);
nor (n409,n410,n583);
xor (n410,n411,n540);
xor (n411,n412,n431);
xor (n412,n413,n418);
xor (n413,n414,n416);
xor (n414,n415,n280);
xor (n415,n271,n275);
xor (n416,n417,n160);
xor (n417,n291,n295);
nand (n418,n419,n429,n430);
nand (n419,n420,n424);
xor (n420,n421,n10);
or (n421,n422,n423);
and (n422,n213,n21);
and (n423,n267,n25);
xor (n424,n425,n14);
or (n425,n426,n427);
and (n426,n299,n8);
and (n427,n428,n12);
nand (n429,n14,n424);
nand (n430,n420,n14);
xor (n431,n432,n502);
xor (n432,n433,n468);
xor (n433,n434,n456);
xor (n434,n14,n435);
nand (n435,n436,n450,n455);
nand (n436,n437,n447);
not (n437,n438);
xor (n438,n439,n166);
or (n439,n440,n444);
and (n440,n7,n441);
xor (n441,n442,n443);
and (n444,n7,n445);
nor (n445,n441,n446);
xnor (n446,n166,n442);
xor (n447,n448,n170);
or (n448,n163,n449);
and (n449,n30,n168);
nand (n450,n451,n447);
xor (n451,n452,n75);
or (n452,n453,n454);
and (n453,n65,n98);
and (n454,n112,n102);
nand (n455,n437,n451);
nand (n456,n457,n462,n467);
nand (n457,n458,n438);
xor (n458,n459,n100);
or (n459,n460,n461);
and (n460,n44,n174);
and (n461,n63,n177);
nand (n462,n463,n438);
xor (n463,n464,n23);
or (n464,n465,n466);
and (n465,n195,n73);
and (n466,n197,n77);
nand (n467,n458,n463);
nand (n468,n469,n488,n501);
nand (n469,n470,n472);
xor (n470,n471,n451);
xor (n471,n437,n447);
nand (n472,n473,n482,n487);
nand (n473,n474,n478);
xor (n474,n475,n170);
or (n475,n476,n477);
and (n476,n30,n164);
and (n477,n44,n168);
xor (n478,n479,n75);
or (n479,n480,n481);
and (n480,n112,n98);
and (n481,n195,n102);
nand (n482,n483,n478);
xor (n483,n484,n100);
or (n484,n485,n486);
and (n485,n63,n174);
and (n486,n65,n177);
nand (n487,n474,n483);
nand (n488,n489,n472);
nand (n489,n490,n495,n500);
nand (n490,n437,n491);
xor (n491,n492,n23);
or (n492,n493,n494);
and (n493,n197,n73);
and (n494,n213,n77);
nand (n495,n496,n491);
xor (n496,n497,n10);
or (n497,n498,n499);
and (n498,n267,n21);
and (n499,n299,n25);
nand (n500,n437,n496);
nand (n501,n470,n489);
nand (n502,n503,n508,n539);
nand (n503,n504,n506);
xor (n504,n505,n14);
xor (n505,n420,n424);
xor (n506,n507,n463);
xor (n507,n458,n438);
nand (n508,n509,n506);
nand (n509,n510,n516,n538);
nand (n510,n511,n14);
xor (n511,n512,n14);
or (n512,n513,n514);
and (n513,n428,n8);
and (n514,n515,n12);
nand (n516,n517,n14);
nand (n517,n518,n532,n537);
nand (n518,n519,n529);
not (n519,n520);
xor (n520,n521,n443);
or (n521,n522,n526);
and (n522,n7,n523);
xor (n523,n524,n525);
and (n526,n7,n527);
nor (n527,n523,n528);
xnor (n528,n443,n524);
xor (n529,n530,n166);
or (n530,n440,n531);
and (n531,n30,n445);
nand (n532,n533,n529);
xor (n533,n534,n170);
or (n534,n535,n536);
and (n535,n44,n164);
and (n536,n63,n168);
nand (n537,n519,n533);
nand (n538,n511,n517);
nand (n539,n504,n509);
nand (n540,n541,n579,n582);
nand (n541,n542,n577);
nand (n542,n543,n563,n576);
nand (n543,n544,n546);
xor (n544,n545,n483);
xor (n545,n474,n478);
nand (n546,n547,n556,n562);
nand (n547,n548,n552);
xor (n548,n549,n100);
or (n549,n550,n551);
and (n550,n65,n174);
and (n551,n112,n177);
xor (n552,n553,n75);
or (n553,n554,n555);
and (n554,n195,n98);
and (n555,n197,n102);
nand (n556,n557,n552);
xor (n557,n558,n14);
or (n558,n559,n560);
and (n559,n515,n8);
and (n560,n561,n12);
nand (n562,n548,n557);
nand (n563,n564,n546);
nand (n564,n565,n570,n575);
nand (n565,n520,n566);
xor (n566,n567,n23);
or (n567,n568,n569);
and (n568,n213,n73);
and (n569,n267,n77);
nand (n570,n571,n566);
xor (n571,n572,n10);
or (n572,n573,n574);
and (n573,n299,n21);
and (n574,n428,n25);
nand (n575,n520,n571);
nand (n576,n544,n564);
xor (n577,n578,n489);
xor (n578,n470,n472);
nand (n579,n580,n577);
xor (n580,n581,n509);
xor (n581,n504,n506);
nand (n582,n542,n580);
nand (n583,n584,n616,n705);
nand (n584,n585,n614);
nand (n585,n586,n590,n613);
nand (n586,n587,n589);
xor (n587,n588,n496);
xor (n588,n437,n491);
xor (n589,n512,n517);
nand (n590,n591,n589);
nand (n591,n592,n595,n612);
nand (n592,n14,n593);
xor (n593,n594,n533);
xor (n594,n519,n529);
nand (n595,n596,n593);
nand (n596,n597,n606,n611);
nand (n597,n598,n602);
xor (n598,n599,n166);
or (n599,n600,n601);
and (n600,n30,n441);
and (n601,n44,n445);
xor (n602,n603,n170);
or (n603,n604,n605);
and (n604,n63,n164);
and (n605,n65,n168);
nand (n606,n607,n602);
xor (n607,n608,n100);
or (n608,n609,n610);
and (n609,n112,n174);
and (n610,n195,n177);
nand (n611,n598,n607);
nand (n612,n14,n596);
nand (n613,n587,n591);
xor (n614,n615,n580);
xor (n615,n542,n577);
nand (n616,n617,n614);
nand (n617,n618,n642,n704);
nand (n618,n619,n621);
xor (n619,n620,n564);
xor (n620,n544,n546);
nand (n621,n622,n638,n641);
nand (n622,n623,n636);
nand (n623,n624,n634,n635);
nand (n624,n625,n629);
xor (n625,n626,n75);
or (n626,n627,n628);
and (n627,n197,n98);
and (n628,n213,n102);
xor (n629,n630,n14);
or (n630,n631,n632);
and (n631,n561,n8);
and (n632,n633,n12);
nand (n634,n519,n629);
nand (n635,n625,n519);
xor (n636,n637,n557);
xor (n637,n548,n552);
nand (n638,n639,n636);
xor (n639,n640,n571);
xor (n640,n520,n566);
nand (n641,n623,n639);
nand (n642,n643,n621);
nand (n643,n644,n700,n703);
nand (n644,n645,n678);
nand (n645,n646,n655,n677);
nand (n646,n647,n651);
xor (n647,n648,n23);
or (n648,n649,n650);
and (n649,n267,n73);
and (n650,n299,n77);
xor (n651,n652,n10);
or (n652,n653,n654);
and (n653,n428,n21);
and (n654,n515,n25);
nand (n655,n656,n651);
nand (n656,n657,n671,n676);
nand (n657,n658,n668);
not (n658,n659);
xor (n659,n660,n525);
or (n660,n661,n665);
and (n661,n7,n662);
xor (n662,n663,n664);
and (n665,n7,n666);
nor (n666,n662,n667);
xnor (n667,n525,n663);
xor (n668,n669,n443);
or (n669,n522,n670);
and (n670,n30,n527);
nand (n671,n672,n668);
xor (n672,n673,n170);
or (n673,n674,n675);
and (n674,n65,n164);
and (n675,n112,n168);
nand (n676,n658,n672);
nand (n677,n647,n656);
nand (n678,n679,n682,n699);
nand (n679,n14,n680);
xor (n680,n681,n607);
xor (n681,n598,n602);
nand (n682,n683,n680);
nand (n683,n684,n693,n698);
nand (n684,n685,n689);
xor (n685,n686,n166);
or (n686,n687,n688);
and (n687,n44,n441);
and (n688,n63,n445);
xor (n689,n690,n100);
or (n690,n691,n692);
and (n691,n195,n174);
and (n692,n197,n177);
nand (n693,n694,n689);
xor (n694,n695,n75);
or (n695,n696,n697);
and (n696,n213,n98);
and (n697,n267,n102);
nand (n698,n685,n694);
nand (n699,n14,n683);
nand (n700,n701,n678);
xor (n701,n702,n596);
xor (n702,n14,n593);
nand (n703,n645,n701);
nand (n704,n619,n643);
nand (n705,n585,n617);
nor (n706,n707,n711);
nand (n707,n708,n709,n710);
nand (n708,n412,n431);
nand (n709,n540,n431);
nand (n710,n412,n540);
xor (n711,n712,n726);
xor (n712,n713,n717);
nand (n713,n714,n715,n716);
nand (n714,n414,n416);
nand (n715,n418,n416);
nand (n716,n414,n418);
xor (n717,n718,n724);
xor (n718,n719,n723);
nand (n719,n720,n721,n722);
nand (n720,n14,n435);
nand (n721,n456,n435);
nand (n722,n14,n456);
xor (n723,n264,n269);
xor (n724,n725,n305);
xor (n725,n289,n302);
nand (n726,n727,n728,n729);
nand (n727,n433,n468);
nand (n728,n502,n468);
nand (n729,n433,n502);
nor (n730,n731,n746);
nor (n731,n732,n736);
nand (n732,n733,n734,n735);
nand (n733,n713,n717);
nand (n734,n726,n717);
nand (n735,n713,n726);
xor (n736,n737,n742);
xor (n737,n738,n740);
xor (n738,n739,n200);
xor (n739,n158,n185);
xor (n740,n741,n287);
xor (n741,n259,n261);
nand (n742,n743,n744,n745);
nand (n743,n719,n723);
nand (n744,n724,n723);
nand (n745,n719,n724);
nor (n746,n747,n751);
nand (n747,n748,n749,n750);
nand (n748,n738,n740);
nand (n749,n742,n740);
nand (n750,n738,n742);
xor (n751,n752,n257);
xor (n752,n156,n215);
nor (n753,n754,n1154);
nor (n754,n755,n1130);
nor (n755,n756,n1128);
nor (n756,n757,n1103);
nand (n757,n758,n1065);
nand (n758,n759,n981,n1064);
nand (n759,n760,n844);
xor (n760,n761,n834);
xor (n761,n762,n784);
xor (n762,n763,n768);
xor (n763,n764,n14);
xor (n764,n765,n23);
or (n765,n766,n767);
and (n766,n299,n73);
and (n767,n428,n77);
nand (n768,n769,n778,n783);
nand (n769,n770,n774);
xor (n770,n771,n170);
or (n771,n772,n773);
and (n772,n112,n164);
and (n773,n195,n168);
xor (n774,n775,n443);
or (n775,n776,n777);
and (n776,n30,n523);
and (n777,n44,n527);
nand (n778,n779,n774);
xor (n779,n780,n166);
or (n780,n781,n782);
and (n781,n63,n441);
and (n782,n65,n445);
nand (n783,n770,n779);
nand (n784,n785,n816,n833);
nand (n785,n786,n802);
nand (n786,n787,n796,n801);
nand (n787,n788,n792);
xor (n788,n789,n170);
or (n789,n790,n791);
and (n790,n195,n164);
and (n791,n197,n168);
xor (n792,n793,n443);
or (n793,n794,n795);
and (n794,n44,n523);
and (n795,n63,n527);
nand (n796,n797,n792);
xor (n797,n798,n100);
or (n798,n799,n800);
and (n799,n213,n174);
and (n800,n267,n177);
nand (n801,n788,n797);
xor (n802,n803,n812);
xor (n803,n804,n808);
xor (n804,n805,n100);
or (n805,n806,n807);
and (n806,n197,n174);
and (n807,n213,n177);
xor (n808,n809,n75);
or (n809,n810,n811);
and (n810,n267,n98);
and (n811,n299,n102);
xor (n812,n813,n10);
or (n813,n814,n815);
and (n814,n561,n21);
and (n815,n633,n25);
nand (n816,n817,n802);
nand (n817,n818,n827,n832);
nand (n818,n819,n823);
xor (n819,n820,n525);
or (n820,n821,n822);
and (n821,n30,n662);
and (n822,n44,n666);
xor (n823,n824,n75);
or (n824,n825,n826);
and (n825,n299,n98);
and (n826,n428,n102);
nand (n827,n828,n823);
xor (n828,n829,n23);
or (n829,n830,n831);
and (n830,n515,n73);
and (n831,n561,n77);
nand (n832,n819,n828);
nand (n833,n786,n817);
xor (n834,n835,n840);
xor (n835,n836,n838);
xor (n836,n837,n672);
xor (n837,n658,n668);
xor (n838,n839,n694);
xor (n839,n685,n689);
nand (n840,n841,n842,n843);
nand (n841,n804,n808);
nand (n842,n812,n808);
nand (n843,n804,n812);
xor (n844,n845,n920);
xor (n845,n846,n900);
nand (n846,n847,n873,n899);
nand (n847,n848,n863);
nand (n848,n849,n861,n862);
nand (n849,n850,n855);
xor (n850,n851,n10);
or (n851,n852,n853);
and (n852,n633,n21);
and (n853,n854,n25);
xor (n855,n856,n14);
or (n856,n857,n859);
and (n857,n858,n8);
and (n859,n860,n12);
nand (n861,n14,n855);
nand (n862,n850,n14);
xor (n863,n864,n869);
xor (n864,n865,n658);
xor (n865,n866,n14);
or (n866,n867,n868);
and (n867,n854,n8);
and (n868,n858,n12);
xor (n869,n870,n23);
or (n870,n871,n872);
and (n871,n428,n73);
and (n872,n515,n77);
nand (n873,n874,n863);
xor (n874,n875,n897);
xor (n875,n14,n876);
nand (n876,n877,n891,n896);
nand (n877,n878,n881);
xor (n878,n879,n525);
or (n879,n661,n880);
and (n880,n30,n666);
not (n881,n882);
xor (n882,n883,n664);
or (n883,n884,n888);
and (n884,n7,n885);
xor (n885,n886,n887);
and (n888,n7,n889);
nor (n889,n885,n890);
xnor (n890,n664,n886);
nand (n891,n892,n881);
xor (n892,n893,n166);
or (n893,n894,n895);
and (n894,n65,n441);
and (n895,n112,n445);
nand (n896,n878,n892);
xor (n897,n898,n779);
xor (n898,n770,n774);
nand (n899,n848,n874);
xor (n900,n901,n916);
xor (n901,n902,n906);
nand (n902,n903,n904,n905);
nand (n903,n865,n658);
nand (n904,n869,n658);
nand (n905,n865,n869);
xor (n906,n907,n659);
xor (n907,n908,n912);
xor (n908,n909,n10);
or (n909,n910,n911);
and (n910,n515,n21);
and (n911,n561,n25);
xor (n912,n913,n14);
or (n913,n914,n915);
and (n914,n633,n8);
and (n915,n854,n12);
nand (n916,n917,n918,n919);
nand (n917,n14,n876);
nand (n918,n897,n876);
nand (n919,n14,n897);
nand (n920,n921,n977,n980);
nand (n921,n922,n942);
nand (n922,n923,n938,n941);
nand (n923,n924,n936);
nand (n924,n925,n930,n935);
nand (n925,n882,n926);
xor (n926,n927,n166);
or (n927,n928,n929);
and (n928,n112,n441);
and (n929,n195,n445);
nand (n930,n931,n926);
xor (n931,n932,n170);
or (n932,n933,n934);
and (n933,n197,n164);
and (n934,n213,n168);
nand (n935,n882,n931);
xor (n936,n937,n797);
xor (n937,n788,n792);
nand (n938,n939,n936);
xor (n939,n940,n892);
xor (n940,n878,n881);
nand (n941,n924,n939);
nand (n942,n943,n973,n976);
nand (n943,n944,n957);
nand (n944,n945,n951,n956);
nand (n945,n946,n950);
xor (n946,n947,n443);
or (n947,n948,n949);
and (n948,n63,n523);
and (n949,n65,n527);
not (n950,n819);
nand (n951,n952,n950);
xor (n952,n953,n100);
or (n953,n954,n955);
and (n954,n267,n174);
and (n955,n299,n177);
nand (n956,n946,n952);
nand (n957,n958,n967,n972);
nand (n958,n959,n963);
xor (n959,n960,n75);
or (n960,n961,n962);
and (n961,n428,n98);
and (n962,n515,n102);
xor (n963,n964,n23);
or (n964,n965,n966);
and (n965,n561,n73);
and (n966,n633,n77);
nand (n967,n968,n963);
xor (n968,n969,n10);
or (n969,n970,n971);
and (n970,n854,n21);
and (n971,n858,n25);
nand (n972,n959,n968);
nand (n973,n974,n957);
xor (n974,n975,n828);
xor (n975,n819,n823);
nand (n976,n944,n974);
nand (n977,n978,n942);
xor (n978,n979,n817);
xor (n979,n786,n802);
nand (n980,n922,n978);
nand (n981,n982,n844);
nand (n982,n983,n1060,n1063);
nand (n983,n984,n986);
xor (n984,n985,n874);
xor (n985,n848,n863);
nand (n986,n987,n1020,n1059);
nand (n987,n988,n1018);
nand (n988,n989,n995,n1017);
nand (n989,n990,n14);
xor (n990,n991,n14);
or (n991,n992,n993);
and (n992,n860,n8);
and (n993,n994,n12);
nand (n995,n996,n14);
nand (n996,n997,n1005,n1016);
nand (n997,n998,n1001);
xor (n998,n999,n664);
or (n999,n884,n1000);
and (n1000,n30,n889);
xor (n1001,n1002,n525);
or (n1002,n1003,n1004);
and (n1003,n44,n662);
and (n1004,n63,n666);
nand (n1005,n1006,n1001);
not (n1006,n1007);
xor (n1007,n1008,n887);
or (n1008,n1009,n1013);
and (n1009,n7,n1010);
xor (n1010,n1011,n1012);
and (n1013,n7,n1014);
nor (n1014,n1010,n1015);
xnor (n1015,n887,n1011);
nand (n1016,n998,n1006);
nand (n1017,n990,n996);
xor (n1018,n1019,n14);
xor (n1019,n850,n855);
nand (n1020,n1021,n1018);
nand (n1021,n1022,n1041,n1058);
nand (n1022,n1023,n1039);
nand (n1023,n1024,n1033,n1038);
nand (n1024,n1025,n1029);
xor (n1025,n1026,n443);
or (n1026,n1027,n1028);
and (n1027,n65,n523);
and (n1028,n112,n527);
xor (n1029,n1030,n166);
or (n1030,n1031,n1032);
and (n1031,n195,n441);
and (n1032,n197,n445);
nand (n1033,n1034,n1029);
xor (n1034,n1035,n170);
or (n1035,n1036,n1037);
and (n1036,n213,n164);
and (n1037,n267,n168);
nand (n1038,n1025,n1034);
xor (n1039,n1040,n931);
xor (n1040,n882,n926);
nand (n1041,n1042,n1039);
nand (n1042,n1043,n1052,n1057);
nand (n1043,n1044,n1048);
xor (n1044,n1045,n75);
or (n1045,n1046,n1047);
and (n1046,n515,n98);
and (n1047,n561,n102);
xor (n1048,n1049,n664);
or (n1049,n1050,n1051);
and (n1050,n30,n885);
and (n1051,n44,n889);
nand (n1052,n1053,n1048);
xor (n1053,n1054,n100);
or (n1054,n1055,n1056);
and (n1055,n299,n174);
and (n1056,n428,n177);
nand (n1057,n1044,n1053);
nand (n1058,n1023,n1042);
nand (n1059,n988,n1021);
nand (n1060,n1061,n986);
xor (n1061,n1062,n978);
xor (n1062,n922,n942);
nand (n1063,n984,n1061);
nand (n1064,n760,n982);
xor (n1065,n1066,n1099);
xor (n1066,n1067,n1071);
nand (n1067,n1068,n1069,n1070);
nand (n1068,n762,n784);
nand (n1069,n834,n784);
nand (n1070,n762,n834);
xor (n1071,n1072,n1087);
xor (n1072,n1073,n1077);
nand (n1073,n1074,n1075,n1076);
nand (n1074,n902,n906);
nand (n1075,n916,n906);
nand (n1076,n902,n916);
xor (n1077,n1078,n1085);
xor (n1078,n1079,n1083);
nand (n1079,n1080,n1081,n1082);
nand (n1080,n908,n912);
nand (n1081,n659,n912);
nand (n1082,n908,n659);
xor (n1083,n1084,n656);
xor (n1084,n647,n651);
xor (n1085,n1086,n519);
xor (n1086,n625,n629);
xor (n1087,n1088,n1095);
xor (n1088,n1089,n1093);
nand (n1089,n1090,n1091,n1092);
nand (n1090,n764,n14);
nand (n1091,n768,n14);
nand (n1092,n764,n768);
xor (n1093,n1094,n683);
xor (n1094,n14,n680);
nand (n1095,n1096,n1097,n1098);
nand (n1096,n836,n838);
nand (n1097,n840,n838);
nand (n1098,n836,n840);
nand (n1099,n1100,n1101,n1102);
nand (n1100,n846,n900);
nand (n1101,n920,n900);
nand (n1102,n846,n920);
nor (n1103,n1104,n1108);
nand (n1104,n1105,n1106,n1107);
nand (n1105,n1067,n1071);
nand (n1106,n1099,n1071);
nand (n1107,n1067,n1099);
xor (n1108,n1109,n1124);
xor (n1109,n1110,n1112);
xor (n1110,n1111,n701);
xor (n1111,n645,n678);
xor (n1112,n1113,n1120);
xor (n1113,n1114,n1116);
xor (n1114,n1115,n639);
xor (n1115,n623,n636);
nand (n1116,n1117,n1118,n1119);
nand (n1117,n1079,n1083);
nand (n1118,n1085,n1083);
nand (n1119,n1079,n1085);
nand (n1120,n1121,n1122,n1123);
nand (n1121,n1089,n1093);
nand (n1122,n1095,n1093);
nand (n1123,n1089,n1095);
nand (n1124,n1125,n1126,n1127);
nand (n1125,n1073,n1077);
nand (n1126,n1087,n1077);
nand (n1127,n1073,n1087);
not (n1128,n1129);
nand (n1129,n1104,n1108);
not (n1130,n1131);
nor (n1131,n1132,n1147);
nor (n1132,n1133,n1137);
nand (n1133,n1134,n1135,n1136);
nand (n1134,n1110,n1112);
nand (n1135,n1124,n1112);
nand (n1136,n1110,n1124);
xor (n1137,n1138,n1143);
xor (n1138,n1139,n1141);
xor (n1139,n1140,n591);
xor (n1140,n587,n589);
xor (n1141,n1142,n643);
xor (n1142,n619,n621);
nand (n1143,n1144,n1145,n1146);
nand (n1144,n1114,n1116);
nand (n1145,n1120,n1116);
nand (n1146,n1114,n1120);
nor (n1147,n1148,n1152);
nand (n1148,n1149,n1150,n1151);
nand (n1149,n1139,n1141);
nand (n1150,n1143,n1141);
nand (n1151,n1139,n1143);
xor (n1152,n1153,n617);
xor (n1153,n585,n614);
not (n1154,n1155);
nor (n1155,n1156,n1158);
nor (n1156,n1157,n1147);
nand (n1157,n1133,n1137);
not (n1158,n1159);
nand (n1159,n1148,n1152);
not (n1160,n1161);
nor (n1161,n1162,n1169);
nor (n1162,n1163,n1168);
nor (n1163,n1164,n1166);
nor (n1164,n1165,n706);
nand (n1165,n410,n583);
not (n1166,n1167);
nand (n1167,n707,n711);
not (n1168,n730);
not (n1169,n1170);
nor (n1170,n1171,n1173);
nor (n1171,n1172,n746);
nand (n1172,n732,n736);
not (n1173,n1174);
nand (n1174,n747,n751);
nand (n1175,n1176,n1180);
nor (n1176,n1177,n407);
nand (n1177,n1178,n1131);
nor (n1178,n1179,n1103);
nor (n1179,n758,n1065);
nand (n1180,n1181,n2711);
nor (n1181,n1182,n2679);
nor (n1182,n1183,n2152);
nor (n1183,n1184,n2137);
nor (n1184,n1185,n1858);
nand (n1185,n1186,n1641);
nor (n1186,n1187,n1540);
nor (n1187,n1188,n1450);
nand (n1188,n1189,n1365,n1449);
nand (n1189,n1190,n1267);
xor (n1190,n1191,n1243);
xor (n1191,n1192,n1217);
xor (n1192,n1193,n1205);
xor (n1193,n1194,n1199);
xor (n1194,n1195,n100);
or (n1195,n1196,n1197);
and (n1196,n994,n174);
and (n1197,n1198,n177);
xor (n1199,n1200,n75);
or (n1200,n1201,n1203);
and (n1201,n1202,n98);
and (n1203,n1204,n102);
xor (n1205,n1206,n1210);
xor (n1206,n1207,n887);
or (n1207,n1208,n1209);
and (n1208,n195,n1010);
and (n1209,n197,n1014);
xnor (n1210,n1211,n1012);
nor (n1211,n1212,n1216);
and (n1212,n112,n1213);
and (n1213,n1214,n1012);
not (n1214,n1215);
and (n1216,n65,n1215);
nand (n1217,n1218,n1228,n1242);
nand (n1218,n1219,n1223);
xor (n1219,n1220,n100);
or (n1220,n1221,n1222);
and (n1221,n1198,n174);
and (n1222,n1202,n177);
xor (n1223,n1224,n75);
or (n1224,n1225,n1226);
and (n1225,n1204,n98);
and (n1226,n1227,n102);
nand (n1228,n1229,n1223);
xor (n1229,n1230,n1239);
xor (n1230,n1231,n1235);
xor (n1231,n1232,n887);
or (n1232,n1233,n1234);
and (n1233,n197,n1010);
and (n1234,n213,n1014);
xor (n1235,n1236,n525);
or (n1236,n1237,n1238);
and (n1237,n428,n662);
and (n1238,n515,n666);
xnor (n1239,n1240,n23);
nand (n1240,n1241,n73);
nand (n1242,n1219,n1229);
xor (n1243,n1244,n1253);
xor (n1244,n1245,n1249);
xor (n1245,n1246,n23);
or (n1246,n1247,n1248);
and (n1247,n1227,n73);
and (n1248,n1241,n77);
nand (n1249,n1250,n1251,n1252);
nand (n1250,n1231,n1235);
nand (n1251,n1239,n1235);
nand (n1252,n1231,n1239);
xor (n1253,n1254,n1263);
xor (n1254,n1255,n1259);
xor (n1255,n1256,n525);
or (n1256,n1257,n1258);
and (n1257,n299,n662);
and (n1258,n428,n666);
xor (n1259,n1260,n664);
or (n1260,n1261,n1262);
and (n1261,n213,n885);
and (n1262,n267,n889);
xor (n1263,n1264,n443);
or (n1264,n1265,n1266);
and (n1265,n515,n523);
and (n1266,n561,n527);
nand (n1267,n1268,n1322,n1364);
nand (n1268,n1269,n1271);
xor (n1269,n1270,n1229);
xor (n1270,n1219,n1223);
xor (n1271,n1272,n1311);
xor (n1272,n1273,n1289);
nand (n1273,n1274,n1283,n1288);
nand (n1274,n1275,n1279);
xor (n1275,n1276,n525);
or (n1276,n1277,n1278);
and (n1277,n515,n662);
and (n1278,n561,n666);
xor (n1279,n1280,n664);
or (n1280,n1281,n1282);
and (n1281,n299,n885);
and (n1282,n428,n889);
nand (n1283,n1284,n1279);
xor (n1284,n1285,n443);
or (n1285,n1286,n1287);
and (n1286,n633,n523);
and (n1287,n854,n527);
nand (n1288,n1275,n1284);
nand (n1289,n1290,n1305,n1310);
nand (n1290,n1291,n1300);
xor (n1291,n1292,n1296);
xnor (n1292,n1293,n1012);
nor (n1293,n1294,n1295);
and (n1294,n197,n1213);
and (n1295,n195,n1215);
xor (n1296,n1297,n887);
or (n1297,n1298,n1299);
and (n1298,n213,n1010);
and (n1299,n267,n1014);
and (n1300,n1301,n75);
xnor (n1301,n1302,n1012);
nor (n1302,n1303,n1304);
and (n1303,n213,n1213);
and (n1304,n197,n1215);
nand (n1305,n1306,n1300);
xor (n1306,n1307,n166);
or (n1307,n1308,n1309);
and (n1308,n858,n441);
and (n1309,n860,n445);
nand (n1310,n1291,n1306);
xor (n1311,n1312,n1318);
xor (n1312,n1313,n1317);
xor (n1313,n1314,n166);
or (n1314,n1315,n1316);
and (n1315,n854,n441);
and (n1316,n858,n445);
and (n1317,n1292,n1296);
xor (n1318,n1319,n170);
or (n1319,n1320,n1321);
and (n1320,n860,n164);
and (n1321,n994,n168);
nand (n1322,n1323,n1271);
nand (n1323,n1324,n1348,n1363);
nand (n1324,n1325,n1346);
nand (n1325,n1326,n1340,n1345);
nand (n1326,n1327,n1336);
and (n1327,n1328,n1332);
xnor (n1328,n1329,n1012);
nor (n1329,n1330,n1331);
and (n1330,n267,n1213);
and (n1331,n213,n1215);
xor (n1332,n1333,n887);
or (n1333,n1334,n1335);
and (n1334,n299,n1010);
and (n1335,n428,n1014);
xor (n1336,n1337,n166);
or (n1337,n1338,n1339);
and (n1338,n860,n441);
and (n1339,n994,n445);
nand (n1340,n1341,n1336);
xor (n1341,n1342,n170);
or (n1342,n1343,n1344);
and (n1343,n1198,n164);
and (n1344,n1202,n168);
nand (n1345,n1327,n1341);
xor (n1346,n1347,n1306);
xor (n1347,n1291,n1300);
nand (n1348,n1349,n1346);
xor (n1349,n1350,n1359);
xor (n1350,n1351,n1355);
xor (n1351,n1352,n170);
or (n1352,n1353,n1354);
and (n1353,n994,n164);
and (n1354,n1198,n168);
xor (n1355,n1356,n100);
or (n1356,n1357,n1358);
and (n1357,n1202,n174);
and (n1358,n1204,n177);
xor (n1359,n1360,n75);
or (n1360,n1361,n1362);
and (n1361,n1227,n98);
and (n1362,n1241,n102);
nand (n1363,n1325,n1349);
nand (n1364,n1269,n1323);
nand (n1365,n1366,n1267);
xor (n1366,n1367,n1406);
xor (n1367,n1368,n1372);
nand (n1368,n1369,n1370,n1371);
nand (n1369,n1273,n1289);
nand (n1370,n1311,n1289);
nand (n1371,n1273,n1311);
xor (n1372,n1373,n1395);
xor (n1373,n1374,n1391);
nand (n1374,n1375,n1385,n1390);
nand (n1375,n1376,n1380);
xor (n1376,n1377,n664);
or (n1377,n1378,n1379);
and (n1378,n267,n885);
and (n1379,n299,n889);
xor (n1380,n1381,n23);
xnor (n1381,n1382,n1012);
nor (n1382,n1383,n1384);
and (n1383,n195,n1213);
and (n1384,n112,n1215);
nand (n1385,n1386,n1380);
xor (n1386,n1387,n443);
or (n1387,n1388,n1389);
and (n1388,n561,n523);
and (n1389,n633,n527);
nand (n1390,n1376,n1386);
nand (n1391,n1392,n1393,n1394);
nand (n1392,n1313,n1317);
nand (n1393,n1318,n1317);
nand (n1394,n1313,n1318);
xor (n1395,n1396,n1402);
xor (n1396,n1397,n1398);
and (n1397,n1381,n23);
xor (n1398,n1399,n166);
or (n1399,n1400,n1401);
and (n1400,n633,n441);
and (n1401,n854,n445);
xor (n1402,n1403,n170);
or (n1403,n1404,n1405);
and (n1404,n858,n164);
and (n1405,n860,n168);
nand (n1406,n1407,n1414,n1448);
nand (n1407,n1408,n1412);
nand (n1408,n1409,n1410,n1411);
nand (n1409,n1351,n1355);
nand (n1410,n1359,n1355);
nand (n1411,n1351,n1359);
xor (n1412,n1413,n1386);
xor (n1413,n1376,n1380);
nand (n1414,n1415,n1412);
nand (n1415,n1416,n1433,n1447);
nand (n1416,n1417,n1431);
nand (n1417,n1418,n1427,n1430);
nand (n1418,n1419,n1423);
xor (n1419,n1420,n887);
or (n1420,n1421,n1422);
and (n1421,n267,n1010);
and (n1422,n299,n1014);
xor (n1423,n1424,n525);
or (n1424,n1425,n1426);
and (n1425,n561,n662);
and (n1426,n633,n666);
nand (n1427,n1428,n1423);
xnor (n1428,n1429,n75);
nand (n1429,n1241,n98);
nand (n1430,n1419,n1428);
xor (n1431,n1432,n1284);
xor (n1432,n1275,n1279);
nand (n1433,n1434,n1431);
nand (n1434,n1435,n1441,n1446);
nand (n1435,n1436,n1440);
xor (n1436,n1437,n664);
or (n1437,n1438,n1439);
and (n1438,n428,n885);
and (n1439,n515,n889);
xor (n1440,n1301,n75);
nand (n1441,n1442,n1440);
xor (n1442,n1443,n443);
or (n1443,n1444,n1445);
and (n1444,n854,n523);
and (n1445,n858,n527);
nand (n1446,n1436,n1442);
nand (n1447,n1417,n1434);
nand (n1448,n1408,n1415);
nand (n1449,n1190,n1366);
xor (n1450,n1451,n1536);
xor (n1451,n1452,n1473);
xor (n1452,n1453,n1469);
xor (n1453,n1454,n1465);
xor (n1454,n1455,n1461);
xor (n1455,n1456,n1460);
xor (n1456,n1457,n75);
or (n1457,n1458,n1459);
and (n1458,n1198,n98);
and (n1459,n1202,n102);
and (n1460,n1206,n1210);
xor (n1461,n1462,n23);
or (n1462,n1463,n1464);
and (n1463,n1204,n73);
and (n1464,n1227,n77);
nand (n1465,n1466,n1467,n1468);
nand (n1466,n1245,n1249);
nand (n1467,n1253,n1249);
nand (n1468,n1245,n1253);
nand (n1469,n1470,n1471,n1472);
nand (n1470,n1374,n1391);
nand (n1471,n1395,n1391);
nand (n1472,n1374,n1395);
xor (n1473,n1474,n1532);
xor (n1474,n1475,n1499);
xor (n1475,n1476,n1495);
xor (n1476,n1477,n1481);
nand (n1477,n1478,n1479,n1480);
nand (n1478,n1397,n1398);
nand (n1479,n1402,n1398);
nand (n1480,n1397,n1402);
xor (n1481,n1482,n1491);
xor (n1482,n1483,n1487);
xnor (n1483,n1484,n1012);
nor (n1484,n1485,n1486);
and (n1485,n65,n1213);
and (n1486,n63,n1215);
xor (n1487,n1488,n525);
or (n1488,n1489,n1490);
and (n1489,n267,n662);
and (n1490,n299,n666);
xor (n1491,n1492,n664);
or (n1492,n1493,n1494);
and (n1493,n197,n885);
and (n1494,n213,n889);
nand (n1495,n1496,n1497,n1498);
nand (n1496,n1255,n1259);
nand (n1497,n1263,n1259);
nand (n1498,n1255,n1263);
xor (n1499,n1500,n1518);
xor (n1500,n1501,n1505);
nand (n1501,n1502,n1503,n1504);
nand (n1502,n1194,n1199);
nand (n1503,n1205,n1199);
nand (n1504,n1194,n1205);
xor (n1505,n1506,n1516);
xor (n1506,n1507,n1511);
xor (n1507,n1508,n443);
or (n1508,n1509,n1510);
and (n1509,n428,n523);
and (n1510,n515,n527);
xor (n1511,n10,n1512);
xor (n1512,n1513,n887);
or (n1513,n1514,n1515);
and (n1514,n112,n1010);
and (n1515,n195,n1014);
xnor (n1516,n1517,n10);
nand (n1517,n1241,n21);
xor (n1518,n1519,n1528);
xor (n1519,n1520,n1524);
xor (n1520,n1521,n166);
or (n1521,n1522,n1523);
and (n1522,n561,n441);
and (n1523,n633,n445);
xor (n1524,n1525,n170);
or (n1525,n1526,n1527);
and (n1526,n854,n164);
and (n1527,n858,n168);
xor (n1528,n1529,n100);
or (n1529,n1530,n1531);
and (n1530,n860,n174);
and (n1531,n994,n177);
nand (n1532,n1533,n1534,n1535);
nand (n1533,n1192,n1217);
nand (n1534,n1243,n1217);
nand (n1535,n1192,n1243);
nand (n1536,n1537,n1538,n1539);
nand (n1537,n1368,n1372);
nand (n1538,n1406,n1372);
nand (n1539,n1368,n1406);
nor (n1540,n1541,n1545);
nand (n1541,n1542,n1543,n1544);
nand (n1542,n1452,n1473);
nand (n1543,n1536,n1473);
nand (n1544,n1452,n1536);
xor (n1545,n1546,n1555);
xor (n1546,n1547,n1551);
nand (n1547,n1548,n1549,n1550);
nand (n1548,n1454,n1465);
nand (n1549,n1469,n1465);
nand (n1550,n1454,n1469);
nand (n1551,n1552,n1553,n1554);
nand (n1552,n1475,n1499);
nand (n1553,n1532,n1499);
nand (n1554,n1475,n1532);
xor (n1555,n1556,n1617);
xor (n1556,n1557,n1588);
xor (n1557,n1558,n1577);
xor (n1558,n1559,n1573);
xor (n1559,n1560,n1569);
xor (n1560,n1561,n1565);
xor (n1561,n1562,n525);
or (n1562,n1563,n1564);
and (n1563,n213,n662);
and (n1564,n267,n666);
xor (n1565,n1566,n664);
or (n1566,n1567,n1568);
and (n1567,n195,n885);
and (n1568,n197,n889);
xor (n1569,n1570,n443);
or (n1570,n1571,n1572);
and (n1571,n299,n523);
and (n1572,n428,n527);
nand (n1573,n1574,n1575,n1576);
nand (n1574,n1507,n1511);
nand (n1575,n1516,n1511);
nand (n1576,n1507,n1516);
xor (n1577,n1578,n1584);
xor (n1578,n1579,n1583);
xor (n1579,n1580,n166);
or (n1580,n1581,n1582);
and (n1581,n515,n441);
and (n1582,n561,n445);
and (n1583,n10,n1512);
xor (n1584,n1585,n170);
or (n1585,n1586,n1587);
and (n1586,n633,n164);
and (n1587,n854,n168);
xor (n1588,n1589,n1613);
xor (n1589,n1590,n1594);
nand (n1590,n1591,n1592,n1593);
nand (n1591,n1520,n1524);
nand (n1592,n1528,n1524);
nand (n1593,n1520,n1528);
xor (n1594,n1595,n1604);
xor (n1595,n1596,n1600);
xor (n1596,n1597,n100);
or (n1597,n1598,n1599);
and (n1598,n858,n174);
and (n1599,n860,n177);
xor (n1600,n1601,n75);
or (n1601,n1602,n1603);
and (n1602,n994,n98);
and (n1603,n1198,n102);
xor (n1604,n1605,n1609);
xnor (n1605,n1606,n1012);
nor (n1606,n1607,n1608);
and (n1607,n63,n1213);
and (n1608,n44,n1215);
xor (n1609,n1610,n887);
or (n1610,n1611,n1612);
and (n1611,n65,n1010);
and (n1612,n112,n1014);
nand (n1613,n1614,n1615,n1616);
nand (n1614,n1456,n1460);
nand (n1615,n1461,n1460);
nand (n1616,n1456,n1461);
xor (n1617,n1618,n1637);
xor (n1618,n1619,n1633);
xor (n1619,n1620,n1629);
xor (n1620,n1621,n1625);
xor (n1621,n1622,n23);
or (n1622,n1623,n1624);
and (n1623,n1202,n73);
and (n1624,n1204,n77);
xor (n1625,n1626,n10);
or (n1626,n1627,n1628);
and (n1627,n1227,n21);
and (n1628,n1241,n25);
nand (n1629,n1630,n1631,n1632);
nand (n1630,n1483,n1487);
nand (n1631,n1491,n1487);
nand (n1632,n1483,n1491);
nand (n1633,n1634,n1635,n1636);
nand (n1634,n1477,n1481);
nand (n1635,n1495,n1481);
nand (n1636,n1477,n1495);
nand (n1637,n1638,n1639,n1640);
nand (n1638,n1501,n1505);
nand (n1639,n1518,n1505);
nand (n1640,n1501,n1518);
nor (n1641,n1642,n1747);
nor (n1642,n1643,n1647);
nand (n1643,n1644,n1645,n1646);
nand (n1644,n1547,n1551);
nand (n1645,n1555,n1551);
nand (n1646,n1547,n1555);
xor (n1647,n1648,n1743);
xor (n1648,n1649,n1683);
xor (n1649,n1650,n1679);
xor (n1650,n1651,n1655);
nand (n1651,n1652,n1653,n1654);
nand (n1652,n1559,n1573);
nand (n1653,n1577,n1573);
nand (n1654,n1559,n1577);
xor (n1655,n1656,n1665);
xor (n1656,n1657,n1661);
xor (n1657,n1658,n10);
or (n1658,n1659,n1660);
and (n1659,n1204,n21);
and (n1660,n1227,n25);
nand (n1661,n1662,n1663,n1664);
nand (n1662,n1579,n1583);
nand (n1663,n1584,n1583);
nand (n1664,n1579,n1584);
xor (n1665,n1666,n1675);
xor (n1666,n1667,n1671);
xor (n1667,n1668,n525);
or (n1668,n1669,n1670);
and (n1669,n197,n662);
and (n1670,n213,n666);
xnor (n1671,n1672,n1012);
nor (n1672,n1673,n1674);
and (n1673,n44,n1213);
and (n1674,n30,n1215);
xor (n1675,n1676,n664);
or (n1676,n1677,n1678);
and (n1677,n112,n885);
and (n1678,n195,n889);
nand (n1679,n1680,n1681,n1682);
nand (n1680,n1590,n1594);
nand (n1681,n1613,n1594);
nand (n1682,n1590,n1613);
xor (n1683,n1684,n1739);
xor (n1684,n1685,n1707);
xor (n1685,n1686,n1695);
xor (n1686,n1687,n1691);
nand (n1687,n1688,n1689,n1690);
nand (n1688,n1561,n1565);
nand (n1689,n1569,n1565);
nand (n1690,n1561,n1569);
nand (n1691,n1692,n1693,n1694);
nand (n1692,n1596,n1600);
nand (n1693,n1604,n1600);
nand (n1694,n1596,n1604);
xor (n1695,n1696,n1703);
xor (n1696,n1697,n1701);
xor (n1697,n1698,n443);
or (n1698,n1699,n1700);
and (n1699,n267,n523);
and (n1700,n299,n527);
xnor (n1701,n1702,n14);
nand (n1702,n1241,n8);
xor (n1703,n1704,n166);
or (n1704,n1705,n1706);
and (n1705,n428,n441);
and (n1706,n515,n445);
xor (n1707,n1708,n1727);
xor (n1708,n1709,n1713);
nand (n1709,n1710,n1711,n1712);
nand (n1710,n1621,n1625);
nand (n1711,n1629,n1625);
nand (n1712,n1621,n1629);
xor (n1713,n1714,n1723);
xor (n1714,n1715,n1719);
xor (n1715,n1716,n170);
or (n1716,n1717,n1718);
and (n1717,n561,n164);
and (n1718,n633,n168);
xor (n1719,n1720,n100);
or (n1720,n1721,n1722);
and (n1721,n854,n174);
and (n1722,n858,n177);
xor (n1723,n1724,n75);
or (n1724,n1725,n1726);
and (n1725,n860,n98);
and (n1726,n994,n102);
xor (n1727,n1728,n1735);
xor (n1728,n1729,n1734);
xor (n1729,n14,n1730);
xor (n1730,n1731,n887);
or (n1731,n1732,n1733);
and (n1732,n63,n1010);
and (n1733,n65,n1014);
and (n1734,n1605,n1609);
xor (n1735,n1736,n23);
or (n1736,n1737,n1738);
and (n1737,n1198,n73);
and (n1738,n1202,n77);
nand (n1739,n1740,n1741,n1742);
nand (n1740,n1619,n1633);
nand (n1741,n1637,n1633);
nand (n1742,n1619,n1637);
nand (n1743,n1744,n1745,n1746);
nand (n1744,n1557,n1588);
nand (n1745,n1617,n1588);
nand (n1746,n1557,n1617);
nor (n1747,n1748,n1752);
nand (n1748,n1749,n1750,n1751);
nand (n1749,n1649,n1683);
nand (n1750,n1743,n1683);
nand (n1751,n1649,n1743);
xor (n1752,n1753,n1762);
xor (n1753,n1754,n1758);
nand (n1754,n1755,n1756,n1757);
nand (n1755,n1651,n1655);
nand (n1756,n1679,n1655);
nand (n1757,n1651,n1679);
nand (n1758,n1759,n1760,n1761);
nand (n1759,n1685,n1707);
nand (n1760,n1739,n1707);
nand (n1761,n1685,n1739);
xor (n1762,n1763,n1824);
xor (n1763,n1764,n1788);
xor (n1764,n1765,n1784);
xor (n1765,n1766,n1770);
nand (n1766,n1767,n1768,n1769);
nand (n1767,n1715,n1719);
nand (n1768,n1723,n1719);
nand (n1769,n1715,n1723);
xor (n1770,n1771,n1780);
xor (n1771,n1772,n1776);
xor (n1772,n1773,n166);
or (n1773,n1774,n1775);
and (n1774,n299,n441);
and (n1775,n428,n445);
xor (n1776,n1777,n170);
or (n1777,n1778,n1779);
and (n1778,n515,n164);
and (n1779,n561,n168);
xor (n1780,n1781,n100);
or (n1781,n1782,n1783);
and (n1782,n633,n174);
and (n1783,n854,n177);
nand (n1784,n1785,n1786,n1787);
nand (n1785,n1729,n1734);
nand (n1786,n1735,n1734);
nand (n1787,n1729,n1735);
xor (n1788,n1789,n1810);
xor (n1789,n1790,n1806);
xor (n1790,n1791,n1805);
xor (n1791,n1792,n1796);
xor (n1792,n1793,n75);
or (n1793,n1794,n1795);
and (n1794,n858,n98);
and (n1795,n860,n102);
xor (n1796,n1797,n1801);
xnor (n1797,n1798,n1012);
nor (n1798,n1799,n1800);
and (n1799,n30,n1213);
and (n1800,n7,n1215);
xor (n1801,n1802,n887);
or (n1802,n1803,n1804);
and (n1803,n44,n1010);
and (n1804,n63,n1014);
and (n1805,n14,n1730);
nand (n1806,n1807,n1808,n1809);
nand (n1807,n1657,n1661);
nand (n1808,n1665,n1661);
nand (n1809,n1657,n1665);
xor (n1810,n1811,n1820);
xor (n1811,n1812,n1816);
xor (n1812,n1813,n23);
or (n1813,n1814,n1815);
and (n1814,n994,n73);
and (n1815,n1198,n77);
xor (n1816,n1817,n14);
or (n1817,n1818,n1819);
and (n1818,n1227,n8);
and (n1819,n1241,n12);
xor (n1820,n1821,n10);
or (n1821,n1822,n1823);
and (n1822,n1202,n21);
and (n1823,n1204,n25);
xor (n1824,n1825,n1854);
xor (n1825,n1826,n1850);
xor (n1826,n1827,n1846);
xor (n1827,n1828,n1832);
nand (n1828,n1829,n1830,n1831);
nand (n1829,n1667,n1671);
nand (n1830,n1675,n1671);
nand (n1831,n1667,n1675);
xor (n1832,n1833,n1842);
xor (n1833,n1834,n1838);
xor (n1834,n1835,n525);
or (n1835,n1836,n1837);
and (n1836,n195,n662);
and (n1837,n197,n666);
xor (n1838,n1839,n664);
or (n1839,n1840,n1841);
and (n1840,n65,n885);
and (n1841,n112,n889);
xor (n1842,n1843,n443);
or (n1843,n1844,n1845);
and (n1844,n213,n523);
and (n1845,n267,n527);
nand (n1846,n1847,n1848,n1849);
nand (n1847,n1697,n1701);
nand (n1848,n1703,n1701);
nand (n1849,n1697,n1703);
nand (n1850,n1851,n1852,n1853);
nand (n1851,n1687,n1691);
nand (n1852,n1695,n1691);
nand (n1853,n1687,n1695);
nand (n1854,n1855,n1856,n1857);
nand (n1855,n1709,n1713);
nand (n1856,n1727,n1713);
nand (n1857,n1709,n1727);
nor (n1858,n1859,n2131);
nor (n1859,n1860,n2107);
nor (n1860,n1861,n2105);
nor (n1861,n1862,n2080);
nand (n1862,n1863,n2042);
nand (n1863,n1864,n1989,n2041);
nand (n1864,n1865,n1916);
xor (n1865,n1866,n1903);
xor (n1866,n1867,n1888);
nand (n1867,n1868,n1882,n1887);
nand (n1868,n1869,n1878);
and (n1869,n1870,n1874);
xnor (n1870,n1871,n1012);
nor (n1871,n1872,n1873);
and (n1872,n428,n1213);
and (n1873,n299,n1215);
xor (n1874,n1875,n887);
or (n1875,n1876,n1877);
and (n1876,n515,n1010);
and (n1877,n561,n1014);
xor (n1878,n1879,n166);
or (n1879,n1880,n1881);
and (n1880,n1198,n441);
and (n1881,n1202,n445);
nand (n1882,n1883,n1878);
xor (n1883,n1884,n170);
or (n1884,n1885,n1886);
and (n1885,n1204,n164);
and (n1886,n1227,n168);
nand (n1887,n1869,n1883);
xor (n1888,n1889,n1898);
xor (n1889,n1890,n1894);
xor (n1890,n1891,n525);
or (n1891,n1892,n1893);
and (n1892,n633,n662);
and (n1893,n854,n666);
xor (n1894,n1895,n664);
or (n1895,n1896,n1897);
and (n1896,n515,n885);
and (n1897,n561,n889);
and (n1898,n1899,n100);
xnor (n1899,n1900,n1012);
nor (n1900,n1901,n1902);
and (n1901,n299,n1213);
and (n1902,n267,n1215);
nand (n1903,n1904,n1910,n1915);
nand (n1904,n1905,n1909);
xor (n1905,n1906,n664);
or (n1906,n1907,n1908);
and (n1907,n561,n885);
and (n1908,n633,n889);
xor (n1909,n1899,n100);
nand (n1910,n1911,n1909);
xor (n1911,n1912,n443);
or (n1912,n1913,n1914);
and (n1913,n860,n523);
and (n1914,n994,n527);
nand (n1915,n1905,n1911);
xor (n1916,n1917,n1953);
xor (n1917,n1918,n1929);
xor (n1918,n1919,n1925);
xor (n1919,n1920,n1924);
xor (n1920,n1921,n443);
or (n1921,n1922,n1923);
and (n1922,n858,n523);
and (n1923,n860,n527);
xor (n1924,n1328,n1332);
xor (n1925,n1926,n166);
or (n1926,n1927,n1928);
and (n1927,n994,n441);
and (n1928,n1198,n445);
xor (n1929,n1930,n1939);
xor (n1930,n1931,n1935);
xor (n1931,n1932,n170);
or (n1932,n1933,n1934);
and (n1933,n1202,n164);
and (n1934,n1204,n168);
xor (n1935,n1936,n100);
or (n1936,n1937,n1938);
and (n1937,n1227,n174);
and (n1938,n1241,n177);
nand (n1939,n1940,n1947,n1952);
nand (n1940,n1941,n1945);
xor (n1941,n1942,n887);
or (n1942,n1943,n1944);
and (n1943,n428,n1010);
and (n1944,n515,n1014);
xnor (n1945,n1946,n100);
nand (n1946,n1241,n174);
nand (n1947,n1948,n1945);
xor (n1948,n1949,n525);
or (n1949,n1950,n1951);
and (n1950,n854,n662);
and (n1951,n858,n666);
nand (n1952,n1941,n1948);
nand (n1953,n1954,n1974,n1988);
nand (n1954,n1955,n1957);
xor (n1955,n1956,n1948);
xor (n1956,n1941,n1945);
nand (n1957,n1958,n1967,n1973);
nand (n1958,n1959,n1963);
xor (n1959,n1960,n525);
or (n1960,n1961,n1962);
and (n1961,n858,n662);
and (n1962,n860,n666);
xor (n1963,n1964,n664);
or (n1964,n1965,n1966);
and (n1965,n633,n885);
and (n1966,n854,n889);
nand (n1967,n1968,n1963);
and (n1968,n1969,n170);
xnor (n1969,n1970,n1012);
nor (n1970,n1971,n1972);
and (n1971,n515,n1213);
and (n1972,n428,n1215);
nand (n1973,n1959,n1968);
nand (n1974,n1975,n1957);
nand (n1975,n1976,n1982,n1987);
nand (n1976,n1977,n1981);
xor (n1977,n1978,n443);
or (n1978,n1979,n1980);
and (n1979,n994,n523);
and (n1980,n1198,n527);
xor (n1981,n1870,n1874);
nand (n1982,n1983,n1981);
xor (n1983,n1984,n166);
or (n1984,n1985,n1986);
and (n1985,n1202,n441);
and (n1986,n1204,n445);
nand (n1987,n1977,n1983);
nand (n1988,n1955,n1975);
nand (n1989,n1990,n1916);
nand (n1990,n1991,n1996,n2040);
nand (n1991,n1992,n1994);
xor (n1992,n1993,n1883);
xor (n1993,n1869,n1878);
xor (n1994,n1995,n1911);
xor (n1995,n1905,n1909);
nand (n1996,n1997,n1994);
nand (n1997,n1998,n2017,n2039);
nand (n1998,n1999,n2003);
xor (n1999,n2000,n170);
or (n2000,n2001,n2002);
and (n2001,n1227,n164);
and (n2002,n1241,n168);
nand (n2003,n2004,n2011,n2016);
nand (n2004,n2005,n2009);
xor (n2005,n2006,n887);
or (n2006,n2007,n2008);
and (n2007,n561,n1010);
and (n2008,n633,n1014);
xnor (n2009,n2010,n170);
nand (n2010,n1241,n164);
nand (n2011,n2012,n2009);
xor (n2012,n2013,n525);
or (n2013,n2014,n2015);
and (n2014,n860,n662);
and (n2015,n994,n666);
nand (n2016,n2005,n2012);
nand (n2017,n2018,n2003);
nand (n2018,n2019,n2033,n2038);
nand (n2019,n2020,n2024);
xor (n2020,n2021,n664);
or (n2021,n2022,n2023);
and (n2022,n854,n885);
and (n2023,n858,n889);
and (n2024,n2025,n2029);
xnor (n2025,n2026,n1012);
nor (n2026,n2027,n2028);
and (n2027,n561,n1213);
and (n2028,n515,n1215);
xor (n2029,n2030,n887);
or (n2030,n2031,n2032);
and (n2031,n633,n1010);
and (n2032,n854,n1014);
nand (n2033,n2034,n2024);
xor (n2034,n2035,n443);
or (n2035,n2036,n2037);
and (n2036,n1198,n523);
and (n2037,n1202,n527);
nand (n2038,n2020,n2034);
nand (n2039,n1999,n2018);
nand (n2040,n1992,n1997);
nand (n2041,n1865,n1990);
xor (n2042,n2043,n2058);
xor (n2043,n2044,n2054);
xor (n2044,n2045,n2052);
xor (n2045,n2046,n2050);
nand (n2046,n2047,n2048,n2049);
nand (n2047,n1890,n1894);
nand (n2048,n1898,n1894);
nand (n2049,n1890,n1898);
xor (n2050,n2051,n1341);
xor (n2051,n1327,n1336);
xor (n2052,n2053,n1442);
xor (n2053,n1436,n1440);
nand (n2054,n2055,n2056,n2057);
nand (n2055,n1918,n1929);
nand (n2056,n1953,n1929);
nand (n2057,n1918,n1953);
xor (n2058,n2059,n2068);
xor (n2059,n2060,n2064);
nand (n2060,n2061,n2062,n2063);
nand (n2061,n1931,n1935);
nand (n2062,n1939,n1935);
nand (n2063,n1931,n1939);
nand (n2064,n2065,n2066,n2067);
nand (n2065,n1867,n1888);
nand (n2066,n1903,n1888);
nand (n2067,n1867,n1903);
xor (n2068,n2069,n2078);
xor (n2069,n2070,n2074);
xor (n2070,n2071,n100);
or (n2071,n2072,n2073);
and (n2072,n1204,n174);
and (n2073,n1227,n177);
nand (n2074,n2075,n2076,n2077);
nand (n2075,n1920,n1924);
nand (n2076,n1925,n1924);
nand (n2077,n1920,n1925);
xor (n2078,n2079,n1428);
xor (n2079,n1419,n1423);
nor (n2080,n2081,n2085);
nand (n2081,n2082,n2083,n2084);
nand (n2082,n2044,n2054);
nand (n2083,n2058,n2054);
nand (n2084,n2044,n2058);
xor (n2085,n2086,n2093);
xor (n2086,n2087,n2089);
xor (n2087,n2088,n1349);
xor (n2088,n1325,n1346);
nand (n2089,n2090,n2091,n2092);
nand (n2090,n2060,n2064);
nand (n2091,n2068,n2064);
nand (n2092,n2060,n2068);
xor (n2093,n2094,n2103);
xor (n2094,n2095,n2099);
nand (n2095,n2096,n2097,n2098);
nand (n2096,n2070,n2074);
nand (n2097,n2078,n2074);
nand (n2098,n2070,n2078);
nand (n2099,n2100,n2101,n2102);
nand (n2100,n2046,n2050);
nand (n2101,n2052,n2050);
nand (n2102,n2046,n2052);
xor (n2103,n2104,n1434);
xor (n2104,n1417,n1431);
not (n2105,n2106);
nand (n2106,n2081,n2085);
not (n2107,n2108);
nor (n2108,n2109,n2124);
nor (n2109,n2110,n2114);
nand (n2110,n2111,n2112,n2113);
nand (n2111,n2087,n2089);
nand (n2112,n2093,n2089);
nand (n2113,n2087,n2093);
xor (n2114,n2115,n2122);
xor (n2115,n2116,n2118);
xor (n2116,n2117,n1415);
xor (n2117,n1408,n1412);
nand (n2118,n2119,n2120,n2121);
nand (n2119,n2095,n2099);
nand (n2120,n2103,n2099);
nand (n2121,n2095,n2103);
xor (n2122,n2123,n1323);
xor (n2123,n1269,n1271);
nor (n2124,n2125,n2129);
nand (n2125,n2126,n2127,n2128);
nand (n2126,n2116,n2118);
nand (n2127,n2122,n2118);
nand (n2128,n2116,n2122);
xor (n2129,n2130,n1366);
xor (n2130,n1190,n1267);
not (n2131,n2132);
nor (n2132,n2133,n2135);
nor (n2133,n2134,n2124);
nand (n2134,n2110,n2114);
not (n2135,n2136);
nand (n2136,n2125,n2129);
not (n2137,n2138);
nor (n2138,n2139,n2146);
nor (n2139,n2140,n2145);
nor (n2140,n2141,n2143);
nor (n2141,n2142,n1540);
nand (n2142,n1188,n1450);
not (n2143,n2144);
nand (n2144,n1541,n1545);
not (n2145,n1641);
not (n2146,n2147);
nor (n2147,n2148,n2150);
nor (n2148,n2149,n1747);
nand (n2149,n1643,n1647);
not (n2150,n2151);
nand (n2151,n1748,n1752);
not (n2152,n2153);
nor (n2153,n2154,n2569);
nand (n2154,n2155,n2382);
nor (n2155,n2156,n2268);
nor (n2156,n2157,n2161);
nand (n2157,n2158,n2159,n2160);
nand (n2158,n1754,n1758);
nand (n2159,n1762,n1758);
nand (n2160,n1754,n1762);
xor (n2161,n2162,n2264);
xor (n2162,n2163,n2196);
xor (n2163,n2164,n2192);
xor (n2164,n2165,n2188);
xor (n2165,n2166,n2184);
xor (n2166,n2167,n2180);
xor (n2167,n2168,n2177);
xor (n2168,n2169,n2173);
xor (n2169,n2170,n887);
or (n2170,n2171,n2172);
and (n2171,n30,n1010);
and (n2172,n44,n1014);
xor (n2173,n2174,n664);
or (n2174,n2175,n2176);
and (n2175,n63,n885);
and (n2176,n65,n889);
xnor (n2177,n2178,n1012);
nor (n2178,n2179,n1800);
and (n2179,n7,n1213);
nand (n2180,n2181,n2182,n2183);
nand (n2181,n1772,n1776);
nand (n2182,n1780,n1776);
nand (n2183,n1772,n1780);
nand (n2184,n2185,n2186,n2187);
nand (n2185,n1792,n1796);
nand (n2186,n1805,n1796);
nand (n2187,n1792,n1805);
nand (n2188,n2189,n2190,n2191);
nand (n2189,n1766,n1770);
nand (n2190,n1784,n1770);
nand (n2191,n1766,n1784);
nand (n2192,n2193,n2194,n2195);
nand (n2193,n1790,n1806);
nand (n2194,n1810,n1806);
nand (n2195,n1790,n1810);
xor (n2196,n2197,n2260);
xor (n2197,n2198,n2236);
xor (n2198,n2199,n2221);
xor (n2199,n2200,n2214);
xor (n2200,n2201,n2210);
xor (n2201,n2202,n2206);
xor (n2202,n2203,n443);
or (n2203,n2204,n2205);
and (n2204,n197,n523);
and (n2205,n213,n527);
xor (n2206,n2207,n166);
or (n2207,n2208,n2209);
and (n2208,n267,n441);
and (n2209,n299,n445);
xor (n2210,n2211,n170);
or (n2211,n2212,n2213);
and (n2212,n428,n164);
and (n2213,n515,n168);
xor (n2214,n2215,n2217);
xor (n2215,n14,n2216);
and (n2216,n1797,n1801);
xor (n2217,n2218,n23);
or (n2218,n2219,n2220);
and (n2219,n860,n73);
and (n2220,n994,n77);
xor (n2221,n2222,n2231);
xor (n2222,n2223,n2227);
xor (n2223,n2224,n100);
or (n2224,n2225,n2226);
and (n2225,n561,n174);
and (n2226,n633,n177);
xor (n2227,n2228,n75);
or (n2228,n2229,n2230);
and (n2229,n854,n98);
and (n2230,n858,n102);
xor (n2231,n14,n2232);
xor (n2232,n2233,n525);
or (n2233,n2234,n2235);
and (n2234,n112,n662);
and (n2235,n195,n666);
xor (n2236,n2237,n2246);
xor (n2237,n2238,n2242);
nand (n2238,n2239,n2240,n2241);
nand (n2239,n1812,n1816);
nand (n2240,n1820,n1816);
nand (n2241,n1812,n1820);
nand (n2242,n2243,n2244,n2245);
nand (n2243,n1828,n1832);
nand (n2244,n1846,n1832);
nand (n2245,n1828,n1846);
xor (n2246,n2247,n2256);
xor (n2247,n2248,n2252);
xor (n2248,n2249,n10);
or (n2249,n2250,n2251);
and (n2250,n1198,n21);
and (n2251,n1202,n25);
xor (n2252,n2253,n14);
or (n2253,n2254,n2255);
and (n2254,n1204,n8);
and (n2255,n1227,n12);
nand (n2256,n2257,n2258,n2259);
nand (n2257,n1834,n1838);
nand (n2258,n1842,n1838);
nand (n2259,n1834,n1842);
nand (n2260,n2261,n2262,n2263);
nand (n2261,n1826,n1850);
nand (n2262,n1854,n1850);
nand (n2263,n1826,n1854);
nand (n2264,n2265,n2266,n2267);
nand (n2265,n1764,n1788);
nand (n2266,n1824,n1788);
nand (n2267,n1764,n1824);
nor (n2268,n2269,n2273);
nand (n2269,n2270,n2271,n2272);
nand (n2270,n2163,n2196);
nand (n2271,n2264,n2196);
nand (n2272,n2163,n2264);
xor (n2273,n2274,n2283);
xor (n2274,n2275,n2279);
nand (n2275,n2276,n2277,n2278);
nand (n2276,n2165,n2188);
nand (n2277,n2192,n2188);
nand (n2278,n2165,n2192);
nand (n2279,n2280,n2281,n2282);
nand (n2280,n2198,n2236);
nand (n2281,n2260,n2236);
nand (n2282,n2198,n2260);
xor (n2283,n2284,n2341);
xor (n2284,n2285,n2316);
xor (n2285,n2286,n2302);
xor (n2286,n2287,n2291);
nand (n2287,n2288,n2289,n2290);
nand (n2288,n14,n2216);
nand (n2289,n2217,n2216);
nand (n2290,n14,n2217);
xor (n2291,n2292,n2298);
xor (n2292,n2293,n2297);
xor (n2293,n2294,n75);
or (n2294,n2295,n2296);
and (n2295,n633,n98);
and (n2296,n854,n102);
and (n2297,n14,n2232);
xor (n2298,n2299,n23);
or (n2299,n2300,n2301);
and (n2300,n858,n73);
and (n2301,n860,n77);
xor (n2302,n2303,n2312);
xor (n2303,n2304,n2308);
xor (n2304,n2305,n10);
or (n2305,n2306,n2307);
and (n2306,n994,n21);
and (n2307,n1198,n25);
xor (n2308,n2309,n14);
or (n2309,n2310,n2311);
and (n2310,n1202,n8);
and (n2311,n1204,n12);
nand (n2312,n2313,n2314,n2315);
nand (n2313,n2169,n2173);
nand (n2314,n2177,n2173);
nand (n2315,n2169,n2177);
xor (n2316,n2317,n2326);
xor (n2317,n2318,n2322);
nand (n2318,n2319,n2320,n2321);
nand (n2319,n2248,n2252);
nand (n2320,n2256,n2252);
nand (n2321,n2248,n2256);
nand (n2322,n2323,n2324,n2325);
nand (n2323,n2167,n2180);
nand (n2324,n2184,n2180);
nand (n2325,n2167,n2184);
xor (n2326,n2327,n14);
xor (n2327,n2328,n2332);
nand (n2328,n2329,n2330,n2331);
nand (n2329,n2202,n2206);
nand (n2330,n2210,n2206);
nand (n2331,n2202,n2210);
xor (n2332,n2333,n2338);
not (n2333,n2334);
xor (n2334,n2335,n525);
or (n2335,n2336,n2337);
and (n2336,n65,n662);
and (n2337,n112,n666);
xor (n2338,n2339,n887);
or (n2339,n1009,n2340);
and (n2340,n30,n1014);
xor (n2341,n2342,n2378);
xor (n2342,n2343,n2347);
nand (n2343,n2344,n2345,n2346);
nand (n2344,n2200,n2214);
nand (n2345,n2221,n2214);
nand (n2346,n2200,n2221);
xor (n2347,n2348,n2367);
xor (n2348,n2349,n2353);
nand (n2349,n2350,n2351,n2352);
nand (n2350,n2223,n2227);
nand (n2351,n2231,n2227);
nand (n2352,n2223,n2231);
xor (n2353,n2354,n2363);
xor (n2354,n2355,n2359);
xor (n2355,n2356,n166);
or (n2356,n2357,n2358);
and (n2357,n213,n441);
and (n2358,n267,n445);
xor (n2359,n2360,n170);
or (n2360,n2361,n2362);
and (n2361,n299,n164);
and (n2362,n428,n168);
xor (n2363,n2364,n100);
or (n2364,n2365,n2366);
and (n2365,n515,n174);
and (n2366,n561,n177);
xor (n2367,n2368,n2374);
xor (n2368,n2369,n2373);
xor (n2369,n2370,n664);
or (n2370,n2371,n2372);
and (n2371,n44,n885);
and (n2372,n63,n889);
not (n2373,n2177);
xor (n2374,n2375,n443);
or (n2375,n2376,n2377);
and (n2376,n195,n523);
and (n2377,n197,n527);
nand (n2378,n2379,n2380,n2381);
nand (n2379,n2238,n2242);
nand (n2380,n2246,n2242);
nand (n2381,n2238,n2246);
nor (n2382,n2383,n2490);
nor (n2383,n2384,n2388);
nand (n2384,n2385,n2386,n2387);
nand (n2385,n2275,n2279);
nand (n2386,n2283,n2279);
nand (n2387,n2275,n2283);
xor (n2388,n2389,n2486);
xor (n2389,n2390,n2430);
xor (n2390,n2391,n2426);
xor (n2391,n2392,n2422);
xor (n2392,n2393,n2418);
xor (n2393,n2394,n2408);
xor (n2394,n2395,n2404);
xor (n2395,n2396,n2400);
xor (n2396,n2397,n166);
or (n2397,n2398,n2399);
and (n2398,n197,n441);
and (n2399,n213,n445);
xor (n2400,n2401,n170);
or (n2401,n2402,n2403);
and (n2402,n267,n164);
and (n2403,n299,n168);
xor (n2404,n2405,n75);
or (n2405,n2406,n2407);
and (n2406,n561,n98);
and (n2407,n633,n102);
xor (n2408,n2409,n2414);
xor (n2409,n2410,n1007);
xor (n2410,n2411,n525);
or (n2411,n2412,n2413);
and (n2412,n63,n662);
and (n2413,n65,n666);
xor (n2414,n2415,n443);
or (n2415,n2416,n2417);
and (n2416,n112,n523);
and (n2417,n195,n527);
nand (n2418,n2419,n2420,n2421);
nand (n2419,n2293,n2297);
nand (n2420,n2298,n2297);
nand (n2421,n2293,n2298);
nand (n2422,n2423,n2424,n2425);
nand (n2423,n2287,n2291);
nand (n2424,n2302,n2291);
nand (n2425,n2287,n2302);
nand (n2426,n2427,n2428,n2429);
nand (n2427,n2318,n2322);
nand (n2428,n2326,n2322);
nand (n2429,n2318,n2326);
xor (n2430,n2431,n2482);
xor (n2431,n2432,n2453);
xor (n2432,n2433,n2449);
xor (n2433,n2434,n2445);
xor (n2434,n2435,n2441);
xor (n2435,n2436,n2437);
not (n2436,n1048);
xor (n2437,n2438,n100);
or (n2438,n2439,n2440);
and (n2439,n428,n174);
and (n2440,n515,n177);
xor (n2441,n2442,n23);
or (n2442,n2443,n2444);
and (n2443,n854,n73);
and (n2444,n858,n77);
nand (n2445,n2446,n2447,n2448);
nand (n2446,n2304,n2308);
nand (n2447,n2312,n2308);
nand (n2448,n2304,n2312);
nand (n2449,n2450,n2451,n2452);
nand (n2450,n2328,n2332);
nand (n2451,n14,n2332);
nand (n2452,n2328,n14);
xor (n2453,n2454,n2478);
xor (n2454,n2455,n2468);
xor (n2455,n2456,n2465);
xor (n2456,n2457,n2461);
xor (n2457,n2458,n10);
or (n2458,n2459,n2460);
and (n2459,n860,n21);
and (n2460,n994,n25);
xor (n2461,n2462,n14);
or (n2462,n2463,n2464);
and (n2463,n1198,n8);
and (n2464,n1202,n12);
nand (n2465,n2333,n2466,n2467);
nand (n2466,n2338,n2334);
not (n2467,n2338);
xor (n2468,n2469,n2474);
xor (n2469,n14,n2470);
nand (n2470,n2471,n2472,n2473);
nand (n2471,n2369,n2373);
nand (n2472,n2374,n2373);
nand (n2473,n2369,n2374);
nand (n2474,n2475,n2476,n2477);
nand (n2475,n2355,n2359);
nand (n2476,n2363,n2359);
nand (n2477,n2355,n2363);
nand (n2478,n2479,n2480,n2481);
nand (n2479,n2349,n2353);
nand (n2480,n2367,n2353);
nand (n2481,n2349,n2367);
nand (n2482,n2483,n2484,n2485);
nand (n2483,n2343,n2347);
nand (n2484,n2378,n2347);
nand (n2485,n2343,n2378);
nand (n2486,n2487,n2488,n2489);
nand (n2487,n2285,n2316);
nand (n2488,n2341,n2316);
nand (n2489,n2285,n2341);
nor (n2490,n2491,n2495);
nand (n2491,n2492,n2493,n2494);
nand (n2492,n2390,n2430);
nand (n2493,n2486,n2430);
nand (n2494,n2390,n2486);
xor (n2495,n2496,n2505);
xor (n2496,n2497,n2501);
nand (n2497,n2498,n2499,n2500);
nand (n2498,n2392,n2422);
nand (n2499,n2426,n2422);
nand (n2500,n2392,n2426);
nand (n2501,n2502,n2503,n2504);
nand (n2502,n2432,n2453);
nand (n2503,n2482,n2453);
nand (n2504,n2432,n2482);
xor (n2505,n2506,n2537);
xor (n2506,n2507,n2511);
nand (n2507,n2508,n2509,n2510);
nand (n2508,n2455,n2468);
nand (n2509,n2478,n2468);
nand (n2510,n2455,n2478);
xor (n2511,n2512,n2525);
xor (n2512,n2513,n2517);
nand (n2513,n2514,n2515,n2516);
nand (n2514,n14,n2470);
nand (n2515,n2474,n2470);
nand (n2516,n14,n2474);
xor (n2517,n2518,n2521);
xor (n2518,n2519,n14);
xor (n2519,n2520,n1006);
xor (n2520,n998,n1001);
nand (n2521,n2522,n2523,n2524);
nand (n2522,n2410,n1007);
nand (n2523,n2414,n1007);
nand (n2524,n2410,n2414);
xor (n2525,n2526,n2533);
xor (n2526,n2527,n2529);
xor (n2527,n2528,n1034);
xor (n2528,n1025,n1029);
nand (n2529,n2530,n2531,n2532);
nand (n2530,n2396,n2400);
nand (n2531,n2404,n2400);
nand (n2532,n2396,n2404);
nand (n2533,n2534,n2535,n2536);
nand (n2534,n2457,n2461);
nand (n2535,n2465,n2461);
nand (n2536,n2457,n2465);
xor (n2537,n2538,n2547);
xor (n2538,n2539,n2543);
nand (n2539,n2540,n2541,n2542);
nand (n2540,n2394,n2408);
nand (n2541,n2418,n2408);
nand (n2542,n2394,n2418);
nand (n2543,n2544,n2545,n2546);
nand (n2544,n2434,n2445);
nand (n2545,n2449,n2445);
nand (n2546,n2434,n2449);
xor (n2547,n2548,n2555);
xor (n2548,n2549,n2553);
nand (n2549,n2550,n2551,n2552);
nand (n2550,n2436,n2437);
nand (n2551,n2441,n2437);
nand (n2552,n2436,n2441);
xor (n2553,n2554,n1053);
xor (n2554,n1044,n1048);
xor (n2555,n2556,n2565);
xor (n2556,n2557,n2561);
xor (n2557,n2558,n23);
or (n2558,n2559,n2560);
and (n2559,n633,n73);
and (n2560,n854,n77);
xor (n2561,n2562,n10);
or (n2562,n2563,n2564);
and (n2563,n858,n21);
and (n2564,n860,n25);
xor (n2565,n2566,n14);
or (n2566,n2567,n2568);
and (n2567,n994,n8);
and (n2568,n1198,n12);
nand (n2569,n2570,n2654);
nor (n2570,n2571,n2621);
nor (n2571,n2572,n2576);
nand (n2572,n2573,n2574,n2575);
nand (n2573,n2497,n2501);
nand (n2574,n2505,n2501);
nand (n2575,n2497,n2505);
xor (n2576,n2577,n2617);
xor (n2577,n2578,n2598);
xor (n2578,n2579,n2586);
xor (n2579,n2580,n2582);
xor (n2580,n2581,n1042);
xor (n2581,n1023,n1039);
nand (n2582,n2583,n2584,n2585);
nand (n2583,n2549,n2553);
nand (n2584,n2555,n2553);
nand (n2585,n2549,n2555);
xor (n2586,n2587,n2594);
xor (n2587,n2588,n2592);
nand (n2588,n2589,n2590,n2591);
nand (n2589,n2557,n2561);
nand (n2590,n2565,n2561);
nand (n2591,n2557,n2565);
xor (n2592,n2593,n952);
xor (n2593,n946,n950);
nand (n2594,n2595,n2596,n2597);
nand (n2595,n2519,n14);
nand (n2596,n2521,n14);
nand (n2597,n2519,n2521);
xor (n2598,n2599,n2613);
xor (n2599,n2600,n2604);
nand (n2600,n2601,n2602,n2603);
nand (n2601,n2513,n2517);
nand (n2602,n2525,n2517);
nand (n2603,n2513,n2525);
xor (n2604,n2605,n2609);
xor (n2605,n2606,n2608);
xor (n2606,n2607,n968);
xor (n2607,n959,n963);
xor (n2608,n991,n996);
nand (n2609,n2610,n2611,n2612);
nand (n2610,n2527,n2529);
nand (n2611,n2533,n2529);
nand (n2612,n2527,n2533);
nand (n2613,n2614,n2615,n2616);
nand (n2614,n2539,n2543);
nand (n2615,n2547,n2543);
nand (n2616,n2539,n2547);
nand (n2617,n2618,n2619,n2620);
nand (n2618,n2507,n2511);
nand (n2619,n2537,n2511);
nand (n2620,n2507,n2537);
nor (n2621,n2622,n2626);
nand (n2622,n2623,n2624,n2625);
nand (n2623,n2578,n2598);
nand (n2624,n2617,n2598);
nand (n2625,n2578,n2617);
xor (n2626,n2627,n2650);
xor (n2627,n2628,n2638);
xor (n2628,n2629,n2636);
xor (n2629,n2630,n2632);
xor (n2630,n2631,n939);
xor (n2631,n924,n936);
nand (n2632,n2633,n2634,n2635);
nand (n2633,n2588,n2592);
nand (n2634,n2594,n2592);
nand (n2635,n2588,n2594);
xor (n2636,n2637,n974);
xor (n2637,n944,n957);
xor (n2638,n2639,n2646);
xor (n2639,n2640,n2642);
xor (n2640,n2641,n1021);
xor (n2641,n988,n1018);
nand (n2642,n2643,n2644,n2645);
nand (n2643,n2606,n2608);
nand (n2644,n2609,n2608);
nand (n2645,n2606,n2609);
nand (n2646,n2647,n2648,n2649);
nand (n2647,n2580,n2582);
nand (n2648,n2586,n2582);
nand (n2649,n2580,n2586);
nand (n2650,n2651,n2652,n2653);
nand (n2651,n2600,n2604);
nand (n2652,n2613,n2604);
nand (n2653,n2600,n2613);
nor (n2654,n2655,n2672);
nor (n2655,n2656,n2660);
nand (n2656,n2657,n2658,n2659);
nand (n2657,n2628,n2638);
nand (n2658,n2650,n2638);
nand (n2659,n2628,n2650);
xor (n2660,n2661,n2668);
xor (n2661,n2662,n2666);
nand (n2662,n2663,n2664,n2665);
nand (n2663,n2630,n2632);
nand (n2664,n2636,n2632);
nand (n2665,n2630,n2636);
xor (n2666,n2667,n1061);
xor (n2667,n984,n986);
nand (n2668,n2669,n2670,n2671);
nand (n2669,n2640,n2642);
nand (n2670,n2646,n2642);
nand (n2671,n2640,n2646);
nor (n2672,n2673,n2677);
nand (n2673,n2674,n2675,n2676);
nand (n2674,n2662,n2666);
nand (n2675,n2668,n2666);
nand (n2676,n2662,n2668);
xor (n2677,n2678,n982);
xor (n2678,n760,n844);
not (n2679,n2680);
nor (n2680,n2681,n2696);
nor (n2681,n2569,n2682);
nor (n2682,n2683,n2690);
nor (n2683,n2684,n2689);
nor (n2684,n2685,n2687);
nor (n2685,n2686,n2268);
nand (n2686,n2157,n2161);
not (n2687,n2688);
nand (n2688,n2269,n2273);
not (n2689,n2382);
not (n2690,n2691);
nor (n2691,n2692,n2694);
nor (n2692,n2693,n2490);
nand (n2693,n2384,n2388);
not (n2694,n2695);
nand (n2695,n2491,n2495);
not (n2696,n2697);
nor (n2697,n2698,n2705);
nor (n2698,n2699,n2704);
nor (n2699,n2700,n2702);
nor (n2700,n2701,n2621);
nand (n2701,n2572,n2576);
not (n2702,n2703);
nand (n2703,n2622,n2626);
not (n2704,n2654);
not (n2705,n2706);
nor (n2706,n2707,n2709);
nor (n2707,n2708,n2672);
nand (n2708,n2656,n2660);
not (n2709,n2710);
nand (n2710,n2673,n2677);
nand (n2711,n2712,n3131);
nand (n2712,n2713,n3024);
nor (n2713,n2714,n3009);
nor (n2714,n2715,n2880);
nand (n2715,n2716,n2857);
nor (n2716,n2717,n2834);
nor (n2717,n2718,n2807);
nand (n2718,n2719,n2764,n2806);
nand (n2719,n2720,n2732);
xor (n2720,n2721,n2727);
xor (n2721,n2722,n2723);
xor (n2722,n2025,n2029);
xor (n2723,n2724,n166);
or (n2724,n2725,n2726);
and (n2725,n1227,n441);
and (n2726,n1241,n445);
and (n2727,n166,n2728);
xor (n2728,n2729,n887);
or (n2729,n2730,n2731);
and (n2730,n854,n1010);
and (n2731,n858,n1014);
nand (n2732,n2733,n2750,n2763);
nand (n2733,n2734,n2735);
xor (n2734,n166,n2728);
nand (n2735,n2736,n2745,n2749);
nand (n2736,n2737,n2741);
xor (n2737,n2738,n525);
or (n2738,n2739,n2740);
and (n2739,n1202,n662);
and (n2740,n1204,n666);
xor (n2741,n2742,n664);
or (n2742,n2743,n2744);
and (n2743,n994,n885);
and (n2744,n1198,n889);
nand (n2745,n2746,n2741);
and (n2746,n443,n2747);
xnor (n2747,n2748,n443);
nand (n2748,n1241,n523);
nand (n2749,n2737,n2746);
nand (n2750,n2751,n2735);
xor (n2751,n2752,n2759);
xor (n2752,n2753,n2757);
xnor (n2753,n2754,n1012);
nor (n2754,n2755,n2756);
and (n2755,n633,n1213);
and (n2756,n561,n1215);
xnor (n2757,n2758,n166);
nand (n2758,n1241,n441);
xor (n2759,n2760,n525);
or (n2760,n2761,n2762);
and (n2761,n1198,n662);
and (n2762,n1202,n666);
nand (n2763,n2734,n2751);
nand (n2764,n2765,n2732);
xor (n2765,n2766,n2785);
xor (n2766,n2767,n2771);
nand (n2767,n2768,n2769,n2770);
nand (n2768,n2753,n2757);
nand (n2769,n2759,n2757);
nand (n2770,n2753,n2759);
xor (n2771,n2772,n2781);
xor (n2772,n2773,n2777);
xor (n2773,n2774,n525);
or (n2774,n2775,n2776);
and (n2775,n994,n662);
and (n2776,n1198,n666);
xor (n2777,n2778,n664);
or (n2778,n2779,n2780);
and (n2779,n858,n885);
and (n2780,n860,n889);
xor (n2781,n2782,n443);
or (n2782,n2783,n2784);
and (n2783,n1202,n523);
and (n2784,n1204,n527);
nand (n2785,n2786,n2800,n2805);
nand (n2786,n2787,n2791);
xor (n2787,n2788,n664);
or (n2788,n2789,n2790);
and (n2789,n860,n885);
and (n2790,n994,n889);
and (n2791,n2792,n2796);
xnor (n2792,n2793,n1012);
nor (n2793,n2794,n2795);
and (n2794,n854,n1213);
and (n2795,n633,n1215);
xor (n2796,n2797,n887);
or (n2797,n2798,n2799);
and (n2798,n858,n1010);
and (n2799,n860,n1014);
nand (n2800,n2801,n2791);
xor (n2801,n2802,n443);
or (n2802,n2803,n2804);
and (n2803,n1204,n523);
and (n2804,n1227,n527);
nand (n2805,n2787,n2801);
nand (n2806,n2720,n2765);
xor (n2807,n2808,n2822);
xor (n2808,n2809,n2818);
xor (n2809,n2810,n2816);
xor (n2810,n2811,n2815);
xor (n2811,n2812,n166);
or (n2812,n2813,n2814);
and (n2813,n1204,n441);
and (n2814,n1227,n445);
xor (n2815,n1969,n170);
xor (n2816,n2817,n2012);
xor (n2817,n2005,n2009);
nand (n2818,n2819,n2820,n2821);
nand (n2819,n2767,n2771);
nand (n2820,n2785,n2771);
nand (n2821,n2767,n2785);
xor (n2822,n2823,n2832);
xor (n2823,n2824,n2828);
nand (n2824,n2825,n2826,n2827);
nand (n2825,n2722,n2723);
nand (n2826,n2727,n2723);
nand (n2827,n2722,n2727);
nand (n2828,n2829,n2830,n2831);
nand (n2829,n2773,n2777);
nand (n2830,n2781,n2777);
nand (n2831,n2773,n2781);
xor (n2832,n2833,n2034);
xor (n2833,n2020,n2024);
nor (n2834,n2835,n2839);
nand (n2835,n2836,n2837,n2838);
nand (n2836,n2809,n2818);
nand (n2837,n2822,n2818);
nand (n2838,n2809,n2822);
xor (n2839,n2840,n2847);
xor (n2840,n2841,n2843);
xor (n2841,n2842,n2018);
xor (n2842,n1999,n2003);
nand (n2843,n2844,n2845,n2846);
nand (n2844,n2824,n2828);
nand (n2845,n2832,n2828);
nand (n2846,n2824,n2832);
xor (n2847,n2848,n2853);
xor (n2848,n2849,n2851);
xor (n2849,n2850,n1968);
xor (n2850,n1959,n1963);
xor (n2851,n2852,n1983);
xor (n2852,n1977,n1981);
nand (n2853,n2854,n2855,n2856);
nand (n2854,n2811,n2815);
nand (n2855,n2816,n2815);
nand (n2856,n2811,n2816);
nor (n2857,n2858,n2873);
nor (n2858,n2859,n2863);
nand (n2859,n2860,n2861,n2862);
nand (n2860,n2841,n2843);
nand (n2861,n2847,n2843);
nand (n2862,n2841,n2847);
xor (n2863,n2864,n2871);
xor (n2864,n2865,n2867);
xor (n2865,n2866,n1975);
xor (n2866,n1955,n1957);
nand (n2867,n2868,n2869,n2870);
nand (n2868,n2849,n2851);
nand (n2869,n2853,n2851);
nand (n2870,n2849,n2853);
xor (n2871,n2872,n1997);
xor (n2872,n1992,n1994);
nor (n2873,n2874,n2878);
nand (n2874,n2875,n2876,n2877);
nand (n2875,n2865,n2867);
nand (n2876,n2871,n2867);
nand (n2877,n2865,n2871);
xor (n2878,n2879,n1990);
xor (n2879,n1865,n1916);
nor (n2880,n2881,n3003);
nor (n2881,n2882,n2979);
nor (n2882,n2883,n2976);
nor (n2883,n2884,n2952);
nand (n2884,n2885,n2924);
or (n2885,n2886,n2910,n2923);
and (n2886,n2887,n2896);
xor (n2887,n2888,n2892);
xnor (n2888,n2889,n1012);
nor (n2889,n2890,n2891);
and (n2890,n860,n1213);
and (n2891,n858,n1215);
xnor (n2892,n2893,n887);
nor (n2893,n2894,n2895);
and (n2894,n1198,n1014);
and (n2895,n994,n1010);
or (n2896,n2897,n2904,n2909);
and (n2897,n2898,n2900);
not (n2898,n2899);
nand (n2899,n1241,n662);
xnor (n2900,n2901,n1012);
nor (n2901,n2902,n2903);
and (n2902,n994,n1213);
and (n2903,n860,n1215);
and (n2904,n2900,n2905);
xnor (n2905,n2906,n887);
nor (n2906,n2907,n2908);
and (n2907,n1202,n1014);
and (n2908,n1198,n1010);
and (n2909,n2898,n2905);
and (n2910,n2896,n2911);
xor (n2911,n2912,n2919);
xor (n2912,n2913,n2915);
and (n2913,n525,n2914);
xnor (n2914,n2899,n525);
xnor (n2915,n2916,n664);
nor (n2916,n2917,n2918);
and (n2917,n1204,n889);
and (n2918,n1202,n885);
xnor (n2919,n2920,n525);
nor (n2920,n2921,n2922);
and (n2921,n1241,n666);
and (n2922,n1227,n662);
and (n2923,n2887,n2911);
xor (n2924,n2925,n2941);
xor (n2925,n2926,n2930);
or (n2926,n2927,n2928,n2929);
and (n2927,n2913,n2915);
and (n2928,n2915,n2919);
and (n2929,n2913,n2919);
xor (n2930,n2931,n2937);
xor (n2931,n2932,n2933);
and (n2932,n2888,n2892);
xnor (n2933,n2934,n664);
nor (n2934,n2935,n2936);
and (n2935,n1202,n889);
and (n2936,n1198,n885);
xnor (n2937,n2938,n525);
nor (n2938,n2939,n2940);
and (n2939,n1227,n666);
and (n2940,n1204,n662);
xor (n2941,n2942,n2948);
xor (n2942,n2943,n2944);
not (n2943,n2748);
xnor (n2944,n2945,n1012);
nor (n2945,n2946,n2947);
and (n2946,n858,n1213);
and (n2947,n854,n1215);
xnor (n2948,n2949,n887);
nor (n2949,n2950,n2951);
and (n2950,n994,n1014);
and (n2951,n860,n1010);
nor (n2952,n2953,n2957);
or (n2953,n2954,n2955,n2956);
and (n2954,n2926,n2930);
and (n2955,n2930,n2941);
and (n2956,n2926,n2941);
xor (n2957,n2958,n2965);
xor (n2958,n2959,n2963);
or (n2959,n2960,n2961,n2962);
and (n2960,n2932,n2933);
and (n2961,n2933,n2937);
and (n2962,n2932,n2937);
xor (n2963,n2964,n2746);
xor (n2964,n2737,n2741);
xor (n2965,n2966,n2972);
xor (n2966,n2967,n2971);
xor (n2967,n2968,n443);
or (n2968,n2969,n2970);
and (n2969,n1227,n523);
and (n2970,n1241,n527);
xor (n2971,n2792,n2796);
or (n2972,n2973,n2974,n2975);
and (n2973,n2943,n2944);
and (n2974,n2944,n2948);
and (n2975,n2943,n2948);
not (n2976,n2977);
not (n2977,n2978);
and (n2978,n2953,n2957);
not (n2979,n2980);
nor (n2980,n2981,n2996);
nor (n2981,n2982,n2986);
nand (n2982,n2983,n2984,n2985);
nand (n2983,n2959,n2963);
nand (n2984,n2965,n2963);
nand (n2985,n2959,n2965);
xor (n2986,n2987,n2994);
xor (n2987,n2988,n2990);
xor (n2988,n2989,n2801);
xor (n2989,n2787,n2791);
nand (n2990,n2991,n2992,n2993);
nand (n2991,n2967,n2971);
nand (n2992,n2972,n2971);
nand (n2993,n2967,n2972);
xor (n2994,n2995,n2751);
xor (n2995,n2734,n2735);
nor (n2996,n2997,n3001);
nand (n2997,n2998,n2999,n3000);
nand (n2998,n2988,n2990);
nand (n2999,n2994,n2990);
nand (n3000,n2988,n2994);
xor (n3001,n3002,n2765);
xor (n3002,n2720,n2732);
not (n3003,n3004);
nor (n3004,n3005,n3007);
nor (n3005,n3006,n2996);
nand (n3006,n2982,n2986);
not (n3007,n3008);
nand (n3008,n2997,n3001);
not (n3009,n3010);
nor (n3010,n3011,n3018);
nor (n3011,n3012,n3017);
nor (n3012,n3013,n3015);
nor (n3013,n3014,n2834);
nand (n3014,n2718,n2807);
not (n3015,n3016);
nand (n3016,n2835,n2839);
not (n3017,n2857);
not (n3018,n3019);
nor (n3019,n3020,n3022);
nor (n3020,n3021,n2873);
nand (n3021,n2859,n2863);
not (n3022,n3023);
nand (n3023,n2874,n2878);
nand (n3024,n3025,n3029);
nor (n3025,n3026,n2715);
nand (n3026,n3027,n2980);
nor (n3027,n3028,n2952);
nor (n3028,n2885,n2924);
or (n3029,n3030,n3052);
and (n3030,n3031,n3033);
xor (n3031,n3032,n2911);
xor (n3032,n2887,n2896);
or (n3033,n3034,n3048,n3051);
and (n3034,n3035,n3044);
and (n3035,n3036,n3040);
xnor (n3036,n3037,n1012);
nor (n3037,n3038,n3039);
and (n3038,n1198,n1213);
and (n3039,n994,n1215);
xnor (n3040,n3041,n887);
nor (n3041,n3042,n3043);
and (n3042,n1204,n1014);
and (n3043,n1202,n1010);
xnor (n3044,n3045,n664);
nor (n3045,n3046,n3047);
and (n3046,n1227,n889);
and (n3047,n1204,n885);
and (n3048,n3044,n3049);
xor (n3049,n3050,n2905);
xor (n3050,n2898,n2900);
and (n3051,n3035,n3049);
and (n3052,n3053,n3054);
xor (n3053,n3031,n3033);
or (n3054,n3055,n3070);
and (n3055,n3056,n3068);
or (n3056,n3057,n3062,n3067);
and (n3057,n3058,n3059);
xor (n3058,n3036,n3040);
and (n3059,n664,n3060);
xnor (n3060,n3061,n664);
nand (n3061,n1241,n885);
and (n3062,n3059,n3063);
xnor (n3063,n3064,n664);
nor (n3064,n3065,n3066);
and (n3065,n1241,n889);
and (n3066,n1227,n885);
and (n3067,n3058,n3063);
xor (n3068,n3069,n3049);
xor (n3069,n3035,n3044);
and (n3070,n3071,n3072);
xor (n3071,n3056,n3068);
or (n3072,n3073,n3089);
and (n3073,n3074,n3076);
xor (n3074,n3075,n3063);
xor (n3075,n3058,n3059);
or (n3076,n3077,n3083,n3088);
and (n3077,n3078,n3079);
not (n3078,n3061);
xnor (n3079,n3080,n1012);
nor (n3080,n3081,n3082);
and (n3081,n1202,n1213);
and (n3082,n1198,n1215);
and (n3083,n3079,n3084);
xnor (n3084,n3085,n887);
nor (n3085,n3086,n3087);
and (n3086,n1227,n1014);
and (n3087,n1204,n1010);
and (n3088,n3078,n3084);
and (n3089,n3090,n3091);
xor (n3090,n3074,n3076);
or (n3091,n3092,n3103);
and (n3092,n3093,n3095);
xor (n3093,n3094,n3084);
xor (n3094,n3078,n3079);
and (n3095,n3096,n3099);
and (n3096,n887,n3097);
xnor (n3097,n3098,n887);
nand (n3098,n1241,n1010);
xnor (n3099,n3100,n1012);
nor (n3100,n3101,n3102);
and (n3101,n1204,n1213);
and (n3102,n1202,n1215);
and (n3103,n3104,n3105);
xor (n3104,n3093,n3095);
or (n3105,n3106,n3112);
and (n3106,n3107,n3111);
xnor (n3107,n3108,n887);
nor (n3108,n3109,n3110);
and (n3109,n1241,n1014);
and (n3110,n1227,n1010);
xor (n3111,n3096,n3099);
and (n3112,n3113,n3114);
xor (n3113,n3107,n3111);
or (n3114,n3115,n3121);
and (n3115,n3116,n3120);
xnor (n3116,n3117,n1012);
nor (n3117,n3118,n3119);
and (n3118,n1227,n1213);
and (n3119,n1204,n1215);
not (n3120,n3098);
and (n3121,n3122,n3123);
xor (n3122,n3116,n3120);
and (n3123,n3124,n3128);
xnor (n3124,n3125,n1012);
nor (n3125,n3126,n3127);
and (n3126,n1241,n1213);
and (n3127,n1227,n1215);
and (n3128,n3129,n1012);
xnor (n3129,n3130,n1012);
nand (n3130,n1241,n1215);
not (n3131,n3132);
nand (n3132,n3133,n2153);
nor (n3133,n3134,n1185);
nand (n3134,n3135,n2108);
nor (n3135,n3136,n2080);
nor (n3136,n1863,n2042);
not (n3137,n3138);
nand (n3138,n3139,n374);
nor (n3139,n3140,n346);
nor (n3140,n154,n310);
not (n3141,n3142);
nor (n3142,n3,n33);
xor (n3143,n3144,n3156);
xor (n3144,n3145,n3147);
not (n3145,n3146);
xnor (n3146,n4,n14);
or (n3147,n3146,n3148);
or (n3148,n3149,n3150,n3155);
not (n3149,n16);
and (n3150,n27,n3151);
or (n3151,n3152,n3153,n3154);
and (n3152,n18,n40);
and (n3153,n40,n127);
and (n3154,n18,n127);
and (n3155,n17,n3151);
and (n3156,n3157,n3158);
xnor (n3157,n3146,n3148);
or (n3158,n3159,n3463);
and (n3159,n3160,n3161);
xor (n3160,n36,n3151);
or (n3161,n3162,n3178,n3462);
and (n3162,n3163,n3165);
xor (n3163,n3164,n127);
xor (n3164,n18,n40);
or (n3165,n3166,n3168,n3177);
and (n3166,n3167,n79);
not (n3167,n55);
and (n3168,n79,n3169);
or (n3169,n3170,n3171,n3176);
and (n3170,n70,n379);
and (n3171,n379,n3172);
or (n3172,n3173,n3174,n3175);
not (n3173,n93);
and (n3174,n104,n117);
and (n3175,n94,n117);
and (n3176,n70,n3172);
and (n3177,n3167,n3169);
and (n3178,n3165,n3179);
or (n3179,n3180,n3220,n3461);
and (n3180,n3181,n3183);
xor (n3181,n3182,n3169);
xor (n3182,n3167,n79);
or (n3183,n3184,n3192,n3219);
and (n3184,n3185,n3190);
or (n3185,n3186,n3187,n3189);
and (n3186,n108,n355);
and (n3187,n355,n3188);
xor (n3188,n360,n117);
and (n3189,n108,n3188);
xor (n3190,n3191,n3172);
xor (n3191,n70,n379);
and (n3192,n3190,n3193);
or (n3193,n3194,n3202,n3218);
and (n3194,n3195,n3200);
or (n3195,n3196,n3197,n3199);
and (n3196,n95,n318);
and (n3197,n318,n3198);
not (n3198,n333);
and (n3199,n95,n3198);
xor (n3200,n3201,n3188);
xor (n3201,n108,n355);
and (n3202,n3200,n3203);
or (n3203,n3204,n3214,n3217);
and (n3204,n3205,n3209);
or (n3205,n3206,n3207,n3208);
and (n3206,n202,n249);
not (n3207,n340);
and (n3208,n202,n252);
or (n3209,n3210,n3211,n3213);
and (n3210,n248,n231);
and (n3211,n231,n3212);
not (n3212,n218);
and (n3213,n248,n3212);
and (n3214,n3209,n3215);
xor (n3215,n3216,n3198);
xor (n3216,n95,n318);
and (n3217,n3205,n3215);
and (n3218,n3195,n3203);
and (n3219,n3185,n3193);
and (n3220,n3183,n3221);
or (n3221,n3222,n3224);
xor (n3222,n3223,n3193);
xor (n3223,n3185,n3190);
or (n3224,n3225,n3256,n3460);
and (n3225,n3226,n3228);
xor (n3226,n3227,n3203);
xor (n3227,n3195,n3200);
or (n3228,n3229,n3241,n3255);
and (n3229,n3230,n3239);
or (n3230,n3231,n3236,n3238);
and (n3231,n3232,n224);
or (n3232,n3233,n3234,n3235);
and (n3233,n248,n205);
not (n3234,n244);
and (n3235,n248,n209);
and (n3236,n224,n3237);
not (n3237,n246);
and (n3238,n3232,n3237);
xor (n3239,n3240,n3215);
xor (n3240,n3205,n3209);
and (n3241,n3239,n3242);
or (n3242,n3243,n3251,n3254);
and (n3243,n3244,n3249);
or (n3244,n3245,n3247,n3248);
and (n3245,n3246,n260);
not (n3246,n200);
and (n3247,n260,n158);
and (n3248,n3246,n158);
xor (n3249,n3250,n3212);
xor (n3250,n248,n231);
and (n3251,n3249,n3252);
xor (n3252,n3253,n3237);
xor (n3253,n3232,n224);
and (n3254,n3244,n3252);
and (n3255,n3230,n3242);
and (n3256,n3228,n3257);
or (n3257,n3258,n3346,n3459);
and (n3258,n3259,n3261);
xor (n3259,n3260,n3242);
xor (n3260,n3230,n3239);
or (n3261,n3262,n3283,n3345);
and (n3262,n3263,n3281);
or (n3263,n3264,n3277,n3280);
and (n3264,n3265,n3269);
or (n3265,n3266,n3267,n3268);
not (n3266,n198);
and (n3267,n192,n263);
and (n3268,n187,n263);
or (n3269,n3270,n3275,n3276);
and (n3270,n269,n3271);
or (n3271,n3272,n3273,n3274);
and (n3272,n161,n291);
not (n3273,n290);
and (n3274,n161,n295);
and (n3275,n3271,n302);
and (n3276,n269,n302);
and (n3277,n3269,n3278);
xor (n3278,n3279,n158);
xor (n3279,n3246,n260);
and (n3280,n3265,n3278);
xor (n3281,n3282,n3252);
xor (n3282,n3244,n3249);
and (n3283,n3281,n3284);
or (n3284,n3285,n3298,n3344);
and (n3285,n3286,n3296);
or (n3286,n3287,n3292,n3295);
and (n3287,n3288,n3290);
xor (n3288,n3289,n263);
xor (n3289,n187,n192);
and (n3290,n414,n3291);
not (n3291,n416);
and (n3292,n3290,n3293);
xor (n3293,n3294,n302);
xor (n3294,n269,n3271);
and (n3295,n3288,n3293);
xor (n3296,n3297,n3278);
xor (n3297,n3265,n3269);
and (n3298,n3296,n3299);
or (n3299,n3300,n3313,n3343);
and (n3300,n3301,n3311);
or (n3301,n3302,n3308,n3310);
and (n3302,n3303,n3304);
not (n3303,n419);
or (n3304,n3305,n3306,n3307);
not (n3305,n436);
and (n3306,n447,n458);
and (n3307,n437,n458);
and (n3308,n3304,n3309);
not (n3309,n413);
and (n3310,n3303,n3309);
xor (n3311,n3312,n3293);
xor (n3312,n3288,n3290);
and (n3313,n3311,n3314);
or (n3314,n3315,n3329,n3342);
and (n3315,n3316,n3320);
or (n3316,n3317,n3318,n3319);
and (n3317,n451,n463);
and (n3318,n463,n505);
and (n3319,n451,n505);
or (n3320,n3321,n3326,n3328);
and (n3321,n472,n3322);
or (n3322,n3323,n3324,n3325);
and (n3323,n438,n491);
not (n3324,n495);
and (n3325,n438,n496);
and (n3326,n3322,n3327);
xor (n3327,n471,n458);
and (n3328,n472,n3327);
and (n3329,n3320,n3330);
or (n3330,n3331,n3338,n3341);
and (n3331,n3332,n3333);
not (n3332,n543);
or (n3333,n3334,n3336,n3337);
and (n3334,n511,n3335);
not (n3335,n587);
and (n3336,n3335,n517);
not (n3337,n538);
and (n3338,n3333,n3339);
xor (n3339,n3340,n505);
xor (n3340,n451,n463);
and (n3341,n3332,n3339);
and (n3342,n3316,n3330);
and (n3343,n3301,n3314);
and (n3344,n3286,n3299);
and (n3345,n3263,n3284);
and (n3346,n3261,n3347);
or (n3347,n3348,n3350);
xor (n3348,n3349,n3284);
xor (n3349,n3263,n3281);
or (n3350,n3351,n3353);
xor (n3351,n3352,n3299);
xor (n3352,n3286,n3296);
or (n3353,n3354,n3386,n3458);
and (n3354,n3355,n3384);
or (n3355,n3356,n3380,n3383);
and (n3356,n3357,n3359);
xor (n3357,n3358,n3309);
xor (n3358,n3303,n3304);
or (n3359,n3360,n3376,n3379);
and (n3360,n3361,n3363);
xor (n3361,n3362,n3327);
xor (n3362,n472,n3322);
or (n3363,n3364,n3370,n3375);
and (n3364,n620,n3365);
and (n3365,n3366,n636);
or (n3366,n3367,n3368,n3369);
and (n3367,n520,n625);
not (n3368,n624);
and (n3369,n520,n629);
and (n3370,n3365,n3371);
or (n3371,n3372,n3373,n3374);
not (n3372,n570);
and (n3373,n571,n596);
and (n3374,n566,n596);
and (n3375,n620,n3371);
and (n3376,n3363,n3377);
xor (n3377,n3378,n3339);
xor (n3378,n3332,n3333);
and (n3379,n3361,n3377);
and (n3380,n3359,n3381);
xor (n3381,n3382,n3330);
xor (n3382,n3316,n3320);
and (n3383,n3357,n3381);
xor (n3384,n3385,n3314);
xor (n3385,n3301,n3311);
and (n3386,n3384,n3387);
or (n3387,n3388,n3390);
xor (n3388,n3389,n3381);
xor (n3389,n3357,n3359);
or (n3390,n3391,n3422,n3457);
and (n3391,n3392,n3420);
or (n3392,n3393,n3402,n3419);
and (n3393,n3394,n3396);
xor (n3394,n3395,n517);
xor (n3395,n511,n3335);
or (n3396,n3397,n3399,n3401);
and (n3397,n3398,n593);
not (n3398,n646);
and (n3399,n593,n3400);
xor (n3400,n3366,n636);
and (n3401,n3398,n3400);
and (n3402,n3396,n3403);
or (n3403,n3404,n3415,n3418);
and (n3404,n3405,n3410);
or (n3405,n3406,n3408,n3409);
and (n3406,n680,n3407);
not (n3407,n1085);
and (n3408,n3407,n1084);
and (n3409,n680,n1084);
or (n3410,n3411,n3413,n3414);
and (n3411,n683,n3412);
not (n3412,n1080);
and (n3413,n3412,n656);
and (n3414,n683,n656);
and (n3415,n3410,n3416);
xor (n3416,n3417,n596);
xor (n3417,n566,n571);
and (n3418,n3405,n3416);
and (n3419,n3394,n3403);
xor (n3420,n3421,n3377);
xor (n3421,n3361,n3363);
and (n3422,n3420,n3423);
or (n3423,n3424,n3453,n3456);
and (n3424,n3425,n3427);
xor (n3425,n3426,n3371);
xor (n3426,n620,n3365);
or (n3427,n3428,n3449,n3452);
and (n3428,n3429,n3447);
or (n3429,n3430,n3443,n3446);
and (n3430,n3431,n3435);
or (n3431,n3432,n3433,n3434);
and (n3432,n764,n838);
and (n3433,n838,n907);
and (n3434,n764,n907);
or (n3435,n3436,n3437,n3442);
and (n3436,n768,n840);
and (n3437,n840,n3438);
or (n3438,n3439,n3440,n3441);
and (n3439,n659,n869);
not (n3440,n905);
and (n3441,n659,n865);
and (n3442,n768,n3438);
and (n3443,n3435,n3444);
xor (n3444,n3445,n1084);
xor (n3445,n680,n3407);
and (n3446,n3431,n3444);
xor (n3447,n3448,n3400);
xor (n3448,n3398,n593);
and (n3449,n3447,n3450);
xor (n3450,n3451,n3416);
xor (n3451,n3405,n3410);
and (n3452,n3429,n3450);
and (n3453,n3427,n3454);
xor (n3454,n3455,n3403);
xor (n3455,n3394,n3396);
and (n3456,n3425,n3454);
and (n3457,n3392,n3423);
and (n3458,n3355,n3387);
and (n3459,n3259,n3347);
and (n3460,n3226,n3257);
and (n3461,n3181,n3221);
and (n3462,n3163,n3179);
and (n3463,n3464,n3465);
xor (n3464,n3160,n3161);
or (n3465,n3466,n3468);
xor (n3466,n3467,n3179);
xor (n3467,n3163,n3165);
and (n3468,n3469,n3470);
not (n3469,n3466);
and (n3470,n3471,n3473);
xor (n3471,n3472,n3221);
xor (n3472,n3181,n3183);
and (n3473,n3474,n3475);
xnor (n3474,n3222,n3224);
and (n3475,n3476,n3478);
xor (n3476,n3477,n3257);
xor (n3477,n3226,n3228);
and (n3478,n3479,n3481);
xor (n3479,n3480,n3347);
xor (n3480,n3259,n3261);
and (n3481,n3482,n3483);
xnor (n3482,n3348,n3350);
and (n3483,n3484,n3485);
xnor (n3484,n3351,n3353);
and (n3485,n3486,n3488);
xor (n3486,n3487,n3387);
xor (n3487,n3355,n3384);
and (n3488,n3489,n3490);
xnor (n3489,n3388,n3390);
or (n3490,n3491,n3571);
and (n3491,n3492,n3494);
xor (n3492,n3493,n3423);
xor (n3493,n3392,n3420);
or (n3494,n3495,n3497);
xor (n3495,n3496,n3454);
xor (n3496,n3425,n3427);
or (n3497,n3498,n3521,n3570);
and (n3498,n3499,n3519);
or (n3499,n3500,n3515,n3518);
and (n3500,n3501,n3503);
xor (n3501,n3502,n656);
xor (n3502,n683,n3412);
or (n3503,n3504,n3511,n3514);
and (n3504,n836,n3505);
or (n3505,n3506,n3508,n3510);
and (n3506,n897,n3507);
not (n3507,n863);
and (n3508,n3507,n3509);
not (n3509,n849);
and (n3510,n897,n3509);
and (n3511,n3505,n3512);
xor (n3512,n3513,n907);
xor (n3513,n764,n838);
and (n3514,n836,n3512);
and (n3515,n3503,n3516);
xor (n3516,n3517,n3444);
xor (n3517,n3431,n3435);
and (n3518,n3501,n3516);
xor (n3519,n3520,n3450);
xor (n3520,n3429,n3447);
and (n3521,n3519,n3522);
or (n3522,n3523,n3534,n3569);
and (n3523,n3524,n3532);
or (n3524,n3525,n3528,n3531);
and (n3525,n3526,n784);
xor (n3526,n3527,n3438);
xor (n3527,n768,n840);
and (n3528,n784,n3529);
xor (n3529,n3530,n3512);
xor (n3530,n836,n3505);
and (n3531,n3526,n3529);
xor (n3532,n3533,n3516);
xor (n3533,n3501,n3503);
and (n3534,n3532,n3535);
or (n3535,n3536,n3565,n3568);
and (n3536,n3537,n3550);
or (n3537,n3538,n3548,n3549);
and (n3538,n3539,n942);
or (n3539,n3540,n3545,n3547);
and (n3540,n3541,n936);
or (n3541,n3542,n3543,n3544);
and (n3542,n881,n926);
not (n3543,n930);
and (n3544,n881,n931);
and (n3545,n936,n3546);
not (n3546,n939);
and (n3547,n3541,n3546);
not (n3548,n977);
and (n3549,n3539,n978);
or (n3550,n3551,n3558,n3564);
and (n3551,n3552,n3556);
or (n3552,n3553,n3554,n3555);
and (n3553,n882,n878);
not (n3554,n896);
and (n3555,n882,n892);
xor (n3556,n3557,n3509);
xor (n3557,n897,n3507);
and (n3558,n3556,n3559);
or (n3559,n3560,n3561,n3563);
and (n3560,n881,n1019);
and (n3561,n1019,n3562);
not (n3562,n2633);
and (n3563,n881,n3562);
and (n3564,n3552,n3559);
and (n3565,n3550,n3566);
xor (n3566,n3567,n3529);
xor (n3567,n3526,n784);
and (n3568,n3537,n3566);
and (n3569,n3524,n3535);
and (n3570,n3499,n3522);
and (n3571,n3572,n3573);
xor (n3572,n3492,n3494);
and (n3573,n3574,n3575);
xnor (n3574,n3495,n3497);
or (n3575,n3576,n3661);
and (n3576,n3577,n3579);
xor (n3577,n3578,n3522);
xor (n3578,n3499,n3519);
or (n3579,n3580,n3582);
xor (n3580,n3581,n3535);
xor (n3581,n3524,n3532);
or (n3582,n3583,n3605,n3660);
and (n3583,n3584,n3603);
or (n3584,n3585,n3599,n3602);
and (n3585,n3586,n3588);
xor (n3586,n3587,n978);
xor (n3587,n3539,n942);
or (n3588,n3589,n3592,n3598);
and (n3589,n3590,n2636);
xor (n3590,n3591,n3546);
xor (n3591,n3541,n936);
and (n3592,n2636,n3593);
or (n3593,n3594,n3595,n3597);
not (n3594,n1058);
and (n3595,n1042,n3596);
not (n3596,n1039);
and (n3597,n1023,n3596);
and (n3598,n3590,n3593);
and (n3599,n3588,n3600);
xor (n3600,n3601,n3559);
xor (n3601,n3552,n3556);
and (n3602,n3586,n3600);
xor (n3603,n3604,n3566);
xor (n3604,n3537,n3550);
and (n3605,n3603,n3606);
or (n3606,n3607,n3622,n3659);
and (n3607,n3608,n3620);
or (n3608,n3609,n3616,n3619);
and (n3609,n3610,n3614);
or (n3610,n3611,n3612,n3613);
and (n3611,n990,n2606);
and (n3612,n2606,n2587);
and (n3613,n990,n2587);
xor (n3614,n3615,n3562);
xor (n3615,n881,n1019);
and (n3616,n3614,n3617);
and (n3617,n2582,n3618);
not (n3618,n2580);
and (n3619,n3610,n3617);
xor (n3620,n3621,n3600);
xor (n3621,n3586,n3588);
and (n3622,n3620,n3623);
or (n3623,n3624,n3644,n3658);
and (n3624,n3625,n3642);
or (n3625,n3626,n3631,n3641);
and (n3626,n3627,n2609);
or (n3627,n3628,n3629,n3630);
and (n3628,n1007,n998);
not (n3629,n997);
and (n3630,n1007,n1001);
and (n3631,n2609,n3632);
or (n3632,n3633,n3638,n3640);
and (n3633,n1006,n3634);
or (n3634,n3635,n3636,n3637);
and (n3635,n1006,n2410);
not (n3636,n2524);
and (n3637,n1006,n2414);
and (n3638,n3634,n3639);
not (n3639,n2519);
and (n3640,n1006,n3639);
and (n3641,n3627,n3632);
xor (n3642,n3643,n3593);
xor (n3643,n3590,n2636);
and (n3644,n3642,n3645);
or (n3645,n3646,n3650,n3657);
and (n3646,n3647,n3649);
xor (n3647,n3648,n2587);
xor (n3648,n990,n2606);
not (n3649,n2579);
and (n3650,n3649,n3651);
or (n3651,n3652,n3655,n3656);
and (n3652,n3653,n2525);
and (n3653,n2394,n3654);
not (n3654,n2408);
and (n3655,n2525,n2547);
and (n3656,n3653,n2547);
and (n3657,n3647,n3651);
and (n3658,n3625,n3645);
and (n3659,n3608,n3623);
and (n3660,n3584,n3606);
and (n3661,n3662,n3663);
xor (n3662,n3577,n3579);
and (n3663,n3664,n3665);
xnor (n3664,n3580,n3582);
or (n3665,n3666,n3870);
and (n3666,n3667,n3669);
xor (n3667,n3668,n3606);
xor (n3668,n3584,n3603);
or (n3669,n3670,n3745,n3869);
and (n3670,n3671,n3743);
or (n3671,n3672,n3739,n3742);
and (n3672,n3673,n3675);
xor (n3673,n3674,n3617);
xor (n3674,n3610,n3614);
or (n3675,n3676,n3710,n3738);
and (n3676,n3677,n3708);
or (n3677,n3678,n3696,n3707);
and (n3678,n3679,n3688);
and (n3679,n3680,n2434);
or (n3680,n3681,n3686,n3687);
and (n3681,n3682,n2304);
or (n3682,n3683,n3684,n3685);
and (n3683,n2373,n2169);
not (n3684,n2313);
and (n3685,n2373,n2173);
not (n3686,n2446);
and (n3687,n3682,n2308);
or (n3688,n3689,n3694,n3695);
and (n3689,n2474,n3690);
or (n3690,n3691,n3692,n3693);
and (n3691,n2373,n2293);
not (n3692,n2421);
and (n3693,n2373,n2298);
and (n3694,n3690,n2455);
and (n3695,n2474,n2455);
and (n3696,n3688,n3697);
or (n3697,n3698,n3704,n3706);
and (n3698,n3699,n3700);
not (n3699,n2393);
or (n3700,n3701,n3702,n3703);
and (n3701,n2177,n2369);
not (n3702,n2473);
and (n3703,n2177,n2374);
and (n3704,n3700,n3705);
not (n3705,n2450);
and (n3706,n3699,n3705);
and (n3707,n3679,n3697);
xor (n3708,n3709,n3632);
xor (n3709,n3627,n2609);
and (n3710,n3708,n3711);
or (n3711,n3712,n3734,n3737);
and (n3712,n3713,n3715);
xor (n3713,n3714,n3639);
xor (n3714,n1006,n3634);
or (n3715,n3716,n3725,n3733);
and (n3716,n3717,n3724);
or (n3717,n3718,n3720,n3723);
and (n3718,n2353,n3719);
not (n3719,n2350);
and (n3720,n3719,n3721);
xor (n3721,n3722,n2298);
xor (n3722,n2373,n2293);
and (n3723,n2353,n3721);
xor (n3724,n3680,n2434);
and (n3725,n3724,n3726);
or (n3726,n3727,n3731,n3732);
and (n3727,n3728,n3729);
not (n3728,n2367);
xor (n3729,n3730,n2308);
xor (n3730,n3682,n2304);
and (n3731,n3729,n2327);
and (n3732,n3728,n2327);
and (n3733,n3717,n3726);
and (n3734,n3715,n3735);
xor (n3735,n3736,n2547);
xor (n3736,n3653,n2525);
and (n3737,n3713,n3735);
and (n3738,n3677,n3711);
and (n3739,n3675,n3740);
xor (n3740,n3741,n3645);
xor (n3741,n3625,n3642);
and (n3742,n3673,n3740);
xor (n3743,n3744,n3623);
xor (n3744,n3608,n3620);
and (n3745,n3743,n3746);
or (n3746,n3747,n3780,n3868);
and (n3747,n3748,n3778);
or (n3748,n3749,n3774,n3777);
and (n3749,n3750,n3752);
xor (n3750,n3751,n3651);
xor (n3751,n3647,n3649);
or (n3752,n3753,n3770,n3773);
and (n3753,n3754,n3756);
xor (n3754,n3755,n3697);
xor (n3755,n3679,n3688);
or (n3756,n3757,n3762,n3769);
and (n3757,n3758,n3760);
xor (n3758,n3759,n2455);
xor (n3759,n2474,n3690);
xor (n3760,n3761,n3705);
xor (n3761,n3699,n3700);
and (n3762,n3760,n3763);
and (n3763,n2318,n3764);
or (n3764,n3765,n3766,n3768);
not (n3765,n2324);
and (n3766,n2184,n3767);
not (n3767,n2167);
and (n3768,n2180,n3767);
and (n3769,n3758,n3763);
and (n3770,n3756,n3771);
xor (n3771,n3772,n3735);
xor (n3772,n3713,n3715);
and (n3773,n3754,n3771);
and (n3774,n3752,n3775);
xor (n3775,n3776,n3711);
xor (n3776,n3677,n3708);
and (n3777,n3750,n3775);
xor (n3778,n3779,n3740);
xor (n3779,n3673,n3675);
and (n3780,n3778,n3781);
or (n3781,n3782,n3839,n3867);
and (n3782,n3783,n3785);
xor (n3783,n3784,n3775);
xor (n3784,n3750,n3752);
or (n3785,n3786,n3818,n3838);
and (n3786,n3787,n3816);
or (n3787,n3788,n3801,n3815);
and (n3788,n3789,n3799);
or (n3789,n3790,n3797,n3798);
and (n3790,n3791,n3795);
or (n3791,n3792,n3793,n3794);
and (n3792,n2232,n2217);
and (n3793,n2217,n2200);
and (n3794,n2232,n2200);
xor (n3795,n3796,n3721);
xor (n3796,n2353,n3719);
and (n3797,n3795,n2378);
and (n3798,n3791,n2378);
xor (n3799,n3800,n3726);
xor (n3800,n3717,n3724);
and (n3801,n3799,n3802);
or (n3802,n3803,n3812,n3814);
and (n3803,n3804,n3810);
or (n3804,n3805,n3806,n3809);
and (n3805,n2222,n2216);
and (n3806,n2216,n3807);
xor (n3807,n3808,n2200);
xor (n3808,n2232,n2217);
and (n3809,n2222,n3807);
xor (n3810,n3811,n2327);
xor (n3811,n3728,n3729);
and (n3812,n3810,n3813);
xor (n3813,n2318,n3764);
and (n3814,n3804,n3813);
and (n3815,n3789,n3802);
xor (n3816,n3817,n3771);
xor (n3817,n3754,n3756);
and (n3818,n3816,n3819);
or (n3819,n3820,n3834,n3837);
and (n3820,n3821,n3823);
xor (n3821,n3822,n3763);
xor (n3822,n3758,n3760);
or (n3823,n3824,n3832,n3833);
and (n3824,n3825,n3827);
xor (n3825,n3826,n2378);
xor (n3826,n3791,n3795);
or (n3827,n3828,n3829,n3831);
not (n3828,n2277);
and (n3829,n2192,n3830);
not (n3830,n2165);
and (n3831,n2188,n3830);
and (n3832,n3827,n2279);
and (n3833,n3825,n2279);
and (n3834,n3823,n3835);
xor (n3835,n3836,n3802);
xor (n3836,n3789,n3799);
and (n3837,n3821,n3835);
and (n3838,n3787,n3819);
and (n3839,n3785,n3840);
or (n3840,n3841,n3843);
xor (n3841,n3842,n3819);
xor (n3842,n3787,n3816);
or (n3843,n3844,n3860,n3866);
and (n3844,n3845,n3858);
or (n3845,n3846,n3854,n3857);
and (n3846,n3847,n3849);
xor (n3847,n3848,n3813);
xor (n3848,n3804,n3810);
or (n3849,n3850,n3852,n3853);
and (n3850,n3851,n2264);
not (n3851,n2163);
not (n3852,n2271);
and (n3853,n3851,n2196);
and (n3854,n3849,n3855);
xor (n3855,n3856,n2279);
xor (n3856,n3825,n3827);
and (n3857,n3847,n3855);
xor (n3858,n3859,n3835);
xor (n3859,n3821,n3823);
and (n3860,n3858,n3861);
or (n3861,n3862,n3864);
or (n3862,n2157,n3863);
not (n3863,n2161);
xor (n3864,n3865,n3855);
xor (n3865,n3847,n3849);
and (n3866,n3845,n3861);
and (n3867,n3783,n3840);
and (n3868,n3748,n3781);
and (n3869,n3671,n3746);
and (n3870,n3871,n3872);
xor (n3871,n3667,n3669);
and (n3872,n3873,n3875);
xor (n3873,n3874,n3746);
xor (n3874,n3671,n3743);
or (n3875,n3876,n3878);
xor (n3876,n3877,n3781);
xor (n3877,n3748,n3778);
and (n3878,n3879,n3880);
not (n3879,n3876);
and (n3880,n3881,n3883);
xor (n3881,n3882,n3840);
xor (n3882,n3783,n3785);
and (n3883,n3884,n3885);
xnor (n3884,n3841,n3843);
and (n3885,n3886,n3888);
xor (n3886,n3887,n3861);
xor (n3887,n3845,n3858);
and (n3888,n3889,n3890);
xnor (n3889,n3862,n3864);
and (n3890,n3891,n3894);
not (n3891,n3892);
nand (n3892,n3893,n2686);
not (n3893,n2156);
nand (n3894,n1183,n3895);
nand (n3895,n3133,n2712);
endmodule
