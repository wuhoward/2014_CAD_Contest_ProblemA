module top (out,n25,n30,n31,n32,n34,n35,n46,n49,n52
        ,n55,n58,n61,n64,n67,n70,n73,n76,n79,n81
        ,n84,n101,n106,n109,n112,n115,n118,n121,n124,n127
        ,n130,n133,n136,n139,n142,n145,n147,n149,n158,n171
        ,n176,n179,n182,n185,n198,n226,n236,n270,n280,n308
        ,n315,n347,n357,n406,n411,n414,n417,n420,n423,n426
        ,n429,n432,n435,n444,n716,n758,n1074,n1101);
output out;
input n25;
input n30;
input n31;
input n32;
input n34;
input n35;
input n46;
input n49;
input n52;
input n55;
input n58;
input n61;
input n64;
input n67;
input n70;
input n73;
input n76;
input n79;
input n81;
input n84;
input n101;
input n106;
input n109;
input n112;
input n115;
input n118;
input n121;
input n124;
input n127;
input n130;
input n133;
input n136;
input n139;
input n142;
input n145;
input n147;
input n149;
input n158;
input n171;
input n176;
input n179;
input n182;
input n185;
input n198;
input n226;
input n236;
input n270;
input n280;
input n308;
input n315;
input n347;
input n357;
input n406;
input n411;
input n414;
input n417;
input n420;
input n423;
input n426;
input n429;
input n432;
input n435;
input n444;
input n716;
input n758;
input n1074;
input n1101;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n26;
wire n27;
wire n28;
wire n29;
wire n33;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n47;
wire n48;
wire n50;
wire n51;
wire n53;
wire n54;
wire n56;
wire n57;
wire n59;
wire n60;
wire n62;
wire n63;
wire n65;
wire n66;
wire n68;
wire n69;
wire n71;
wire n72;
wire n74;
wire n75;
wire n77;
wire n78;
wire n80;
wire n82;
wire n83;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n102;
wire n103;
wire n104;
wire n105;
wire n107;
wire n108;
wire n110;
wire n111;
wire n113;
wire n114;
wire n116;
wire n117;
wire n119;
wire n120;
wire n122;
wire n123;
wire n125;
wire n126;
wire n128;
wire n129;
wire n131;
wire n132;
wire n134;
wire n135;
wire n137;
wire n138;
wire n140;
wire n141;
wire n143;
wire n144;
wire n146;
wire n148;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n172;
wire n173;
wire n174;
wire n175;
wire n177;
wire n178;
wire n180;
wire n181;
wire n183;
wire n184;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n407;
wire n408;
wire n409;
wire n410;
wire n412;
wire n413;
wire n415;
wire n416;
wire n418;
wire n419;
wire n421;
wire n422;
wire n424;
wire n425;
wire n427;
wire n428;
wire n430;
wire n431;
wire n433;
wire n434;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2988;
wire n2989;
wire n2990;
wire n2991;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2996;
wire n2997;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3003;
wire n3004;
wire n3005;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3010;
wire n3011;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3038;
wire n3039;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
wire n3056;
wire n3057;
wire n3058;
wire n3059;
wire n3060;
wire n3061;
wire n3062;
wire n3063;
wire n3064;
wire n3065;
wire n3066;
wire n3067;
wire n3068;
wire n3069;
wire n3070;
wire n3071;
wire n3072;
wire n3073;
wire n3074;
wire n3075;
wire n3076;
wire n3077;
wire n3078;
wire n3079;
wire n3080;
wire n3081;
wire n3082;
wire n3083;
wire n3084;
wire n3085;
wire n3086;
wire n3087;
wire n3088;
wire n3089;
wire n3090;
wire n3091;
wire n3092;
wire n3093;
wire n3094;
wire n3095;
wire n3096;
wire n3097;
wire n3098;
wire n3099;
wire n3100;
wire n3101;
wire n3102;
wire n3103;
wire n3104;
wire n3105;
wire n3106;
wire n3107;
wire n3108;
wire n3109;
wire n3110;
wire n3111;
wire n3112;
wire n3113;
wire n3114;
wire n3115;
wire n3116;
wire n3117;
wire n3118;
wire n3119;
wire n3120;
wire n3121;
wire n3122;
wire n3123;
wire n3124;
wire n3125;
wire n3126;
wire n3127;
wire n3128;
wire n3129;
wire n3130;
wire n3131;
wire n3132;
wire n3133;
wire n3134;
wire n3135;
wire n3136;
wire n3137;
wire n3138;
wire n3139;
wire n3140;
wire n3141;
wire n3142;
wire n3143;
wire n3144;
wire n3145;
wire n3146;
wire n3147;
wire n3148;
wire n3149;
wire n3150;
wire n3151;
wire n3152;
wire n3153;
wire n3154;
wire n3155;
wire n3156;
wire n3157;
wire n3158;
wire n3159;
wire n3160;
wire n3161;
wire n3162;
wire n3163;
wire n3164;
wire n3165;
wire n3166;
wire n3167;
wire n3168;
wire n3169;
wire n3170;
wire n3171;
wire n3172;
wire n3173;
wire n3174;
wire n3175;
wire n3176;
wire n3177;
wire n3178;
wire n3179;
wire n3180;
wire n3181;
wire n3182;
wire n3183;
wire n3184;
wire n3185;
wire n3186;
wire n3187;
wire n3188;
wire n3189;
wire n3190;
wire n3191;
wire n3192;
wire n3193;
wire n3194;
wire n3195;
wire n3196;
wire n3197;
wire n3198;
wire n3199;
wire n3200;
wire n3201;
wire n3202;
wire n3203;
wire n3204;
wire n3205;
wire n3206;
wire n3207;
wire n3208;
wire n3209;
wire n3210;
wire n3211;
wire n3212;
wire n3213;
wire n3214;
wire n3215;
wire n3216;
wire n3217;
wire n3218;
wire n3219;
wire n3220;
wire n3221;
wire n3222;
wire n3223;
wire n3224;
wire n3225;
wire n3226;
wire n3227;
wire n3228;
wire n3229;
wire n3230;
wire n3231;
wire n3232;
wire n3233;
wire n3234;
wire n3235;
wire n3236;
wire n3237;
wire n3238;
wire n3239;
wire n3240;
wire n3241;
wire n3242;
wire n3243;
wire n3244;
wire n3245;
wire n3246;
wire n3247;
wire n3248;
wire n3249;
wire n3250;
wire n3251;
wire n3252;
wire n3253;
wire n3254;
wire n3255;
wire n3256;
wire n3257;
wire n3258;
wire n3259;
wire n3260;
wire n3261;
wire n3262;
wire n3263;
wire n3264;
wire n3265;
wire n3266;
wire n3267;
wire n3268;
wire n3269;
wire n3270;
wire n3271;
wire n3272;
wire n3273;
wire n3274;
wire n3275;
wire n3276;
wire n3277;
wire n3278;
wire n3279;
wire n3280;
wire n3281;
wire n3282;
wire n3283;
wire n3284;
wire n3285;
wire n3286;
wire n3287;
wire n3288;
wire n3289;
wire n3290;
wire n3291;
wire n3292;
wire n3293;
wire n3294;
wire n3295;
wire n3296;
wire n3297;
wire n3298;
wire n3299;
wire n3300;
wire n3301;
wire n3302;
wire n3303;
wire n3304;
wire n3305;
wire n3306;
wire n3307;
wire n3308;
wire n3309;
wire n3310;
wire n3311;
wire n3312;
wire n3313;
wire n3314;
wire n3315;
wire n3316;
wire n3317;
wire n3318;
wire n3319;
wire n3320;
wire n3321;
wire n3322;
wire n3323;
wire n3324;
wire n3325;
wire n3326;
wire n3327;
wire n3328;
wire n3329;
wire n3330;
wire n3331;
wire n3332;
wire n3333;
wire n3334;
wire n3335;
wire n3336;
wire n3337;
wire n3338;
wire n3339;
wire n3340;
wire n3341;
wire n3342;
wire n3343;
wire n3344;
wire n3345;
wire n3346;
wire n3347;
wire n3348;
wire n3349;
wire n3350;
wire n3351;
wire n3352;
wire n3353;
wire n3354;
wire n3355;
wire n3356;
wire n3357;
wire n3358;
wire n3359;
wire n3360;
wire n3361;
wire n3362;
wire n3363;
wire n3364;
wire n3365;
wire n3366;
wire n3367;
wire n3368;
wire n3369;
wire n3370;
wire n3371;
wire n3372;
wire n3373;
wire n3374;
wire n3375;
wire n3376;
wire n3377;
wire n3378;
wire n3379;
wire n3380;
wire n3381;
wire n3382;
wire n3383;
wire n3384;
wire n3385;
wire n3386;
wire n3387;
wire n3388;
wire n3389;
wire n3390;
wire n3391;
wire n3392;
wire n3393;
wire n3394;
wire n3395;
wire n3396;
wire n3397;
wire n3398;
wire n3399;
wire n3400;
wire n3401;
wire n3402;
wire n3403;
wire n3404;
wire n3405;
wire n3406;
wire n3407;
wire n3408;
wire n3409;
wire n3410;
wire n3411;
wire n3412;
wire n3413;
wire n3414;
wire n3415;
wire n3416;
wire n3417;
wire n3418;
wire n3419;
wire n3420;
wire n3421;
wire n3422;
wire n3423;
wire n3424;
wire n3425;
wire n3426;
wire n3427;
wire n3428;
wire n3429;
wire n3430;
wire n3431;
wire n3432;
wire n3433;
wire n3434;
wire n3435;
wire n3436;
wire n3437;
wire n3438;
wire n3439;
wire n3440;
wire n3441;
wire n3442;
wire n3443;
wire n3444;
wire n3445;
wire n3446;
wire n3447;
wire n3448;
wire n3449;
wire n3450;
wire n3451;
wire n3452;
wire n3453;
wire n3454;
wire n3455;
wire n3456;
wire n3457;
wire n3458;
wire n3459;
wire n3460;
wire n3461;
wire n3462;
wire n3463;
wire n3464;
wire n3465;
wire n3466;
wire n3467;
wire n3468;
wire n3469;
wire n3470;
wire n3471;
wire n3472;
wire n3473;
wire n3474;
wire n3475;
wire n3476;
wire n3477;
wire n3478;
wire n3479;
wire n3480;
wire n3481;
wire n3482;
wire n3483;
wire n3484;
wire n3485;
wire n3486;
wire n3487;
wire n3488;
wire n3489;
wire n3490;
wire n3491;
wire n3492;
wire n3493;
wire n3494;
wire n3495;
wire n3496;
wire n3497;
wire n3498;
wire n3499;
wire n3500;
wire n3501;
wire n3502;
wire n3503;
wire n3504;
wire n3505;
wire n3506;
wire n3507;
wire n3508;
wire n3509;
wire n3510;
wire n3511;
wire n3512;
wire n3513;
wire n3514;
wire n3515;
wire n3516;
wire n3517;
wire n3518;
wire n3519;
wire n3520;
wire n3521;
wire n3522;
wire n3523;
wire n3524;
wire n3525;
wire n3526;
wire n3527;
wire n3528;
wire n3529;
wire n3530;
wire n3531;
wire n3532;
wire n3533;
wire n3534;
wire n3535;
wire n3536;
wire n3537;
wire n3538;
wire n3539;
wire n3540;
wire n3541;
wire n3542;
wire n3543;
wire n3544;
wire n3545;
wire n3546;
wire n3547;
wire n3548;
wire n3549;
wire n3550;
wire n3551;
wire n3552;
wire n3553;
wire n3554;
wire n3555;
wire n3556;
wire n3557;
wire n3558;
wire n3559;
wire n3560;
wire n3561;
wire n3562;
wire n3563;
wire n3564;
wire n3565;
wire n3566;
wire n3567;
wire n3568;
wire n3569;
wire n3570;
wire n3571;
wire n3572;
wire n3573;
wire n3574;
wire n3575;
wire n3576;
wire n3577;
wire n3578;
wire n3579;
wire n3580;
wire n3581;
wire n3582;
wire n3583;
wire n3584;
wire n3585;
wire n3586;
wire n3587;
wire n3588;
wire n3589;
wire n3590;
wire n3591;
wire n3592;
wire n3593;
wire n3594;
wire n3595;
wire n3596;
wire n3597;
wire n3598;
wire n3599;
wire n3600;
wire n3601;
wire n3602;
wire n3603;
wire n3604;
wire n3605;
wire n3606;
wire n3607;
wire n3608;
wire n3609;
wire n3610;
wire n3611;
wire n3612;
wire n3613;
wire n3614;
wire n3615;
wire n3616;
wire n3617;
wire n3618;
wire n3619;
wire n3620;
wire n3621;
wire n3622;
wire n3623;
wire n3624;
wire n3625;
wire n3626;
wire n3627;
wire n3628;
wire n3629;
wire n3630;
wire n3631;
wire n3632;
wire n3633;
wire n3634;
wire n3635;
wire n3636;
wire n3637;
wire n3638;
wire n3639;
wire n3640;
wire n3641;
wire n3642;
wire n3643;
wire n3644;
wire n3645;
wire n3646;
wire n3647;
wire n3648;
wire n3649;
wire n3650;
wire n3651;
wire n3652;
wire n3653;
wire n3654;
wire n3655;
wire n3656;
wire n3657;
wire n3658;
wire n3659;
wire n3660;
wire n3661;
wire n3662;
wire n3663;
wire n3664;
wire n3665;
wire n3666;
wire n3667;
wire n3668;
wire n3669;
wire n3670;
wire n3671;
wire n3672;
wire n3673;
wire n3674;
wire n3675;
wire n3676;
wire n3677;
wire n3678;
wire n3679;
wire n3680;
wire n3681;
wire n3682;
wire n3683;
wire n3684;
wire n3685;
wire n3686;
wire n3687;
wire n3688;
wire n3689;
wire n3690;
wire n3691;
wire n3692;
wire n3693;
wire n3694;
wire n3695;
wire n3696;
wire n3697;
wire n3698;
wire n3699;
wire n3700;
wire n3701;
wire n3702;
wire n3703;
wire n3704;
wire n3705;
wire n3706;
wire n3707;
wire n3708;
wire n3709;
wire n3710;
wire n3711;
wire n3712;
wire n3713;
wire n3714;
wire n3715;
wire n3716;
wire n3717;
wire n3718;
wire n3719;
wire n3720;
wire n3721;
wire n3722;
wire n3723;
wire n3724;
wire n3725;
wire n3726;
wire n3727;
wire n3728;
wire n3729;
wire n3730;
wire n3731;
wire n3732;
wire n3733;
wire n3734;
wire n3735;
wire n3736;
wire n3737;
wire n3738;
wire n3739;
wire n3740;
wire n3741;
wire n3742;
wire n3743;
wire n3744;
wire n3745;
wire n3746;
wire n3747;
wire n3748;
wire n3749;
wire n3750;
wire n3751;
wire n3752;
wire n3753;
wire n3754;
wire n3755;
wire n3756;
wire n3757;
wire n3758;
wire n3759;
wire n3760;
wire n3761;
wire n3762;
wire n3763;
wire n3764;
wire n3765;
wire n3766;
wire n3767;
wire n3768;
wire n3769;
wire n3770;
wire n3771;
wire n3772;
wire n3773;
wire n3774;
wire n3775;
wire n3776;
wire n3777;
wire n3778;
wire n3779;
wire n3780;
wire n3781;
wire n3782;
wire n3783;
wire n3784;
wire n3785;
wire n3786;
wire n3787;
wire n3788;
wire n3789;
wire n3790;
wire n3791;
wire n3792;
wire n3793;
wire n3794;
wire n3795;
wire n3796;
wire n3797;
wire n3798;
wire n3799;
wire n3800;
wire n3801;
wire n3802;
wire n3803;
wire n3804;
wire n3805;
wire n3806;
wire n3807;
wire n3808;
wire n3809;
wire n3810;
wire n3811;
wire n3812;
wire n3813;
wire n3814;
wire n3815;
wire n3816;
wire n3817;
wire n3818;
wire n3819;
wire n3820;
wire n3821;
wire n3822;
wire n3823;
wire n3824;
wire n3825;
wire n3826;
wire n3827;
wire n3828;
wire n3829;
wire n3830;
wire n3831;
wire n3832;
wire n3833;
wire n3834;
wire n3835;
wire n3836;
wire n3837;
wire n3838;
wire n3839;
wire n3840;
wire n3841;
wire n3842;
wire n3843;
wire n3844;
wire n3845;
wire n3846;
wire n3847;
wire n3848;
wire n3849;
wire n3850;
wire n3851;
wire n3852;
wire n3853;
wire n3854;
wire n3855;
wire n3856;
wire n3857;
wire n3858;
wire n3859;
wire n3860;
wire n3861;
wire n3862;
wire n3863;
wire n3864;
wire n3865;
wire n3866;
wire n3867;
wire n3868;
wire n3869;
wire n3870;
wire n3871;
wire n3872;
wire n3873;
wire n3874;
wire n3875;
wire n3876;
wire n3877;
wire n3878;
wire n3879;
wire n3880;
wire n3881;
wire n3882;
wire n3883;
wire n3884;
wire n3885;
wire n3886;
wire n3887;
wire n3888;
wire n3889;
wire n3890;
wire n3891;
wire n3892;
wire n3893;
wire n3894;
wire n3895;
wire n3896;
wire n3897;
wire n3898;
wire n3899;
wire n3900;
wire n3901;
wire n3902;
wire n3903;
wire n3904;
wire n3905;
wire n3906;
wire n3907;
wire n3908;
wire n3909;
wire n3910;
wire n3911;
wire n3912;
wire n3913;
wire n3914;
wire n3915;
wire n3916;
wire n3917;
wire n3918;
wire n3919;
wire n3920;
wire n3921;
wire n3922;
wire n3923;
wire n3924;
wire n3925;
wire n3926;
wire n3927;
wire n3928;
wire n3929;
wire n3930;
wire n3931;
wire n3932;
wire n3933;
wire n3934;
wire n3935;
wire n3936;
wire n3937;
wire n3938;
wire n3939;
wire n3940;
wire n3941;
wire n3942;
wire n3943;
wire n3944;
wire n3945;
wire n3946;
wire n3947;
wire n3948;
wire n3949;
wire n3950;
wire n3951;
wire n3952;
wire n3953;
wire n3954;
wire n3955;
wire n3956;
wire n3957;
wire n3958;
wire n3959;
wire n3960;
wire n3961;
wire n3962;
wire n3963;
wire n3964;
wire n3965;
wire n3966;
wire n3967;
wire n3968;
wire n3969;
wire n3970;
wire n3971;
wire n3972;
wire n3973;
wire n3974;
wire n3975;
wire n3976;
wire n3977;
wire n3978;
wire n3979;
wire n3980;
wire n3981;
wire n3982;
wire n3983;
wire n3984;
wire n3985;
wire n3986;
wire n3987;
wire n3988;
wire n3989;
wire n3990;
wire n3991;
wire n3992;
wire n3993;
wire n3994;
wire n3995;
wire n3996;
wire n3997;
wire n3998;
wire n3999;
wire n4000;
wire n4001;
wire n4002;
wire n4003;
wire n4004;
wire n4005;
wire n4006;
wire n4007;
wire n4008;
wire n4009;
wire n4010;
wire n4011;
wire n4012;
wire n4013;
wire n4014;
wire n4015;
wire n4016;
wire n4017;
wire n4018;
wire n4019;
wire n4020;
wire n4021;
wire n4022;
wire n4023;
wire n4024;
wire n4025;
wire n4026;
wire n4027;
wire n4028;
wire n4029;
wire n4030;
wire n4031;
wire n4032;
wire n4033;
wire n4034;
wire n4035;
wire n4036;
wire n4037;
wire n4038;
wire n4039;
wire n4040;
wire n4041;
wire n4042;
wire n4043;
wire n4044;
wire n4045;
wire n4046;
wire n4047;
wire n4048;
wire n4049;
wire n4050;
wire n4051;
wire n4052;
wire n4053;
wire n4054;
wire n4055;
wire n4056;
wire n4057;
wire n4058;
wire n4059;
wire n4060;
wire n4061;
wire n4062;
wire n4063;
wire n4064;
wire n4065;
wire n4066;
wire n4067;
wire n4068;
wire n4069;
wire n4070;
wire n4071;
wire n4072;
wire n4073;
wire n4074;
wire n4075;
wire n4076;
wire n4077;
wire n4078;
wire n4079;
wire n4080;
wire n4081;
wire n4082;
wire n4083;
wire n4084;
wire n4085;
wire n4086;
wire n4087;
wire n4088;
wire n4089;
wire n4090;
wire n4091;
wire n4092;
wire n4093;
wire n4094;
wire n4095;
wire n4096;
wire n4097;
wire n4098;
wire n4099;
wire n4100;
wire n4101;
wire n4102;
wire n4103;
wire n4104;
wire n4105;
wire n4106;
wire n4107;
wire n4108;
wire n4109;
wire n4110;
wire n4111;
wire n4112;
wire n4113;
wire n4114;
wire n4115;
wire n4116;
wire n4117;
wire n4118;
wire n4119;
wire n4120;
wire n4121;
wire n4122;
wire n4123;
wire n4124;
wire n4125;
wire n4126;
wire n4127;
wire n4128;
wire n4129;
wire n4130;
wire n4131;
wire n4132;
wire n4133;
wire n4134;
wire n4135;
wire n4136;
wire n4137;
wire n4138;
wire n4139;
wire n4140;
wire n4141;
wire n4142;
wire n4143;
wire n4144;
wire n4145;
wire n4146;
wire n4147;
wire n4148;
wire n4149;
wire n4150;
wire n4151;
wire n4152;
wire n4153;
wire n4154;
wire n4155;
wire n4156;
wire n4157;
wire n4158;
wire n4159;
wire n4160;
wire n4161;
wire n4162;
wire n4163;
wire n4164;
wire n4165;
wire n4166;
wire n4167;
wire n4168;
wire n4169;
wire n4170;
wire n4171;
wire n4172;
wire n4173;
wire n4174;
wire n4175;
wire n4176;
wire n4177;
wire n4178;
wire n4179;
wire n4180;
wire n4181;
wire n4182;
wire n4183;
wire n4184;
wire n4185;
wire n4186;
wire n4187;
wire n4188;
wire n4189;
wire n4190;
wire n4191;
wire n4192;
wire n4193;
wire n4194;
wire n4195;
wire n4196;
wire n4197;
wire n4198;
wire n4199;
wire n4200;
wire n4201;
wire n4202;
wire n4203;
wire n4204;
wire n4205;
wire n4206;
wire n4207;
wire n4208;
wire n4209;
wire n4210;
wire n4211;
wire n4212;
wire n4213;
wire n4214;
wire n4215;
wire n4216;
wire n4217;
wire n4218;
wire n4219;
wire n4220;
wire n4221;
wire n4222;
wire n4223;
wire n4224;
wire n4225;
wire n4226;
wire n4227;
wire n4228;
wire n4229;
wire n4230;
wire n4231;
wire n4232;
wire n4233;
wire n4234;
wire n4235;
wire n4236;
wire n4237;
wire n4238;
wire n4239;
wire n4240;
wire n4241;
wire n4242;
wire n4243;
wire n4244;
wire n4245;
wire n4246;
wire n4247;
wire n4248;
wire n4249;
wire n4250;
wire n4251;
wire n4252;
wire n4253;
wire n4254;
wire n4255;
wire n4256;
wire n4257;
wire n4258;
wire n4259;
wire n4260;
wire n4261;
wire n4262;
wire n4263;
wire n4264;
wire n4265;
wire n4266;
wire n4267;
wire n4268;
wire n4269;
wire n4270;
wire n4271;
wire n4272;
wire n4273;
wire n4274;
wire n4275;
wire n4276;
wire n4277;
wire n4278;
wire n4279;
wire n4280;
wire n4281;
wire n4282;
wire n4283;
wire n4284;
wire n4285;
wire n4286;
wire n4287;
wire n4288;
wire n4289;
wire n4290;
wire n4291;
wire n4292;
wire n4293;
wire n4294;
wire n4295;
wire n4296;
wire n4297;
wire n4298;
wire n4299;
wire n4300;
wire n4301;
wire n4302;
wire n4303;
wire n4304;
wire n4305;
wire n4306;
wire n4307;
wire n4308;
wire n4309;
wire n4310;
wire n4311;
wire n4312;
wire n4313;
wire n4314;
wire n4315;
wire n4316;
wire n4317;
wire n4318;
wire n4319;
wire n4320;
wire n4321;
wire n4322;
wire n4323;
wire n4324;
wire n4325;
wire n4326;
wire n4327;
wire n4328;
wire n4329;
wire n4330;
wire n4331;
wire n4332;
wire n4333;
wire n4334;
wire n4335;
wire n4336;
wire n4337;
wire n4338;
wire n4339;
wire n4340;
wire n4341;
wire n4342;
wire n4343;
wire n4344;
wire n4345;
wire n4346;
wire n4347;
wire n4348;
wire n4349;
wire n4350;
wire n4351;
wire n4352;
wire n4353;
wire n4354;
wire n4355;
wire n4356;
wire n4357;
wire n4358;
wire n4359;
wire n4360;
wire n4361;
wire n4362;
wire n4363;
wire n4364;
wire n4365;
wire n4366;
wire n4367;
wire n4368;
wire n4369;
wire n4370;
wire n4371;
wire n4372;
wire n4373;
wire n4374;
wire n4375;
wire n4376;
wire n4377;
wire n4378;
wire n4379;
wire n4380;
wire n4381;
wire n4382;
wire n4383;
wire n4384;
wire n4385;
wire n4386;
wire n4387;
wire n4388;
wire n4389;
wire n4390;
wire n4391;
wire n4392;
wire n4393;
wire n4394;
wire n4395;
wire n4396;
wire n4397;
wire n4398;
wire n4399;
wire n4400;
wire n4401;
wire n4402;
wire n4403;
wire n4404;
wire n4405;
wire n4406;
wire n4407;
wire n4408;
wire n4409;
wire n4410;
wire n4411;
wire n4412;
wire n4413;
wire n4414;
wire n4415;
wire n4416;
wire n4417;
wire n4418;
wire n4419;
wire n4420;
wire n4421;
wire n4422;
wire n4423;
wire n4424;
wire n4425;
wire n4426;
wire n4427;
wire n4428;
wire n4429;
wire n4430;
wire n4431;
wire n4432;
wire n4433;
wire n4434;
wire n4435;
wire n4436;
wire n4437;
wire n4438;
wire n4439;
wire n4440;
wire n4441;
wire n4442;
wire n4443;
wire n4444;
wire n4445;
wire n4446;
wire n4447;
wire n4448;
wire n4449;
wire n4450;
wire n4451;
wire n4452;
wire n4453;
wire n4454;
wire n4455;
wire n4456;
wire n4457;
wire n4458;
wire n4459;
wire n4460;
wire n4461;
wire n4462;
wire n4463;
wire n4464;
wire n4465;
wire n4466;
wire n4467;
wire n4468;
wire n4469;
wire n4470;
wire n4471;
wire n4472;
wire n4473;
wire n4474;
wire n4475;
wire n4476;
wire n4477;
wire n4478;
wire n4479;
wire n4480;
wire n4481;
wire n4482;
wire n4483;
wire n4484;
wire n4485;
wire n4486;
wire n4487;
wire n4488;
wire n4489;
wire n4490;
wire n4491;
wire n4492;
wire n4493;
wire n4494;
wire n4495;
wire n4496;
wire n4497;
wire n4498;
wire n4499;
wire n4500;
wire n4501;
wire n4502;
wire n4503;
wire n4504;
wire n4505;
wire n4506;
wire n4507;
wire n4508;
wire n4509;
wire n4510;
wire n4511;
wire n4512;
wire n4513;
wire n4514;
wire n4515;
wire n4516;
wire n4517;
wire n4518;
wire n4519;
wire n4520;
wire n4521;
wire n4522;
wire n4523;
wire n4524;
wire n4525;
wire n4526;
wire n4527;
wire n4528;
wire n4529;
wire n4530;
wire n4531;
wire n4532;
wire n4533;
wire n4534;
wire n4535;
wire n4536;
wire n4537;
wire n4538;
wire n4539;
wire n4540;
wire n4541;
wire n4542;
wire n4543;
wire n4544;
wire n4545;
wire n4546;
wire n4547;
wire n4548;
wire n4549;
wire n4550;
wire n4551;
wire n4552;
wire n4553;
wire n4554;
wire n4555;
wire n4556;
wire n4557;
wire n4558;
wire n4559;
wire n4560;
wire n4561;
wire n4562;
wire n4563;
wire n4564;
wire n4565;
wire n4566;
wire n4567;
wire n4568;
wire n4569;
wire n4570;
wire n4571;
wire n4572;
wire n4573;
wire n4574;
wire n4575;
wire n4576;
wire n4577;
wire n4578;
wire n4579;
wire n4580;
wire n4581;
wire n4582;
wire n4583;
wire n4584;
wire n4585;
wire n4586;
wire n4587;
wire n4588;
wire n4589;
wire n4590;
wire n4591;
wire n4592;
wire n4593;
wire n4594;
wire n4595;
wire n4596;
wire n4597;
wire n4598;
wire n4599;
wire n4600;
wire n4601;
wire n4602;
wire n4603;
wire n4604;
wire n4605;
wire n4606;
wire n4607;
wire n4608;
wire n4609;
wire n4610;
wire n4611;
wire n4612;
wire n4613;
wire n4614;
wire n4615;
wire n4616;
wire n4617;
wire n4618;
wire n4619;
wire n4620;
wire n4621;
wire n4622;
wire n4623;
wire n4624;
wire n4625;
wire n4626;
wire n4627;
wire n4628;
wire n4629;
wire n4630;
wire n4631;
wire n4632;
wire n4633;
wire n4634;
wire n4635;
wire n4636;
wire n4637;
wire n4638;
wire n4639;
wire n4640;
wire n4641;
wire n4642;
wire n4643;
wire n4644;
wire n4645;
wire n4646;
wire n4647;
wire n4648;
wire n4649;
wire n4650;
wire n4651;
wire n4652;
wire n4653;
wire n4654;
wire n4655;
wire n4656;
wire n4657;
wire n4658;
wire n4659;
wire n4660;
wire n4661;
wire n4662;
wire n4663;
wire n4664;
wire n4665;
wire n4666;
wire n4667;
wire n4668;
wire n4669;
wire n4670;
wire n4671;
wire n4672;
wire n4673;
wire n4674;
wire n4675;
wire n4676;
wire n4677;
wire n4678;
wire n4679;
wire n4680;
wire n4681;
wire n4682;
wire n4683;
wire n4684;
wire n4685;
wire n4686;
wire n4687;
wire n4688;
wire n4689;
wire n4690;
wire n4691;
wire n4692;
wire n4693;
wire n4694;
wire n4695;
wire n4696;
wire n4697;
wire n4698;
wire n4699;
wire n4700;
wire n4701;
wire n4702;
wire n4703;
wire n4704;
wire n4705;
wire n4706;
wire n4707;
wire n4708;
wire n4709;
wire n4710;
wire n4711;
wire n4712;
wire n4713;
wire n4714;
wire n4715;
wire n4716;
wire n4717;
wire n4718;
wire n4719;
wire n4720;
wire n4721;
wire n4722;
wire n4723;
wire n4724;
wire n4725;
wire n4726;
wire n4727;
wire n4728;
wire n4729;
wire n4730;
wire n4731;
wire n4732;
wire n4733;
wire n4734;
wire n4735;
wire n4736;
wire n4737;
wire n4738;
wire n4739;
wire n4740;
wire n4741;
wire n4742;
wire n4743;
wire n4744;
wire n4745;
wire n4746;
wire n4747;
wire n4748;
wire n4749;
wire n4750;
wire n4751;
wire n4752;
wire n4753;
wire n4754;
wire n4755;
wire n4756;
wire n4757;
wire n4758;
wire n4759;
wire n4760;
wire n4761;
wire n4762;
wire n4763;
wire n4764;
wire n4765;
wire n4766;
wire n4767;
wire n4768;
wire n4769;
wire n4770;
wire n4771;
wire n4772;
wire n4773;
wire n4774;
wire n4775;
wire n4776;
wire n4777;
wire n4778;
wire n4779;
wire n4780;
wire n4781;
wire n4782;
wire n4783;
wire n4784;
wire n4785;
wire n4786;
wire n4787;
wire n4788;
wire n4789;
wire n4790;
wire n4791;
wire n4792;
wire n4793;
wire n4794;
wire n4795;
wire n4796;
wire n4797;
wire n4798;
wire n4799;
wire n4800;
wire n4801;
wire n4802;
wire n4803;
wire n4804;
wire n4805;
wire n4806;
wire n4807;
wire n4808;
wire n4809;
wire n4810;
wire n4811;
wire n4812;
wire n4813;
wire n4814;
wire n4815;
wire n4816;
wire n4817;
wire n4818;
wire n4819;
wire n4820;
wire n4821;
wire n4822;
wire n4823;
wire n4824;
wire n4825;
wire n4826;
wire n4827;
wire n4828;
wire n4829;
wire n4830;
wire n4831;
wire n4832;
wire n4833;
wire n4834;
wire n4835;
wire n4836;
wire n4837;
wire n4838;
wire n4839;
wire n4840;
wire n4841;
wire n4842;
wire n4843;
wire n4844;
wire n4845;
wire n4846;
wire n4847;
wire n4848;
wire n4849;
wire n4850;
wire n4851;
wire n4852;
wire n4853;
wire n4854;
wire n4855;
wire n4856;
wire n4857;
wire n4858;
wire n4859;
wire n4860;
wire n4861;
wire n4862;
wire n4863;
wire n4864;
wire n4865;
wire n4866;
wire n4867;
wire n4868;
wire n4869;
wire n4870;
wire n4871;
wire n4872;
wire n4873;
wire n4874;
wire n4875;
wire n4876;
wire n4877;
wire n4878;
wire n4879;
wire n4880;
wire n4881;
wire n4882;
wire n4883;
wire n4884;
wire n4885;
wire n4886;
wire n4887;
wire n4888;
wire n4889;
wire n4890;
wire n4891;
wire n4892;
wire n4893;
wire n4894;
wire n4895;
wire n4896;
wire n4897;
wire n4898;
wire n4899;
wire n4900;
wire n4901;
wire n4902;
wire n4903;
wire n4904;
wire n4905;
wire n4906;
wire n4907;
wire n4908;
wire n4909;
wire n4910;
wire n4911;
wire n4912;
wire n4913;
wire n4914;
wire n4915;
wire n4916;
wire n4917;
wire n4918;
wire n4919;
wire n4920;
wire n4921;
wire n4922;
wire n4923;
wire n4924;
wire n4925;
wire n4926;
wire n4927;
wire n4928;
wire n4929;
wire n4930;
wire n4931;
wire n4932;
wire n4933;
wire n4934;
wire n4935;
wire n4936;
wire n4937;
wire n4938;
wire n4939;
wire n4940;
wire n4941;
wire n4942;
wire n4943;
wire n4944;
wire n4945;
wire n4946;
wire n4947;
wire n4948;
wire n4949;
wire n4950;
wire n4951;
wire n4952;
wire n4953;
wire n4954;
wire n4955;
wire n4956;
wire n4957;
wire n4958;
wire n4959;
wire n4960;
wire n4961;
wire n4962;
wire n4963;
wire n4964;
wire n4965;
wire n4966;
wire n4967;
wire n4968;
wire n4969;
wire n4970;
wire n4971;
wire n4972;
wire n4973;
wire n4974;
wire n4975;
wire n4976;
wire n4977;
wire n4978;
wire n4979;
wire n4980;
wire n4981;
wire n4982;
wire n4983;
wire n4984;
wire n4985;
wire n4986;
wire n4987;
wire n4988;
wire n4989;
wire n4990;
wire n4991;
wire n4992;
wire n4993;
wire n4994;
wire n4995;
wire n4996;
wire n4997;
wire n4998;
wire n4999;
wire n5000;
wire n5001;
wire n5002;
wire n5003;
wire n5004;
wire n5005;
wire n5006;
wire n5007;
wire n5008;
wire n5009;
wire n5010;
wire n5011;
wire n5012;
wire n5013;
wire n5014;
wire n5015;
wire n5016;
wire n5017;
wire n5018;
wire n5019;
wire n5020;
wire n5021;
wire n5022;
wire n5023;
wire n5024;
wire n5025;
wire n5026;
wire n5027;
wire n5028;
wire n5029;
wire n5030;
wire n5031;
wire n5032;
wire n5033;
wire n5034;
wire n5035;
wire n5036;
wire n5037;
wire n5038;
wire n5039;
wire n5040;
wire n5041;
wire n5042;
wire n5043;
wire n5044;
wire n5045;
wire n5046;
wire n5047;
wire n5048;
wire n5049;
wire n5050;
wire n5051;
wire n5052;
wire n5053;
wire n5054;
wire n5055;
wire n5056;
wire n5057;
wire n5058;
wire n5059;
wire n5060;
wire n5061;
wire n5062;
wire n5063;
wire n5064;
wire n5065;
wire n5066;
wire n5067;
wire n5068;
wire n5069;
wire n5070;
wire n5071;
wire n5072;
wire n5073;
wire n5074;
wire n5075;
wire n5076;
wire n5077;
wire n5078;
wire n5079;
wire n5080;
wire n5081;
wire n5082;
wire n5083;
wire n5084;
wire n5085;
wire n5086;
wire n5087;
wire n5088;
wire n5089;
wire n5090;
wire n5091;
wire n5092;
wire n5093;
wire n5094;
wire n5095;
wire n5096;
wire n5097;
wire n5098;
wire n5099;
wire n5100;
wire n5101;
wire n5102;
wire n5103;
wire n5104;
wire n5105;
wire n5106;
wire n5107;
wire n5108;
wire n5109;
wire n5110;
wire n5111;
wire n5112;
wire n5113;
wire n5114;
wire n5115;
wire n5116;
wire n5117;
wire n5118;
wire n5119;
wire n5120;
wire n5121;
wire n5122;
wire n5123;
wire n5124;
wire n5125;
wire n5126;
wire n5127;
wire n5128;
wire n5129;
wire n5130;
wire n5131;
wire n5132;
wire n5133;
wire n5134;
wire n5135;
wire n5136;
wire n5137;
wire n5138;
wire n5139;
wire n5140;
wire n5141;
wire n5142;
wire n5143;
wire n5144;
wire n5145;
wire n5146;
wire n5147;
wire n5148;
wire n5149;
wire n5150;
wire n5151;
wire n5152;
wire n5153;
wire n5154;
wire n5155;
wire n5156;
wire n5157;
wire n5158;
wire n5159;
wire n5160;
wire n5161;
wire n5162;
wire n5163;
wire n5164;
wire n5165;
wire n5166;
wire n5167;
wire n5168;
wire n5169;
wire n5170;
wire n5171;
wire n5172;
wire n5173;
wire n5174;
wire n5175;
wire n5176;
wire n5177;
wire n5178;
wire n5179;
wire n5180;
wire n5181;
wire n5182;
wire n5183;
wire n5184;
wire n5185;
wire n5186;
wire n5187;
wire n5188;
wire n5189;
wire n5190;
wire n5191;
wire n5192;
wire n5193;
wire n5194;
wire n5195;
wire n5196;
wire n5197;
wire n5198;
wire n5199;
wire n5200;
wire n5201;
wire n5202;
wire n5203;
wire n5204;
wire n5205;
wire n5206;
wire n5207;
wire n5208;
wire n5209;
wire n5210;
wire n5211;
wire n5212;
wire n5213;
wire n5214;
wire n5215;
wire n5216;
wire n5217;
wire n5218;
wire n5219;
wire n5220;
wire n5221;
wire n5222;
wire n5223;
wire n5224;
wire n5225;
wire n5226;
wire n5227;
wire n5228;
wire n5229;
wire n5230;
wire n5231;
wire n5232;
wire n5233;
wire n5234;
wire n5235;
wire n5236;
wire n5237;
wire n5238;
wire n5239;
wire n5240;
wire n5241;
wire n5242;
wire n5243;
wire n5244;
wire n5245;
wire n5246;
wire n5247;
wire n5248;
wire n5249;
wire n5250;
wire n5251;
wire n5252;
wire n5253;
wire n5254;
wire n5255;
wire n5256;
wire n5257;
wire n5258;
wire n5259;
wire n5260;
wire n5261;
wire n5262;
wire n5263;
wire n5264;
wire n5265;
wire n5266;
wire n5267;
wire n5268;
wire n5269;
wire n5270;
wire n5271;
wire n5272;
wire n5273;
wire n5274;
wire n5275;
wire n5276;
wire n5277;
wire n5278;
wire n5279;
wire n5280;
wire n5281;
wire n5282;
wire n5283;
wire n5284;
wire n5285;
wire n5286;
wire n5287;
wire n5288;
wire n5289;
wire n5290;
wire n5291;
wire n5292;
wire n5293;
wire n5294;
wire n5295;
wire n5296;
wire n5297;
wire n5298;
wire n5299;
wire n5300;
wire n5301;
wire n5302;
wire n5303;
wire n5304;
wire n5305;
wire n5306;
wire n5307;
wire n5308;
wire n5309;
wire n5310;
wire n5311;
wire n5312;
wire n5313;
wire n5314;
wire n5315;
wire n5316;
wire n5317;
wire n5318;
wire n5319;
wire n5320;
wire n5321;
wire n5322;
wire n5323;
wire n5324;
wire n5325;
wire n5326;
wire n5327;
wire n5328;
wire n5329;
wire n5330;
wire n5331;
wire n5332;
wire n5333;
wire n5334;
wire n5335;
wire n5336;
wire n5337;
wire n5338;
wire n5339;
wire n5340;
wire n5341;
wire n5342;
wire n5343;
wire n5344;
wire n5345;
wire n5346;
wire n5347;
wire n5348;
wire n5349;
wire n5350;
wire n5351;
wire n5352;
wire n5353;
wire n5354;
wire n5355;
wire n5356;
wire n5357;
wire n5358;
wire n5359;
wire n5360;
wire n5361;
wire n5362;
wire n5363;
wire n5364;
wire n5365;
wire n5366;
wire n5367;
wire n5368;
wire n5369;
wire n5370;
wire n5371;
wire n5372;
wire n5373;
wire n5374;
wire n5375;
wire n5376;
wire n5377;
wire n5378;
wire n5379;
wire n5380;
wire n5381;
wire n5382;
wire n5383;
wire n5384;
wire n5385;
wire n5386;
wire n5387;
wire n5388;
wire n5389;
wire n5390;
wire n5391;
wire n5392;
wire n5393;
wire n5394;
wire n5395;
wire n5396;
wire n5397;
wire n5398;
wire n5399;
wire n5400;
wire n5401;
wire n5402;
wire n5403;
wire n5404;
wire n5405;
wire n5406;
wire n5407;
wire n5408;
wire n5409;
wire n5410;
wire n5411;
wire n5412;
wire n5413;
wire n5414;
wire n5415;
wire n5416;
wire n5417;
wire n5418;
wire n5419;
wire n5420;
wire n5421;
wire n5422;
wire n5423;
wire n5424;
wire n5425;
wire n5426;
wire n5427;
wire n5428;
wire n5429;
wire n5430;
wire n5431;
wire n5432;
wire n5433;
wire n5434;
wire n5435;
wire n5436;
wire n5437;
wire n5438;
wire n5439;
wire n5440;
wire n5441;
wire n5442;
wire n5443;
wire n5444;
wire n5445;
wire n5446;
wire n5447;
wire n5448;
wire n5449;
wire n5450;
wire n5451;
wire n5452;
wire n5453;
wire n5454;
wire n5455;
wire n5456;
wire n5457;
wire n5458;
wire n5459;
wire n5460;
wire n5461;
wire n5462;
wire n5463;
wire n5464;
wire n5465;
wire n5466;
wire n5467;
wire n5468;
wire n5469;
wire n5470;
wire n5471;
wire n5472;
wire n5473;
wire n5474;
wire n5475;
wire n5476;
wire n5477;
wire n5478;
wire n5479;
wire n5480;
wire n5481;
wire n5482;
wire n5483;
wire n5484;
wire n5485;
wire n5486;
wire n5487;
wire n5488;
wire n5489;
wire n5490;
wire n5491;
wire n5492;
wire n5493;
wire n5494;
wire n5495;
wire n5496;
wire n5497;
wire n5498;
wire n5499;
wire n5500;
wire n5501;
wire n5502;
wire n5503;
wire n5504;
wire n5505;
wire n5506;
wire n5507;
xor (out,n0,n3085);
nand (n0,n1,n3084);
or (n1,n2,n1342);
not (n2,n3);
nor (n3,n4,n1341);
not (n4,n5);
nand (n5,n6,n1218);
not (n6,n7);
xor (n7,n8,n998);
xor (n8,n9,n824);
xor (n9,n10,n790);
xor (n10,n11,n516);
xor (n11,n12,n379);
xor (n12,n13,n258);
or (n13,n14,n257);
and (n14,n15,n219);
xor (n15,n16,n164);
nand (n16,n17,n152);
or (n17,n18,n97);
or (n18,n19,n90);
nor (n19,n20,n88);
and (n20,n21,n85);
not (n21,n22);
wire s0n22,s1n22,notn22;
or (n22,s0n22,s1n22);
not(notn22,n82);
and (s0n22,notn22,n23);
and (s1n22,n82,n42);
wire s0n23,s1n23,notn23;
or (n23,s0n23,s1n23);
not(notn23,n26);
and (s0n23,notn23,1'b0);
and (s1n23,n26,n25);
or (n26,n27,n38);
or (n27,n28,n36);
nor (n28,n29,n31,n32,n33,n35);
not (n29,n30);
not (n33,n34);
nor (n36,n30,n37,n32,n33,n35);
not (n37,n31);
or (n38,n39,n41);
and (n39,n29,n31,n32,n33,n40);
not (n40,n35);
nor (n41,n29,n37,n32,n33,n35);
xor (n42,n43,n44);
not (n43,n25);
and (n44,n45,n47);
not (n45,n46);
and (n47,n48,n50);
not (n48,n49);
and (n50,n51,n53);
not (n51,n52);
and (n53,n54,n56);
not (n54,n55);
and (n56,n57,n59);
not (n57,n58);
and (n59,n60,n62);
not (n60,n61);
and (n62,n63,n65);
not (n63,n64);
and (n65,n66,n68);
not (n66,n67);
and (n68,n69,n71);
not (n69,n70);
and (n71,n72,n74);
not (n72,n73);
and (n74,n75,n77);
not (n75,n76);
and (n77,n78,n80);
not (n78,n79);
not (n80,n81);
and (n82,n83,n84);
or (n83,n28,n39);
wire s0n85,s1n85,notn85;
or (n85,s0n85,s1n85);
not(notn85,n82);
and (s0n85,notn85,n86);
and (s1n85,n82,n87);
wire s0n86,s1n86,notn86;
or (n86,s0n86,s1n86);
not(notn86,n26);
and (s0n86,notn86,1'b0);
and (s1n86,n26,n46);
xor (n87,n45,n47);
and (n88,n89,n22);
not (n89,n85);
nor (n90,n91,n95);
and (n91,n85,n92);
wire s0n92,s1n92,notn92;
or (n92,s0n92,s1n92);
not(notn92,n82);
and (s0n92,notn92,n93);
and (s1n92,n82,n94);
wire s0n93,s1n93,notn93;
or (n93,s0n93,s1n93);
not(notn93,n26);
and (s0n93,notn93,1'b0);
and (s1n93,n26,n49);
xor (n94,n48,n50);
and (n95,n89,n96);
not (n96,n92);
nor (n97,n98,n150);
and (n98,n21,n99);
wire s0n99,s1n99,notn99;
or (n99,s0n99,s1n99);
not(notn99,n148);
and (s0n99,notn99,n100);
and (s1n99,n148,n102);
wire s0n100,s1n100,notn100;
or (n100,s0n100,s1n100);
not(notn100,n26);
and (s0n100,notn100,1'b0);
and (s1n100,n26,n101);
xor (n102,n103,n104);
not (n103,n101);
and (n104,n105,n107);
not (n105,n106);
and (n107,n108,n110);
not (n108,n109);
and (n110,n111,n113);
not (n111,n112);
and (n113,n114,n116);
not (n114,n115);
and (n116,n117,n119);
not (n117,n118);
and (n119,n120,n122);
not (n120,n121);
and (n122,n123,n125);
not (n123,n124);
and (n125,n126,n128);
not (n126,n127);
and (n128,n129,n131);
not (n129,n130);
and (n131,n132,n134);
not (n132,n133);
and (n134,n135,n137);
not (n135,n136);
and (n137,n138,n140);
not (n138,n139);
and (n140,n141,n143);
not (n141,n142);
and (n143,n144,n146);
not (n144,n145);
not (n146,n147);
and (n148,n83,n149);
and (n150,n22,n151);
not (n151,n99);
or (n152,n153,n154);
not (n153,n90);
nor (n154,n155,n162);
and (n155,n21,n156);
wire s0n156,s1n156,notn156;
or (n156,s0n156,s1n156);
not(notn156,n148);
and (s0n156,notn156,n157);
and (s1n156,n148,n159);
wire s0n157,s1n157,notn157;
or (n157,s0n157,s1n157);
not(notn157,n26);
and (s0n157,notn157,1'b0);
and (s1n157,n26,n158);
xor (n159,n160,n161);
not (n160,n158);
and (n161,n103,n104);
and (n162,n22,n163);
not (n163,n156);
nand (n164,n165,n210);
or (n165,n166,n203);
or (n166,n167,n193);
nor (n167,n168,n190);
and (n168,n169,n187);
wire s0n169,s1n169,notn169;
or (n169,s0n169,s1n169);
not(notn169,n82);
and (s0n169,notn169,n170);
and (s1n169,n82,n172);
wire s0n170,s1n170,notn170;
or (n170,s0n170,s1n170);
not(notn170,n26);
and (s0n170,notn170,1'b0);
and (s1n170,n26,n171);
xor (n172,n173,n174);
not (n173,n171);
and (n174,n175,n177);
not (n175,n176);
and (n177,n178,n180);
not (n178,n179);
and (n180,n181,n183);
not (n181,n182);
and (n183,n184,n186);
not (n184,n185);
and (n186,n43,n44);
wire s0n187,s1n187,notn187;
or (n187,s0n187,s1n187);
not(notn187,n82);
and (s0n187,notn187,n188);
and (s1n187,n82,n189);
wire s0n188,s1n188,notn188;
or (n188,s0n188,s1n188);
not(notn188,n26);
and (s0n188,notn188,1'b0);
and (s1n188,n26,n176);
xor (n189,n175,n177);
and (n190,n191,n192);
not (n191,n169);
not (n192,n187);
nor (n193,n194,n202);
and (n194,n169,n195);
not (n195,n196);
wire s0n196,s1n196,notn196;
or (n196,s0n196,s1n196);
not(notn196,n82);
and (s0n196,notn196,n197);
and (s1n196,n82,n199);
wire s0n197,s1n197,notn197;
or (n197,s0n197,s1n197);
not(notn197,n26);
and (s0n197,notn197,1'b0);
and (s1n197,n26,n198);
xor (n199,n200,n201);
not (n200,n198);
and (n201,n173,n174);
and (n202,n191,n196);
nor (n203,n204,n208);
and (n204,n195,n205);
wire s0n205,s1n205,notn205;
or (n205,s0n205,s1n205);
not(notn205,n148);
and (s0n205,notn205,n206);
and (s1n205,n148,n207);
wire s0n206,s1n206,notn206;
or (n206,s0n206,s1n206);
not(notn206,n26);
and (s0n206,notn206,1'b0);
and (s1n206,n26,n121);
xor (n207,n120,n122);
and (n208,n196,n209);
not (n209,n205);
or (n210,n211,n212);
not (n211,n167);
nor (n212,n213,n217);
and (n213,n195,n214);
wire s0n214,s1n214,notn214;
or (n214,s0n214,s1n214);
not(notn214,n148);
and (s0n214,notn214,n215);
and (s1n214,n148,n216);
wire s0n215,s1n215,notn215;
or (n215,s0n215,s1n215);
not(notn215,n26);
and (s0n215,notn215,1'b0);
and (s1n215,n26,n118);
xor (n216,n117,n119);
and (n217,n196,n218);
not (n218,n214);
nand (n219,n220,n249);
or (n220,n221,n242);
nand (n221,n222,n232);
nor (n222,n223,n230);
and (n223,n195,n224);
wire s0n224,s1n224,notn224;
or (n224,s0n224,s1n224);
not(notn224,n82);
and (s0n224,notn224,n225);
and (s1n224,n82,n227);
wire s0n225,s1n225,notn225;
or (n225,s0n225,s1n225);
not(notn225,n26);
and (s0n225,notn225,1'b0);
and (s1n225,n26,n226);
xor (n227,n228,n229);
not (n228,n226);
and (n229,n200,n201);
and (n230,n196,n231);
not (n231,n224);
nand (n232,n233,n240);
or (n233,n231,n234);
wire s0n234,s1n234,notn234;
or (n234,s0n234,s1n234);
not(notn234,n82);
and (s0n234,notn234,n235);
and (s1n234,n82,n237);
wire s0n235,s1n235,notn235;
or (n235,s0n235,s1n235);
not(notn235,n26);
and (s0n235,notn235,1'b0);
and (s1n235,n26,n236);
xor (n237,n238,n239);
not (n238,n236);
and (n239,n228,n229);
or (n240,n224,n241);
not (n241,n234);
nor (n242,n243,n247);
and (n243,n241,n244);
wire s0n244,s1n244,notn244;
or (n244,s0n244,s1n244);
not(notn244,n148);
and (s0n244,notn244,n245);
and (s1n244,n148,n246);
wire s0n245,s1n245,notn245;
or (n245,s0n245,s1n245);
not(notn245,n26);
and (s0n245,notn245,1'b0);
and (s1n245,n26,n127);
xor (n246,n126,n128);
and (n247,n248,n234);
not (n248,n244);
or (n249,n222,n250);
nor (n250,n251,n255);
and (n251,n241,n252);
wire s0n252,s1n252,notn252;
or (n252,s0n252,s1n252);
not(notn252,n148);
and (s0n252,notn252,n253);
and (s1n252,n148,n254);
wire s0n253,s1n253,notn253;
or (n253,s0n253,s1n253);
not(notn253,n26);
and (s0n253,notn253,1'b0);
and (s1n253,n26,n124);
xor (n254,n123,n125);
and (n255,n256,n234);
not (n256,n252);
and (n257,n16,n164);
or (n258,n259,n378);
and (n259,n260,n340);
xor (n260,n261,n300);
nand (n261,n262,n292);
or (n262,n263,n285);
or (n263,n264,n275);
not (n264,n265);
and (n265,n266,n274);
nand (n266,n267,n234);
not (n267,n268);
wire s0n268,s1n268,notn268;
or (n268,s0n268,s1n268);
not(notn268,n82);
and (s0n268,notn268,n269);
and (s1n268,n82,n271);
wire s0n269,s1n269,notn269;
or (n269,s0n269,s1n269);
not(notn269,n26);
and (s0n269,notn269,1'b0);
and (s1n269,n26,n270);
xor (n271,n272,n273);
not (n272,n270);
and (n273,n238,n239);
nand (n274,n268,n241);
nor (n275,n276,n284);
and (n276,n268,n277);
not (n277,n278);
wire s0n278,s1n278,notn278;
or (n278,s0n278,s1n278);
not(notn278,n82);
and (s0n278,notn278,n279);
and (s1n278,n82,n281);
wire s0n279,s1n279,notn279;
or (n279,s0n279,s1n279);
not(notn279,n26);
and (s0n279,notn279,1'b0);
and (s1n279,n26,n280);
xor (n281,n282,n283);
not (n282,n280);
and (n283,n272,n273);
and (n284,n267,n278);
nor (n285,n286,n290);
and (n286,n277,n287);
wire s0n287,s1n287,notn287;
or (n287,s0n287,s1n287);
not(notn287,n148);
and (s0n287,notn287,n288);
and (s1n287,n148,n289);
wire s0n288,s1n288,notn288;
or (n288,s0n288,s1n288);
not(notn288,n26);
and (s0n288,notn288,1'b0);
and (s1n288,n26,n133);
xor (n289,n132,n134);
and (n290,n291,n278);
not (n291,n287);
or (n292,n265,n293);
nor (n293,n294,n298);
and (n294,n277,n295);
wire s0n295,s1n295,notn295;
or (n295,s0n295,s1n295);
not(notn295,n148);
and (s0n295,notn295,n296);
and (s1n295,n148,n297);
wire s0n296,s1n296,notn296;
or (n296,s0n296,s1n296);
not(notn296,n26);
and (s0n296,notn296,1'b0);
and (s1n296,n26,n130);
xor (n297,n129,n131);
and (n298,n299,n278);
not (n299,n295);
nand (n300,n301,n332);
or (n301,n302,n325);
nand (n302,n303,n322);
or (n303,n304,n319);
not (n304,n305);
nand (n305,n306,n312);
wire s0n306,s1n306,notn306;
or (n306,s0n306,s1n306);
not(notn306,n82);
and (s0n306,notn306,n307);
and (s1n306,n82,n309);
wire s0n307,s1n307,notn307;
or (n307,s0n307,s1n307);
not(notn307,n26);
and (s0n307,notn307,1'b0);
and (s1n307,n26,n308);
xor (n309,n310,n311);
not (n310,n308);
and (n311,n282,n283);
not (n312,n313);
wire s0n313,s1n313,notn313;
or (n313,s0n313,s1n313);
not(notn313,n82);
and (s0n313,notn313,n314);
and (s1n313,n82,n316);
wire s0n314,s1n314,notn314;
or (n314,s0n314,s1n314);
not(notn314,n26);
and (s0n314,notn314,1'b0);
and (s1n314,n26,n315);
xor (n316,n317,n318);
not (n317,n315);
and (n318,n310,n311);
not (n319,n320);
nand (n320,n321,n313);
not (n321,n306);
and (n322,n323,n324);
nand (n323,n321,n278);
nand (n324,n306,n277);
nor (n325,n326,n330);
and (n326,n327,n312);
wire s0n327,s1n327,notn327;
or (n327,s0n327,s1n327);
not(notn327,n148);
and (s0n327,notn327,n328);
and (s1n327,n148,n329);
wire s0n328,s1n328,notn328;
or (n328,s0n328,s1n328);
not(notn328,n26);
and (s0n328,notn328,1'b0);
and (s1n328,n26,n139);
xor (n329,n138,n140);
and (n330,n331,n313);
not (n331,n327);
or (n332,n322,n333);
nor (n333,n334,n338);
and (n334,n312,n335);
wire s0n335,s1n335,notn335;
or (n335,s0n335,s1n335);
not(notn335,n148);
and (s0n335,notn335,n336);
and (s1n335,n148,n337);
wire s0n336,s1n336,notn336;
or (n336,s0n336,s1n336);
not(notn336,n26);
and (s0n336,notn336,1'b0);
and (s1n336,n26,n136);
xor (n337,n135,n137);
and (n338,n339,n313);
not (n339,n335);
nand (n340,n341,n370);
or (n341,n342,n363);
nand (n342,n343,n353);
nor (n343,n344,n351);
and (n344,n312,n345);
wire s0n345,s1n345,notn345;
or (n345,s0n345,s1n345);
not(notn345,n82);
and (s0n345,notn345,n346);
and (s1n345,n82,n348);
wire s0n346,s1n346,notn346;
or (n346,s0n346,s1n346);
not(notn346,n26);
and (s0n346,notn346,1'b0);
and (s1n346,n26,n347);
xor (n348,n349,n350);
not (n349,n347);
and (n350,n317,n318);
and (n351,n313,n352);
not (n352,n345);
nand (n353,n354,n361);
or (n354,n352,n355);
wire s0n355,s1n355,notn355;
or (n355,s0n355,s1n355);
not(notn355,n82);
and (s0n355,notn355,n356);
and (s1n355,n82,n358);
wire s0n356,s1n356,notn356;
or (n356,s0n356,s1n356);
not(notn356,n26);
and (s0n356,notn356,1'b0);
and (s1n356,n26,n357);
xor (n358,n359,n360);
not (n359,n357);
and (n360,n349,n350);
or (n361,n345,n362);
not (n362,n355);
nor (n363,n364,n368);
and (n364,n362,n365);
wire s0n365,s1n365,notn365;
or (n365,s0n365,s1n365);
not(notn365,n148);
and (s0n365,notn365,n366);
and (s1n365,n148,n367);
wire s0n366,s1n366,notn366;
or (n366,s0n366,s1n366);
not(notn366,n26);
and (s0n366,notn366,1'b0);
and (s1n366,n26,n145);
xor (n367,n144,n146);
and (n368,n369,n355);
not (n369,n365);
or (n370,n343,n371);
nor (n371,n372,n376);
and (n372,n373,n362);
wire s0n373,s1n373,notn373;
or (n373,s0n373,s1n373);
not(notn373,n148);
and (s0n373,notn373,n374);
and (s1n373,n148,n375);
wire s0n374,s1n374,notn374;
or (n374,s0n374,s1n374);
not(notn374,n26);
and (s0n374,notn374,1'b0);
and (s1n374,n26,n142);
xor (n375,n141,n143);
and (n376,n377,n355);
not (n377,n373);
and (n378,n261,n300);
xor (n379,n380,n486);
xor (n380,n381,n450);
nand (n381,n382,n439);
or (n382,n383,n402);
nand (n383,n384,n395);
nor (n384,n385,n393);
and (n385,n386,n390);
not (n386,n387);
wire s0n387,s1n387,notn387;
or (n387,s0n387,s1n387);
not(notn387,n82);
and (s0n387,notn387,n388);
and (s1n387,n82,n389);
wire s0n388,s1n388,notn388;
or (n388,s0n388,s1n388);
not(notn388,n26);
and (s0n388,notn388,1'b0);
and (s1n388,n26,n79);
xor (n389,n78,n80);
wire s0n390,s1n390,notn390;
or (n390,s0n390,s1n390);
not(notn390,n82);
and (s0n390,notn390,n391);
and (s1n390,n82,n392);
wire s0n391,s1n391,notn391;
or (n391,s0n391,s1n391);
not(notn391,n26);
and (s0n391,notn391,1'b0);
and (s1n391,n26,n76);
xor (n392,n75,n77);
and (n393,n387,n394);
not (n394,n390);
nand (n395,n396,n401);
or (n396,n397,n390);
not (n397,n398);
wire s0n398,s1n398,notn398;
or (n398,s0n398,s1n398);
not(notn398,n82);
and (s0n398,notn398,n399);
and (s1n398,n82,n400);
wire s0n399,s1n399,notn399;
or (n399,s0n399,s1n399);
not(notn399,n26);
and (s0n399,notn399,1'b0);
and (s1n399,n26,n73);
xor (n400,n72,n74);
nand (n401,n397,n390);
nor (n402,n403,n437);
and (n403,n404,n397);
wire s0n404,s1n404,notn404;
or (n404,s0n404,s1n404);
not(notn404,n148);
and (s0n404,notn404,n405);
and (s1n404,n148,n407);
wire s0n405,s1n405,notn405;
or (n405,s0n405,s1n405);
not(notn405,n26);
and (s0n405,notn405,1'b0);
and (s1n405,n26,n406);
xor (n407,n408,n409);
not (n408,n406);
and (n409,n410,n412);
not (n410,n411);
and (n412,n413,n415);
not (n413,n414);
and (n415,n416,n418);
not (n416,n417);
and (n418,n419,n421);
not (n419,n420);
and (n421,n422,n424);
not (n422,n423);
and (n424,n425,n427);
not (n425,n426);
and (n427,n428,n430);
not (n428,n429);
and (n430,n431,n433);
not (n431,n432);
and (n433,n434,n436);
not (n434,n435);
and (n436,n160,n161);
and (n437,n438,n398);
not (n438,n404);
or (n439,n440,n384);
nor (n440,n441,n448);
and (n441,n442,n397);
wire s0n442,s1n442,notn442;
or (n442,s0n442,s1n442);
not(notn442,n148);
and (s0n442,notn442,n443);
and (s1n442,n148,n445);
wire s0n443,s1n443,notn443;
or (n443,s0n443,s1n443);
not(notn443,n26);
and (s0n443,notn443,1'b0);
and (s1n443,n26,n444);
xor (n445,n446,n447);
not (n446,n444);
and (n447,n408,n409);
and (n448,n449,n398);
not (n449,n442);
nand (n450,n451,n478);
or (n451,n452,n471);
nand (n452,n453,n464);
or (n453,n454,n461);
and (n454,n455,n458);
wire s0n455,s1n455,notn455;
or (n455,s0n455,s1n455);
not(notn455,n82);
and (s0n455,notn455,n456);
and (s1n455,n82,n457);
wire s0n456,s1n456,notn456;
or (n456,s0n456,s1n456);
not(notn456,n26);
and (s0n456,notn456,1'b0);
and (s1n456,n26,n67);
xor (n457,n66,n68);
wire s0n458,s1n458,notn458;
or (n458,s0n458,s1n458);
not(notn458,n82);
and (s0n458,notn458,n459);
and (s1n458,n82,n460);
wire s0n459,s1n459,notn459;
or (n459,s0n459,s1n459);
not(notn459,n26);
and (s0n459,notn459,1'b0);
and (s1n459,n26,n64);
xor (n460,n63,n65);
and (n461,n462,n463);
not (n462,n455);
not (n463,n458);
nor (n464,n465,n469);
and (n465,n466,n458);
wire s0n466,s1n466,notn466;
or (n466,s0n466,s1n466);
not(notn466,n82);
and (s0n466,notn466,n467);
and (s1n466,n82,n468);
wire s0n467,s1n467,notn467;
or (n467,s0n467,s1n467);
not(notn467,n26);
and (s0n467,notn467,1'b0);
and (s1n467,n26,n61);
xor (n468,n60,n62);
and (n469,n470,n463);
not (n470,n466);
nor (n471,n472,n476);
and (n472,n473,n470);
wire s0n473,s1n473,notn473;
or (n473,s0n473,s1n473);
not(notn473,n148);
and (s0n473,notn473,n474);
and (s1n473,n148,n475);
wire s0n474,s1n474,notn474;
or (n474,s0n474,s1n474);
not(notn474,n26);
and (s0n474,notn474,1'b0);
and (s1n474,n26,n420);
xor (n475,n419,n421);
and (n476,n477,n466);
not (n477,n473);
or (n478,n479,n453);
nor (n479,n480,n484);
and (n480,n481,n470);
wire s0n481,s1n481,notn481;
or (n481,s0n481,s1n481);
not(notn481,n148);
and (s0n481,notn481,n482);
and (s1n481,n148,n483);
wire s0n482,s1n482,notn482;
or (n482,s0n482,s1n482);
not(notn482,n26);
and (s0n482,notn482,1'b0);
and (s1n482,n26,n417);
xor (n483,n416,n418);
and (n484,n485,n466);
not (n485,n481);
nand (n486,n487,n511);
or (n487,n488,n504);
not (n488,n489);
nor (n489,n490,n496);
nand (n490,n491,n495);
or (n491,n21,n492);
wire s0n492,s1n492,notn492;
or (n492,s0n492,s1n492);
not(notn492,n82);
and (s0n492,notn492,n493);
and (s1n492,n82,n494);
wire s0n493,s1n493,notn493;
or (n493,s0n493,s1n493);
not(notn493,n26);
and (s0n493,notn493,1'b0);
and (s1n493,n26,n185);
xor (n494,n184,n186);
nand (n495,n21,n492);
nor (n496,n497,n502);
and (n497,n498,n492);
not (n498,n499);
wire s0n499,s1n499,notn499;
or (n499,s0n499,s1n499);
not(notn499,n82);
and (s0n499,notn499,n500);
and (s1n499,n82,n501);
wire s0n500,s1n500,notn500;
or (n500,s0n500,s1n500);
not(notn500,n26);
and (s0n500,notn500,1'b0);
and (s1n500,n26,n182);
xor (n501,n181,n183);
and (n502,n503,n499);
not (n503,n492);
nor (n504,n505,n509);
and (n505,n498,n506);
wire s0n506,s1n506,notn506;
or (n506,s0n506,s1n506);
not(notn506,n148);
and (s0n506,notn506,n507);
and (s1n506,n148,n508);
wire s0n507,s1n507,notn507;
or (n507,s0n507,s1n507);
not(notn507,n26);
and (s0n507,notn507,1'b0);
and (s1n507,n26,n106);
xor (n508,n105,n107);
and (n509,n499,n510);
not (n510,n506);
or (n511,n512,n513);
not (n512,n490);
nor (n513,n514,n515);
and (n514,n498,n99);
and (n515,n499,n151);
xor (n516,n517,n704);
xor (n517,n518,n538);
xor (n518,n519,n532);
xor (n519,n520,n526);
nand (n520,n521,n522);
or (n521,n221,n250);
or (n522,n222,n523);
nor (n523,n524,n525);
and (n524,n241,n205);
and (n525,n234,n209);
nand (n526,n527,n528);
or (n527,n263,n293);
or (n528,n265,n529);
nor (n529,n530,n531);
and (n530,n244,n277);
and (n531,n248,n278);
nand (n532,n533,n534);
or (n533,n302,n333);
or (n534,n322,n535);
nor (n535,n536,n537);
and (n536,n287,n312);
and (n537,n291,n313);
or (n538,n539,n703);
and (n539,n540,n630);
xor (n540,n541,n567);
and (n541,n542,n550);
nor (n542,n543,n362);
nor (n543,n544,n548);
and (n544,n312,n545);
not (n545,n546);
and (n546,n547,n345);
wire s0n547,s1n547,notn547;
or (n547,s0n547,s1n547);
not(notn547,n26);
and (s0n547,notn547,1'b0);
and (s1n547,n26,n147);
and (n548,n352,n549);
not (n549,n547);
nand (n550,n551,n559);
or (n551,n383,n552);
nor (n552,n553,n557);
and (n553,n554,n397);
wire s0n554,s1n554,notn554;
or (n554,s0n554,s1n554);
not(notn554,n148);
and (s0n554,notn554,n555);
and (s1n554,n148,n556);
wire s0n555,s1n555,notn555;
or (n555,s0n555,s1n555);
not(notn555,n26);
and (s0n555,notn555,1'b0);
and (s1n555,n26,n414);
xor (n556,n413,n415);
and (n557,n558,n398);
not (n558,n554);
or (n559,n560,n384);
nor (n560,n561,n565);
and (n561,n562,n397);
wire s0n562,s1n562,notn562;
or (n562,s0n562,s1n562);
not(notn562,n148);
and (s0n562,notn562,n563);
and (s1n562,n148,n564);
wire s0n563,s1n563,notn563;
or (n563,s0n563,s1n563);
not(notn563,n26);
and (s0n563,notn563,1'b0);
and (s1n563,n26,n411);
xor (n564,n410,n412);
and (n565,n566,n398);
not (n566,n562);
or (n567,n568,n629);
and (n568,n569,n604);
xor (n569,n570,n587);
nand (n570,n571,n579);
or (n571,n452,n572);
nor (n572,n573,n577);
and (n573,n574,n470);
wire s0n574,s1n574,notn574;
or (n574,s0n574,s1n574);
not(notn574,n148);
and (s0n574,notn574,n575);
and (s1n574,n148,n576);
wire s0n575,s1n575,notn575;
or (n575,s0n575,s1n575);
not(notn575,n26);
and (s0n575,notn575,1'b0);
and (s1n575,n26,n426);
xor (n576,n425,n427);
and (n577,n578,n466);
not (n578,n574);
or (n579,n580,n453);
nor (n580,n581,n585);
and (n581,n582,n470);
wire s0n582,s1n582,notn582;
or (n582,s0n582,s1n582);
not(notn582,n148);
and (s0n582,notn582,n583);
and (s1n582,n148,n584);
wire s0n583,s1n583,notn583;
or (n583,s0n583,s1n583);
not(notn583,n26);
and (s0n583,notn583,1'b0);
and (s1n583,n26,n423);
xor (n584,n422,n424);
and (n585,n586,n466);
not (n586,n582);
nand (n587,n588,n596);
or (n588,n488,n589);
nor (n589,n590,n594);
and (n590,n498,n591);
wire s0n591,s1n591,notn591;
or (n591,s0n591,s1n591);
not(notn591,n148);
and (s0n591,notn591,n592);
and (s1n591,n148,n593);
wire s0n592,s1n592,notn592;
or (n592,s0n592,s1n592);
not(notn592,n26);
and (s0n592,notn592,1'b0);
and (s1n592,n26,n112);
xor (n593,n111,n113);
and (n594,n499,n595);
not (n595,n591);
or (n596,n512,n597);
nor (n597,n598,n602);
and (n598,n498,n599);
wire s0n599,s1n599,notn599;
or (n599,s0n599,s1n599);
not(notn599,n148);
and (s0n599,notn599,n600);
and (s1n599,n148,n601);
wire s0n600,s1n600,notn600;
or (n600,s0n600,s1n600);
not(notn600,n26);
and (s0n600,notn600,1'b0);
and (s1n600,n26,n109);
xor (n601,n108,n110);
and (n602,n499,n603);
not (n603,n599);
nand (n604,n605,n621);
or (n605,n606,n618);
not (n606,n607);
and (n607,n608,n615);
nor (n608,n609,n614);
and (n609,n499,n610);
not (n610,n611);
wire s0n611,s1n611,notn611;
or (n611,s0n611,s1n611);
not(notn611,n82);
and (s0n611,notn611,n612);
and (s1n611,n82,n613);
wire s0n612,s1n612,notn612;
or (n612,s0n612,s1n612);
not(notn612,n26);
and (s0n612,notn612,1'b0);
and (s1n612,n26,n179);
xor (n613,n178,n180);
and (n614,n498,n611);
nand (n615,n616,n617);
or (n616,n610,n187);
or (n617,n192,n611);
nor (n618,n619,n620);
and (n619,n192,n214);
and (n620,n187,n218);
or (n621,n608,n622);
nor (n622,n623,n627);
and (n623,n192,n624);
wire s0n624,s1n624,notn624;
or (n624,s0n624,s1n624);
not(notn624,n148);
and (s0n624,notn624,n625);
and (s1n624,n148,n626);
wire s0n625,s1n625,notn625;
or (n625,s0n625,s1n625);
not(notn625,n26);
and (s0n625,notn625,1'b0);
and (s1n625,n26,n115);
xor (n626,n114,n116);
and (n627,n187,n628);
not (n628,n624);
and (n629,n570,n587);
or (n630,n631,n702);
and (n631,n632,n678);
xor (n632,n633,n666);
nand (n633,n634,n658);
or (n634,n635,n651);
nand (n635,n636,n647);
nor (n636,n637,n644);
and (n637,n638,n641);
wire s0n638,s1n638,notn638;
or (n638,s0n638,s1n638);
not(notn638,n82);
and (s0n638,notn638,n639);
and (s1n638,n82,n640);
wire s0n639,s1n639,notn639;
or (n639,s0n639,s1n639);
not(notn639,n26);
and (s0n639,notn639,1'b0);
and (s1n639,n26,n58);
xor (n640,n57,n59);
wire s0n641,s1n641,notn641;
or (n641,s0n641,s1n641);
not(notn641,n82);
and (s0n641,notn641,n642);
and (s1n641,n82,n643);
wire s0n642,s1n642,notn642;
or (n642,s0n642,s1n642);
not(notn642,n26);
and (s0n642,notn642,1'b0);
and (s1n642,n26,n55);
xor (n643,n54,n56);
and (n644,n645,n646);
not (n645,n638);
not (n646,n641);
not (n647,n648);
nor (n648,n649,n650);
and (n649,n466,n638);
and (n650,n470,n645);
nor (n651,n652,n656);
and (n652,n653,n646);
wire s0n653,s1n653,notn653;
or (n653,s0n653,s1n653);
not(notn653,n148);
and (s0n653,notn653,n654);
and (s1n653,n148,n655);
wire s0n654,s1n654,notn654;
or (n654,s0n654,s1n654);
not(notn654,n26);
and (s0n654,notn654,1'b0);
and (s1n654,n26,n432);
xor (n655,n431,n433);
and (n656,n657,n641);
not (n657,n653);
or (n658,n659,n647);
nor (n659,n660,n664);
and (n660,n661,n646);
wire s0n661,s1n661,notn661;
or (n661,s0n661,s1n661);
not(notn661,n148);
and (s0n661,notn661,n662);
and (s1n661,n148,n663);
wire s0n662,s1n662,notn662;
or (n662,s0n662,s1n662);
not(notn662,n26);
and (s0n662,notn662,1'b0);
and (s1n662,n26,n429);
xor (n663,n428,n430);
and (n664,n665,n641);
not (n665,n661);
nand (n666,n667,n674);
or (n667,n668,n671);
nor (n668,n669,n670);
and (n669,n404,n386);
and (n670,n438,n387);
nand (n671,n387,n672);
not (n672,n673);
wire s0n673,s1n673,notn673;
or (n673,s0n673,s1n673);
not(notn673,n26);
and (s0n673,notn673,1'b0);
and (s1n673,n26,n81);
or (n674,n675,n672);
nor (n675,n676,n677);
and (n676,n442,n386);
and (n677,n449,n387);
nand (n678,n679,n694);
or (n679,n680,n691);
nand (n680,n681,n688);
or (n681,n682,n686);
and (n682,n683,n641);
wire s0n683,s1n683,notn683;
or (n683,s0n683,s1n683);
not(notn683,n82);
and (s0n683,notn683,n684);
and (s1n683,n82,n685);
wire s0n684,s1n684,notn684;
or (n684,s0n684,s1n684);
not(notn684,n26);
and (s0n684,notn684,1'b0);
and (s1n684,n26,n52);
xor (n685,n51,n53);
and (n686,n687,n646);
not (n687,n683);
nand (n688,n689,n690);
or (n689,n687,n92);
or (n690,n96,n683);
nor (n691,n692,n693);
and (n692,n96,n156);
and (n693,n92,n163);
or (n694,n681,n695);
nor (n695,n696,n700);
and (n696,n697,n96);
wire s0n697,s1n697,notn697;
or (n697,s0n697,s1n697);
not(notn697,n148);
and (s0n697,notn697,n698);
and (s1n697,n148,n699);
wire s0n698,s1n698,notn698;
or (n698,s0n698,s1n698);
not(notn698,n26);
and (s0n698,notn698,1'b0);
and (s1n698,n26,n435);
xor (n699,n434,n436);
and (n700,n701,n92);
not (n701,n697);
and (n702,n633,n666);
and (n703,n541,n567);
xor (n704,n705,n771);
xor (n705,n706,n750);
or (n706,n707,n749);
and (n707,n708,n728);
xor (n708,n709,n722);
nand (n709,n710,n711);
or (n710,n675,n671);
or (n711,n712,n672);
nor (n712,n713,n720);
and (n713,n714,n386);
wire s0n714,s1n714,notn714;
or (n714,s0n714,s1n714);
not(notn714,n148);
and (s0n714,notn714,n715);
and (s1n714,n148,n717);
wire s0n715,s1n715,notn715;
or (n715,s0n715,s1n715);
not(notn715,n26);
and (s0n715,notn715,1'b0);
and (s1n715,n26,n716);
xor (n717,n718,n719);
not (n718,n716);
and (n719,n446,n447);
and (n720,n721,n387);
not (n721,n714);
nand (n722,n723,n724);
or (n723,n680,n695);
or (n724,n681,n725);
nor (n725,n726,n727);
and (n726,n96,n653);
and (n727,n657,n92);
nand (n728,n729,n745);
or (n729,n730,n742);
nand (n730,n731,n738);
not (n731,n732);
nand (n732,n733,n737);
or (n733,n397,n734);
wire s0n734,s1n734,notn734;
or (n734,s0n734,s1n734);
not(notn734,n82);
and (s0n734,notn734,n735);
and (s1n734,n82,n736);
wire s0n735,s1n735,notn735;
or (n735,s0n735,s1n735);
not(notn735,n26);
and (s0n735,notn735,1'b0);
and (s1n735,n26,n70);
xor (n736,n69,n71);
nand (n737,n734,n397);
nor (n738,n739,n741);
and (n739,n462,n740);
not (n740,n734);
and (n741,n455,n734);
nor (n742,n743,n744);
and (n743,n481,n462);
and (n744,n485,n455);
or (n745,n746,n731);
nor (n746,n747,n748);
and (n747,n554,n462);
and (n748,n558,n455);
and (n749,n709,n722);
or (n750,n751,n770);
and (n751,n752,n767);
xor (n752,n753,n764);
nor (n753,n754,n549);
nor (n754,n755,n762);
and (n755,n362,n756);
wire s0n756,s1n756,notn756;
or (n756,s0n756,s1n756);
not(notn756,n82);
and (s0n756,notn756,n757);
and (s1n756,n82,n759);
wire s0n757,s1n757,notn757;
or (n757,s0n757,s1n757);
not(notn757,n26);
and (s0n757,notn757,1'b0);
and (s1n757,n26,n758);
xor (n759,n760,n761);
not (n760,n758);
and (n761,n359,n360);
and (n762,n355,n763);
not (n763,n756);
nand (n764,n765,n766);
or (n765,n383,n560);
or (n766,n402,n384);
nand (n767,n768,n769);
or (n768,n452,n580);
or (n769,n471,n453);
and (n770,n753,n764);
or (n771,n772,n789);
and (n772,n773,n783);
xor (n773,n774,n777);
nand (n774,n775,n776);
or (n775,n488,n597);
or (n776,n512,n504);
nand (n777,n778,n779);
or (n778,n606,n622);
or (n779,n608,n780);
nor (n780,n781,n782);
and (n781,n192,n591);
and (n782,n187,n595);
nand (n783,n784,n785);
or (n784,n635,n659);
or (n785,n786,n647);
nor (n786,n787,n788);
and (n787,n646,n574);
and (n788,n578,n641);
and (n789,n774,n777);
or (n790,n791,n823);
and (n791,n792,n822);
xor (n792,n793,n794);
xor (n793,n15,n219);
or (n794,n795,n821);
and (n795,n796,n804);
xor (n796,n797,n803);
nand (n797,n798,n802);
or (n798,n342,n799);
nor (n799,n800,n801);
and (n800,n355,n549);
and (n801,n362,n547);
or (n802,n343,n363);
xor (n803,n542,n550);
or (n804,n805,n820);
and (n805,n806,n814);
xor (n806,n807,n808);
nor (n807,n343,n549);
nand (n808,n809,n813);
or (n809,n383,n810);
nor (n810,n811,n812);
and (n811,n481,n397);
and (n812,n485,n398);
or (n813,n552,n384);
nand (n814,n815,n819);
or (n815,n452,n816);
nor (n816,n817,n818);
and (n817,n661,n470);
and (n818,n665,n466);
or (n819,n572,n453);
and (n820,n807,n808);
and (n821,n797,n803);
xor (n822,n540,n630);
and (n823,n793,n794);
or (n824,n825,n997);
and (n825,n826,n936);
xor (n826,n827,n828);
xor (n827,n792,n822);
xor (n828,n829,n929);
xor (n829,n830,n882);
or (n830,n831,n881);
and (n831,n832,n880);
xor (n832,n833,n855);
or (n833,n834,n854);
and (n834,n835,n848);
xor (n835,n836,n842);
nand (n836,n837,n841);
or (n837,n488,n838);
nor (n838,n839,n840);
and (n839,n498,n624);
and (n840,n499,n628);
or (n841,n512,n589);
nand (n842,n843,n847);
or (n843,n606,n844);
nor (n844,n845,n846);
and (n845,n192,n205);
and (n846,n187,n209);
or (n847,n608,n618);
nand (n848,n849,n853);
or (n849,n635,n850);
nor (n850,n851,n852);
and (n851,n697,n646);
and (n852,n701,n641);
or (n853,n651,n647);
and (n854,n836,n842);
or (n855,n856,n879);
and (n856,n857,n870);
xor (n857,n858,n864);
nand (n858,n859,n863);
or (n859,n860,n671);
nor (n860,n861,n862);
and (n861,n562,n386);
and (n862,n566,n387);
or (n863,n668,n672);
nand (n864,n865,n869);
or (n865,n680,n866);
nor (n866,n867,n868);
and (n867,n96,n99);
and (n868,n92,n151);
or (n869,n681,n691);
nand (n870,n871,n875);
or (n871,n730,n872);
nor (n872,n873,n874);
and (n873,n582,n462);
and (n874,n586,n455);
or (n875,n876,n731);
nor (n876,n877,n878);
and (n877,n473,n462);
and (n878,n477,n455);
and (n879,n858,n864);
xor (n880,n632,n678);
and (n881,n833,n855);
or (n882,n883,n928);
and (n883,n884,n903);
xor (n884,n885,n902);
xor (n885,n886,n896);
xor (n886,n887,n890);
nand (n887,n888,n889);
or (n888,n730,n876);
or (n889,n742,n731);
nand (n890,n891,n895);
or (n891,n18,n892);
nor (n892,n893,n894);
and (n893,n21,n506);
and (n894,n22,n510);
or (n895,n153,n97);
nand (n896,n897,n901);
or (n897,n166,n898);
nor (n898,n899,n900);
and (n899,n195,n252);
and (n900,n196,n256);
or (n901,n211,n203);
xor (n902,n569,n604);
or (n903,n904,n927);
and (n904,n905,n918);
xor (n905,n906,n912);
nand (n906,n907,n911);
or (n907,n18,n908);
nor (n908,n909,n910);
and (n909,n21,n599);
and (n910,n22,n603);
or (n911,n153,n892);
nand (n912,n913,n917);
or (n913,n166,n914);
nor (n914,n915,n916);
and (n915,n195,n244);
and (n916,n196,n248);
or (n917,n211,n898);
nand (n918,n919,n923);
or (n919,n221,n920);
nor (n920,n921,n922);
and (n921,n241,n287);
and (n922,n291,n234);
or (n923,n222,n924);
nor (n924,n925,n926);
and (n925,n241,n295);
and (n926,n299,n234);
and (n927,n906,n912);
and (n928,n885,n902);
xor (n929,n930,n935);
xor (n930,n931,n934);
or (n931,n932,n933);
and (n932,n886,n896);
and (n933,n887,n890);
xor (n934,n773,n783);
xor (n935,n260,n340);
or (n936,n937,n996);
and (n937,n938,n979);
xor (n938,n939,n978);
or (n939,n940,n977);
and (n940,n941,n976);
xor (n941,n942,n943);
xor (n942,n835,n848);
xor (n943,n944,n963);
xor (n944,n945,n954);
nand (n945,n946,n950);
or (n946,n263,n947);
nor (n947,n948,n949);
and (n948,n327,n277);
and (n949,n331,n278);
or (n950,n265,n951);
nor (n951,n952,n953);
and (n952,n277,n335);
and (n953,n339,n278);
nand (n954,n955,n959);
or (n955,n302,n956);
nor (n956,n957,n958);
and (n957,n365,n312);
and (n958,n369,n313);
or (n959,n960,n322);
nor (n960,n961,n962);
and (n961,n373,n312);
and (n962,n377,n313);
and (n963,n964,n970);
nor (n964,n965,n312);
nor (n965,n966,n969);
and (n966,n967,n277);
not (n967,n968);
and (n968,n547,n306);
and (n969,n321,n549);
nand (n970,n971,n975);
or (n971,n383,n972);
nor (n972,n973,n974);
and (n973,n473,n397);
and (n974,n477,n398);
or (n975,n384,n810);
xor (n976,n905,n918);
and (n977,n942,n943);
xor (n978,n884,n903);
xor (n979,n980,n995);
xor (n980,n981,n992);
xor (n981,n982,n989);
xor (n982,n983,n986);
nand (n983,n984,n985);
or (n984,n221,n924);
or (n985,n222,n242);
nand (n986,n987,n988);
or (n987,n263,n951);
or (n988,n265,n285);
nand (n989,n990,n991);
or (n990,n302,n960);
or (n991,n322,n325);
or (n992,n993,n994);
and (n993,n944,n963);
and (n994,n945,n954);
xor (n995,n796,n804);
and (n996,n939,n978);
and (n997,n827,n828);
xor (n998,n999,n1107);
xor (n999,n1000,n1003);
or (n1000,n1001,n1002);
and (n1001,n829,n929);
and (n1002,n830,n882);
xor (n1003,n1004,n1017);
xor (n1004,n1005,n1014);
or (n1005,n1006,n1013);
and (n1006,n1007,n1012);
xor (n1007,n1008,n1009);
xor (n1008,n752,n767);
or (n1009,n1010,n1011);
and (n1010,n982,n989);
and (n1011,n983,n986);
xor (n1012,n708,n728);
and (n1013,n1008,n1009);
or (n1014,n1015,n1016);
and (n1015,n930,n935);
and (n1016,n931,n934);
xor (n1017,n1018,n1059);
xor (n1018,n1019,n1039);
xor (n1019,n1020,n1033);
xor (n1020,n1021,n1027);
nand (n1021,n1022,n1023);
or (n1022,n680,n725);
or (n1023,n681,n1024);
nor (n1024,n1025,n1026);
and (n1025,n96,n661);
and (n1026,n665,n92);
nand (n1027,n1028,n1029);
or (n1028,n18,n154);
or (n1029,n153,n1030);
nor (n1030,n1031,n1032);
and (n1031,n697,n21);
and (n1032,n701,n22);
nand (n1033,n1034,n1035);
or (n1034,n166,n212);
or (n1035,n211,n1036);
nor (n1036,n1037,n1038);
and (n1037,n195,n624);
and (n1038,n196,n628);
xor (n1039,n1040,n1053);
xor (n1040,n1041,n1047);
nand (n1041,n1042,n1043);
or (n1042,n606,n780);
or (n1043,n1044,n608);
nor (n1044,n1045,n1046);
and (n1045,n192,n599);
and (n1046,n187,n603);
nand (n1047,n1048,n1049);
or (n1048,n635,n786);
or (n1049,n1050,n647);
nor (n1050,n1051,n1052);
and (n1051,n646,n582);
and (n1052,n586,n641);
nand (n1053,n1054,n1055);
or (n1054,n730,n746);
or (n1055,n731,n1056);
nor (n1056,n1057,n1058);
and (n1057,n562,n462);
and (n1058,n566,n455);
xor (n1059,n1060,n1087);
xor (n1060,n1061,n1067);
nand (n1061,n1062,n1063);
or (n1062,n342,n371);
or (n1063,n1064,n343);
nor (n1064,n1065,n1066);
and (n1065,n327,n362);
and (n1066,n331,n355);
nand (n1067,n1068,n1083);
or (n1068,n1069,n1080);
nand (n1069,n754,n1070);
nand (n1070,n1071,n1078);
or (n1071,n763,n1072);
wire s0n1072,s1n1072,notn1072;
or (n1072,s0n1072,s1n1072);
not(notn1072,n82);
and (s0n1072,notn1072,n1073);
and (s1n1072,n82,n1075);
wire s0n1073,s1n1073,notn1073;
or (n1073,s0n1073,s1n1073);
not(notn1073,n26);
and (s0n1073,notn1073,1'b0);
and (s1n1073,n26,n1074);
xor (n1075,n1076,n1077);
not (n1076,n1074);
and (n1077,n760,n761);
or (n1078,n756,n1079);
not (n1079,n1072);
nor (n1080,n1081,n1082);
and (n1081,n1072,n549);
and (n1082,n1079,n547);
or (n1083,n1084,n754);
nor (n1084,n1085,n1086);
and (n1085,n365,n1079);
and (n1086,n369,n1072);
xor (n1087,n1088,n1094);
nor (n1088,n1089,n1079);
nor (n1089,n1090,n1093);
and (n1090,n1091,n362);
not (n1091,n1092);
and (n1092,n547,n756);
and (n1093,n763,n549);
nand (n1094,n1095,n1096);
or (n1095,n712,n671);
or (n1096,n1097,n672);
nor (n1097,n1098,n1105);
and (n1098,n1099,n386);
wire s0n1099,s1n1099,notn1099;
or (n1099,s0n1099,s1n1099);
not(notn1099,n148);
and (s0n1099,notn1099,n1100);
and (s1n1099,n148,n1102);
wire s0n1100,s1n1100,notn1100;
or (n1100,s0n1100,s1n1100);
not(notn1100,n26);
and (s0n1100,notn1100,1'b0);
and (s1n1100,n26,n1101);
xor (n1102,n1103,n1104);
not (n1103,n1101);
and (n1104,n718,n719);
and (n1105,n1106,n387);
not (n1106,n1099);
or (n1107,n1108,n1217);
and (n1108,n1109,n1114);
xor (n1109,n1110,n1111);
xor (n1110,n1007,n1012);
or (n1111,n1112,n1113);
and (n1112,n980,n995);
and (n1113,n981,n992);
or (n1114,n1115,n1216);
and (n1115,n1116,n1215);
xor (n1116,n1117,n1187);
or (n1117,n1118,n1186);
and (n1118,n1119,n1164);
xor (n1119,n1120,n1142);
or (n1120,n1121,n1141);
and (n1121,n1122,n1135);
xor (n1122,n1123,n1129);
nand (n1123,n1124,n1128);
or (n1124,n452,n1125);
nor (n1125,n1126,n1127);
and (n1126,n653,n470);
and (n1127,n657,n466);
or (n1128,n816,n453);
nand (n1129,n1130,n1134);
or (n1130,n488,n1131);
nor (n1131,n1132,n1133);
and (n1132,n498,n214);
and (n1133,n499,n218);
or (n1134,n512,n838);
nand (n1135,n1136,n1140);
or (n1136,n606,n1137);
nor (n1137,n1138,n1139);
and (n1138,n192,n252);
and (n1139,n187,n256);
or (n1140,n844,n608);
and (n1141,n1123,n1129);
or (n1142,n1143,n1163);
and (n1143,n1144,n1157);
xor (n1144,n1145,n1151);
nand (n1145,n1146,n1150);
or (n1146,n635,n1147);
nor (n1147,n1148,n1149);
and (n1148,n646,n156);
and (n1149,n641,n163);
or (n1150,n850,n647);
nand (n1151,n1152,n1156);
or (n1152,n1153,n671);
nor (n1153,n1154,n1155);
and (n1154,n554,n386);
and (n1155,n558,n387);
or (n1156,n860,n672);
nand (n1157,n1158,n1162);
or (n1158,n680,n1159);
nor (n1159,n1160,n1161);
and (n1160,n96,n506);
and (n1161,n92,n510);
or (n1162,n681,n866);
and (n1163,n1145,n1151);
or (n1164,n1165,n1185);
and (n1165,n1166,n1179);
xor (n1166,n1167,n1173);
nand (n1167,n1168,n1172);
or (n1168,n221,n1169);
nor (n1169,n1170,n1171);
and (n1170,n241,n335);
and (n1171,n234,n339);
or (n1172,n222,n920);
nand (n1173,n1174,n1178);
or (n1174,n263,n1175);
nor (n1175,n1176,n1177);
and (n1176,n373,n277);
and (n1177,n377,n278);
or (n1178,n265,n947);
nand (n1179,n1180,n1184);
or (n1180,n302,n1181);
nor (n1181,n1182,n1183);
and (n1182,n313,n549);
and (n1183,n312,n547);
or (n1184,n322,n956);
and (n1185,n1167,n1173);
and (n1186,n1120,n1142);
or (n1187,n1188,n1214);
and (n1188,n1189,n1213);
xor (n1189,n1190,n1212);
or (n1190,n1191,n1211);
and (n1191,n1192,n1205);
xor (n1192,n1193,n1199);
nand (n1193,n1194,n1198);
or (n1194,n730,n1195);
nor (n1195,n1196,n1197);
and (n1196,n574,n462);
and (n1197,n578,n455);
or (n1198,n872,n731);
nand (n1199,n1200,n1204);
or (n1200,n18,n1201);
nor (n1201,n1202,n1203);
and (n1202,n21,n591);
and (n1203,n22,n595);
or (n1204,n153,n908);
nand (n1205,n1206,n1210);
or (n1206,n166,n1207);
nor (n1207,n1208,n1209);
and (n1208,n195,n295);
and (n1209,n196,n299);
or (n1210,n211,n914);
and (n1211,n1193,n1199);
xor (n1212,n857,n870);
xor (n1213,n806,n814);
and (n1214,n1190,n1212);
xor (n1215,n832,n880);
and (n1216,n1117,n1187);
and (n1217,n1110,n1111);
not (n1218,n1219);
or (n1219,n1220,n1340);
and (n1220,n1221,n1224);
xor (n1221,n1222,n1223);
xor (n1222,n1109,n1114);
xor (n1223,n826,n936);
or (n1224,n1225,n1339);
and (n1225,n1226,n1326);
xor (n1226,n1227,n1325);
or (n1227,n1228,n1324);
and (n1228,n1229,n1280);
xor (n1229,n1230,n1279);
or (n1230,n1231,n1278);
and (n1231,n1232,n1256);
xor (n1232,n1233,n1234);
xor (n1233,n964,n970);
or (n1234,n1235,n1255);
and (n1235,n1236,n1249);
xor (n1236,n1237,n1243);
nand (n1237,n1238,n1242);
or (n1238,n488,n1239);
nor (n1239,n1240,n1241);
and (n1240,n498,n205);
and (n1241,n499,n209);
or (n1242,n512,n1131);
nand (n1243,n1244,n1248);
or (n1244,n606,n1245);
nor (n1245,n1246,n1247);
and (n1246,n192,n244);
and (n1247,n187,n248);
or (n1248,n1137,n608);
nand (n1249,n1250,n1254);
or (n1250,n635,n1251);
nor (n1251,n1252,n1253);
and (n1252,n646,n99);
and (n1253,n641,n151);
or (n1254,n1147,n647);
and (n1255,n1237,n1243);
or (n1256,n1257,n1277);
and (n1257,n1258,n1271);
xor (n1258,n1259,n1265);
nand (n1259,n1260,n1264);
or (n1260,n1261,n671);
nor (n1261,n1262,n1263);
and (n1262,n481,n386);
and (n1263,n485,n387);
or (n1264,n1153,n672);
nand (n1265,n1266,n1270);
or (n1266,n730,n1267);
nor (n1267,n1268,n1269);
and (n1268,n661,n462);
and (n1269,n665,n455);
or (n1270,n731,n1195);
nand (n1271,n1272,n1276);
or (n1272,n680,n1273);
nor (n1273,n1274,n1275);
and (n1274,n96,n599);
and (n1275,n92,n603);
or (n1276,n681,n1159);
and (n1277,n1259,n1265);
and (n1278,n1233,n1234);
xor (n1279,n1119,n1164);
or (n1280,n1281,n1323);
and (n1281,n1282,n1322);
xor (n1282,n1283,n1300);
or (n1283,n1284,n1299);
and (n1284,n1285,n1293);
xor (n1285,n1286,n1287);
nor (n1286,n322,n549);
nand (n1287,n1288,n1292);
or (n1288,n383,n1289);
nor (n1289,n1290,n1291);
and (n1290,n582,n397);
and (n1291,n586,n398);
or (n1292,n384,n972);
nand (n1293,n1294,n1298);
or (n1294,n452,n1295);
nor (n1295,n1296,n1297);
and (n1296,n697,n470);
and (n1297,n701,n466);
or (n1298,n1125,n453);
and (n1299,n1286,n1287);
or (n1300,n1301,n1321);
and (n1301,n1302,n1315);
xor (n1302,n1303,n1309);
nand (n1303,n1304,n1308);
or (n1304,n18,n1305);
nor (n1305,n1306,n1307);
and (n1306,n21,n624);
and (n1307,n22,n628);
or (n1308,n153,n1201);
nand (n1309,n1310,n1314);
or (n1310,n166,n1311);
nor (n1311,n1312,n1313);
and (n1312,n287,n195);
and (n1313,n291,n196);
or (n1314,n211,n1207);
nand (n1315,n1316,n1320);
or (n1316,n221,n1317);
nor (n1317,n1318,n1319);
and (n1318,n327,n241);
and (n1319,n331,n234);
or (n1320,n222,n1169);
and (n1321,n1303,n1309);
xor (n1322,n1144,n1157);
and (n1323,n1283,n1300);
and (n1324,n1230,n1279);
xor (n1325,n1116,n1215);
or (n1326,n1327,n1338);
and (n1327,n1328,n1337);
xor (n1328,n1329,n1330);
xor (n1329,n1189,n1213);
or (n1330,n1331,n1336);
and (n1331,n1332,n1335);
xor (n1332,n1333,n1334);
xor (n1333,n1122,n1135);
xor (n1334,n1192,n1205);
xor (n1335,n1166,n1179);
and (n1336,n1333,n1334);
xor (n1337,n941,n976);
and (n1338,n1329,n1330);
and (n1339,n1227,n1325);
and (n1340,n1222,n1223);
nor (n1341,n6,n1218);
not (n1342,n1343);
nor (n1343,n1344,n3083);
nor (n1344,n1345,n3078);
nor (n1345,n1346,n3077);
and (n1346,n1347,n3064);
or (n1347,n1348,n3063);
and (n1348,n1349,n1706);
xor (n1349,n1350,n1691);
or (n1350,n1351,n1690);
and (n1351,n1352,n1659);
xor (n1352,n1353,n1364);
xor (n1353,n1354,n1363);
xor (n1354,n1355,n1362);
or (n1355,n1356,n1361);
and (n1356,n1357,n1360);
xor (n1357,n1358,n1359);
xor (n1358,n1285,n1293);
xor (n1359,n1236,n1249);
xor (n1360,n1302,n1315);
and (n1361,n1358,n1359);
xor (n1362,n1332,n1335);
xor (n1363,n1282,n1322);
or (n1364,n1365,n1658);
and (n1365,n1366,n1583);
xor (n1366,n1367,n1503);
or (n1367,n1368,n1502);
and (n1368,n1369,n1420);
xor (n1369,n1370,n1390);
xor (n1370,n1371,n1384);
xor (n1371,n1372,n1378);
nand (n1372,n1373,n1377);
or (n1373,n452,n1374);
nor (n1374,n1375,n1376);
and (n1375,n156,n470);
and (n1376,n163,n466);
or (n1377,n1295,n453);
nand (n1378,n1379,n1383);
or (n1379,n488,n1380);
nor (n1380,n1381,n1382);
and (n1381,n498,n252);
and (n1382,n499,n256);
or (n1383,n512,n1239);
nand (n1384,n1385,n1389);
or (n1385,n606,n1386);
nor (n1386,n1387,n1388);
and (n1387,n192,n295);
and (n1388,n187,n299);
or (n1389,n1245,n608);
xor (n1390,n1391,n1407);
xor (n1391,n1392,n1398);
nand (n1392,n1393,n1397);
or (n1393,n221,n1394);
nor (n1394,n1395,n1396);
and (n1395,n373,n241);
and (n1396,n377,n234);
or (n1397,n222,n1317);
nand (n1398,n1399,n1403);
or (n1399,n263,n1400);
nor (n1400,n1401,n1402);
and (n1401,n278,n549);
and (n1402,n277,n547);
or (n1403,n265,n1404);
nor (n1404,n1405,n1406);
and (n1405,n365,n277);
and (n1406,n369,n278);
xor (n1407,n1408,n1414);
nor (n1408,n1409,n277);
nor (n1409,n1410,n1413);
and (n1410,n1411,n241);
not (n1411,n1412);
and (n1412,n547,n268);
and (n1413,n267,n549);
nand (n1414,n1415,n1419);
or (n1415,n383,n1416);
nor (n1416,n1417,n1418);
and (n1417,n574,n397);
and (n1418,n578,n398);
or (n1419,n1289,n384);
or (n1420,n1421,n1501);
and (n1421,n1422,n1470);
xor (n1422,n1423,n1439);
and (n1423,n1424,n1430);
nor (n1424,n1425,n241);
nor (n1425,n1426,n1429);
and (n1426,n1427,n195);
not (n1427,n1428);
and (n1428,n547,n224);
and (n1429,n231,n549);
nand (n1430,n1431,n1435);
or (n1431,n383,n1432);
nor (n1432,n1433,n1434);
and (n1433,n653,n397);
and (n1434,n657,n398);
or (n1435,n384,n1436);
nor (n1436,n1437,n1438);
and (n1437,n661,n397);
and (n1438,n665,n398);
or (n1439,n1440,n1469);
and (n1440,n1441,n1460);
xor (n1441,n1442,n1451);
nand (n1442,n1443,n1447);
or (n1443,n635,n1444);
nor (n1444,n1445,n1446);
and (n1445,n646,n591);
and (n1446,n641,n595);
or (n1447,n1448,n647);
nor (n1448,n1449,n1450);
and (n1449,n646,n599);
and (n1450,n641,n603);
nand (n1451,n1452,n1456);
or (n1452,n1453,n671);
nor (n1453,n1454,n1455);
and (n1454,n574,n386);
and (n1455,n578,n387);
or (n1456,n1457,n672);
nor (n1457,n1458,n1459);
and (n1458,n582,n386);
and (n1459,n586,n387);
nand (n1460,n1461,n1465);
or (n1461,n730,n1462);
nor (n1462,n1463,n1464);
and (n1463,n156,n462);
and (n1464,n163,n455);
or (n1465,n1466,n731);
nor (n1466,n1467,n1468);
and (n1467,n697,n462);
and (n1468,n701,n455);
and (n1469,n1442,n1451);
or (n1470,n1471,n1500);
and (n1471,n1472,n1491);
xor (n1472,n1473,n1482);
nand (n1473,n1474,n1478);
or (n1474,n452,n1475);
nor (n1475,n1476,n1477);
and (n1476,n506,n470);
and (n1477,n510,n466);
or (n1478,n453,n1479);
nor (n1479,n1480,n1481);
and (n1480,n99,n470);
and (n1481,n151,n466);
nand (n1482,n1483,n1487);
or (n1483,n488,n1484);
nor (n1484,n1485,n1486);
and (n1485,n498,n295);
and (n1486,n499,n299);
or (n1487,n1488,n512);
nor (n1488,n1489,n1490);
and (n1489,n498,n244);
and (n1490,n499,n248);
nand (n1491,n1492,n1496);
or (n1492,n606,n1493);
nor (n1493,n1494,n1495);
and (n1494,n192,n335);
and (n1495,n187,n339);
or (n1496,n1497,n608);
nor (n1497,n1498,n1499);
and (n1498,n192,n287);
and (n1499,n187,n291);
and (n1500,n1473,n1482);
and (n1501,n1423,n1439);
and (n1502,n1370,n1390);
xor (n1503,n1504,n1536);
xor (n1504,n1505,n1508);
or (n1505,n1506,n1507);
and (n1506,n1391,n1407);
and (n1507,n1392,n1398);
xor (n1508,n1509,n1514);
xor (n1509,n1510,n1513);
nand (n1510,n1511,n1512);
or (n1511,n263,n1404);
or (n1512,n265,n1175);
and (n1513,n1408,n1414);
or (n1514,n1515,n1535);
and (n1515,n1516,n1529);
xor (n1516,n1517,n1523);
nand (n1517,n1518,n1522);
or (n1518,n635,n1519);
nor (n1519,n1520,n1521);
and (n1520,n646,n506);
and (n1521,n641,n510);
or (n1522,n1251,n647);
nand (n1523,n1524,n1528);
or (n1524,n1525,n671);
nor (n1525,n1526,n1527);
and (n1526,n473,n386);
and (n1527,n477,n387);
or (n1528,n1261,n672);
nand (n1529,n1530,n1534);
or (n1530,n730,n1531);
nor (n1531,n1532,n1533);
and (n1532,n653,n462);
and (n1533,n657,n455);
or (n1534,n1267,n731);
and (n1535,n1517,n1523);
or (n1536,n1537,n1582);
and (n1537,n1538,n1569);
xor (n1538,n1539,n1558);
or (n1539,n1540,n1557);
and (n1540,n1541,n1548);
xor (n1541,n1542,n1545);
nand (n1542,n1543,n1544);
or (n1543,n1457,n671);
or (n1544,n1525,n672);
nand (n1545,n1546,n1547);
or (n1546,n730,n1466);
or (n1547,n1531,n731);
nand (n1548,n1549,n1553);
or (n1549,n680,n1550);
nor (n1550,n1551,n1552);
and (n1551,n96,n624);
and (n1552,n92,n628);
or (n1553,n681,n1554);
nor (n1554,n1555,n1556);
and (n1555,n96,n591);
and (n1556,n92,n595);
and (n1557,n1542,n1545);
or (n1558,n1559,n1568);
and (n1559,n1560,n1565);
xor (n1560,n1561,n1562);
nor (n1561,n265,n549);
nand (n1562,n1563,n1564);
or (n1563,n383,n1436);
or (n1564,n384,n1416);
nand (n1565,n1566,n1567);
or (n1566,n452,n1479);
or (n1567,n453,n1374);
and (n1568,n1561,n1562);
or (n1569,n1570,n1581);
and (n1570,n1571,n1578);
xor (n1571,n1572,n1575);
nand (n1572,n1573,n1574);
or (n1573,n488,n1488);
or (n1574,n512,n1380);
nand (n1575,n1576,n1577);
or (n1576,n606,n1497);
or (n1577,n1386,n608);
nand (n1578,n1579,n1580);
or (n1579,n635,n1448);
or (n1580,n1519,n647);
and (n1581,n1572,n1575);
and (n1582,n1539,n1558);
or (n1583,n1584,n1657);
and (n1584,n1585,n1621);
xor (n1585,n1586,n1620);
or (n1586,n1587,n1619);
and (n1587,n1588,n1618);
xor (n1588,n1589,n1617);
or (n1589,n1590,n1616);
and (n1590,n1591,n1607);
xor (n1591,n1592,n1598);
nand (n1592,n1593,n1597);
or (n1593,n680,n1594);
nor (n1594,n1595,n1596);
and (n1595,n96,n214);
and (n1596,n92,n218);
or (n1597,n681,n1550);
nand (n1598,n1599,n1603);
or (n1599,n18,n1600);
nor (n1600,n1601,n1602);
and (n1601,n21,n252);
and (n1602,n22,n256);
or (n1603,n153,n1604);
nor (n1604,n1605,n1606);
and (n1605,n21,n205);
and (n1606,n22,n209);
nand (n1607,n1608,n1612);
or (n1608,n166,n1609);
nor (n1609,n1610,n1611);
and (n1610,n373,n195);
and (n1611,n377,n196);
or (n1612,n211,n1613);
nor (n1613,n1614,n1615);
and (n1614,n327,n195);
and (n1615,n331,n196);
and (n1616,n1592,n1598);
xor (n1617,n1541,n1548);
xor (n1618,n1571,n1578);
and (n1619,n1589,n1617);
xor (n1620,n1538,n1569);
xor (n1621,n1622,n1641);
xor (n1622,n1623,n1640);
xor (n1623,n1624,n1634);
xor (n1624,n1625,n1628);
nand (n1625,n1626,n1627);
or (n1626,n680,n1554);
or (n1627,n681,n1273);
nand (n1628,n1629,n1633);
or (n1629,n18,n1630);
nor (n1630,n1631,n1632);
and (n1631,n21,n214);
and (n1632,n22,n218);
or (n1633,n153,n1305);
nand (n1634,n1635,n1639);
or (n1635,n166,n1636);
nor (n1636,n1637,n1638);
and (n1637,n195,n335);
and (n1638,n196,n339);
or (n1639,n211,n1311);
xor (n1640,n1516,n1529);
or (n1641,n1642,n1656);
and (n1642,n1643,n1650);
xor (n1643,n1644,n1647);
nand (n1644,n1645,n1646);
or (n1645,n18,n1604);
or (n1646,n153,n1630);
nand (n1647,n1648,n1649);
or (n1648,n166,n1613);
or (n1649,n211,n1636);
nand (n1650,n1651,n1655);
or (n1651,n221,n1652);
nor (n1652,n1653,n1654);
and (n1653,n365,n241);
and (n1654,n369,n234);
or (n1655,n222,n1394);
and (n1656,n1644,n1647);
and (n1657,n1586,n1620);
and (n1658,n1367,n1503);
xor (n1659,n1660,n1681);
xor (n1660,n1661,n1664);
or (n1661,n1662,n1663);
and (n1662,n1504,n1536);
and (n1663,n1505,n1508);
xor (n1664,n1665,n1680);
xor (n1665,n1666,n1669);
or (n1666,n1667,n1668);
and (n1667,n1509,n1514);
and (n1668,n1510,n1513);
or (n1669,n1670,n1679);
and (n1670,n1671,n1678);
xor (n1671,n1672,n1675);
or (n1672,n1673,n1674);
and (n1673,n1371,n1384);
and (n1674,n1372,n1378);
or (n1675,n1676,n1677);
and (n1676,n1624,n1634);
and (n1677,n1625,n1628);
xor (n1678,n1258,n1271);
and (n1679,n1672,n1675);
xor (n1680,n1232,n1256);
or (n1681,n1682,n1689);
and (n1682,n1683,n1688);
xor (n1683,n1684,n1687);
or (n1684,n1685,n1686);
and (n1685,n1622,n1641);
and (n1686,n1623,n1640);
xor (n1687,n1357,n1360);
xor (n1688,n1671,n1678);
and (n1689,n1684,n1687);
and (n1690,n1353,n1364);
xor (n1691,n1692,n1697);
xor (n1692,n1693,n1694);
xor (n1693,n1328,n1337);
or (n1694,n1695,n1696);
and (n1695,n1660,n1681);
and (n1696,n1661,n1664);
xor (n1697,n1698,n1705);
xor (n1698,n1699,n1702);
or (n1699,n1700,n1701);
and (n1700,n1665,n1680);
and (n1701,n1666,n1669);
or (n1702,n1703,n1704);
and (n1703,n1354,n1363);
and (n1704,n1355,n1362);
xor (n1705,n1229,n1280);
nand (n1706,n1707,n3057);
or (n1707,n1708,n3039,n3052);
nor (n1708,n1709,n3038);
and (n1709,n1710,n3017);
or (n1710,n1711,n3016);
and (n1711,n1712,n2066);
xor (n1712,n1713,n2039);
or (n1713,n1714,n2038);
and (n1714,n1715,n1953);
xor (n1715,n1716,n1840);
xor (n1716,n1717,n1810);
xor (n1717,n1718,n1749);
xor (n1718,n1719,n1727);
xor (n1719,n1720,n1726);
nand (n1720,n1721,n1725);
or (n1721,n221,n1722);
nor (n1722,n1723,n1724);
and (n1723,n234,n549);
and (n1724,n241,n547);
or (n1725,n222,n1652);
xor (n1726,n1424,n1430);
or (n1727,n1728,n1748);
and (n1728,n1729,n1742);
xor (n1729,n1730,n1736);
nand (n1730,n1731,n1735);
or (n1731,n635,n1732);
nor (n1732,n1733,n1734);
and (n1733,n646,n624);
and (n1734,n641,n628);
or (n1735,n1444,n647);
nand (n1736,n1737,n1741);
or (n1737,n730,n1738);
nor (n1738,n1739,n1740);
and (n1739,n99,n462);
and (n1740,n151,n455);
or (n1741,n731,n1462);
nand (n1742,n1743,n1747);
or (n1743,n680,n1744);
nor (n1744,n1745,n1746);
and (n1745,n96,n205);
and (n1746,n92,n209);
or (n1747,n681,n1594);
and (n1748,n1730,n1736);
or (n1749,n1750,n1809);
and (n1750,n1751,n1808);
xor (n1751,n1752,n1783);
or (n1752,n1753,n1782);
and (n1753,n1754,n1773);
xor (n1754,n1755,n1764);
nand (n1755,n1756,n1760);
or (n1756,n452,n1757);
nor (n1757,n1758,n1759);
and (n1758,n591,n470);
and (n1759,n595,n466);
or (n1760,n453,n1761);
nor (n1761,n1762,n1763);
and (n1762,n599,n470);
and (n1763,n603,n466);
nand (n1764,n1765,n1769);
or (n1765,n488,n1766);
nor (n1766,n1767,n1768);
and (n1767,n498,n335);
and (n1768,n339,n499);
or (n1769,n512,n1770);
nor (n1770,n1771,n1772);
and (n1771,n287,n498);
and (n1772,n291,n499);
nand (n1773,n1774,n1778);
or (n1774,n606,n1775);
nor (n1775,n1776,n1777);
and (n1776,n373,n192);
and (n1777,n377,n187);
or (n1778,n1779,n608);
nor (n1779,n1780,n1781);
and (n1780,n327,n192);
and (n1781,n331,n187);
and (n1782,n1755,n1764);
or (n1783,n1784,n1807);
and (n1784,n1785,n1801);
xor (n1785,n1786,n1795);
nand (n1786,n1787,n1791);
or (n1787,n383,n1788);
nor (n1788,n1789,n1790);
and (n1789,n397,n156);
and (n1790,n163,n398);
or (n1791,n1792,n384);
nor (n1792,n1793,n1794);
and (n1793,n697,n397);
and (n1794,n701,n398);
nand (n1795,n1796,n1800);
or (n1796,n635,n1797);
nor (n1797,n1798,n1799);
and (n1798,n646,n214);
and (n1799,n641,n218);
or (n1800,n1732,n647);
nand (n1801,n1802,n1806);
or (n1802,n730,n1803);
nor (n1803,n1804,n1805);
and (n1804,n506,n462);
and (n1805,n510,n455);
or (n1806,n731,n1738);
and (n1807,n1786,n1795);
xor (n1808,n1729,n1742);
and (n1809,n1752,n1783);
xor (n1810,n1811,n1839);
xor (n1811,n1812,n1826);
or (n1812,n1813,n1825);
and (n1813,n1814,n1822);
xor (n1814,n1815,n1816);
nor (n1815,n222,n549);
nand (n1816,n1817,n1821);
or (n1817,n1818,n671);
nor (n1818,n1819,n1820);
and (n1819,n661,n386);
and (n1820,n665,n387);
or (n1821,n1453,n672);
nand (n1822,n1823,n1824);
or (n1823,n452,n1761);
or (n1824,n453,n1475);
and (n1825,n1815,n1816);
or (n1826,n1827,n1838);
and (n1827,n1828,n1835);
xor (n1828,n1829,n1832);
nand (n1829,n1830,n1831);
or (n1830,n488,n1770);
or (n1831,n1484,n512);
nand (n1832,n1833,n1834);
or (n1833,n606,n1779);
or (n1834,n1493,n608);
nand (n1835,n1836,n1837);
or (n1836,n383,n1792);
or (n1837,n384,n1432);
and (n1838,n1829,n1832);
xor (n1839,n1441,n1460);
xor (n1840,n1841,n1903);
xor (n1841,n1842,n1876);
or (n1842,n1843,n1875);
and (n1843,n1844,n1847);
xor (n1844,n1845,n1846);
xor (n1845,n1814,n1822);
xor (n1846,n1828,n1835);
or (n1847,n1848,n1874);
and (n1848,n1849,n1865);
xor (n1849,n1850,n1856);
nand (n1850,n1851,n1855);
or (n1851,n680,n1852);
nor (n1852,n1853,n1854);
and (n1853,n96,n252);
and (n1854,n92,n256);
or (n1855,n681,n1744);
nand (n1856,n1857,n1861);
or (n1857,n18,n1858);
nor (n1858,n1859,n1860);
and (n1859,n21,n295);
and (n1860,n22,n299);
or (n1861,n1862,n153);
nor (n1862,n1863,n1864);
and (n1863,n21,n244);
and (n1864,n22,n248);
nand (n1865,n1866,n1870);
or (n1866,n166,n1867);
nor (n1867,n1868,n1869);
and (n1868,n196,n549);
and (n1869,n195,n547);
or (n1870,n211,n1871);
nor (n1871,n1872,n1873);
and (n1872,n365,n195);
and (n1873,n369,n196);
and (n1874,n1850,n1856);
and (n1875,n1845,n1846);
xor (n1876,n1877,n1880);
xor (n1877,n1878,n1879);
xor (n1878,n1472,n1491);
xor (n1879,n1591,n1607);
or (n1880,n1881,n1902);
and (n1881,n1882,n1889);
xor (n1882,n1883,n1886);
nand (n1883,n1884,n1885);
or (n1884,n18,n1862);
or (n1885,n153,n1600);
nand (n1886,n1887,n1888);
or (n1887,n166,n1871);
or (n1888,n211,n1609);
and (n1889,n1890,n1896);
nor (n1890,n1891,n195);
nor (n1891,n1892,n1895);
and (n1892,n1893,n192);
not (n1893,n1894);
and (n1894,n547,n169);
and (n1895,n191,n549);
nand (n1896,n1897,n1901);
or (n1897,n1898,n671);
nor (n1898,n1899,n1900);
and (n1899,n653,n386);
and (n1900,n657,n387);
or (n1901,n1818,n672);
and (n1902,n1883,n1886);
or (n1903,n1904,n1952);
and (n1904,n1905,n1951);
xor (n1905,n1906,n1907);
xor (n1906,n1882,n1889);
or (n1907,n1908,n1950);
and (n1908,n1909,n1928);
xor (n1909,n1910,n1911);
xor (n1910,n1890,n1896);
or (n1911,n1912,n1927);
and (n1912,n1913,n1921);
xor (n1913,n1914,n1915);
nor (n1914,n211,n549);
nand (n1915,n1916,n1920);
or (n1916,n1917,n671);
nor (n1917,n1918,n1919);
and (n1918,n697,n386);
and (n1919,n701,n387);
or (n1920,n1898,n672);
nand (n1921,n1922,n1923);
or (n1922,n1757,n453);
or (n1923,n452,n1924);
nor (n1924,n1925,n1926);
and (n1925,n624,n470);
and (n1926,n628,n466);
and (n1927,n1914,n1915);
or (n1928,n1929,n1949);
and (n1929,n1930,n1943);
xor (n1930,n1931,n1937);
nand (n1931,n1932,n1936);
or (n1932,n488,n1933);
nor (n1933,n1934,n1935);
and (n1934,n327,n498);
and (n1935,n331,n499);
or (n1936,n1766,n512);
nand (n1937,n1938,n1942);
or (n1938,n606,n1939);
nor (n1939,n1940,n1941);
and (n1940,n365,n192);
and (n1941,n369,n187);
or (n1942,n1775,n608);
nand (n1943,n1944,n1948);
or (n1944,n383,n1945);
nor (n1945,n1946,n1947);
and (n1946,n397,n99);
and (n1947,n151,n398);
or (n1948,n384,n1788);
and (n1949,n1931,n1937);
and (n1950,n1910,n1911);
xor (n1951,n1751,n1808);
and (n1952,n1906,n1907);
or (n1953,n1954,n2037);
and (n1954,n1955,n1985);
xor (n1955,n1956,n1984);
or (n1956,n1957,n1983);
and (n1957,n1958,n1982);
xor (n1958,n1959,n1981);
or (n1959,n1960,n1980);
and (n1960,n1961,n1974);
xor (n1961,n1962,n1968);
nand (n1962,n1963,n1967);
or (n1963,n635,n1964);
nor (n1964,n1965,n1966);
and (n1965,n646,n205);
and (n1966,n641,n209);
or (n1967,n1797,n647);
nand (n1968,n1969,n1973);
or (n1969,n730,n1970);
nor (n1970,n1971,n1972);
and (n1971,n599,n462);
and (n1972,n603,n455);
or (n1973,n731,n1803);
nand (n1974,n1975,n1979);
or (n1975,n680,n1976);
nor (n1976,n1977,n1978);
and (n1977,n96,n244);
and (n1978,n92,n248);
or (n1979,n681,n1852);
and (n1980,n1962,n1968);
xor (n1981,n1785,n1801);
xor (n1982,n1754,n1773);
and (n1983,n1959,n1981);
xor (n1984,n1844,n1847);
or (n1985,n1986,n2036);
and (n1986,n1987,n2035);
xor (n1987,n1988,n1989);
xor (n1988,n1849,n1865);
or (n1989,n1990,n2034);
and (n1990,n1991,n2011);
xor (n1991,n1992,n1998);
nand (n1992,n1993,n1997);
or (n1993,n18,n1994);
nor (n1994,n1995,n1996);
and (n1995,n21,n287);
and (n1996,n22,n291);
or (n1997,n1858,n153);
and (n1998,n1999,n2005);
nor (n1999,n2000,n192);
nor (n2000,n2001,n2004);
and (n2001,n498,n2002);
not (n2002,n2003);
and (n2003,n547,n611);
and (n2004,n610,n549);
nand (n2005,n2006,n2010);
or (n2006,n2007,n671);
nor (n2007,n2008,n2009);
and (n2008,n156,n386);
and (n2009,n163,n387);
or (n2010,n1917,n672);
or (n2011,n2012,n2033);
and (n2012,n2013,n2026);
xor (n2013,n2014,n2020);
nand (n2014,n2015,n2019);
or (n2015,n452,n2016);
nor (n2016,n2017,n2018);
and (n2017,n214,n470);
and (n2018,n218,n466);
or (n2019,n1924,n453);
nand (n2020,n2021,n2025);
or (n2021,n488,n2022);
nor (n2022,n2023,n2024);
and (n2023,n373,n498);
and (n2024,n377,n499);
or (n2025,n512,n1933);
nand (n2026,n2027,n2032);
or (n2027,n2028,n606);
not (n2028,n2029);
nand (n2029,n2030,n2031);
or (n2030,n192,n547);
or (n2031,n187,n549);
or (n2032,n1939,n608);
and (n2033,n2014,n2020);
and (n2034,n1992,n1998);
xor (n2035,n1909,n1928);
and (n2036,n1988,n1989);
and (n2037,n1956,n1984);
and (n2038,n1716,n1840);
xor (n2039,n2040,n2063);
xor (n2040,n2041,n2050);
xor (n2041,n2042,n2047);
xor (n2042,n2043,n2044);
xor (n2043,n1422,n1470);
or (n2044,n2045,n2046);
and (n2045,n1811,n1839);
and (n2046,n1812,n1826);
or (n2047,n2048,n2049);
and (n2048,n1877,n1880);
and (n2049,n1878,n1879);
xor (n2050,n2051,n2060);
xor (n2051,n2052,n2053);
xor (n2052,n1588,n1618);
xor (n2053,n2054,n2057);
xor (n2054,n2055,n2056);
xor (n2055,n1560,n1565);
xor (n2056,n1643,n1650);
or (n2057,n2058,n2059);
and (n2058,n1719,n1727);
and (n2059,n1720,n1726);
or (n2060,n2061,n2062);
and (n2061,n1717,n1810);
and (n2062,n1718,n1749);
or (n2063,n2064,n2065);
and (n2064,n1841,n1903);
and (n2065,n1842,n1876);
nand (n2066,n2067,n3010);
or (n2067,n2068,n3003);
nand (n2068,n2069,n2992);
not (n2069,n2070);
nor (n2070,n2071,n2981);
nor (n2071,n2072,n2930);
nand (n2072,n2073,n2804);
or (n2073,n2074,n2803);
and (n2074,n2075,n2393);
xor (n2075,n2076,n2307);
or (n2076,n2077,n2306);
and (n2077,n2078,n2255);
xor (n2078,n2079,n2162);
xor (n2079,n2080,n2131);
xor (n2080,n2081,n2102);
xor (n2081,n2082,n2093);
xor (n2082,n2083,n2084);
nor (n2083,n512,n549);
nand (n2084,n2085,n2089);
or (n2085,n2086,n671);
nor (n2086,n2087,n2088);
and (n2087,n386,n599);
and (n2088,n603,n387);
or (n2089,n2090,n672);
nor (n2090,n2091,n2092);
and (n2091,n506,n386);
and (n2092,n510,n387);
nand (n2093,n2094,n2098);
or (n2094,n383,n2095);
nor (n2095,n2096,n2097);
and (n2096,n397,n624);
and (n2097,n628,n398);
or (n2098,n384,n2099);
nor (n2099,n2100,n2101);
and (n2100,n591,n397);
and (n2101,n595,n398);
or (n2102,n2103,n2130);
and (n2103,n2104,n2120);
xor (n2104,n2105,n2111);
nand (n2105,n2106,n2110);
or (n2106,n383,n2107);
nor (n2107,n2108,n2109);
and (n2108,n397,n214);
and (n2109,n218,n398);
or (n2110,n384,n2095);
nand (n2111,n2112,n2116);
or (n2112,n452,n2113);
nor (n2113,n2114,n2115);
and (n2114,n295,n470);
and (n2115,n299,n466);
or (n2116,n453,n2117);
nor (n2117,n2118,n2119);
and (n2118,n244,n470);
and (n2119,n248,n466);
nand (n2120,n2121,n2126);
or (n2121,n2122,n635);
not (n2122,n2123);
nand (n2123,n2124,n2125);
or (n2124,n641,n339);
or (n2125,n646,n335);
or (n2126,n2127,n647);
nor (n2127,n2128,n2129);
and (n2128,n646,n287);
and (n2129,n641,n291);
and (n2130,n2105,n2111);
or (n2131,n2132,n2161);
and (n2132,n2133,n2152);
xor (n2133,n2134,n2143);
nand (n2134,n2135,n2139);
or (n2135,n730,n2136);
nor (n2136,n2137,n2138);
and (n2137,n252,n462);
and (n2138,n256,n455);
or (n2139,n2140,n731);
nor (n2140,n2141,n2142);
and (n2141,n205,n462);
and (n2142,n209,n455);
nand (n2143,n2144,n2148);
or (n2144,n680,n2145);
nor (n2145,n2146,n2147);
and (n2146,n373,n96);
and (n2147,n377,n92);
or (n2148,n2149,n681);
nor (n2149,n2150,n2151);
and (n2150,n327,n96);
and (n2151,n331,n92);
nand (n2152,n2153,n2157);
or (n2153,n153,n2154);
nor (n2154,n2155,n2156);
and (n2155,n365,n21);
and (n2156,n369,n22);
or (n2157,n18,n2158);
nor (n2158,n2159,n2160);
and (n2159,n22,n549);
and (n2160,n21,n547);
and (n2161,n2134,n2143);
xor (n2162,n2163,n2211);
xor (n2163,n2164,n2191);
xor (n2164,n2165,n2178);
xor (n2165,n2166,n2172);
nand (n2166,n2167,n2168);
or (n2167,n680,n2149);
or (n2168,n2169,n681);
nor (n2169,n2170,n2171);
and (n2170,n96,n335);
and (n2171,n92,n339);
nand (n2172,n2173,n2174);
or (n2173,n18,n2154);
or (n2174,n2175,n153);
nor (n2175,n2176,n2177);
and (n2176,n373,n21);
and (n2177,n377,n22);
and (n2178,n2179,n2185);
nand (n2179,n2180,n2184);
or (n2180,n2181,n671);
nor (n2181,n2182,n2183);
and (n2182,n386,n591);
and (n2183,n595,n387);
or (n2184,n2086,n672);
nor (n2185,n2186,n21);
nor (n2186,n2187,n2190);
and (n2187,n96,n2188);
not (n2188,n2189);
and (n2189,n547,n85);
and (n2190,n89,n549);
xor (n2191,n2192,n2205);
xor (n2192,n2193,n2199);
nand (n2193,n2194,n2195);
or (n2194,n452,n2117);
or (n2195,n2196,n453);
nor (n2196,n2197,n2198);
and (n2197,n252,n470);
and (n2198,n256,n466);
nand (n2199,n2200,n2201);
or (n2200,n635,n2127);
or (n2201,n2202,n647);
nor (n2202,n2203,n2204);
and (n2203,n646,n295);
and (n2204,n641,n299);
nand (n2205,n2206,n2210);
or (n2206,n731,n2207);
nor (n2207,n2208,n2209);
and (n2208,n214,n462);
and (n2209,n218,n455);
or (n2210,n730,n2140);
or (n2211,n2212,n2254);
and (n2212,n2213,n2232);
xor (n2213,n2214,n2215);
xor (n2214,n2179,n2185);
or (n2215,n2216,n2231);
and (n2216,n2217,n2225);
xor (n2217,n2218,n2219);
nor (n2218,n153,n549);
nand (n2219,n2220,n2224);
or (n2220,n2221,n671);
nor (n2221,n2222,n2223);
and (n2222,n386,n624);
and (n2223,n628,n387);
or (n2224,n2181,n672);
nand (n2225,n2226,n2227);
or (n2226,n384,n2107);
or (n2227,n383,n2228);
nor (n2228,n2229,n2230);
and (n2229,n205,n397);
and (n2230,n209,n398);
and (n2231,n2218,n2219);
or (n2232,n2233,n2253);
and (n2233,n2234,n2247);
xor (n2234,n2235,n2241);
nand (n2235,n2236,n2240);
or (n2236,n452,n2237);
nor (n2237,n2238,n2239);
and (n2238,n287,n470);
and (n2239,n291,n466);
or (n2240,n2113,n453);
nand (n2241,n2242,n2243);
or (n2242,n647,n2122);
or (n2243,n635,n2244);
nor (n2244,n2245,n2246);
and (n2245,n646,n327);
and (n2246,n641,n331);
nand (n2247,n2248,n2249);
or (n2248,n681,n2145);
or (n2249,n680,n2250);
nor (n2250,n2251,n2252);
and (n2251,n365,n96);
and (n2252,n369,n92);
and (n2253,n2235,n2241);
and (n2254,n2214,n2215);
or (n2255,n2256,n2305);
and (n2256,n2257,n2260);
xor (n2257,n2258,n2259);
xor (n2258,n2133,n2152);
xor (n2259,n2104,n2120);
or (n2260,n2261,n2304);
and (n2261,n2262,n2282);
xor (n2262,n2263,n2269);
nand (n2263,n2264,n2268);
or (n2264,n730,n2265);
nor (n2265,n2266,n2267);
and (n2266,n244,n462);
and (n2267,n248,n455);
or (n2268,n731,n2136);
and (n2269,n2270,n2276);
nand (n2270,n2271,n2275);
or (n2271,n2272,n671);
nor (n2272,n2273,n2274);
and (n2273,n214,n386);
and (n2274,n218,n387);
or (n2275,n2221,n672);
nor (n2276,n2277,n96);
nor (n2277,n2278,n2281);
and (n2278,n646,n2279);
not (n2279,n2280);
and (n2280,n547,n683);
and (n2281,n687,n549);
or (n2282,n2283,n2303);
and (n2283,n2284,n2297);
xor (n2284,n2285,n2291);
nand (n2285,n2286,n2290);
or (n2286,n383,n2287);
nor (n2287,n2288,n2289);
and (n2288,n252,n397);
and (n2289,n256,n398);
or (n2290,n384,n2228);
nand (n2291,n2292,n2296);
or (n2292,n452,n2293);
nor (n2293,n2294,n2295);
and (n2294,n335,n470);
and (n2295,n339,n466);
or (n2296,n2237,n453);
nand (n2297,n2298,n2302);
or (n2298,n635,n2299);
nor (n2299,n2300,n2301);
and (n2300,n373,n646);
and (n2301,n377,n641);
or (n2302,n2244,n647);
and (n2303,n2285,n2291);
and (n2304,n2263,n2269);
and (n2305,n2258,n2259);
and (n2306,n2079,n2162);
xor (n2307,n2308,n2341);
xor (n2308,n2309,n2338);
xor (n2309,n2310,n2317);
xor (n2310,n2311,n2314);
or (n2311,n2312,n2313);
and (n2312,n2192,n2205);
and (n2313,n2193,n2199);
or (n2314,n2315,n2316);
and (n2315,n2165,n2178);
and (n2316,n2166,n2172);
xor (n2317,n2318,n2331);
xor (n2318,n2319,n2325);
nand (n2319,n2320,n2321);
or (n2320,n635,n2202);
or (n2321,n2322,n647);
nor (n2322,n2323,n2324);
and (n2323,n646,n244);
and (n2324,n641,n248);
nand (n2325,n2326,n2327);
or (n2326,n730,n2207);
or (n2327,n731,n2328);
nor (n2328,n2329,n2330);
and (n2329,n624,n462);
and (n2330,n628,n455);
nand (n2331,n2332,n2337);
or (n2332,n681,n2333);
not (n2333,n2334);
nand (n2334,n2335,n2336);
or (n2335,n291,n92);
or (n2336,n96,n287);
or (n2337,n680,n2169);
or (n2338,n2339,n2340);
and (n2339,n2163,n2211);
and (n2340,n2164,n2191);
xor (n2341,n2342,n2369);
xor (n2342,n2343,n2366);
xor (n2343,n2344,n2360);
xor (n2344,n2345,n2351);
nand (n2345,n2346,n2347);
or (n2346,n383,n2099);
or (n2347,n384,n2348);
nor (n2348,n2349,n2350);
and (n2349,n397,n599);
and (n2350,n603,n398);
nand (n2351,n2352,n2356);
or (n2352,n488,n2353);
nor (n2353,n2354,n2355);
and (n2354,n499,n549);
and (n2355,n498,n547);
or (n2356,n2357,n512);
nor (n2357,n2358,n2359);
and (n2358,n365,n498);
and (n2359,n369,n499);
nand (n2360,n2361,n2365);
or (n2361,n2362,n453);
nor (n2362,n2363,n2364);
and (n2363,n205,n470);
and (n2364,n209,n466);
or (n2365,n452,n2196);
or (n2366,n2367,n2368);
and (n2367,n2080,n2131);
and (n2368,n2081,n2102);
xor (n2369,n2370,n2390);
xor (n2370,n2371,n2377);
nand (n2371,n2372,n2373);
or (n2372,n18,n2175);
or (n2373,n2374,n153);
nor (n2374,n2375,n2376);
and (n2375,n327,n21);
and (n2376,n331,n22);
xor (n2377,n2378,n2384);
nand (n2378,n2379,n2380);
or (n2379,n2090,n671);
or (n2380,n2381,n672);
nor (n2381,n2382,n2383);
and (n2382,n99,n386);
and (n2383,n151,n387);
nor (n2384,n2385,n498);
nor (n2385,n2386,n2389);
and (n2386,n21,n2387);
not (n2387,n2388);
and (n2388,n547,n492);
and (n2389,n503,n549);
or (n2390,n2391,n2392);
and (n2391,n2082,n2093);
and (n2392,n2083,n2084);
or (n2393,n2394,n2802);
and (n2394,n2395,n2426);
xor (n2395,n2396,n2425);
or (n2396,n2397,n2424);
and (n2397,n2398,n2423);
xor (n2398,n2399,n2422);
or (n2399,n2400,n2421);
and (n2400,n2401,n2404);
xor (n2401,n2402,n2403);
xor (n2402,n2217,n2225);
xor (n2403,n2234,n2247);
or (n2404,n2405,n2420);
and (n2405,n2406,n2419);
xor (n2406,n2407,n2413);
nand (n2407,n2408,n2412);
or (n2408,n680,n2409);
nor (n2409,n2410,n2411);
and (n2410,n92,n549);
and (n2411,n96,n547);
or (n2412,n2250,n681);
nand (n2413,n2414,n2418);
or (n2414,n730,n2415);
nor (n2415,n2416,n2417);
and (n2416,n295,n462);
and (n2417,n299,n455);
or (n2418,n2265,n731);
xor (n2419,n2270,n2276);
and (n2420,n2407,n2413);
and (n2421,n2402,n2403);
xor (n2422,n2213,n2232);
xor (n2423,n2257,n2260);
and (n2424,n2399,n2422);
xor (n2425,n2078,n2255);
nand (n2426,n2427,n2799,n2801);
or (n2427,n2428,n2794);
nand (n2428,n2429,n2783);
or (n2429,n2430,n2782);
and (n2430,n2431,n2552);
xor (n2431,n2432,n2537);
or (n2432,n2433,n2536);
and (n2433,n2434,n2502);
xor (n2434,n2435,n2457);
xor (n2435,n2436,n2451);
xor (n2436,n2437,n2444);
nand (n2437,n2438,n2443);
or (n2438,n452,n2439);
not (n2439,n2440);
nor (n2440,n2441,n2442);
and (n2441,n470,n331);
and (n2442,n327,n466);
or (n2443,n2293,n453);
nand (n2444,n2445,n2450);
or (n2445,n2446,n635);
not (n2446,n2447);
nand (n2447,n2448,n2449);
or (n2448,n369,n641);
or (n2449,n365,n646);
or (n2450,n2299,n647);
nand (n2451,n2452,n2456);
or (n2452,n730,n2453);
nor (n2453,n2454,n2455);
and (n2454,n287,n462);
and (n2455,n291,n455);
or (n2456,n731,n2415);
or (n2457,n2458,n2501);
and (n2458,n2459,n2481);
xor (n2459,n2460,n2466);
nand (n2460,n2461,n2465);
or (n2461,n730,n2462);
nor (n2462,n2463,n2464);
and (n2463,n335,n462);
and (n2464,n339,n455);
or (n2465,n2453,n731);
xor (n2466,n2467,n2473);
nor (n2467,n2468,n646);
nor (n2468,n2469,n2472);
and (n2469,n2470,n470);
not (n2470,n2471);
and (n2471,n547,n638);
and (n2472,n645,n549);
nand (n2473,n2474,n2477);
or (n2474,n671,n2475);
not (n2475,n2476);
xnor (n2476,n252,n386);
or (n2477,n2478,n672);
nor (n2478,n2479,n2480);
and (n2479,n386,n205);
and (n2480,n209,n387);
or (n2481,n2482,n2500);
and (n2482,n2483,n2491);
xor (n2483,n2484,n2485);
nor (n2484,n647,n549);
nand (n2485,n2486,n2487);
or (n2486,n672,n2475);
or (n2487,n2488,n671);
nor (n2488,n2489,n2490);
and (n2489,n386,n244);
and (n2490,n248,n387);
nand (n2491,n2492,n2496);
or (n2492,n452,n2493);
nor (n2493,n2494,n2495);
and (n2494,n365,n470);
and (n2495,n369,n466);
or (n2496,n2497,n453);
nor (n2497,n2498,n2499);
and (n2498,n373,n470);
and (n2499,n377,n466);
and (n2500,n2484,n2485);
and (n2501,n2460,n2466);
xor (n2502,n2503,n2517);
xor (n2503,n2504,n2505);
and (n2504,n2467,n2473);
xor (n2505,n2506,n2511);
xor (n2506,n2507,n2508);
nor (n2507,n681,n549);
nand (n2508,n2509,n2510);
or (n2509,n2478,n671);
or (n2510,n2272,n672);
nand (n2511,n2512,n2516);
or (n2512,n383,n2513);
nor (n2513,n2514,n2515);
and (n2514,n244,n397);
and (n2515,n248,n398);
or (n2516,n384,n2287);
or (n2517,n2518,n2535);
and (n2518,n2519,n2529);
xor (n2519,n2520,n2526);
nand (n2520,n2521,n2525);
or (n2521,n383,n2522);
nor (n2522,n2523,n2524);
and (n2523,n397,n295);
and (n2524,n299,n398);
or (n2525,n2513,n384);
nand (n2526,n2527,n2528);
or (n2527,n453,n2439);
or (n2528,n2497,n452);
nand (n2529,n2530,n2531);
or (n2530,n647,n2446);
or (n2531,n635,n2532);
nor (n2532,n2533,n2534);
and (n2533,n641,n549);
and (n2534,n646,n547);
and (n2535,n2520,n2526);
and (n2536,n2435,n2457);
xor (n2537,n2538,n2543);
xor (n2538,n2539,n2540);
xor (n2539,n2284,n2297);
or (n2540,n2541,n2542);
and (n2541,n2503,n2517);
and (n2542,n2504,n2505);
xor (n2543,n2544,n2551);
xor (n2544,n2545,n2548);
or (n2545,n2546,n2547);
and (n2546,n2506,n2511);
and (n2547,n2507,n2508);
or (n2548,n2549,n2550);
and (n2549,n2436,n2451);
and (n2550,n2437,n2444);
xor (n2551,n2406,n2419);
or (n2552,n2553,n2781);
and (n2553,n2554,n2591);
xor (n2554,n2555,n2590);
or (n2555,n2556,n2589);
and (n2556,n2557,n2588);
xor (n2557,n2558,n2587);
or (n2558,n2559,n2586);
and (n2559,n2560,n2573);
xor (n2560,n2561,n2567);
nand (n2561,n2562,n2566);
or (n2562,n383,n2563);
nor (n2563,n2564,n2565);
and (n2564,n287,n397);
and (n2565,n398,n291);
or (n2566,n2522,n384);
nand (n2567,n2568,n2572);
or (n2568,n730,n2569);
nor (n2569,n2570,n2571);
and (n2570,n327,n462);
and (n2571,n331,n455);
or (n2572,n2462,n731);
and (n2573,n2574,n2580);
nor (n2574,n2575,n470);
nor (n2575,n2576,n2579);
and (n2576,n2577,n462);
not (n2577,n2578);
and (n2578,n547,n458);
and (n2579,n463,n549);
nand (n2580,n2581,n2585);
or (n2581,n2582,n671);
nor (n2582,n2583,n2584);
and (n2583,n386,n295);
and (n2584,n299,n387);
or (n2585,n2488,n672);
and (n2586,n2561,n2567);
xor (n2587,n2519,n2529);
xor (n2588,n2459,n2481);
and (n2589,n2558,n2587);
xor (n2590,n2434,n2502);
nand (n2591,n2592,n2778,n2780);
or (n2592,n2593,n2651);
nand (n2593,n2594,n2646);
not (n2594,n2595);
nor (n2595,n2596,n2622);
xor (n2596,n2597,n2621);
xor (n2597,n2598,n2620);
or (n2598,n2599,n2619);
and (n2599,n2600,n2613);
xor (n2600,n2601,n2607);
nand (n2601,n2602,n2606);
or (n2602,n452,n2603);
nor (n2603,n2604,n2605);
and (n2604,n466,n549);
and (n2605,n470,n547);
or (n2606,n2493,n453);
nand (n2607,n2608,n2612);
or (n2608,n2609,n383);
nor (n2609,n2610,n2611);
and (n2610,n398,n339);
and (n2611,n397,n335);
or (n2612,n2563,n384);
nand (n2613,n2614,n2618);
or (n2614,n730,n2615);
nor (n2615,n2616,n2617);
and (n2616,n373,n462);
and (n2617,n377,n455);
or (n2618,n2569,n731);
and (n2619,n2601,n2607);
xor (n2620,n2483,n2491);
xor (n2621,n2560,n2573);
or (n2622,n2623,n2645);
and (n2623,n2624,n2644);
xor (n2624,n2625,n2626);
xor (n2625,n2574,n2580);
or (n2626,n2627,n2643);
and (n2627,n2628,n2637);
xor (n2628,n2629,n2630);
nor (n2629,n453,n549);
nand (n2630,n2631,n2636);
or (n2631,n2632,n671);
not (n2632,n2633);
nand (n2633,n2634,n2635);
or (n2634,n387,n291);
nand (n2635,n291,n387);
or (n2636,n2582,n672);
nand (n2637,n2638,n2642);
or (n2638,n383,n2639);
nor (n2639,n2640,n2641);
and (n2640,n397,n327);
and (n2641,n398,n331);
or (n2642,n2609,n384);
and (n2643,n2629,n2630);
xor (n2644,n2600,n2613);
and (n2645,n2625,n2626);
or (n2646,n2647,n2648);
xor (n2647,n2557,n2588);
or (n2648,n2649,n2650);
and (n2649,n2597,n2621);
and (n2650,n2598,n2620);
nor (n2651,n2652,n2777);
and (n2652,n2653,n2772);
or (n2653,n2654,n2771);
and (n2654,n2655,n2696);
xor (n2655,n2656,n2689);
or (n2656,n2657,n2688);
and (n2657,n2658,n2674);
xor (n2658,n2659,n2665);
nand (n2659,n2660,n2664);
or (n2660,n383,n2661);
nor (n2661,n2662,n2663);
and (n2662,n398,n377);
and (n2663,n397,n373);
or (n2664,n2639,n384);
or (n2665,n2666,n2670);
nor (n2666,n2667,n731);
nor (n2667,n2668,n2669);
and (n2668,n462,n365);
and (n2669,n455,n369);
nor (n2670,n730,n2671);
nor (n2671,n2672,n2673);
and (n2672,n455,n549);
and (n2673,n462,n547);
xor (n2674,n2675,n2681);
nor (n2675,n2676,n462);
nor (n2676,n2677,n2680);
and (n2677,n2678,n397);
not (n2678,n2679);
and (n2679,n547,n734);
and (n2680,n740,n549);
nand (n2681,n2682,n2687);
or (n2682,n671,n2683);
not (n2683,n2684);
nand (n2684,n2685,n2686);
or (n2685,n386,n335);
nand (n2686,n335,n386);
nand (n2687,n2633,n673);
and (n2688,n2659,n2665);
xor (n2689,n2690,n2695);
xor (n2690,n2691,n2694);
nand (n2691,n2692,n2693);
or (n2692,n730,n2667);
or (n2693,n2615,n731);
and (n2694,n2675,n2681);
xor (n2695,n2628,n2637);
or (n2696,n2697,n2770);
and (n2697,n2698,n2718);
xor (n2698,n2699,n2717);
or (n2699,n2700,n2716);
and (n2700,n2701,n2710);
xor (n2701,n2702,n2703);
and (n2702,n732,n547);
nand (n2703,n2704,n2709);
or (n2704,n671,n2705);
not (n2705,n2706);
nand (n2706,n2707,n2708);
or (n2707,n387,n331);
nand (n2708,n331,n387);
nand (n2709,n2684,n673);
nand (n2710,n2711,n2715);
or (n2711,n383,n2712);
nor (n2712,n2713,n2714);
and (n2713,n397,n365);
and (n2714,n398,n369);
or (n2715,n2661,n384);
and (n2716,n2702,n2703);
xor (n2717,n2658,n2674);
or (n2718,n2719,n2769);
and (n2719,n2720,n2737);
xor (n2720,n2721,n2736);
and (n2721,n2722,n2728);
and (n2722,n2723,n398);
nand (n2723,n2724,n2727);
nand (n2724,n2725,n386);
not (n2725,n2726);
and (n2726,n547,n390);
nand (n2727,n394,n549);
nand (n2728,n2729,n2730);
or (n2729,n672,n2705);
nand (n2730,n2731,n2735);
not (n2731,n2732);
nor (n2732,n2733,n2734);
and (n2733,n377,n387);
and (n2734,n373,n386);
not (n2735,n671);
xor (n2736,n2701,n2710);
or (n2737,n2738,n2768);
and (n2738,n2739,n2747);
xor (n2739,n2740,n2746);
nand (n2740,n2741,n2745);
or (n2741,n383,n2742);
nor (n2742,n2743,n2744);
and (n2743,n398,n549);
and (n2744,n397,n547);
or (n2745,n2712,n384);
xor (n2746,n2722,n2728);
or (n2747,n2748,n2767);
and (n2748,n2749,n2757);
xor (n2749,n2750,n2751);
nor (n2750,n384,n549);
nand (n2751,n2752,n2756);
or (n2752,n2753,n671);
or (n2753,n2754,n2755);
and (n2754,n386,n369);
and (n2755,n365,n387);
or (n2756,n2732,n672);
nor (n2757,n2758,n2765);
nor (n2758,n2759,n2761);
and (n2759,n2760,n673);
not (n2760,n2753);
and (n2761,n2762,n2735);
nand (n2762,n2763,n2764);
or (n2763,n386,n547);
or (n2764,n387,n549);
or (n2765,n386,n2766);
and (n2766,n547,n673);
and (n2767,n2750,n2751);
and (n2768,n2740,n2746);
and (n2769,n2721,n2736);
and (n2770,n2699,n2717);
and (n2771,n2656,n2689);
or (n2772,n2773,n2774);
xor (n2773,n2624,n2644);
or (n2774,n2775,n2776);
and (n2775,n2690,n2695);
and (n2776,n2691,n2694);
and (n2777,n2773,n2774);
nand (n2778,n2646,n2779);
and (n2779,n2596,n2622);
nand (n2780,n2647,n2648);
and (n2781,n2555,n2590);
and (n2782,n2432,n2537);
or (n2783,n2784,n2791);
xor (n2784,n2785,n2790);
xor (n2785,n2786,n2787);
xor (n2786,n2262,n2282);
or (n2787,n2788,n2789);
and (n2788,n2544,n2551);
and (n2789,n2545,n2548);
xor (n2790,n2401,n2404);
or (n2791,n2792,n2793);
and (n2792,n2538,n2543);
and (n2793,n2539,n2540);
nor (n2794,n2795,n2796);
xor (n2795,n2398,n2423);
or (n2796,n2797,n2798);
and (n2797,n2785,n2790);
and (n2798,n2786,n2787);
or (n2799,n2794,n2800);
nand (n2800,n2784,n2791);
nand (n2801,n2795,n2796);
and (n2802,n2396,n2425);
and (n2803,n2076,n2307);
nor (n2804,n2805,n2925);
nor (n2805,n2806,n2916);
xor (n2806,n2807,n2871);
xor (n2807,n2808,n2846);
xor (n2808,n2809,n2831);
xor (n2809,n2810,n2811);
xor (n2810,n2013,n2026);
xor (n2811,n2812,n2825);
xor (n2812,n2813,n2819);
nand (n2813,n2814,n2818);
or (n2814,n383,n2815);
nor (n2815,n2816,n2817);
and (n2816,n397,n506);
and (n2817,n510,n398);
or (n2818,n384,n1945);
nand (n2819,n2820,n2824);
or (n2820,n635,n2821);
nor (n2821,n2822,n2823);
and (n2822,n646,n252);
and (n2823,n641,n256);
or (n2824,n1964,n647);
nand (n2825,n2826,n2830);
or (n2826,n2827,n730);
nor (n2827,n2828,n2829);
and (n2828,n591,n462);
and (n2829,n595,n455);
or (n2830,n731,n1970);
xor (n2831,n2832,n2845);
xor (n2832,n2833,n2839);
nand (n2833,n2834,n2838);
or (n2834,n680,n2835);
nor (n2835,n2836,n2837);
and (n2836,n96,n295);
and (n2837,n92,n299);
or (n2838,n1976,n681);
nand (n2839,n2840,n2844);
or (n2840,n18,n2841);
nor (n2841,n2842,n2843);
and (n2842,n21,n335);
and (n2843,n339,n22);
or (n2844,n153,n1994);
xor (n2845,n1999,n2005);
or (n2846,n2847,n2870);
and (n2847,n2848,n2855);
xor (n2848,n2849,n2852);
or (n2849,n2850,n2851);
and (n2850,n2370,n2390);
and (n2851,n2371,n2377);
or (n2852,n2853,n2854);
and (n2853,n2310,n2317);
and (n2854,n2311,n2314);
xor (n2855,n2856,n2867);
xor (n2856,n2857,n2858);
and (n2857,n2378,n2384);
xor (n2858,n2859,n2864);
xor (n2859,n2860,n2861);
nor (n2860,n608,n549);
nand (n2861,n2862,n2863);
or (n2862,n2381,n671);
or (n2863,n2007,n672);
nand (n2864,n2865,n2866);
or (n2865,n383,n2348);
or (n2866,n384,n2815);
or (n2867,n2868,n2869);
and (n2868,n2344,n2360);
and (n2869,n2345,n2351);
and (n2870,n2849,n2852);
xor (n2871,n2872,n2907);
xor (n2872,n2873,n2876);
or (n2873,n2874,n2875);
and (n2874,n2856,n2867);
and (n2875,n2857,n2858);
xor (n2876,n2877,n2894);
xor (n2877,n2878,n2881);
or (n2878,n2879,n2880);
and (n2879,n2859,n2864);
and (n2880,n2860,n2861);
or (n2881,n2882,n2893);
and (n2882,n2883,n2890);
xor (n2883,n2884,n2887);
nand (n2884,n2885,n2886);
or (n2885,n730,n2328);
or (n2886,n731,n2827);
nand (n2887,n2888,n2889);
or (n2888,n2333,n680);
or (n2889,n2835,n681);
nand (n2890,n2891,n2892);
or (n2891,n18,n2374);
or (n2892,n2841,n153);
and (n2893,n2884,n2887);
or (n2894,n2895,n2906);
and (n2895,n2896,n2903);
xor (n2896,n2897,n2900);
nand (n2897,n2898,n2899);
or (n2898,n488,n2357);
or (n2899,n2022,n512);
nand (n2900,n2901,n2902);
or (n2901,n452,n2362);
or (n2902,n2016,n453);
nand (n2903,n2904,n2905);
or (n2904,n635,n2322);
or (n2905,n2821,n647);
and (n2906,n2897,n2900);
or (n2907,n2908,n2915);
and (n2908,n2909,n2914);
xor (n2909,n2910,n2913);
or (n2910,n2911,n2912);
and (n2911,n2318,n2331);
and (n2912,n2319,n2325);
xor (n2913,n2883,n2890);
xor (n2914,n2896,n2903);
and (n2915,n2910,n2913);
or (n2916,n2917,n2924);
and (n2917,n2918,n2923);
xor (n2918,n2919,n2920);
xor (n2919,n2909,n2914);
or (n2920,n2921,n2922);
and (n2921,n2342,n2369);
and (n2922,n2343,n2366);
xor (n2923,n2848,n2855);
and (n2924,n2919,n2920);
nor (n2925,n2926,n2927);
xor (n2926,n2918,n2923);
or (n2927,n2928,n2929);
and (n2928,n2308,n2341);
and (n2929,n2309,n2338);
or (n2930,n2931,n2976);
nor (n2931,n2932,n2967);
xor (n2932,n2933,n2952);
xor (n2933,n2934,n2935);
xor (n2934,n1987,n2035);
or (n2935,n2936,n2951);
and (n2936,n2937,n2944);
xor (n2937,n2938,n2941);
or (n2938,n2939,n2940);
and (n2939,n2877,n2894);
and (n2940,n2878,n2881);
or (n2941,n2942,n2943);
and (n2942,n2809,n2831);
and (n2943,n2810,n2811);
xor (n2944,n2945,n2950);
xor (n2945,n2946,n2949);
or (n2946,n2947,n2948);
and (n2947,n2812,n2825);
and (n2948,n2813,n2819);
xor (n2949,n1961,n1974);
xor (n2950,n1913,n1921);
and (n2951,n2938,n2941);
xor (n2952,n2953,n2958);
xor (n2953,n2954,n2957);
or (n2954,n2955,n2956);
and (n2955,n2945,n2950);
and (n2956,n2946,n2949);
xor (n2957,n1958,n1982);
or (n2958,n2959,n2966);
and (n2959,n2960,n2965);
xor (n2960,n2961,n2962);
xor (n2961,n1930,n1943);
or (n2962,n2963,n2964);
and (n2963,n2832,n2845);
and (n2964,n2833,n2839);
xor (n2965,n1991,n2011);
and (n2966,n2961,n2962);
or (n2967,n2968,n2975);
and (n2968,n2969,n2974);
xor (n2969,n2970,n2971);
xor (n2970,n2960,n2965);
or (n2971,n2972,n2973);
and (n2972,n2872,n2907);
and (n2973,n2873,n2876);
xor (n2974,n2937,n2944);
and (n2975,n2970,n2971);
nor (n2976,n2977,n2980);
or (n2977,n2978,n2979);
and (n2978,n2807,n2871);
and (n2979,n2808,n2846);
xor (n2980,n2969,n2974);
nand (n2981,n2982,n2991);
or (n2982,n2983,n2931);
nor (n2983,n2984,n2990);
and (n2984,n2985,n2989);
nand (n2985,n2986,n2988);
or (n2986,n2805,n2987);
nand (n2987,n2926,n2927);
nand (n2988,n2806,n2916);
not (n2989,n2976);
and (n2990,n2977,n2980);
nand (n2991,n2932,n2967);
or (n2992,n2993,n3000);
xor (n2993,n2994,n2999);
xor (n2994,n2995,n2996);
xor (n2995,n1905,n1951);
or (n2996,n2997,n2998);
and (n2997,n2953,n2958);
and (n2998,n2954,n2957);
xor (n2999,n1955,n1985);
or (n3000,n3001,n3002);
and (n3001,n2933,n2952);
and (n3002,n2934,n2935);
and (n3003,n3004,n3006);
not (n3004,n3005);
xor (n3005,n1715,n1953);
not (n3006,n3007);
or (n3007,n3008,n3009);
and (n3008,n2994,n2999);
and (n3009,n2995,n2996);
nor (n3010,n3011,n3015);
and (n3011,n3012,n3013);
not (n3012,n3003);
not (n3013,n3014);
nand (n3014,n2993,n3000);
nor (n3015,n3004,n3006);
and (n3016,n1713,n2039);
nand (n3017,n3018,n3022);
not (n3018,n3019);
or (n3019,n3020,n3021);
and (n3020,n2040,n2063);
and (n3021,n2041,n2050);
not (n3022,n3023);
xor (n3023,n3024,n3029);
xor (n3024,n3025,n3026);
xor (n3025,n1585,n1621);
or (n3026,n3027,n3028);
and (n3027,n2051,n2060);
and (n3028,n2052,n2053);
xor (n3029,n3030,n3035);
xor (n3030,n3031,n3032);
xor (n3031,n1369,n1420);
or (n3032,n3033,n3034);
and (n3033,n2054,n2057);
and (n3034,n2055,n2056);
or (n3035,n3036,n3037);
and (n3036,n2042,n2047);
and (n3037,n2043,n2044);
nor (n3038,n3022,n3018);
and (n3039,n3040,n3050);
not (n3040,n3041);
or (n3041,n3042,n3049);
and (n3042,n3043,n3046);
xor (n3043,n3044,n3045);
xor (n3044,n1683,n1688);
xor (n3045,n1366,n1583);
or (n3046,n3047,n3048);
and (n3047,n3030,n3035);
and (n3048,n3031,n3032);
and (n3049,n3044,n3045);
not (n3050,n3051);
xor (n3051,n1352,n1659);
nor (n3052,n3053,n3054);
xor (n3053,n3043,n3046);
or (n3054,n3055,n3056);
and (n3055,n3024,n3029);
and (n3056,n3025,n3026);
nor (n3057,n3058,n3062);
and (n3058,n3059,n3060);
not (n3059,n3039);
not (n3060,n3061);
nand (n3061,n3053,n3054);
nor (n3062,n3040,n3050);
and (n3063,n1350,n1691);
nand (n3064,n3065,n3073);
not (n3065,n3066);
xor (n3066,n3067,n3072);
xor (n3067,n3068,n3069);
xor (n3068,n938,n979);
or (n3069,n3070,n3071);
and (n3070,n1698,n1705);
and (n3071,n1699,n1702);
xor (n3072,n1226,n1326);
not (n3073,n3074);
or (n3074,n3075,n3076);
and (n3075,n1692,n1697);
and (n3076,n1693,n1694);
nor (n3077,n3065,n3073);
nor (n3078,n3079,n3080);
xor (n3079,n1221,n1224);
or (n3080,n3081,n3082);
and (n3081,n3067,n3072);
and (n3082,n3068,n3069);
and (n3083,n3079,n3080);
or (n3084,n1343,n3);
xor (n3085,n3086,n5507);
xor (n3086,n3087,n5505);
xor (n3087,n3088,n5504);
xor (n3088,n3089,n5495);
xor (n3089,n3090,n5494);
xor (n3090,n3091,n5480);
xor (n3091,n3092,n5479);
xor (n3092,n3093,n5458);
xor (n3093,n3094,n5457);
xor (n3094,n3095,n5431);
xor (n3095,n3096,n5430);
xor (n3096,n3097,n5397);
xor (n3097,n3098,n5396);
xor (n3098,n3099,n5358);
xor (n3099,n3100,n5357);
xor (n3100,n3101,n5312);
xor (n3101,n3102,n5311);
xor (n3102,n3103,n5261);
xor (n3103,n3104,n5260);
xor (n3104,n3105,n5203);
xor (n3105,n3106,n5202);
xor (n3106,n3107,n5140);
xor (n3107,n3108,n5139);
xor (n3108,n3109,n5070);
xor (n3109,n3110,n5069);
xor (n3110,n3111,n4995);
xor (n3111,n3112,n4994);
xor (n3112,n3113,n4913);
xor (n3113,n3114,n4912);
xor (n3114,n3115,n4826);
xor (n3115,n3116,n4825);
xor (n3116,n3117,n4732);
xor (n3117,n3118,n4731);
xor (n3118,n3119,n4633);
xor (n3119,n3120,n4632);
xor (n3120,n3121,n4527);
xor (n3121,n3122,n4526);
xor (n3122,n3123,n4416);
xor (n3123,n3124,n4415);
xor (n3124,n3125,n4298);
xor (n3125,n3126,n4297);
xor (n3126,n3127,n4175);
xor (n3127,n3128,n4174);
xor (n3128,n3129,n4046);
xor (n3129,n3130,n4045);
xor (n3130,n3131,n3911);
xor (n3131,n3132,n3910);
xor (n3132,n3133,n3769);
xor (n3133,n3134,n3768);
xor (n3134,n3135,n3622);
xor (n3135,n3136,n3621);
xor (n3136,n3137,n3468);
xor (n3137,n3138,n3467);
xor (n3138,n3139,n3309);
xor (n3139,n3140,n3308);
xor (n3140,n3141,n3144);
xor (n3141,n3142,n3143);
and (n3142,n1099,n673);
and (n3143,n714,n387);
or (n3144,n3145,n3148);
and (n3145,n3146,n3147);
and (n3146,n714,n673);
and (n3147,n442,n387);
and (n3148,n3149,n3150);
xor (n3149,n3146,n3147);
or (n3150,n3151,n3154);
and (n3151,n3152,n3153);
and (n3152,n442,n673);
and (n3153,n404,n387);
and (n3154,n3155,n3156);
xor (n3155,n3152,n3153);
or (n3156,n3157,n3160);
and (n3157,n3158,n3159);
and (n3158,n404,n673);
and (n3159,n562,n387);
and (n3160,n3161,n3162);
xor (n3161,n3158,n3159);
or (n3162,n3163,n3166);
and (n3163,n3164,n3165);
and (n3164,n562,n673);
and (n3165,n554,n387);
and (n3166,n3167,n3168);
xor (n3167,n3164,n3165);
or (n3168,n3169,n3172);
and (n3169,n3170,n3171);
and (n3170,n554,n673);
and (n3171,n481,n387);
and (n3172,n3173,n3174);
xor (n3173,n3170,n3171);
or (n3174,n3175,n3178);
and (n3175,n3176,n3177);
and (n3176,n481,n673);
and (n3177,n473,n387);
and (n3178,n3179,n3180);
xor (n3179,n3176,n3177);
or (n3180,n3181,n3184);
and (n3181,n3182,n3183);
and (n3182,n473,n673);
and (n3183,n582,n387);
and (n3184,n3185,n3186);
xor (n3185,n3182,n3183);
or (n3186,n3187,n3190);
and (n3187,n3188,n3189);
and (n3188,n582,n673);
and (n3189,n574,n387);
and (n3190,n3191,n3192);
xor (n3191,n3188,n3189);
or (n3192,n3193,n3196);
and (n3193,n3194,n3195);
and (n3194,n574,n673);
and (n3195,n661,n387);
and (n3196,n3197,n3198);
xor (n3197,n3194,n3195);
or (n3198,n3199,n3202);
and (n3199,n3200,n3201);
and (n3200,n661,n673);
and (n3201,n653,n387);
and (n3202,n3203,n3204);
xor (n3203,n3200,n3201);
or (n3204,n3205,n3208);
and (n3205,n3206,n3207);
and (n3206,n653,n673);
and (n3207,n697,n387);
and (n3208,n3209,n3210);
xor (n3209,n3206,n3207);
or (n3210,n3211,n3214);
and (n3211,n3212,n3213);
and (n3212,n697,n673);
and (n3213,n156,n387);
and (n3214,n3215,n3216);
xor (n3215,n3212,n3213);
or (n3216,n3217,n3220);
and (n3217,n3218,n3219);
and (n3218,n156,n673);
and (n3219,n99,n387);
and (n3220,n3221,n3222);
xor (n3221,n3218,n3219);
or (n3222,n3223,n3226);
and (n3223,n3224,n3225);
and (n3224,n99,n673);
and (n3225,n506,n387);
and (n3226,n3227,n3228);
xor (n3227,n3224,n3225);
or (n3228,n3229,n3232);
and (n3229,n3230,n3231);
and (n3230,n506,n673);
and (n3231,n599,n387);
and (n3232,n3233,n3234);
xor (n3233,n3230,n3231);
or (n3234,n3235,n3238);
and (n3235,n3236,n3237);
and (n3236,n599,n673);
and (n3237,n591,n387);
and (n3238,n3239,n3240);
xor (n3239,n3236,n3237);
or (n3240,n3241,n3244);
and (n3241,n3242,n3243);
and (n3242,n591,n673);
and (n3243,n624,n387);
and (n3244,n3245,n3246);
xor (n3245,n3242,n3243);
or (n3246,n3247,n3250);
and (n3247,n3248,n3249);
and (n3248,n624,n673);
and (n3249,n214,n387);
and (n3250,n3251,n3252);
xor (n3251,n3248,n3249);
or (n3252,n3253,n3256);
and (n3253,n3254,n3255);
and (n3254,n214,n673);
and (n3255,n205,n387);
and (n3256,n3257,n3258);
xor (n3257,n3254,n3255);
or (n3258,n3259,n3262);
and (n3259,n3260,n3261);
and (n3260,n205,n673);
and (n3261,n252,n387);
and (n3262,n3263,n3264);
xor (n3263,n3260,n3261);
or (n3264,n3265,n3268);
and (n3265,n3266,n3267);
and (n3266,n252,n673);
and (n3267,n244,n387);
and (n3268,n3269,n3270);
xor (n3269,n3266,n3267);
or (n3270,n3271,n3274);
and (n3271,n3272,n3273);
and (n3272,n244,n673);
and (n3273,n295,n387);
and (n3274,n3275,n3276);
xor (n3275,n3272,n3273);
or (n3276,n3277,n3280);
and (n3277,n3278,n3279);
and (n3278,n295,n673);
and (n3279,n287,n387);
and (n3280,n3281,n3282);
xor (n3281,n3278,n3279);
or (n3282,n3283,n3286);
and (n3283,n3284,n3285);
and (n3284,n287,n673);
and (n3285,n335,n387);
and (n3286,n3287,n3288);
xor (n3287,n3284,n3285);
or (n3288,n3289,n3292);
and (n3289,n3290,n3291);
and (n3290,n335,n673);
and (n3291,n327,n387);
and (n3292,n3293,n3294);
xor (n3293,n3290,n3291);
or (n3294,n3295,n3298);
and (n3295,n3296,n3297);
and (n3296,n327,n673);
and (n3297,n373,n387);
and (n3298,n3299,n3300);
xor (n3299,n3296,n3297);
or (n3300,n3301,n3303);
and (n3301,n3302,n2755);
and (n3302,n373,n673);
and (n3303,n3304,n3305);
xor (n3304,n3302,n2755);
and (n3305,n3306,n3307);
and (n3306,n365,n673);
and (n3307,n547,n387);
and (n3308,n442,n390);
or (n3309,n3310,n3313);
and (n3310,n3311,n3312);
xor (n3311,n3149,n3150);
and (n3312,n404,n390);
and (n3313,n3314,n3315);
xor (n3314,n3311,n3312);
or (n3315,n3316,n3319);
and (n3316,n3317,n3318);
xor (n3317,n3155,n3156);
and (n3318,n562,n390);
and (n3319,n3320,n3321);
xor (n3320,n3317,n3318);
or (n3321,n3322,n3325);
and (n3322,n3323,n3324);
xor (n3323,n3161,n3162);
and (n3324,n554,n390);
and (n3325,n3326,n3327);
xor (n3326,n3323,n3324);
or (n3327,n3328,n3331);
and (n3328,n3329,n3330);
xor (n3329,n3167,n3168);
and (n3330,n481,n390);
and (n3331,n3332,n3333);
xor (n3332,n3329,n3330);
or (n3333,n3334,n3337);
and (n3334,n3335,n3336);
xor (n3335,n3173,n3174);
and (n3336,n473,n390);
and (n3337,n3338,n3339);
xor (n3338,n3335,n3336);
or (n3339,n3340,n3343);
and (n3340,n3341,n3342);
xor (n3341,n3179,n3180);
and (n3342,n582,n390);
and (n3343,n3344,n3345);
xor (n3344,n3341,n3342);
or (n3345,n3346,n3349);
and (n3346,n3347,n3348);
xor (n3347,n3185,n3186);
and (n3348,n574,n390);
and (n3349,n3350,n3351);
xor (n3350,n3347,n3348);
or (n3351,n3352,n3355);
and (n3352,n3353,n3354);
xor (n3353,n3191,n3192);
and (n3354,n661,n390);
and (n3355,n3356,n3357);
xor (n3356,n3353,n3354);
or (n3357,n3358,n3361);
and (n3358,n3359,n3360);
xor (n3359,n3197,n3198);
and (n3360,n653,n390);
and (n3361,n3362,n3363);
xor (n3362,n3359,n3360);
or (n3363,n3364,n3367);
and (n3364,n3365,n3366);
xor (n3365,n3203,n3204);
and (n3366,n697,n390);
and (n3367,n3368,n3369);
xor (n3368,n3365,n3366);
or (n3369,n3370,n3373);
and (n3370,n3371,n3372);
xor (n3371,n3209,n3210);
and (n3372,n156,n390);
and (n3373,n3374,n3375);
xor (n3374,n3371,n3372);
or (n3375,n3376,n3379);
and (n3376,n3377,n3378);
xor (n3377,n3215,n3216);
and (n3378,n99,n390);
and (n3379,n3380,n3381);
xor (n3380,n3377,n3378);
or (n3381,n3382,n3385);
and (n3382,n3383,n3384);
xor (n3383,n3221,n3222);
and (n3384,n506,n390);
and (n3385,n3386,n3387);
xor (n3386,n3383,n3384);
or (n3387,n3388,n3391);
and (n3388,n3389,n3390);
xor (n3389,n3227,n3228);
and (n3390,n599,n390);
and (n3391,n3392,n3393);
xor (n3392,n3389,n3390);
or (n3393,n3394,n3397);
and (n3394,n3395,n3396);
xor (n3395,n3233,n3234);
and (n3396,n591,n390);
and (n3397,n3398,n3399);
xor (n3398,n3395,n3396);
or (n3399,n3400,n3403);
and (n3400,n3401,n3402);
xor (n3401,n3239,n3240);
and (n3402,n624,n390);
and (n3403,n3404,n3405);
xor (n3404,n3401,n3402);
or (n3405,n3406,n3409);
and (n3406,n3407,n3408);
xor (n3407,n3245,n3246);
and (n3408,n214,n390);
and (n3409,n3410,n3411);
xor (n3410,n3407,n3408);
or (n3411,n3412,n3415);
and (n3412,n3413,n3414);
xor (n3413,n3251,n3252);
and (n3414,n205,n390);
and (n3415,n3416,n3417);
xor (n3416,n3413,n3414);
or (n3417,n3418,n3421);
and (n3418,n3419,n3420);
xor (n3419,n3257,n3258);
and (n3420,n252,n390);
and (n3421,n3422,n3423);
xor (n3422,n3419,n3420);
or (n3423,n3424,n3427);
and (n3424,n3425,n3426);
xor (n3425,n3263,n3264);
and (n3426,n244,n390);
and (n3427,n3428,n3429);
xor (n3428,n3425,n3426);
or (n3429,n3430,n3433);
and (n3430,n3431,n3432);
xor (n3431,n3269,n3270);
and (n3432,n295,n390);
and (n3433,n3434,n3435);
xor (n3434,n3431,n3432);
or (n3435,n3436,n3439);
and (n3436,n3437,n3438);
xor (n3437,n3275,n3276);
and (n3438,n287,n390);
and (n3439,n3440,n3441);
xor (n3440,n3437,n3438);
or (n3441,n3442,n3445);
and (n3442,n3443,n3444);
xor (n3443,n3281,n3282);
and (n3444,n335,n390);
and (n3445,n3446,n3447);
xor (n3446,n3443,n3444);
or (n3447,n3448,n3451);
and (n3448,n3449,n3450);
xor (n3449,n3287,n3288);
and (n3450,n327,n390);
and (n3451,n3452,n3453);
xor (n3452,n3449,n3450);
or (n3453,n3454,n3457);
and (n3454,n3455,n3456);
xor (n3455,n3293,n3294);
and (n3456,n373,n390);
and (n3457,n3458,n3459);
xor (n3458,n3455,n3456);
or (n3459,n3460,n3463);
and (n3460,n3461,n3462);
xor (n3461,n3299,n3300);
and (n3462,n365,n390);
and (n3463,n3464,n3465);
xor (n3464,n3461,n3462);
and (n3465,n3466,n2726);
xor (n3466,n3304,n3305);
and (n3467,n404,n398);
or (n3468,n3469,n3472);
and (n3469,n3470,n3471);
xor (n3470,n3314,n3315);
and (n3471,n562,n398);
and (n3472,n3473,n3474);
xor (n3473,n3470,n3471);
or (n3474,n3475,n3478);
and (n3475,n3476,n3477);
xor (n3476,n3320,n3321);
and (n3477,n554,n398);
and (n3478,n3479,n3480);
xor (n3479,n3476,n3477);
or (n3480,n3481,n3484);
and (n3481,n3482,n3483);
xor (n3482,n3326,n3327);
and (n3483,n481,n398);
and (n3484,n3485,n3486);
xor (n3485,n3482,n3483);
or (n3486,n3487,n3490);
and (n3487,n3488,n3489);
xor (n3488,n3332,n3333);
and (n3489,n473,n398);
and (n3490,n3491,n3492);
xor (n3491,n3488,n3489);
or (n3492,n3493,n3496);
and (n3493,n3494,n3495);
xor (n3494,n3338,n3339);
and (n3495,n582,n398);
and (n3496,n3497,n3498);
xor (n3497,n3494,n3495);
or (n3498,n3499,n3502);
and (n3499,n3500,n3501);
xor (n3500,n3344,n3345);
and (n3501,n574,n398);
and (n3502,n3503,n3504);
xor (n3503,n3500,n3501);
or (n3504,n3505,n3508);
and (n3505,n3506,n3507);
xor (n3506,n3350,n3351);
and (n3507,n661,n398);
and (n3508,n3509,n3510);
xor (n3509,n3506,n3507);
or (n3510,n3511,n3514);
and (n3511,n3512,n3513);
xor (n3512,n3356,n3357);
and (n3513,n653,n398);
and (n3514,n3515,n3516);
xor (n3515,n3512,n3513);
or (n3516,n3517,n3520);
and (n3517,n3518,n3519);
xor (n3518,n3362,n3363);
and (n3519,n697,n398);
and (n3520,n3521,n3522);
xor (n3521,n3518,n3519);
or (n3522,n3523,n3526);
and (n3523,n3524,n3525);
xor (n3524,n3368,n3369);
and (n3525,n156,n398);
and (n3526,n3527,n3528);
xor (n3527,n3524,n3525);
or (n3528,n3529,n3532);
and (n3529,n3530,n3531);
xor (n3530,n3374,n3375);
and (n3531,n99,n398);
and (n3532,n3533,n3534);
xor (n3533,n3530,n3531);
or (n3534,n3535,n3538);
and (n3535,n3536,n3537);
xor (n3536,n3380,n3381);
and (n3537,n506,n398);
and (n3538,n3539,n3540);
xor (n3539,n3536,n3537);
or (n3540,n3541,n3544);
and (n3541,n3542,n3543);
xor (n3542,n3386,n3387);
and (n3543,n599,n398);
and (n3544,n3545,n3546);
xor (n3545,n3542,n3543);
or (n3546,n3547,n3550);
and (n3547,n3548,n3549);
xor (n3548,n3392,n3393);
and (n3549,n591,n398);
and (n3550,n3551,n3552);
xor (n3551,n3548,n3549);
or (n3552,n3553,n3556);
and (n3553,n3554,n3555);
xor (n3554,n3398,n3399);
and (n3555,n624,n398);
and (n3556,n3557,n3558);
xor (n3557,n3554,n3555);
or (n3558,n3559,n3562);
and (n3559,n3560,n3561);
xor (n3560,n3404,n3405);
and (n3561,n214,n398);
and (n3562,n3563,n3564);
xor (n3563,n3560,n3561);
or (n3564,n3565,n3568);
and (n3565,n3566,n3567);
xor (n3566,n3410,n3411);
and (n3567,n205,n398);
and (n3568,n3569,n3570);
xor (n3569,n3566,n3567);
or (n3570,n3571,n3574);
and (n3571,n3572,n3573);
xor (n3572,n3416,n3417);
and (n3573,n252,n398);
and (n3574,n3575,n3576);
xor (n3575,n3572,n3573);
or (n3576,n3577,n3580);
and (n3577,n3578,n3579);
xor (n3578,n3422,n3423);
and (n3579,n244,n398);
and (n3580,n3581,n3582);
xor (n3581,n3578,n3579);
or (n3582,n3583,n3586);
and (n3583,n3584,n3585);
xor (n3584,n3428,n3429);
and (n3585,n295,n398);
and (n3586,n3587,n3588);
xor (n3587,n3584,n3585);
or (n3588,n3589,n3592);
and (n3589,n3590,n3591);
xor (n3590,n3434,n3435);
and (n3591,n287,n398);
and (n3592,n3593,n3594);
xor (n3593,n3590,n3591);
or (n3594,n3595,n3598);
and (n3595,n3596,n3597);
xor (n3596,n3440,n3441);
and (n3597,n335,n398);
and (n3598,n3599,n3600);
xor (n3599,n3596,n3597);
or (n3600,n3601,n3604);
and (n3601,n3602,n3603);
xor (n3602,n3446,n3447);
and (n3603,n327,n398);
and (n3604,n3605,n3606);
xor (n3605,n3602,n3603);
or (n3606,n3607,n3610);
and (n3607,n3608,n3609);
xor (n3608,n3452,n3453);
and (n3609,n373,n398);
and (n3610,n3611,n3612);
xor (n3611,n3608,n3609);
or (n3612,n3613,n3616);
and (n3613,n3614,n3615);
xor (n3614,n3458,n3459);
and (n3615,n365,n398);
and (n3616,n3617,n3618);
xor (n3617,n3614,n3615);
and (n3618,n3619,n3620);
xor (n3619,n3464,n3465);
and (n3620,n547,n398);
and (n3621,n562,n734);
or (n3622,n3623,n3626);
and (n3623,n3624,n3625);
xor (n3624,n3473,n3474);
and (n3625,n554,n734);
and (n3626,n3627,n3628);
xor (n3627,n3624,n3625);
or (n3628,n3629,n3632);
and (n3629,n3630,n3631);
xor (n3630,n3479,n3480);
and (n3631,n481,n734);
and (n3632,n3633,n3634);
xor (n3633,n3630,n3631);
or (n3634,n3635,n3638);
and (n3635,n3636,n3637);
xor (n3636,n3485,n3486);
and (n3637,n473,n734);
and (n3638,n3639,n3640);
xor (n3639,n3636,n3637);
or (n3640,n3641,n3644);
and (n3641,n3642,n3643);
xor (n3642,n3491,n3492);
and (n3643,n582,n734);
and (n3644,n3645,n3646);
xor (n3645,n3642,n3643);
or (n3646,n3647,n3650);
and (n3647,n3648,n3649);
xor (n3648,n3497,n3498);
and (n3649,n574,n734);
and (n3650,n3651,n3652);
xor (n3651,n3648,n3649);
or (n3652,n3653,n3656);
and (n3653,n3654,n3655);
xor (n3654,n3503,n3504);
and (n3655,n661,n734);
and (n3656,n3657,n3658);
xor (n3657,n3654,n3655);
or (n3658,n3659,n3662);
and (n3659,n3660,n3661);
xor (n3660,n3509,n3510);
and (n3661,n653,n734);
and (n3662,n3663,n3664);
xor (n3663,n3660,n3661);
or (n3664,n3665,n3668);
and (n3665,n3666,n3667);
xor (n3666,n3515,n3516);
and (n3667,n697,n734);
and (n3668,n3669,n3670);
xor (n3669,n3666,n3667);
or (n3670,n3671,n3674);
and (n3671,n3672,n3673);
xor (n3672,n3521,n3522);
and (n3673,n156,n734);
and (n3674,n3675,n3676);
xor (n3675,n3672,n3673);
or (n3676,n3677,n3680);
and (n3677,n3678,n3679);
xor (n3678,n3527,n3528);
and (n3679,n99,n734);
and (n3680,n3681,n3682);
xor (n3681,n3678,n3679);
or (n3682,n3683,n3686);
and (n3683,n3684,n3685);
xor (n3684,n3533,n3534);
and (n3685,n506,n734);
and (n3686,n3687,n3688);
xor (n3687,n3684,n3685);
or (n3688,n3689,n3692);
and (n3689,n3690,n3691);
xor (n3690,n3539,n3540);
and (n3691,n599,n734);
and (n3692,n3693,n3694);
xor (n3693,n3690,n3691);
or (n3694,n3695,n3698);
and (n3695,n3696,n3697);
xor (n3696,n3545,n3546);
and (n3697,n591,n734);
and (n3698,n3699,n3700);
xor (n3699,n3696,n3697);
or (n3700,n3701,n3704);
and (n3701,n3702,n3703);
xor (n3702,n3551,n3552);
and (n3703,n624,n734);
and (n3704,n3705,n3706);
xor (n3705,n3702,n3703);
or (n3706,n3707,n3710);
and (n3707,n3708,n3709);
xor (n3708,n3557,n3558);
and (n3709,n214,n734);
and (n3710,n3711,n3712);
xor (n3711,n3708,n3709);
or (n3712,n3713,n3716);
and (n3713,n3714,n3715);
xor (n3714,n3563,n3564);
and (n3715,n205,n734);
and (n3716,n3717,n3718);
xor (n3717,n3714,n3715);
or (n3718,n3719,n3722);
and (n3719,n3720,n3721);
xor (n3720,n3569,n3570);
and (n3721,n252,n734);
and (n3722,n3723,n3724);
xor (n3723,n3720,n3721);
or (n3724,n3725,n3728);
and (n3725,n3726,n3727);
xor (n3726,n3575,n3576);
and (n3727,n244,n734);
and (n3728,n3729,n3730);
xor (n3729,n3726,n3727);
or (n3730,n3731,n3734);
and (n3731,n3732,n3733);
xor (n3732,n3581,n3582);
and (n3733,n295,n734);
and (n3734,n3735,n3736);
xor (n3735,n3732,n3733);
or (n3736,n3737,n3740);
and (n3737,n3738,n3739);
xor (n3738,n3587,n3588);
and (n3739,n287,n734);
and (n3740,n3741,n3742);
xor (n3741,n3738,n3739);
or (n3742,n3743,n3746);
and (n3743,n3744,n3745);
xor (n3744,n3593,n3594);
and (n3745,n335,n734);
and (n3746,n3747,n3748);
xor (n3747,n3744,n3745);
or (n3748,n3749,n3752);
and (n3749,n3750,n3751);
xor (n3750,n3599,n3600);
and (n3751,n327,n734);
and (n3752,n3753,n3754);
xor (n3753,n3750,n3751);
or (n3754,n3755,n3758);
and (n3755,n3756,n3757);
xor (n3756,n3605,n3606);
and (n3757,n373,n734);
and (n3758,n3759,n3760);
xor (n3759,n3756,n3757);
or (n3760,n3761,n3764);
and (n3761,n3762,n3763);
xor (n3762,n3611,n3612);
and (n3763,n365,n734);
and (n3764,n3765,n3766);
xor (n3765,n3762,n3763);
and (n3766,n3767,n2679);
xor (n3767,n3617,n3618);
and (n3768,n554,n455);
or (n3769,n3770,n3773);
and (n3770,n3771,n3772);
xor (n3771,n3627,n3628);
and (n3772,n481,n455);
and (n3773,n3774,n3775);
xor (n3774,n3771,n3772);
or (n3775,n3776,n3779);
and (n3776,n3777,n3778);
xor (n3777,n3633,n3634);
and (n3778,n473,n455);
and (n3779,n3780,n3781);
xor (n3780,n3777,n3778);
or (n3781,n3782,n3785);
and (n3782,n3783,n3784);
xor (n3783,n3639,n3640);
and (n3784,n582,n455);
and (n3785,n3786,n3787);
xor (n3786,n3783,n3784);
or (n3787,n3788,n3791);
and (n3788,n3789,n3790);
xor (n3789,n3645,n3646);
and (n3790,n574,n455);
and (n3791,n3792,n3793);
xor (n3792,n3789,n3790);
or (n3793,n3794,n3797);
and (n3794,n3795,n3796);
xor (n3795,n3651,n3652);
and (n3796,n661,n455);
and (n3797,n3798,n3799);
xor (n3798,n3795,n3796);
or (n3799,n3800,n3803);
and (n3800,n3801,n3802);
xor (n3801,n3657,n3658);
and (n3802,n653,n455);
and (n3803,n3804,n3805);
xor (n3804,n3801,n3802);
or (n3805,n3806,n3809);
and (n3806,n3807,n3808);
xor (n3807,n3663,n3664);
and (n3808,n697,n455);
and (n3809,n3810,n3811);
xor (n3810,n3807,n3808);
or (n3811,n3812,n3815);
and (n3812,n3813,n3814);
xor (n3813,n3669,n3670);
and (n3814,n156,n455);
and (n3815,n3816,n3817);
xor (n3816,n3813,n3814);
or (n3817,n3818,n3821);
and (n3818,n3819,n3820);
xor (n3819,n3675,n3676);
and (n3820,n99,n455);
and (n3821,n3822,n3823);
xor (n3822,n3819,n3820);
or (n3823,n3824,n3827);
and (n3824,n3825,n3826);
xor (n3825,n3681,n3682);
and (n3826,n506,n455);
and (n3827,n3828,n3829);
xor (n3828,n3825,n3826);
or (n3829,n3830,n3833);
and (n3830,n3831,n3832);
xor (n3831,n3687,n3688);
and (n3832,n599,n455);
and (n3833,n3834,n3835);
xor (n3834,n3831,n3832);
or (n3835,n3836,n3839);
and (n3836,n3837,n3838);
xor (n3837,n3693,n3694);
and (n3838,n591,n455);
and (n3839,n3840,n3841);
xor (n3840,n3837,n3838);
or (n3841,n3842,n3845);
and (n3842,n3843,n3844);
xor (n3843,n3699,n3700);
and (n3844,n624,n455);
and (n3845,n3846,n3847);
xor (n3846,n3843,n3844);
or (n3847,n3848,n3851);
and (n3848,n3849,n3850);
xor (n3849,n3705,n3706);
and (n3850,n214,n455);
and (n3851,n3852,n3853);
xor (n3852,n3849,n3850);
or (n3853,n3854,n3857);
and (n3854,n3855,n3856);
xor (n3855,n3711,n3712);
and (n3856,n205,n455);
and (n3857,n3858,n3859);
xor (n3858,n3855,n3856);
or (n3859,n3860,n3863);
and (n3860,n3861,n3862);
xor (n3861,n3717,n3718);
and (n3862,n252,n455);
and (n3863,n3864,n3865);
xor (n3864,n3861,n3862);
or (n3865,n3866,n3869);
and (n3866,n3867,n3868);
xor (n3867,n3723,n3724);
and (n3868,n244,n455);
and (n3869,n3870,n3871);
xor (n3870,n3867,n3868);
or (n3871,n3872,n3875);
and (n3872,n3873,n3874);
xor (n3873,n3729,n3730);
and (n3874,n295,n455);
and (n3875,n3876,n3877);
xor (n3876,n3873,n3874);
or (n3877,n3878,n3881);
and (n3878,n3879,n3880);
xor (n3879,n3735,n3736);
and (n3880,n287,n455);
and (n3881,n3882,n3883);
xor (n3882,n3879,n3880);
or (n3883,n3884,n3887);
and (n3884,n3885,n3886);
xor (n3885,n3741,n3742);
and (n3886,n335,n455);
and (n3887,n3888,n3889);
xor (n3888,n3885,n3886);
or (n3889,n3890,n3893);
and (n3890,n3891,n3892);
xor (n3891,n3747,n3748);
and (n3892,n327,n455);
and (n3893,n3894,n3895);
xor (n3894,n3891,n3892);
or (n3895,n3896,n3899);
and (n3896,n3897,n3898);
xor (n3897,n3753,n3754);
and (n3898,n373,n455);
and (n3899,n3900,n3901);
xor (n3900,n3897,n3898);
or (n3901,n3902,n3905);
and (n3902,n3903,n3904);
xor (n3903,n3759,n3760);
and (n3904,n365,n455);
and (n3905,n3906,n3907);
xor (n3906,n3903,n3904);
and (n3907,n3908,n3909);
xor (n3908,n3765,n3766);
and (n3909,n547,n455);
and (n3910,n481,n458);
or (n3911,n3912,n3915);
and (n3912,n3913,n3914);
xor (n3913,n3774,n3775);
and (n3914,n473,n458);
and (n3915,n3916,n3917);
xor (n3916,n3913,n3914);
or (n3917,n3918,n3921);
and (n3918,n3919,n3920);
xor (n3919,n3780,n3781);
and (n3920,n582,n458);
and (n3921,n3922,n3923);
xor (n3922,n3919,n3920);
or (n3923,n3924,n3927);
and (n3924,n3925,n3926);
xor (n3925,n3786,n3787);
and (n3926,n574,n458);
and (n3927,n3928,n3929);
xor (n3928,n3925,n3926);
or (n3929,n3930,n3933);
and (n3930,n3931,n3932);
xor (n3931,n3792,n3793);
and (n3932,n661,n458);
and (n3933,n3934,n3935);
xor (n3934,n3931,n3932);
or (n3935,n3936,n3939);
and (n3936,n3937,n3938);
xor (n3937,n3798,n3799);
and (n3938,n653,n458);
and (n3939,n3940,n3941);
xor (n3940,n3937,n3938);
or (n3941,n3942,n3945);
and (n3942,n3943,n3944);
xor (n3943,n3804,n3805);
and (n3944,n697,n458);
and (n3945,n3946,n3947);
xor (n3946,n3943,n3944);
or (n3947,n3948,n3951);
and (n3948,n3949,n3950);
xor (n3949,n3810,n3811);
and (n3950,n156,n458);
and (n3951,n3952,n3953);
xor (n3952,n3949,n3950);
or (n3953,n3954,n3957);
and (n3954,n3955,n3956);
xor (n3955,n3816,n3817);
and (n3956,n99,n458);
and (n3957,n3958,n3959);
xor (n3958,n3955,n3956);
or (n3959,n3960,n3963);
and (n3960,n3961,n3962);
xor (n3961,n3822,n3823);
and (n3962,n506,n458);
and (n3963,n3964,n3965);
xor (n3964,n3961,n3962);
or (n3965,n3966,n3969);
and (n3966,n3967,n3968);
xor (n3967,n3828,n3829);
and (n3968,n599,n458);
and (n3969,n3970,n3971);
xor (n3970,n3967,n3968);
or (n3971,n3972,n3975);
and (n3972,n3973,n3974);
xor (n3973,n3834,n3835);
and (n3974,n591,n458);
and (n3975,n3976,n3977);
xor (n3976,n3973,n3974);
or (n3977,n3978,n3981);
and (n3978,n3979,n3980);
xor (n3979,n3840,n3841);
and (n3980,n624,n458);
and (n3981,n3982,n3983);
xor (n3982,n3979,n3980);
or (n3983,n3984,n3987);
and (n3984,n3985,n3986);
xor (n3985,n3846,n3847);
and (n3986,n214,n458);
and (n3987,n3988,n3989);
xor (n3988,n3985,n3986);
or (n3989,n3990,n3993);
and (n3990,n3991,n3992);
xor (n3991,n3852,n3853);
and (n3992,n205,n458);
and (n3993,n3994,n3995);
xor (n3994,n3991,n3992);
or (n3995,n3996,n3999);
and (n3996,n3997,n3998);
xor (n3997,n3858,n3859);
and (n3998,n252,n458);
and (n3999,n4000,n4001);
xor (n4000,n3997,n3998);
or (n4001,n4002,n4005);
and (n4002,n4003,n4004);
xor (n4003,n3864,n3865);
and (n4004,n244,n458);
and (n4005,n4006,n4007);
xor (n4006,n4003,n4004);
or (n4007,n4008,n4011);
and (n4008,n4009,n4010);
xor (n4009,n3870,n3871);
and (n4010,n295,n458);
and (n4011,n4012,n4013);
xor (n4012,n4009,n4010);
or (n4013,n4014,n4017);
and (n4014,n4015,n4016);
xor (n4015,n3876,n3877);
and (n4016,n287,n458);
and (n4017,n4018,n4019);
xor (n4018,n4015,n4016);
or (n4019,n4020,n4023);
and (n4020,n4021,n4022);
xor (n4021,n3882,n3883);
and (n4022,n335,n458);
and (n4023,n4024,n4025);
xor (n4024,n4021,n4022);
or (n4025,n4026,n4029);
and (n4026,n4027,n4028);
xor (n4027,n3888,n3889);
and (n4028,n327,n458);
and (n4029,n4030,n4031);
xor (n4030,n4027,n4028);
or (n4031,n4032,n4035);
and (n4032,n4033,n4034);
xor (n4033,n3894,n3895);
and (n4034,n373,n458);
and (n4035,n4036,n4037);
xor (n4036,n4033,n4034);
or (n4037,n4038,n4041);
and (n4038,n4039,n4040);
xor (n4039,n3900,n3901);
and (n4040,n365,n458);
and (n4041,n4042,n4043);
xor (n4042,n4039,n4040);
and (n4043,n4044,n2578);
xor (n4044,n3906,n3907);
and (n4045,n473,n466);
or (n4046,n4047,n4050);
and (n4047,n4048,n4049);
xor (n4048,n3916,n3917);
and (n4049,n582,n466);
and (n4050,n4051,n4052);
xor (n4051,n4048,n4049);
or (n4052,n4053,n4056);
and (n4053,n4054,n4055);
xor (n4054,n3922,n3923);
and (n4055,n574,n466);
and (n4056,n4057,n4058);
xor (n4057,n4054,n4055);
or (n4058,n4059,n4062);
and (n4059,n4060,n4061);
xor (n4060,n3928,n3929);
and (n4061,n661,n466);
and (n4062,n4063,n4064);
xor (n4063,n4060,n4061);
or (n4064,n4065,n4068);
and (n4065,n4066,n4067);
xor (n4066,n3934,n3935);
and (n4067,n653,n466);
and (n4068,n4069,n4070);
xor (n4069,n4066,n4067);
or (n4070,n4071,n4074);
and (n4071,n4072,n4073);
xor (n4072,n3940,n3941);
and (n4073,n697,n466);
and (n4074,n4075,n4076);
xor (n4075,n4072,n4073);
or (n4076,n4077,n4080);
and (n4077,n4078,n4079);
xor (n4078,n3946,n3947);
and (n4079,n156,n466);
and (n4080,n4081,n4082);
xor (n4081,n4078,n4079);
or (n4082,n4083,n4086);
and (n4083,n4084,n4085);
xor (n4084,n3952,n3953);
and (n4085,n99,n466);
and (n4086,n4087,n4088);
xor (n4087,n4084,n4085);
or (n4088,n4089,n4092);
and (n4089,n4090,n4091);
xor (n4090,n3958,n3959);
and (n4091,n506,n466);
and (n4092,n4093,n4094);
xor (n4093,n4090,n4091);
or (n4094,n4095,n4098);
and (n4095,n4096,n4097);
xor (n4096,n3964,n3965);
and (n4097,n599,n466);
and (n4098,n4099,n4100);
xor (n4099,n4096,n4097);
or (n4100,n4101,n4104);
and (n4101,n4102,n4103);
xor (n4102,n3970,n3971);
and (n4103,n591,n466);
and (n4104,n4105,n4106);
xor (n4105,n4102,n4103);
or (n4106,n4107,n4110);
and (n4107,n4108,n4109);
xor (n4108,n3976,n3977);
and (n4109,n624,n466);
and (n4110,n4111,n4112);
xor (n4111,n4108,n4109);
or (n4112,n4113,n4116);
and (n4113,n4114,n4115);
xor (n4114,n3982,n3983);
and (n4115,n214,n466);
and (n4116,n4117,n4118);
xor (n4117,n4114,n4115);
or (n4118,n4119,n4122);
and (n4119,n4120,n4121);
xor (n4120,n3988,n3989);
and (n4121,n205,n466);
and (n4122,n4123,n4124);
xor (n4123,n4120,n4121);
or (n4124,n4125,n4128);
and (n4125,n4126,n4127);
xor (n4126,n3994,n3995);
and (n4127,n252,n466);
and (n4128,n4129,n4130);
xor (n4129,n4126,n4127);
or (n4130,n4131,n4134);
and (n4131,n4132,n4133);
xor (n4132,n4000,n4001);
and (n4133,n244,n466);
and (n4134,n4135,n4136);
xor (n4135,n4132,n4133);
or (n4136,n4137,n4140);
and (n4137,n4138,n4139);
xor (n4138,n4006,n4007);
and (n4139,n295,n466);
and (n4140,n4141,n4142);
xor (n4141,n4138,n4139);
or (n4142,n4143,n4146);
and (n4143,n4144,n4145);
xor (n4144,n4012,n4013);
and (n4145,n287,n466);
and (n4146,n4147,n4148);
xor (n4147,n4144,n4145);
or (n4148,n4149,n4152);
and (n4149,n4150,n4151);
xor (n4150,n4018,n4019);
and (n4151,n335,n466);
and (n4152,n4153,n4154);
xor (n4153,n4150,n4151);
or (n4154,n4155,n4157);
and (n4155,n4156,n2442);
xor (n4156,n4024,n4025);
and (n4157,n4158,n4159);
xor (n4158,n4156,n2442);
or (n4159,n4160,n4163);
and (n4160,n4161,n4162);
xor (n4161,n4030,n4031);
and (n4162,n373,n466);
and (n4163,n4164,n4165);
xor (n4164,n4161,n4162);
or (n4165,n4166,n4169);
and (n4166,n4167,n4168);
xor (n4167,n4036,n4037);
and (n4168,n365,n466);
and (n4169,n4170,n4171);
xor (n4170,n4167,n4168);
and (n4171,n4172,n4173);
xor (n4172,n4042,n4043);
and (n4173,n547,n466);
and (n4174,n582,n638);
or (n4175,n4176,n4179);
and (n4176,n4177,n4178);
xor (n4177,n4051,n4052);
and (n4178,n574,n638);
and (n4179,n4180,n4181);
xor (n4180,n4177,n4178);
or (n4181,n4182,n4185);
and (n4182,n4183,n4184);
xor (n4183,n4057,n4058);
and (n4184,n661,n638);
and (n4185,n4186,n4187);
xor (n4186,n4183,n4184);
or (n4187,n4188,n4191);
and (n4188,n4189,n4190);
xor (n4189,n4063,n4064);
and (n4190,n653,n638);
and (n4191,n4192,n4193);
xor (n4192,n4189,n4190);
or (n4193,n4194,n4197);
and (n4194,n4195,n4196);
xor (n4195,n4069,n4070);
and (n4196,n697,n638);
and (n4197,n4198,n4199);
xor (n4198,n4195,n4196);
or (n4199,n4200,n4203);
and (n4200,n4201,n4202);
xor (n4201,n4075,n4076);
and (n4202,n156,n638);
and (n4203,n4204,n4205);
xor (n4204,n4201,n4202);
or (n4205,n4206,n4209);
and (n4206,n4207,n4208);
xor (n4207,n4081,n4082);
and (n4208,n99,n638);
and (n4209,n4210,n4211);
xor (n4210,n4207,n4208);
or (n4211,n4212,n4215);
and (n4212,n4213,n4214);
xor (n4213,n4087,n4088);
and (n4214,n506,n638);
and (n4215,n4216,n4217);
xor (n4216,n4213,n4214);
or (n4217,n4218,n4221);
and (n4218,n4219,n4220);
xor (n4219,n4093,n4094);
and (n4220,n599,n638);
and (n4221,n4222,n4223);
xor (n4222,n4219,n4220);
or (n4223,n4224,n4227);
and (n4224,n4225,n4226);
xor (n4225,n4099,n4100);
and (n4226,n591,n638);
and (n4227,n4228,n4229);
xor (n4228,n4225,n4226);
or (n4229,n4230,n4233);
and (n4230,n4231,n4232);
xor (n4231,n4105,n4106);
and (n4232,n624,n638);
and (n4233,n4234,n4235);
xor (n4234,n4231,n4232);
or (n4235,n4236,n4239);
and (n4236,n4237,n4238);
xor (n4237,n4111,n4112);
and (n4238,n214,n638);
and (n4239,n4240,n4241);
xor (n4240,n4237,n4238);
or (n4241,n4242,n4245);
and (n4242,n4243,n4244);
xor (n4243,n4117,n4118);
and (n4244,n205,n638);
and (n4245,n4246,n4247);
xor (n4246,n4243,n4244);
or (n4247,n4248,n4251);
and (n4248,n4249,n4250);
xor (n4249,n4123,n4124);
and (n4250,n252,n638);
and (n4251,n4252,n4253);
xor (n4252,n4249,n4250);
or (n4253,n4254,n4257);
and (n4254,n4255,n4256);
xor (n4255,n4129,n4130);
and (n4256,n244,n638);
and (n4257,n4258,n4259);
xor (n4258,n4255,n4256);
or (n4259,n4260,n4263);
and (n4260,n4261,n4262);
xor (n4261,n4135,n4136);
and (n4262,n295,n638);
and (n4263,n4264,n4265);
xor (n4264,n4261,n4262);
or (n4265,n4266,n4269);
and (n4266,n4267,n4268);
xor (n4267,n4141,n4142);
and (n4268,n287,n638);
and (n4269,n4270,n4271);
xor (n4270,n4267,n4268);
or (n4271,n4272,n4275);
and (n4272,n4273,n4274);
xor (n4273,n4147,n4148);
and (n4274,n335,n638);
and (n4275,n4276,n4277);
xor (n4276,n4273,n4274);
or (n4277,n4278,n4281);
and (n4278,n4279,n4280);
xor (n4279,n4153,n4154);
and (n4280,n327,n638);
and (n4281,n4282,n4283);
xor (n4282,n4279,n4280);
or (n4283,n4284,n4287);
and (n4284,n4285,n4286);
xor (n4285,n4158,n4159);
and (n4286,n373,n638);
and (n4287,n4288,n4289);
xor (n4288,n4285,n4286);
or (n4289,n4290,n4293);
and (n4290,n4291,n4292);
xor (n4291,n4164,n4165);
and (n4292,n365,n638);
and (n4293,n4294,n4295);
xor (n4294,n4291,n4292);
and (n4295,n4296,n2471);
xor (n4296,n4170,n4171);
and (n4297,n574,n641);
or (n4298,n4299,n4302);
and (n4299,n4300,n4301);
xor (n4300,n4180,n4181);
and (n4301,n661,n641);
and (n4302,n4303,n4304);
xor (n4303,n4300,n4301);
or (n4304,n4305,n4308);
and (n4305,n4306,n4307);
xor (n4306,n4186,n4187);
and (n4307,n653,n641);
and (n4308,n4309,n4310);
xor (n4309,n4306,n4307);
or (n4310,n4311,n4314);
and (n4311,n4312,n4313);
xor (n4312,n4192,n4193);
and (n4313,n697,n641);
and (n4314,n4315,n4316);
xor (n4315,n4312,n4313);
or (n4316,n4317,n4320);
and (n4317,n4318,n4319);
xor (n4318,n4198,n4199);
and (n4319,n156,n641);
and (n4320,n4321,n4322);
xor (n4321,n4318,n4319);
or (n4322,n4323,n4326);
and (n4323,n4324,n4325);
xor (n4324,n4204,n4205);
and (n4325,n99,n641);
and (n4326,n4327,n4328);
xor (n4327,n4324,n4325);
or (n4328,n4329,n4332);
and (n4329,n4330,n4331);
xor (n4330,n4210,n4211);
and (n4331,n506,n641);
and (n4332,n4333,n4334);
xor (n4333,n4330,n4331);
or (n4334,n4335,n4338);
and (n4335,n4336,n4337);
xor (n4336,n4216,n4217);
and (n4337,n599,n641);
and (n4338,n4339,n4340);
xor (n4339,n4336,n4337);
or (n4340,n4341,n4344);
and (n4341,n4342,n4343);
xor (n4342,n4222,n4223);
and (n4343,n591,n641);
and (n4344,n4345,n4346);
xor (n4345,n4342,n4343);
or (n4346,n4347,n4350);
and (n4347,n4348,n4349);
xor (n4348,n4228,n4229);
and (n4349,n624,n641);
and (n4350,n4351,n4352);
xor (n4351,n4348,n4349);
or (n4352,n4353,n4356);
and (n4353,n4354,n4355);
xor (n4354,n4234,n4235);
and (n4355,n214,n641);
and (n4356,n4357,n4358);
xor (n4357,n4354,n4355);
or (n4358,n4359,n4362);
and (n4359,n4360,n4361);
xor (n4360,n4240,n4241);
and (n4361,n205,n641);
and (n4362,n4363,n4364);
xor (n4363,n4360,n4361);
or (n4364,n4365,n4368);
and (n4365,n4366,n4367);
xor (n4366,n4246,n4247);
and (n4367,n252,n641);
and (n4368,n4369,n4370);
xor (n4369,n4366,n4367);
or (n4370,n4371,n4374);
and (n4371,n4372,n4373);
xor (n4372,n4252,n4253);
and (n4373,n244,n641);
and (n4374,n4375,n4376);
xor (n4375,n4372,n4373);
or (n4376,n4377,n4380);
and (n4377,n4378,n4379);
xor (n4378,n4258,n4259);
and (n4379,n295,n641);
and (n4380,n4381,n4382);
xor (n4381,n4378,n4379);
or (n4382,n4383,n4386);
and (n4383,n4384,n4385);
xor (n4384,n4264,n4265);
and (n4385,n287,n641);
and (n4386,n4387,n4388);
xor (n4387,n4384,n4385);
or (n4388,n4389,n4392);
and (n4389,n4390,n4391);
xor (n4390,n4270,n4271);
and (n4391,n335,n641);
and (n4392,n4393,n4394);
xor (n4393,n4390,n4391);
or (n4394,n4395,n4398);
and (n4395,n4396,n4397);
xor (n4396,n4276,n4277);
and (n4397,n327,n641);
and (n4398,n4399,n4400);
xor (n4399,n4396,n4397);
or (n4400,n4401,n4404);
and (n4401,n4402,n4403);
xor (n4402,n4282,n4283);
and (n4403,n373,n641);
and (n4404,n4405,n4406);
xor (n4405,n4402,n4403);
or (n4406,n4407,n4410);
and (n4407,n4408,n4409);
xor (n4408,n4288,n4289);
and (n4409,n365,n641);
and (n4410,n4411,n4412);
xor (n4411,n4408,n4409);
and (n4412,n4413,n4414);
xor (n4413,n4294,n4295);
and (n4414,n547,n641);
and (n4415,n661,n683);
or (n4416,n4417,n4420);
and (n4417,n4418,n4419);
xor (n4418,n4303,n4304);
and (n4419,n653,n683);
and (n4420,n4421,n4422);
xor (n4421,n4418,n4419);
or (n4422,n4423,n4426);
and (n4423,n4424,n4425);
xor (n4424,n4309,n4310);
and (n4425,n697,n683);
and (n4426,n4427,n4428);
xor (n4427,n4424,n4425);
or (n4428,n4429,n4432);
and (n4429,n4430,n4431);
xor (n4430,n4315,n4316);
and (n4431,n156,n683);
and (n4432,n4433,n4434);
xor (n4433,n4430,n4431);
or (n4434,n4435,n4438);
and (n4435,n4436,n4437);
xor (n4436,n4321,n4322);
and (n4437,n99,n683);
and (n4438,n4439,n4440);
xor (n4439,n4436,n4437);
or (n4440,n4441,n4444);
and (n4441,n4442,n4443);
xor (n4442,n4327,n4328);
and (n4443,n506,n683);
and (n4444,n4445,n4446);
xor (n4445,n4442,n4443);
or (n4446,n4447,n4450);
and (n4447,n4448,n4449);
xor (n4448,n4333,n4334);
and (n4449,n599,n683);
and (n4450,n4451,n4452);
xor (n4451,n4448,n4449);
or (n4452,n4453,n4456);
and (n4453,n4454,n4455);
xor (n4454,n4339,n4340);
and (n4455,n591,n683);
and (n4456,n4457,n4458);
xor (n4457,n4454,n4455);
or (n4458,n4459,n4462);
and (n4459,n4460,n4461);
xor (n4460,n4345,n4346);
and (n4461,n624,n683);
and (n4462,n4463,n4464);
xor (n4463,n4460,n4461);
or (n4464,n4465,n4468);
and (n4465,n4466,n4467);
xor (n4466,n4351,n4352);
and (n4467,n214,n683);
and (n4468,n4469,n4470);
xor (n4469,n4466,n4467);
or (n4470,n4471,n4474);
and (n4471,n4472,n4473);
xor (n4472,n4357,n4358);
and (n4473,n205,n683);
and (n4474,n4475,n4476);
xor (n4475,n4472,n4473);
or (n4476,n4477,n4480);
and (n4477,n4478,n4479);
xor (n4478,n4363,n4364);
and (n4479,n252,n683);
and (n4480,n4481,n4482);
xor (n4481,n4478,n4479);
or (n4482,n4483,n4486);
and (n4483,n4484,n4485);
xor (n4484,n4369,n4370);
and (n4485,n244,n683);
and (n4486,n4487,n4488);
xor (n4487,n4484,n4485);
or (n4488,n4489,n4492);
and (n4489,n4490,n4491);
xor (n4490,n4375,n4376);
and (n4491,n295,n683);
and (n4492,n4493,n4494);
xor (n4493,n4490,n4491);
or (n4494,n4495,n4498);
and (n4495,n4496,n4497);
xor (n4496,n4381,n4382);
and (n4497,n287,n683);
and (n4498,n4499,n4500);
xor (n4499,n4496,n4497);
or (n4500,n4501,n4504);
and (n4501,n4502,n4503);
xor (n4502,n4387,n4388);
and (n4503,n335,n683);
and (n4504,n4505,n4506);
xor (n4505,n4502,n4503);
or (n4506,n4507,n4510);
and (n4507,n4508,n4509);
xor (n4508,n4393,n4394);
and (n4509,n327,n683);
and (n4510,n4511,n4512);
xor (n4511,n4508,n4509);
or (n4512,n4513,n4516);
and (n4513,n4514,n4515);
xor (n4514,n4399,n4400);
and (n4515,n373,n683);
and (n4516,n4517,n4518);
xor (n4517,n4514,n4515);
or (n4518,n4519,n4522);
and (n4519,n4520,n4521);
xor (n4520,n4405,n4406);
and (n4521,n365,n683);
and (n4522,n4523,n4524);
xor (n4523,n4520,n4521);
and (n4524,n4525,n2280);
xor (n4525,n4411,n4412);
and (n4526,n653,n92);
or (n4527,n4528,n4531);
and (n4528,n4529,n4530);
xor (n4529,n4421,n4422);
and (n4530,n697,n92);
and (n4531,n4532,n4533);
xor (n4532,n4529,n4530);
or (n4533,n4534,n4537);
and (n4534,n4535,n4536);
xor (n4535,n4427,n4428);
and (n4536,n156,n92);
and (n4537,n4538,n4539);
xor (n4538,n4535,n4536);
or (n4539,n4540,n4543);
and (n4540,n4541,n4542);
xor (n4541,n4433,n4434);
and (n4542,n99,n92);
and (n4543,n4544,n4545);
xor (n4544,n4541,n4542);
or (n4545,n4546,n4549);
and (n4546,n4547,n4548);
xor (n4547,n4439,n4440);
and (n4548,n506,n92);
and (n4549,n4550,n4551);
xor (n4550,n4547,n4548);
or (n4551,n4552,n4555);
and (n4552,n4553,n4554);
xor (n4553,n4445,n4446);
and (n4554,n599,n92);
and (n4555,n4556,n4557);
xor (n4556,n4553,n4554);
or (n4557,n4558,n4561);
and (n4558,n4559,n4560);
xor (n4559,n4451,n4452);
and (n4560,n591,n92);
and (n4561,n4562,n4563);
xor (n4562,n4559,n4560);
or (n4563,n4564,n4567);
and (n4564,n4565,n4566);
xor (n4565,n4457,n4458);
and (n4566,n624,n92);
and (n4567,n4568,n4569);
xor (n4568,n4565,n4566);
or (n4569,n4570,n4573);
and (n4570,n4571,n4572);
xor (n4571,n4463,n4464);
and (n4572,n214,n92);
and (n4573,n4574,n4575);
xor (n4574,n4571,n4572);
or (n4575,n4576,n4579);
and (n4576,n4577,n4578);
xor (n4577,n4469,n4470);
and (n4578,n205,n92);
and (n4579,n4580,n4581);
xor (n4580,n4577,n4578);
or (n4581,n4582,n4585);
and (n4582,n4583,n4584);
xor (n4583,n4475,n4476);
and (n4584,n252,n92);
and (n4585,n4586,n4587);
xor (n4586,n4583,n4584);
or (n4587,n4588,n4591);
and (n4588,n4589,n4590);
xor (n4589,n4481,n4482);
and (n4590,n244,n92);
and (n4591,n4592,n4593);
xor (n4592,n4589,n4590);
or (n4593,n4594,n4597);
and (n4594,n4595,n4596);
xor (n4595,n4487,n4488);
and (n4596,n295,n92);
and (n4597,n4598,n4599);
xor (n4598,n4595,n4596);
or (n4599,n4600,n4603);
and (n4600,n4601,n4602);
xor (n4601,n4493,n4494);
and (n4602,n287,n92);
and (n4603,n4604,n4605);
xor (n4604,n4601,n4602);
or (n4605,n4606,n4609);
and (n4606,n4607,n4608);
xor (n4607,n4499,n4500);
and (n4608,n335,n92);
and (n4609,n4610,n4611);
xor (n4610,n4607,n4608);
or (n4611,n4612,n4615);
and (n4612,n4613,n4614);
xor (n4613,n4505,n4506);
and (n4614,n327,n92);
and (n4615,n4616,n4617);
xor (n4616,n4613,n4614);
or (n4617,n4618,n4621);
and (n4618,n4619,n4620);
xor (n4619,n4511,n4512);
and (n4620,n373,n92);
and (n4621,n4622,n4623);
xor (n4622,n4619,n4620);
or (n4623,n4624,n4627);
and (n4624,n4625,n4626);
xor (n4625,n4517,n4518);
and (n4626,n365,n92);
and (n4627,n4628,n4629);
xor (n4628,n4625,n4626);
and (n4629,n4630,n4631);
xor (n4630,n4523,n4524);
and (n4631,n547,n92);
and (n4632,n697,n85);
or (n4633,n4634,n4637);
and (n4634,n4635,n4636);
xor (n4635,n4532,n4533);
and (n4636,n156,n85);
and (n4637,n4638,n4639);
xor (n4638,n4635,n4636);
or (n4639,n4640,n4643);
and (n4640,n4641,n4642);
xor (n4641,n4538,n4539);
and (n4642,n99,n85);
and (n4643,n4644,n4645);
xor (n4644,n4641,n4642);
or (n4645,n4646,n4649);
and (n4646,n4647,n4648);
xor (n4647,n4544,n4545);
and (n4648,n506,n85);
and (n4649,n4650,n4651);
xor (n4650,n4647,n4648);
or (n4651,n4652,n4655);
and (n4652,n4653,n4654);
xor (n4653,n4550,n4551);
and (n4654,n599,n85);
and (n4655,n4656,n4657);
xor (n4656,n4653,n4654);
or (n4657,n4658,n4661);
and (n4658,n4659,n4660);
xor (n4659,n4556,n4557);
and (n4660,n591,n85);
and (n4661,n4662,n4663);
xor (n4662,n4659,n4660);
or (n4663,n4664,n4667);
and (n4664,n4665,n4666);
xor (n4665,n4562,n4563);
and (n4666,n624,n85);
and (n4667,n4668,n4669);
xor (n4668,n4665,n4666);
or (n4669,n4670,n4673);
and (n4670,n4671,n4672);
xor (n4671,n4568,n4569);
and (n4672,n214,n85);
and (n4673,n4674,n4675);
xor (n4674,n4671,n4672);
or (n4675,n4676,n4679);
and (n4676,n4677,n4678);
xor (n4677,n4574,n4575);
and (n4678,n205,n85);
and (n4679,n4680,n4681);
xor (n4680,n4677,n4678);
or (n4681,n4682,n4685);
and (n4682,n4683,n4684);
xor (n4683,n4580,n4581);
and (n4684,n252,n85);
and (n4685,n4686,n4687);
xor (n4686,n4683,n4684);
or (n4687,n4688,n4691);
and (n4688,n4689,n4690);
xor (n4689,n4586,n4587);
and (n4690,n244,n85);
and (n4691,n4692,n4693);
xor (n4692,n4689,n4690);
or (n4693,n4694,n4697);
and (n4694,n4695,n4696);
xor (n4695,n4592,n4593);
and (n4696,n295,n85);
and (n4697,n4698,n4699);
xor (n4698,n4695,n4696);
or (n4699,n4700,n4703);
and (n4700,n4701,n4702);
xor (n4701,n4598,n4599);
and (n4702,n287,n85);
and (n4703,n4704,n4705);
xor (n4704,n4701,n4702);
or (n4705,n4706,n4709);
and (n4706,n4707,n4708);
xor (n4707,n4604,n4605);
and (n4708,n335,n85);
and (n4709,n4710,n4711);
xor (n4710,n4707,n4708);
or (n4711,n4712,n4715);
and (n4712,n4713,n4714);
xor (n4713,n4610,n4611);
and (n4714,n327,n85);
and (n4715,n4716,n4717);
xor (n4716,n4713,n4714);
or (n4717,n4718,n4721);
and (n4718,n4719,n4720);
xor (n4719,n4616,n4617);
and (n4720,n373,n85);
and (n4721,n4722,n4723);
xor (n4722,n4719,n4720);
or (n4723,n4724,n4727);
and (n4724,n4725,n4726);
xor (n4725,n4622,n4623);
and (n4726,n365,n85);
and (n4727,n4728,n4729);
xor (n4728,n4725,n4726);
and (n4729,n4730,n2189);
xor (n4730,n4628,n4629);
and (n4731,n156,n22);
or (n4732,n4733,n4736);
and (n4733,n4734,n4735);
xor (n4734,n4638,n4639);
and (n4735,n99,n22);
and (n4736,n4737,n4738);
xor (n4737,n4734,n4735);
or (n4738,n4739,n4742);
and (n4739,n4740,n4741);
xor (n4740,n4644,n4645);
and (n4741,n506,n22);
and (n4742,n4743,n4744);
xor (n4743,n4740,n4741);
or (n4744,n4745,n4748);
and (n4745,n4746,n4747);
xor (n4746,n4650,n4651);
and (n4747,n599,n22);
and (n4748,n4749,n4750);
xor (n4749,n4746,n4747);
or (n4750,n4751,n4754);
and (n4751,n4752,n4753);
xor (n4752,n4656,n4657);
and (n4753,n591,n22);
and (n4754,n4755,n4756);
xor (n4755,n4752,n4753);
or (n4756,n4757,n4760);
and (n4757,n4758,n4759);
xor (n4758,n4662,n4663);
and (n4759,n624,n22);
and (n4760,n4761,n4762);
xor (n4761,n4758,n4759);
or (n4762,n4763,n4766);
and (n4763,n4764,n4765);
xor (n4764,n4668,n4669);
and (n4765,n214,n22);
and (n4766,n4767,n4768);
xor (n4767,n4764,n4765);
or (n4768,n4769,n4772);
and (n4769,n4770,n4771);
xor (n4770,n4674,n4675);
and (n4771,n205,n22);
and (n4772,n4773,n4774);
xor (n4773,n4770,n4771);
or (n4774,n4775,n4778);
and (n4775,n4776,n4777);
xor (n4776,n4680,n4681);
and (n4777,n252,n22);
and (n4778,n4779,n4780);
xor (n4779,n4776,n4777);
or (n4780,n4781,n4784);
and (n4781,n4782,n4783);
xor (n4782,n4686,n4687);
and (n4783,n244,n22);
and (n4784,n4785,n4786);
xor (n4785,n4782,n4783);
or (n4786,n4787,n4790);
and (n4787,n4788,n4789);
xor (n4788,n4692,n4693);
and (n4789,n295,n22);
and (n4790,n4791,n4792);
xor (n4791,n4788,n4789);
or (n4792,n4793,n4796);
and (n4793,n4794,n4795);
xor (n4794,n4698,n4699);
and (n4795,n287,n22);
and (n4796,n4797,n4798);
xor (n4797,n4794,n4795);
or (n4798,n4799,n4802);
and (n4799,n4800,n4801);
xor (n4800,n4704,n4705);
and (n4801,n335,n22);
and (n4802,n4803,n4804);
xor (n4803,n4800,n4801);
or (n4804,n4805,n4808);
and (n4805,n4806,n4807);
xor (n4806,n4710,n4711);
and (n4807,n327,n22);
and (n4808,n4809,n4810);
xor (n4809,n4806,n4807);
or (n4810,n4811,n4814);
and (n4811,n4812,n4813);
xor (n4812,n4716,n4717);
and (n4813,n373,n22);
and (n4814,n4815,n4816);
xor (n4815,n4812,n4813);
or (n4816,n4817,n4820);
and (n4817,n4818,n4819);
xor (n4818,n4722,n4723);
and (n4819,n365,n22);
and (n4820,n4821,n4822);
xor (n4821,n4818,n4819);
and (n4822,n4823,n4824);
xor (n4823,n4728,n4729);
and (n4824,n547,n22);
and (n4825,n99,n492);
or (n4826,n4827,n4830);
and (n4827,n4828,n4829);
xor (n4828,n4737,n4738);
and (n4829,n506,n492);
and (n4830,n4831,n4832);
xor (n4831,n4828,n4829);
or (n4832,n4833,n4836);
and (n4833,n4834,n4835);
xor (n4834,n4743,n4744);
and (n4835,n599,n492);
and (n4836,n4837,n4838);
xor (n4837,n4834,n4835);
or (n4838,n4839,n4842);
and (n4839,n4840,n4841);
xor (n4840,n4749,n4750);
and (n4841,n591,n492);
and (n4842,n4843,n4844);
xor (n4843,n4840,n4841);
or (n4844,n4845,n4848);
and (n4845,n4846,n4847);
xor (n4846,n4755,n4756);
and (n4847,n624,n492);
and (n4848,n4849,n4850);
xor (n4849,n4846,n4847);
or (n4850,n4851,n4854);
and (n4851,n4852,n4853);
xor (n4852,n4761,n4762);
and (n4853,n214,n492);
and (n4854,n4855,n4856);
xor (n4855,n4852,n4853);
or (n4856,n4857,n4860);
and (n4857,n4858,n4859);
xor (n4858,n4767,n4768);
and (n4859,n205,n492);
and (n4860,n4861,n4862);
xor (n4861,n4858,n4859);
or (n4862,n4863,n4866);
and (n4863,n4864,n4865);
xor (n4864,n4773,n4774);
and (n4865,n252,n492);
and (n4866,n4867,n4868);
xor (n4867,n4864,n4865);
or (n4868,n4869,n4872);
and (n4869,n4870,n4871);
xor (n4870,n4779,n4780);
and (n4871,n244,n492);
and (n4872,n4873,n4874);
xor (n4873,n4870,n4871);
or (n4874,n4875,n4878);
and (n4875,n4876,n4877);
xor (n4876,n4785,n4786);
and (n4877,n295,n492);
and (n4878,n4879,n4880);
xor (n4879,n4876,n4877);
or (n4880,n4881,n4884);
and (n4881,n4882,n4883);
xor (n4882,n4791,n4792);
and (n4883,n287,n492);
and (n4884,n4885,n4886);
xor (n4885,n4882,n4883);
or (n4886,n4887,n4890);
and (n4887,n4888,n4889);
xor (n4888,n4797,n4798);
and (n4889,n335,n492);
and (n4890,n4891,n4892);
xor (n4891,n4888,n4889);
or (n4892,n4893,n4896);
and (n4893,n4894,n4895);
xor (n4894,n4803,n4804);
and (n4895,n327,n492);
and (n4896,n4897,n4898);
xor (n4897,n4894,n4895);
or (n4898,n4899,n4902);
and (n4899,n4900,n4901);
xor (n4900,n4809,n4810);
and (n4901,n373,n492);
and (n4902,n4903,n4904);
xor (n4903,n4900,n4901);
or (n4904,n4905,n4908);
and (n4905,n4906,n4907);
xor (n4906,n4815,n4816);
and (n4907,n365,n492);
and (n4908,n4909,n4910);
xor (n4909,n4906,n4907);
and (n4910,n4911,n2388);
xor (n4911,n4821,n4822);
and (n4912,n506,n499);
or (n4913,n4914,n4917);
and (n4914,n4915,n4916);
xor (n4915,n4831,n4832);
and (n4916,n599,n499);
and (n4917,n4918,n4919);
xor (n4918,n4915,n4916);
or (n4919,n4920,n4923);
and (n4920,n4921,n4922);
xor (n4921,n4837,n4838);
and (n4922,n591,n499);
and (n4923,n4924,n4925);
xor (n4924,n4921,n4922);
or (n4925,n4926,n4929);
and (n4926,n4927,n4928);
xor (n4927,n4843,n4844);
and (n4928,n624,n499);
and (n4929,n4930,n4931);
xor (n4930,n4927,n4928);
or (n4931,n4932,n4935);
and (n4932,n4933,n4934);
xor (n4933,n4849,n4850);
and (n4934,n214,n499);
and (n4935,n4936,n4937);
xor (n4936,n4933,n4934);
or (n4937,n4938,n4941);
and (n4938,n4939,n4940);
xor (n4939,n4855,n4856);
and (n4940,n205,n499);
and (n4941,n4942,n4943);
xor (n4942,n4939,n4940);
or (n4943,n4944,n4947);
and (n4944,n4945,n4946);
xor (n4945,n4861,n4862);
and (n4946,n252,n499);
and (n4947,n4948,n4949);
xor (n4948,n4945,n4946);
or (n4949,n4950,n4953);
and (n4950,n4951,n4952);
xor (n4951,n4867,n4868);
and (n4952,n244,n499);
and (n4953,n4954,n4955);
xor (n4954,n4951,n4952);
or (n4955,n4956,n4959);
and (n4956,n4957,n4958);
xor (n4957,n4873,n4874);
and (n4958,n295,n499);
and (n4959,n4960,n4961);
xor (n4960,n4957,n4958);
or (n4961,n4962,n4965);
and (n4962,n4963,n4964);
xor (n4963,n4879,n4880);
and (n4964,n287,n499);
and (n4965,n4966,n4967);
xor (n4966,n4963,n4964);
or (n4967,n4968,n4971);
and (n4968,n4969,n4970);
xor (n4969,n4885,n4886);
and (n4970,n335,n499);
and (n4971,n4972,n4973);
xor (n4972,n4969,n4970);
or (n4973,n4974,n4977);
and (n4974,n4975,n4976);
xor (n4975,n4891,n4892);
and (n4976,n327,n499);
and (n4977,n4978,n4979);
xor (n4978,n4975,n4976);
or (n4979,n4980,n4983);
and (n4980,n4981,n4982);
xor (n4981,n4897,n4898);
and (n4982,n373,n499);
and (n4983,n4984,n4985);
xor (n4984,n4981,n4982);
or (n4985,n4986,n4989);
and (n4986,n4987,n4988);
xor (n4987,n4903,n4904);
and (n4988,n365,n499);
and (n4989,n4990,n4991);
xor (n4990,n4987,n4988);
and (n4991,n4992,n4993);
xor (n4992,n4909,n4910);
and (n4993,n547,n499);
and (n4994,n599,n611);
or (n4995,n4996,n4999);
and (n4996,n4997,n4998);
xor (n4997,n4918,n4919);
and (n4998,n591,n611);
and (n4999,n5000,n5001);
xor (n5000,n4997,n4998);
or (n5001,n5002,n5005);
and (n5002,n5003,n5004);
xor (n5003,n4924,n4925);
and (n5004,n624,n611);
and (n5005,n5006,n5007);
xor (n5006,n5003,n5004);
or (n5007,n5008,n5011);
and (n5008,n5009,n5010);
xor (n5009,n4930,n4931);
and (n5010,n214,n611);
and (n5011,n5012,n5013);
xor (n5012,n5009,n5010);
or (n5013,n5014,n5017);
and (n5014,n5015,n5016);
xor (n5015,n4936,n4937);
and (n5016,n205,n611);
and (n5017,n5018,n5019);
xor (n5018,n5015,n5016);
or (n5019,n5020,n5023);
and (n5020,n5021,n5022);
xor (n5021,n4942,n4943);
and (n5022,n252,n611);
and (n5023,n5024,n5025);
xor (n5024,n5021,n5022);
or (n5025,n5026,n5029);
and (n5026,n5027,n5028);
xor (n5027,n4948,n4949);
and (n5028,n244,n611);
and (n5029,n5030,n5031);
xor (n5030,n5027,n5028);
or (n5031,n5032,n5035);
and (n5032,n5033,n5034);
xor (n5033,n4954,n4955);
and (n5034,n295,n611);
and (n5035,n5036,n5037);
xor (n5036,n5033,n5034);
or (n5037,n5038,n5041);
and (n5038,n5039,n5040);
xor (n5039,n4960,n4961);
and (n5040,n287,n611);
and (n5041,n5042,n5043);
xor (n5042,n5039,n5040);
or (n5043,n5044,n5047);
and (n5044,n5045,n5046);
xor (n5045,n4966,n4967);
and (n5046,n335,n611);
and (n5047,n5048,n5049);
xor (n5048,n5045,n5046);
or (n5049,n5050,n5053);
and (n5050,n5051,n5052);
xor (n5051,n4972,n4973);
and (n5052,n327,n611);
and (n5053,n5054,n5055);
xor (n5054,n5051,n5052);
or (n5055,n5056,n5059);
and (n5056,n5057,n5058);
xor (n5057,n4978,n4979);
and (n5058,n373,n611);
and (n5059,n5060,n5061);
xor (n5060,n5057,n5058);
or (n5061,n5062,n5065);
and (n5062,n5063,n5064);
xor (n5063,n4984,n4985);
and (n5064,n365,n611);
and (n5065,n5066,n5067);
xor (n5066,n5063,n5064);
and (n5067,n5068,n2003);
xor (n5068,n4990,n4991);
and (n5069,n591,n187);
or (n5070,n5071,n5074);
and (n5071,n5072,n5073);
xor (n5072,n5000,n5001);
and (n5073,n624,n187);
and (n5074,n5075,n5076);
xor (n5075,n5072,n5073);
or (n5076,n5077,n5080);
and (n5077,n5078,n5079);
xor (n5078,n5006,n5007);
and (n5079,n214,n187);
and (n5080,n5081,n5082);
xor (n5081,n5078,n5079);
or (n5082,n5083,n5086);
and (n5083,n5084,n5085);
xor (n5084,n5012,n5013);
and (n5085,n205,n187);
and (n5086,n5087,n5088);
xor (n5087,n5084,n5085);
or (n5088,n5089,n5092);
and (n5089,n5090,n5091);
xor (n5090,n5018,n5019);
and (n5091,n252,n187);
and (n5092,n5093,n5094);
xor (n5093,n5090,n5091);
or (n5094,n5095,n5098);
and (n5095,n5096,n5097);
xor (n5096,n5024,n5025);
and (n5097,n244,n187);
and (n5098,n5099,n5100);
xor (n5099,n5096,n5097);
or (n5100,n5101,n5104);
and (n5101,n5102,n5103);
xor (n5102,n5030,n5031);
and (n5103,n295,n187);
and (n5104,n5105,n5106);
xor (n5105,n5102,n5103);
or (n5106,n5107,n5110);
and (n5107,n5108,n5109);
xor (n5108,n5036,n5037);
and (n5109,n287,n187);
and (n5110,n5111,n5112);
xor (n5111,n5108,n5109);
or (n5112,n5113,n5116);
and (n5113,n5114,n5115);
xor (n5114,n5042,n5043);
and (n5115,n335,n187);
and (n5116,n5117,n5118);
xor (n5117,n5114,n5115);
or (n5118,n5119,n5122);
and (n5119,n5120,n5121);
xor (n5120,n5048,n5049);
and (n5121,n327,n187);
and (n5122,n5123,n5124);
xor (n5123,n5120,n5121);
or (n5124,n5125,n5128);
and (n5125,n5126,n5127);
xor (n5126,n5054,n5055);
and (n5127,n373,n187);
and (n5128,n5129,n5130);
xor (n5129,n5126,n5127);
or (n5130,n5131,n5134);
and (n5131,n5132,n5133);
xor (n5132,n5060,n5061);
and (n5133,n365,n187);
and (n5134,n5135,n5136);
xor (n5135,n5132,n5133);
and (n5136,n5137,n5138);
xor (n5137,n5066,n5067);
and (n5138,n547,n187);
and (n5139,n624,n169);
or (n5140,n5141,n5144);
and (n5141,n5142,n5143);
xor (n5142,n5075,n5076);
and (n5143,n214,n169);
and (n5144,n5145,n5146);
xor (n5145,n5142,n5143);
or (n5146,n5147,n5150);
and (n5147,n5148,n5149);
xor (n5148,n5081,n5082);
and (n5149,n205,n169);
and (n5150,n5151,n5152);
xor (n5151,n5148,n5149);
or (n5152,n5153,n5156);
and (n5153,n5154,n5155);
xor (n5154,n5087,n5088);
and (n5155,n252,n169);
and (n5156,n5157,n5158);
xor (n5157,n5154,n5155);
or (n5158,n5159,n5162);
and (n5159,n5160,n5161);
xor (n5160,n5093,n5094);
and (n5161,n244,n169);
and (n5162,n5163,n5164);
xor (n5163,n5160,n5161);
or (n5164,n5165,n5168);
and (n5165,n5166,n5167);
xor (n5166,n5099,n5100);
and (n5167,n295,n169);
and (n5168,n5169,n5170);
xor (n5169,n5166,n5167);
or (n5170,n5171,n5174);
and (n5171,n5172,n5173);
xor (n5172,n5105,n5106);
and (n5173,n287,n169);
and (n5174,n5175,n5176);
xor (n5175,n5172,n5173);
or (n5176,n5177,n5180);
and (n5177,n5178,n5179);
xor (n5178,n5111,n5112);
and (n5179,n335,n169);
and (n5180,n5181,n5182);
xor (n5181,n5178,n5179);
or (n5182,n5183,n5186);
and (n5183,n5184,n5185);
xor (n5184,n5117,n5118);
and (n5185,n327,n169);
and (n5186,n5187,n5188);
xor (n5187,n5184,n5185);
or (n5188,n5189,n5192);
and (n5189,n5190,n5191);
xor (n5190,n5123,n5124);
and (n5191,n373,n169);
and (n5192,n5193,n5194);
xor (n5193,n5190,n5191);
or (n5194,n5195,n5198);
and (n5195,n5196,n5197);
xor (n5196,n5129,n5130);
and (n5197,n365,n169);
and (n5198,n5199,n5200);
xor (n5199,n5196,n5197);
and (n5200,n5201,n1894);
xor (n5201,n5135,n5136);
and (n5202,n214,n196);
or (n5203,n5204,n5207);
and (n5204,n5205,n5206);
xor (n5205,n5145,n5146);
and (n5206,n205,n196);
and (n5207,n5208,n5209);
xor (n5208,n5205,n5206);
or (n5209,n5210,n5213);
and (n5210,n5211,n5212);
xor (n5211,n5151,n5152);
and (n5212,n252,n196);
and (n5213,n5214,n5215);
xor (n5214,n5211,n5212);
or (n5215,n5216,n5219);
and (n5216,n5217,n5218);
xor (n5217,n5157,n5158);
and (n5218,n244,n196);
and (n5219,n5220,n5221);
xor (n5220,n5217,n5218);
or (n5221,n5222,n5225);
and (n5222,n5223,n5224);
xor (n5223,n5163,n5164);
and (n5224,n295,n196);
and (n5225,n5226,n5227);
xor (n5226,n5223,n5224);
or (n5227,n5228,n5231);
and (n5228,n5229,n5230);
xor (n5229,n5169,n5170);
and (n5230,n287,n196);
and (n5231,n5232,n5233);
xor (n5232,n5229,n5230);
or (n5233,n5234,n5237);
and (n5234,n5235,n5236);
xor (n5235,n5175,n5176);
and (n5236,n335,n196);
and (n5237,n5238,n5239);
xor (n5238,n5235,n5236);
or (n5239,n5240,n5243);
and (n5240,n5241,n5242);
xor (n5241,n5181,n5182);
and (n5242,n327,n196);
and (n5243,n5244,n5245);
xor (n5244,n5241,n5242);
or (n5245,n5246,n5249);
and (n5246,n5247,n5248);
xor (n5247,n5187,n5188);
and (n5248,n373,n196);
and (n5249,n5250,n5251);
xor (n5250,n5247,n5248);
or (n5251,n5252,n5255);
and (n5252,n5253,n5254);
xor (n5253,n5193,n5194);
and (n5254,n365,n196);
and (n5255,n5256,n5257);
xor (n5256,n5253,n5254);
and (n5257,n5258,n5259);
xor (n5258,n5199,n5200);
and (n5259,n547,n196);
and (n5260,n205,n224);
or (n5261,n5262,n5265);
and (n5262,n5263,n5264);
xor (n5263,n5208,n5209);
and (n5264,n252,n224);
and (n5265,n5266,n5267);
xor (n5266,n5263,n5264);
or (n5267,n5268,n5271);
and (n5268,n5269,n5270);
xor (n5269,n5214,n5215);
and (n5270,n244,n224);
and (n5271,n5272,n5273);
xor (n5272,n5269,n5270);
or (n5273,n5274,n5277);
and (n5274,n5275,n5276);
xor (n5275,n5220,n5221);
and (n5276,n295,n224);
and (n5277,n5278,n5279);
xor (n5278,n5275,n5276);
or (n5279,n5280,n5283);
and (n5280,n5281,n5282);
xor (n5281,n5226,n5227);
and (n5282,n287,n224);
and (n5283,n5284,n5285);
xor (n5284,n5281,n5282);
or (n5285,n5286,n5289);
and (n5286,n5287,n5288);
xor (n5287,n5232,n5233);
and (n5288,n335,n224);
and (n5289,n5290,n5291);
xor (n5290,n5287,n5288);
or (n5291,n5292,n5295);
and (n5292,n5293,n5294);
xor (n5293,n5238,n5239);
and (n5294,n327,n224);
and (n5295,n5296,n5297);
xor (n5296,n5293,n5294);
or (n5297,n5298,n5301);
and (n5298,n5299,n5300);
xor (n5299,n5244,n5245);
and (n5300,n373,n224);
and (n5301,n5302,n5303);
xor (n5302,n5299,n5300);
or (n5303,n5304,n5307);
and (n5304,n5305,n5306);
xor (n5305,n5250,n5251);
and (n5306,n365,n224);
and (n5307,n5308,n5309);
xor (n5308,n5305,n5306);
and (n5309,n5310,n1428);
xor (n5310,n5256,n5257);
and (n5311,n252,n234);
or (n5312,n5313,n5316);
and (n5313,n5314,n5315);
xor (n5314,n5266,n5267);
and (n5315,n244,n234);
and (n5316,n5317,n5318);
xor (n5317,n5314,n5315);
or (n5318,n5319,n5322);
and (n5319,n5320,n5321);
xor (n5320,n5272,n5273);
and (n5321,n295,n234);
and (n5322,n5323,n5324);
xor (n5323,n5320,n5321);
or (n5324,n5325,n5328);
and (n5325,n5326,n5327);
xor (n5326,n5278,n5279);
and (n5327,n287,n234);
and (n5328,n5329,n5330);
xor (n5329,n5326,n5327);
or (n5330,n5331,n5334);
and (n5331,n5332,n5333);
xor (n5332,n5284,n5285);
and (n5333,n335,n234);
and (n5334,n5335,n5336);
xor (n5335,n5332,n5333);
or (n5336,n5337,n5340);
and (n5337,n5338,n5339);
xor (n5338,n5290,n5291);
and (n5339,n327,n234);
and (n5340,n5341,n5342);
xor (n5341,n5338,n5339);
or (n5342,n5343,n5346);
and (n5343,n5344,n5345);
xor (n5344,n5296,n5297);
and (n5345,n373,n234);
and (n5346,n5347,n5348);
xor (n5347,n5344,n5345);
or (n5348,n5349,n5352);
and (n5349,n5350,n5351);
xor (n5350,n5302,n5303);
and (n5351,n365,n234);
and (n5352,n5353,n5354);
xor (n5353,n5350,n5351);
and (n5354,n5355,n5356);
xor (n5355,n5308,n5309);
and (n5356,n547,n234);
and (n5357,n244,n268);
or (n5358,n5359,n5362);
and (n5359,n5360,n5361);
xor (n5360,n5317,n5318);
and (n5361,n295,n268);
and (n5362,n5363,n5364);
xor (n5363,n5360,n5361);
or (n5364,n5365,n5368);
and (n5365,n5366,n5367);
xor (n5366,n5323,n5324);
and (n5367,n287,n268);
and (n5368,n5369,n5370);
xor (n5369,n5366,n5367);
or (n5370,n5371,n5374);
and (n5371,n5372,n5373);
xor (n5372,n5329,n5330);
and (n5373,n335,n268);
and (n5374,n5375,n5376);
xor (n5375,n5372,n5373);
or (n5376,n5377,n5380);
and (n5377,n5378,n5379);
xor (n5378,n5335,n5336);
and (n5379,n327,n268);
and (n5380,n5381,n5382);
xor (n5381,n5378,n5379);
or (n5382,n5383,n5386);
and (n5383,n5384,n5385);
xor (n5384,n5341,n5342);
and (n5385,n373,n268);
and (n5386,n5387,n5388);
xor (n5387,n5384,n5385);
or (n5388,n5389,n5392);
and (n5389,n5390,n5391);
xor (n5390,n5347,n5348);
and (n5391,n365,n268);
and (n5392,n5393,n5394);
xor (n5393,n5390,n5391);
and (n5394,n5395,n1412);
xor (n5395,n5353,n5354);
and (n5396,n295,n278);
or (n5397,n5398,n5401);
and (n5398,n5399,n5400);
xor (n5399,n5363,n5364);
and (n5400,n287,n278);
and (n5401,n5402,n5403);
xor (n5402,n5399,n5400);
or (n5403,n5404,n5407);
and (n5404,n5405,n5406);
xor (n5405,n5369,n5370);
and (n5406,n335,n278);
and (n5407,n5408,n5409);
xor (n5408,n5405,n5406);
or (n5409,n5410,n5413);
and (n5410,n5411,n5412);
xor (n5411,n5375,n5376);
and (n5412,n327,n278);
and (n5413,n5414,n5415);
xor (n5414,n5411,n5412);
or (n5415,n5416,n5419);
and (n5416,n5417,n5418);
xor (n5417,n5381,n5382);
and (n5418,n373,n278);
and (n5419,n5420,n5421);
xor (n5420,n5417,n5418);
or (n5421,n5422,n5425);
and (n5422,n5423,n5424);
xor (n5423,n5387,n5388);
and (n5424,n365,n278);
and (n5425,n5426,n5427);
xor (n5426,n5423,n5424);
and (n5427,n5428,n5429);
xor (n5428,n5393,n5394);
and (n5429,n547,n278);
and (n5430,n287,n306);
or (n5431,n5432,n5435);
and (n5432,n5433,n5434);
xor (n5433,n5402,n5403);
and (n5434,n335,n306);
and (n5435,n5436,n5437);
xor (n5436,n5433,n5434);
or (n5437,n5438,n5441);
and (n5438,n5439,n5440);
xor (n5439,n5408,n5409);
and (n5440,n327,n306);
and (n5441,n5442,n5443);
xor (n5442,n5439,n5440);
or (n5443,n5444,n5447);
and (n5444,n5445,n5446);
xor (n5445,n5414,n5415);
and (n5446,n373,n306);
and (n5447,n5448,n5449);
xor (n5448,n5445,n5446);
or (n5449,n5450,n5453);
and (n5450,n5451,n5452);
xor (n5451,n5420,n5421);
and (n5452,n365,n306);
and (n5453,n5454,n5455);
xor (n5454,n5451,n5452);
and (n5455,n5456,n968);
xor (n5456,n5426,n5427);
and (n5457,n335,n313);
or (n5458,n5459,n5462);
and (n5459,n5460,n5461);
xor (n5460,n5436,n5437);
and (n5461,n327,n313);
and (n5462,n5463,n5464);
xor (n5463,n5460,n5461);
or (n5464,n5465,n5468);
and (n5465,n5466,n5467);
xor (n5466,n5442,n5443);
and (n5467,n373,n313);
and (n5468,n5469,n5470);
xor (n5469,n5466,n5467);
or (n5470,n5471,n5474);
and (n5471,n5472,n5473);
xor (n5472,n5448,n5449);
and (n5473,n365,n313);
and (n5474,n5475,n5476);
xor (n5475,n5472,n5473);
and (n5476,n5477,n5478);
xor (n5477,n5454,n5455);
and (n5478,n547,n313);
and (n5479,n327,n345);
or (n5480,n5481,n5484);
and (n5481,n5482,n5483);
xor (n5482,n5463,n5464);
and (n5483,n373,n345);
and (n5484,n5485,n5486);
xor (n5485,n5482,n5483);
or (n5486,n5487,n5490);
and (n5487,n5488,n5489);
xor (n5488,n5469,n5470);
and (n5489,n365,n345);
and (n5490,n5491,n5492);
xor (n5491,n5488,n5489);
and (n5492,n5493,n546);
xor (n5493,n5475,n5476);
and (n5494,n373,n355);
or (n5495,n5496,n5499);
and (n5496,n5497,n5498);
xor (n5497,n5485,n5486);
and (n5498,n365,n355);
and (n5499,n5500,n5501);
xor (n5500,n5497,n5498);
and (n5501,n5502,n5503);
xor (n5502,n5491,n5492);
and (n5503,n547,n355);
and (n5504,n365,n756);
and (n5505,n5506,n1092);
xor (n5506,n5500,n5501);
and (n5507,n547,n1072);
endmodule
