module top (out,n11,n12,n14,n15,n18,n19,n25,n30,n31
        ,n40,n41,n43,n50,n53,n111,n217,n219,n222,n231
        ,n239,n241,n250,n307);
output out;
input n11;
input n12;
input n14;
input n15;
input n18;
input n19;
input n25;
input n30;
input n31;
input n40;
input n41;
input n43;
input n50;
input n53;
input n111;
input n217;
input n219;
input n222;
input n231;
input n239;
input n241;
input n250;
input n307;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n13;
wire n16;
wire n17;
wire n20;
wire n21;
wire n22;
wire n23;
wire n24;
wire n26;
wire n27;
wire n28;
wire n29;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n42;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n51;
wire n52;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n218;
wire n220;
wire n221;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n240;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
xor (out,n0,n453);
xor (n0,n1,n404);
xor (n1,n2,n208);
xor (n2,n3,n116);
xor (n3,n4,n100);
xor (n4,n5,n73);
xor (n5,n6,n34);
or (n6,n7,n26,n33);
and (n7,n8,n21);
or (n8,n9,n16,n20);
and (n9,n10,n13);
and (n10,n11,n12);
and (n13,n14,n15);
and (n16,n13,n17);
and (n17,n18,n19);
and (n20,n10,n17);
nor (n21,n22,n23);
not (n22,n11);
and (n23,n24,n11);
not (n24,n25);
and (n26,n21,n27);
nor (n27,n28,n32);
and (n28,n29,n31);
not (n29,n30);
not (n32,n31);
and (n33,n8,n27);
or (n34,n35,n57,n72);
and (n35,n36,n55);
or (n36,n37,n46,n54);
and (n37,n38,n44);
and (n38,n39,n42);
and (n39,n40,n41);
and (n42,n43,n31);
xor (n44,n45,n17);
xor (n45,n10,n13);
and (n46,n44,n47);
xor (n47,n48,n52);
xor (n48,n49,n51);
and (n49,n40,n50);
and (n51,n43,n41);
and (n52,n53,n31);
and (n54,n38,n47);
xor (n55,n56,n27);
xor (n56,n8,n21);
and (n57,n55,n58);
xor (n58,n59,n69);
xor (n59,n60,n64);
or (n60,n61,n62,n63);
and (n61,n49,n51);
and (n62,n51,n52);
and (n63,n49,n52);
xor (n64,n65,n68);
xor (n65,n66,n67);
and (n66,n40,n19);
and (n67,n43,n50);
and (n68,n53,n41);
xor (n69,n70,n71);
and (n70,n14,n12);
and (n71,n18,n15);
and (n72,n36,n58);
xor (n73,n74,n88);
xor (n74,n75,n79);
or (n75,n76,n77,n78);
and (n76,n60,n64);
and (n77,n64,n69);
and (n78,n60,n69);
xor (n79,n80,n85);
xor (n80,n81,n84);
nor (n81,n82,n83);
not (n82,n14);
and (n83,n24,n14);
and (n84,n18,n12);
nor (n85,n86,n87);
and (n86,n29,n41);
not (n87,n41);
xor (n88,n89,n95);
xor (n89,n90,n94);
or (n90,n91,n92,n93);
and (n91,n66,n67);
and (n92,n67,n68);
and (n93,n66,n68);
and (n94,n70,n71);
xor (n95,n96,n99);
xor (n96,n97,n98);
and (n97,n40,n15);
and (n98,n43,n19);
and (n99,n53,n50);
and (n100,n101,n114);
or (n101,n102,n108,n113);
and (n102,n103,n106);
and (n103,n104,n105);
and (n104,n18,n50);
xor (n105,n39,n42);
xor (n106,n107,n47);
xor (n107,n38,n44);
and (n108,n106,n109);
nor (n109,n110,n112);
not (n110,n111);
and (n112,n24,n111);
and (n113,n103,n109);
xor (n114,n115,n58);
xor (n115,n36,n55);
or (n116,n117,n147);
and (n117,n118,n119);
xor (n118,n101,n114);
or (n119,n120,n143,n146);
and (n120,n121,n128);
or (n121,n122,n125,n127);
and (n122,n123,n124);
and (n123,n111,n12);
and (n124,n11,n15);
and (n125,n124,n126);
and (n126,n14,n19);
and (n127,n123,n126);
or (n128,n129,n140,n142);
and (n129,n130,n138);
or (n130,n131,n134,n137);
and (n131,n132,n133);
and (n132,n14,n41);
and (n133,n18,n31);
and (n134,n135,n136);
and (n135,n18,n41);
and (n136,n40,n31);
and (n137,n131,n136);
xor (n138,n139,n126);
xor (n139,n123,n124);
and (n140,n138,n141);
xor (n141,n104,n105);
and (n142,n130,n141);
and (n143,n128,n144);
xor (n144,n145,n109);
xor (n145,n103,n106);
and (n146,n121,n144);
and (n147,n148,n149);
xor (n148,n118,n119);
or (n149,n150,n178);
and (n150,n151,n153);
xor (n151,n152,n144);
xor (n152,n121,n128);
or (n153,n154,n174,n177);
and (n154,n155,n158);
and (n155,n156,n157);
and (n156,n11,n19);
and (n157,n14,n50);
or (n158,n159,n170,n173);
and (n159,n160,n169);
or (n160,n161,n166,n168);
and (n161,n162,n165);
and (n162,n163,n164);
and (n163,n11,n41);
and (n164,n14,n31);
and (n165,n11,n50);
and (n166,n165,n167);
xor (n167,n132,n133);
and (n168,n162,n167);
xor (n169,n156,n157);
and (n170,n169,n171);
xor (n171,n172,n136);
xor (n172,n131,n135);
and (n173,n160,n171);
and (n174,n158,n175);
xor (n175,n176,n141);
xor (n176,n130,n138);
and (n177,n155,n175);
and (n178,n179,n180);
xor (n179,n151,n153);
or (n180,n181,n203);
and (n181,n182,n184);
xor (n182,n183,n175);
xor (n183,n155,n158);
and (n184,n185,n201);
or (n185,n186,n197,n200);
and (n186,n187,n196);
or (n187,n188,n193,n195);
and (n188,n189,n192);
and (n189,n190,n191);
and (n190,n111,n41);
and (n191,n11,n31);
and (n192,n111,n50);
and (n193,n192,n194);
xor (n194,n163,n164);
and (n195,n189,n194);
and (n196,n111,n19);
and (n197,n196,n198);
xor (n198,n199,n167);
xor (n199,n162,n165);
and (n200,n187,n198);
xor (n201,n202,n171);
xor (n202,n160,n169);
and (n203,n204,n205);
xor (n204,n182,n184);
and (n205,n206,n207);
and (n206,n111,n15);
xor (n207,n185,n201);
xor (n208,n209,n312);
xor (n209,n210,n296);
xor (n210,n211,n270);
xor (n211,n212,n233);
or (n212,n213,n227,n232);
and (n213,n214,n224);
or (n214,n215,n220,n223);
and (n215,n216,n218);
and (n216,n217,n12);
and (n218,n219,n15);
and (n220,n218,n221);
and (n221,n222,n19);
and (n223,n216,n221);
nor (n224,n225,n226);
not (n225,n217);
and (n226,n24,n217);
and (n227,n224,n228);
nor (n228,n229,n32);
and (n229,n230,n31);
not (n230,n231);
and (n232,n214,n228);
or (n233,n234,n254,n269);
and (n234,n235,n252);
or (n235,n236,n244,n251);
and (n236,n237,n242);
and (n237,n238,n240);
and (n238,n239,n41);
and (n240,n241,n31);
xor (n242,n243,n221);
xor (n243,n216,n218);
and (n244,n242,n245);
xor (n245,n246,n249);
xor (n246,n247,n248);
and (n247,n239,n50);
and (n248,n241,n41);
and (n249,n250,n31);
and (n251,n237,n245);
xor (n252,n253,n228);
xor (n253,n214,n224);
and (n254,n252,n255);
xor (n255,n256,n266);
xor (n256,n257,n261);
or (n257,n258,n259,n260);
and (n258,n247,n248);
and (n259,n248,n249);
and (n260,n247,n249);
xor (n261,n262,n265);
xor (n262,n263,n264);
and (n263,n239,n19);
and (n264,n241,n50);
and (n265,n250,n41);
xor (n266,n267,n268);
and (n267,n219,n12);
and (n268,n222,n15);
and (n269,n235,n255);
xor (n270,n271,n284);
xor (n271,n272,n276);
or (n272,n273,n274,n275);
and (n273,n257,n261);
and (n274,n261,n266);
and (n275,n257,n266);
xor (n276,n277,n282);
xor (n277,n278,n281);
nor (n278,n279,n280);
not (n279,n219);
and (n280,n24,n219);
and (n281,n222,n12);
nor (n282,n283,n87);
and (n283,n230,n41);
xor (n284,n285,n291);
xor (n285,n286,n290);
or (n286,n287,n288,n289);
and (n287,n263,n264);
and (n288,n264,n265);
and (n289,n263,n265);
and (n290,n267,n268);
xor (n291,n292,n295);
xor (n292,n293,n294);
and (n293,n239,n15);
and (n294,n241,n19);
and (n295,n250,n50);
and (n296,n297,n310);
or (n297,n298,n304,n309);
and (n298,n299,n302);
and (n299,n300,n301);
and (n300,n222,n50);
xor (n301,n238,n240);
xor (n302,n303,n245);
xor (n303,n237,n242);
and (n304,n302,n305);
nor (n305,n306,n308);
not (n306,n307);
and (n308,n24,n307);
and (n309,n299,n305);
xor (n310,n311,n255);
xor (n311,n235,n252);
or (n312,n313,n343);
and (n313,n314,n315);
xor (n314,n297,n310);
or (n315,n316,n339,n342);
and (n316,n317,n324);
or (n317,n318,n321,n323);
and (n318,n319,n320);
and (n319,n307,n12);
and (n320,n217,n15);
and (n321,n320,n322);
and (n322,n219,n19);
and (n323,n319,n322);
or (n324,n325,n336,n338);
and (n325,n326,n334);
or (n326,n327,n330,n333);
and (n327,n328,n329);
and (n328,n219,n41);
and (n329,n222,n31);
and (n330,n331,n332);
and (n331,n222,n41);
and (n332,n239,n31);
and (n333,n327,n332);
xor (n334,n335,n322);
xor (n335,n319,n320);
and (n336,n334,n337);
xor (n337,n300,n301);
and (n338,n326,n337);
and (n339,n324,n340);
xor (n340,n341,n305);
xor (n341,n299,n302);
and (n342,n317,n340);
and (n343,n344,n345);
xor (n344,n314,n315);
or (n345,n346,n374);
and (n346,n347,n349);
xor (n347,n348,n340);
xor (n348,n317,n324);
or (n349,n350,n370,n373);
and (n350,n351,n354);
and (n351,n352,n353);
and (n352,n217,n19);
and (n353,n219,n50);
or (n354,n355,n366,n369);
and (n355,n356,n365);
or (n356,n357,n362,n364);
and (n357,n358,n361);
and (n358,n359,n360);
and (n359,n217,n41);
and (n360,n219,n31);
and (n361,n217,n50);
and (n362,n361,n363);
xor (n363,n328,n329);
and (n364,n358,n363);
xor (n365,n352,n353);
and (n366,n365,n367);
xor (n367,n368,n332);
xor (n368,n327,n331);
and (n369,n356,n367);
and (n370,n354,n371);
xor (n371,n372,n337);
xor (n372,n326,n334);
and (n373,n351,n371);
and (n374,n375,n376);
xor (n375,n347,n349);
or (n376,n377,n399);
and (n377,n378,n380);
xor (n378,n379,n371);
xor (n379,n351,n354);
and (n380,n381,n397);
or (n381,n382,n393,n396);
and (n382,n383,n392);
or (n383,n384,n389,n391);
and (n384,n385,n388);
and (n385,n386,n387);
and (n386,n307,n41);
and (n387,n217,n31);
and (n388,n307,n50);
and (n389,n388,n390);
xor (n390,n359,n360);
and (n391,n385,n390);
and (n392,n307,n19);
and (n393,n392,n394);
xor (n394,n395,n363);
xor (n395,n358,n361);
and (n396,n383,n394);
xor (n397,n398,n367);
xor (n398,n356,n365);
and (n399,n400,n401);
xor (n400,n378,n380);
and (n401,n402,n403);
and (n402,n307,n15);
xor (n403,n381,n397);
or (n404,n405,n408,n452);
and (n405,n406,n407);
xor (n406,n148,n149);
xor (n407,n344,n345);
and (n408,n407,n409);
or (n409,n410,n413,n451);
and (n410,n411,n412);
xor (n411,n179,n180);
xor (n412,n375,n376);
and (n413,n412,n414);
or (n414,n415,n418,n450);
and (n415,n416,n417);
xor (n416,n204,n205);
xor (n417,n400,n401);
and (n418,n417,n419);
or (n419,n420,n423,n449);
and (n420,n421,n422);
xor (n421,n206,n207);
xor (n422,n402,n403);
and (n423,n422,n424);
or (n424,n425,n430,n448);
and (n425,n426,n428);
xor (n426,n427,n198);
xor (n427,n187,n196);
xor (n428,n429,n394);
xor (n429,n383,n392);
and (n430,n428,n431);
or (n431,n432,n437,n447);
and (n432,n433,n435);
xor (n433,n434,n194);
xor (n434,n189,n192);
xor (n435,n436,n390);
xor (n436,n385,n388);
and (n437,n435,n438);
or (n438,n439,n442,n446);
and (n439,n440,n441);
xor (n440,n190,n191);
xor (n441,n386,n387);
and (n442,n441,n443);
and (n443,n444,n445);
and (n444,n111,n31);
and (n445,n307,n31);
and (n446,n440,n443);
and (n447,n433,n438);
and (n448,n426,n431);
and (n449,n421,n424);
and (n450,n416,n419);
and (n451,n411,n414);
and (n452,n406,n409);
xor (n453,n454,n595);
xor (n454,n455,n573);
xor (n455,n456,n537);
xor (n456,n457,n499);
and (n457,n458,n484);
or (n458,n459,n475,n483);
and (n459,n460,n468);
and (n460,n461,n15);
xor (n461,n462,n463);
xor (n462,n14,n219);
or (n463,n464,n465,n467);
and (n464,n11,n217);
and (n465,n217,n466);
and (n466,n111,n307);
and (n467,n11,n466);
and (n468,n469,n19);
xor (n469,n470,n471);
xor (n470,n18,n222);
or (n471,n472,n473,n474);
and (n472,n14,n219);
and (n473,n219,n463);
and (n474,n14,n463);
and (n475,n468,n476);
and (n476,n477,n50);
xor (n477,n478,n479);
xor (n478,n40,n239);
or (n479,n480,n481,n482);
and (n480,n18,n222);
and (n481,n222,n471);
and (n482,n18,n471);
and (n483,n460,n476);
and (n484,n485,n492);
and (n485,n486,n41);
xor (n486,n487,n488);
xor (n487,n43,n241);
or (n488,n489,n490,n491);
and (n489,n40,n239);
and (n490,n239,n479);
and (n491,n40,n479);
and (n492,n493,n31);
xor (n493,n494,n495);
xor (n494,n53,n250);
or (n495,n496,n497,n498);
and (n496,n43,n241);
and (n497,n241,n488);
and (n498,n43,n488);
or (n499,n500,n512,n536);
and (n500,n501,n511);
or (n501,n502,n508,n510);
and (n502,n503,n506);
and (n503,n504,n505);
and (n504,n477,n41);
and (n505,n486,n31);
xor (n506,n507,n476);
xor (n507,n460,n468);
and (n508,n506,n509);
xor (n509,n485,n492);
and (n510,n503,n509);
xor (n511,n458,n484);
and (n512,n511,n513);
xor (n513,n514,n531);
xor (n514,n515,n520);
nor (n515,n516,n519);
not (n516,n517);
xor (n517,n518,n466);
xor (n518,n11,n217);
and (n519,n24,n517);
xor (n520,n521,n524);
xor (n521,n522,n523);
and (n522,n486,n50);
and (n523,n493,n41);
and (n524,n525,n31);
xor (n525,n526,n527);
xor (n526,n30,n231);
or (n527,n528,n529,n530);
and (n528,n53,n250);
and (n529,n250,n495);
and (n530,n53,n495);
xor (n531,n532,n535);
xor (n532,n533,n534);
and (n533,n461,n12);
and (n534,n469,n15);
and (n535,n477,n19);
and (n536,n501,n513);
xor (n537,n538,n561);
xor (n538,n539,n543);
or (n539,n540,n541,n542);
and (n540,n515,n520);
and (n541,n520,n531);
and (n542,n515,n531);
xor (n543,n544,n554);
xor (n544,n545,n549);
or (n545,n546,n547,n548);
and (n546,n522,n523);
and (n547,n523,n524);
and (n548,n522,n524);
xor (n549,n550,n553);
xor (n550,n551,n552);
and (n551,n486,n19);
and (n552,n493,n50);
and (n553,n525,n41);
xor (n554,n555,n560);
xor (n555,n556,n559);
nor (n556,n557,n558);
not (n557,n461);
and (n558,n24,n461);
and (n559,n469,n12);
and (n560,n477,n15);
xor (n561,n562,n566);
or (n562,n563,n564,n565);
and (n563,n533,n534);
and (n564,n534,n535);
and (n565,n533,n535);
nor (n566,n567,n32);
and (n567,n568,n31);
not (n568,n569);
or (n569,n570,n571,n572);
and (n570,n30,n231);
and (n571,n231,n527);
and (n572,n30,n527);
or (n573,n574,n591,n594);
and (n574,n575,n581);
and (n575,n576,n580);
nor (n576,n577,n579);
not (n577,n578);
xor (n578,n111,n307);
and (n579,n24,n578);
and (n580,n517,n12);
or (n581,n582,n588,n590);
and (n582,n583,n586);
and (n583,n584,n585);
and (n584,n469,n50);
xor (n585,n504,n505);
xor (n586,n587,n509);
xor (n587,n503,n506);
and (n588,n586,n589);
xor (n589,n576,n580);
and (n590,n583,n589);
and (n591,n581,n592);
xor (n592,n593,n513);
xor (n593,n501,n511);
and (n594,n575,n592);
or (n595,n596,n627);
and (n596,n597,n599);
xor (n597,n598,n592);
xor (n598,n575,n581);
or (n599,n600,n623,n626);
and (n600,n601,n608);
or (n601,n602,n605,n607);
and (n602,n603,n604);
and (n603,n578,n12);
and (n604,n517,n15);
and (n605,n604,n606);
and (n606,n461,n19);
and (n607,n603,n606);
or (n608,n609,n620,n622);
and (n609,n610,n618);
or (n610,n611,n614,n617);
and (n611,n612,n613);
and (n612,n461,n41);
and (n613,n469,n31);
and (n614,n615,n616);
and (n615,n469,n41);
and (n616,n477,n31);
and (n617,n611,n616);
xor (n618,n619,n606);
xor (n619,n603,n604);
and (n620,n618,n621);
xor (n621,n584,n585);
and (n622,n610,n621);
and (n623,n608,n624);
xor (n624,n625,n589);
xor (n625,n583,n586);
and (n626,n601,n624);
and (n627,n628,n629);
xor (n628,n597,n599);
or (n629,n630,n658);
and (n630,n631,n633);
xor (n631,n632,n624);
xor (n632,n601,n608);
or (n633,n634,n654,n657);
and (n634,n635,n638);
and (n635,n636,n637);
and (n636,n517,n19);
and (n637,n461,n50);
or (n638,n639,n650,n653);
and (n639,n640,n649);
or (n640,n641,n646,n648);
and (n641,n642,n645);
and (n642,n643,n644);
and (n643,n517,n41);
and (n644,n461,n31);
and (n645,n517,n50);
and (n646,n645,n647);
xor (n647,n612,n613);
and (n648,n642,n647);
xor (n649,n636,n637);
and (n650,n649,n651);
xor (n651,n652,n616);
xor (n652,n611,n615);
and (n653,n640,n651);
and (n654,n638,n655);
xor (n655,n656,n621);
xor (n656,n610,n618);
and (n657,n635,n655);
and (n658,n659,n660);
xor (n659,n631,n633);
or (n660,n661,n683);
and (n661,n662,n664);
xor (n662,n663,n655);
xor (n663,n635,n638);
and (n664,n665,n681);
or (n665,n666,n677,n680);
and (n666,n667,n676);
or (n667,n668,n673,n675);
and (n668,n669,n672);
and (n669,n670,n671);
and (n670,n578,n41);
and (n671,n517,n31);
and (n672,n578,n50);
and (n673,n672,n674);
xor (n674,n643,n644);
and (n675,n669,n674);
and (n676,n578,n19);
and (n677,n676,n678);
xor (n678,n679,n647);
xor (n679,n642,n645);
and (n680,n667,n678);
xor (n681,n682,n651);
xor (n682,n640,n649);
and (n683,n684,n685);
xor (n684,n662,n664);
and (n685,n686,n687);
and (n686,n578,n15);
xor (n687,n665,n681);
endmodule
