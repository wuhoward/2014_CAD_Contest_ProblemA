module top (out,n13,n15,n20,n22,n32,n41,n47,n51,n57
        ,n70,n71,n91,n128,n134,n152,n153,n188,n189,n210
        ,n215,n255,n382,n388,n395,n401,n435,n436,n443,n456
        ,n528,n548,n608);
output out;
input n13;
input n15;
input n20;
input n22;
input n32;
input n41;
input n47;
input n51;
input n57;
input n70;
input n71;
input n91;
input n128;
input n134;
input n152;
input n153;
input n188;
input n189;
input n210;
input n215;
input n255;
input n382;
input n388;
input n395;
input n401;
input n435;
input n436;
input n443;
input n456;
input n528;
input n548;
input n608;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n14;
wire n16;
wire n17;
wire n18;
wire n19;
wire n21;
wire n23;
wire n24;
wire n25;
wire n26;
wire n27;
wire n28;
wire n29;
wire n30;
wire n31;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n48;
wire n49;
wire n50;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n211;
wire n212;
wire n213;
wire n214;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2988;
wire n2989;
wire n2990;
wire n2991;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2996;
wire n2997;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3003;
wire n3004;
wire n3005;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3010;
wire n3011;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3038;
wire n3039;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
wire n3056;
wire n3057;
wire n3058;
wire n3059;
wire n3060;
wire n3061;
wire n3062;
wire n3063;
wire n3064;
wire n3065;
wire n3066;
wire n3067;
wire n3068;
wire n3069;
wire n3070;
wire n3071;
wire n3072;
wire n3073;
wire n3074;
wire n3075;
wire n3076;
wire n3077;
wire n3078;
wire n3079;
wire n3080;
wire n3081;
wire n3082;
wire n3083;
wire n3084;
wire n3085;
wire n3086;
wire n3087;
wire n3088;
wire n3089;
wire n3090;
wire n3091;
wire n3092;
wire n3093;
wire n3094;
wire n3095;
wire n3096;
wire n3097;
wire n3098;
wire n3099;
wire n3100;
wire n3101;
wire n3102;
wire n3103;
wire n3104;
wire n3105;
wire n3106;
wire n3107;
wire n3108;
wire n3109;
wire n3110;
wire n3111;
wire n3112;
wire n3113;
wire n3114;
wire n3115;
wire n3116;
wire n3117;
wire n3118;
wire n3119;
wire n3120;
wire n3121;
wire n3122;
wire n3123;
wire n3124;
wire n3125;
wire n3126;
wire n3127;
wire n3128;
wire n3129;
wire n3130;
wire n3131;
wire n3132;
wire n3133;
wire n3134;
wire n3135;
wire n3136;
wire n3137;
wire n3138;
wire n3139;
wire n3140;
wire n3141;
wire n3142;
wire n3143;
wire n3144;
wire n3145;
wire n3146;
wire n3147;
wire n3148;
wire n3149;
wire n3150;
wire n3151;
wire n3152;
wire n3153;
wire n3154;
wire n3155;
wire n3156;
wire n3157;
wire n3158;
wire n3159;
wire n3160;
wire n3161;
wire n3162;
wire n3163;
wire n3164;
wire n3165;
wire n3166;
wire n3167;
wire n3168;
wire n3169;
wire n3170;
wire n3171;
wire n3172;
wire n3173;
wire n3174;
wire n3175;
wire n3176;
wire n3177;
wire n3178;
wire n3179;
wire n3180;
wire n3181;
wire n3182;
wire n3183;
wire n3184;
wire n3185;
wire n3186;
wire n3187;
wire n3188;
wire n3189;
wire n3190;
wire n3191;
wire n3192;
wire n3193;
wire n3194;
wire n3195;
wire n3196;
wire n3197;
wire n3198;
wire n3199;
wire n3200;
wire n3201;
wire n3202;
wire n3203;
wire n3204;
wire n3205;
wire n3206;
wire n3207;
wire n3208;
wire n3209;
wire n3210;
wire n3211;
wire n3212;
wire n3213;
wire n3214;
wire n3215;
wire n3216;
wire n3217;
wire n3218;
wire n3219;
wire n3220;
wire n3221;
wire n3222;
wire n3223;
wire n3224;
wire n3225;
wire n3226;
wire n3227;
wire n3228;
wire n3229;
wire n3230;
wire n3231;
wire n3232;
wire n3233;
wire n3234;
wire n3235;
wire n3236;
wire n3237;
wire n3238;
wire n3239;
wire n3240;
wire n3241;
wire n3242;
wire n3243;
wire n3244;
wire n3245;
wire n3246;
wire n3247;
wire n3248;
wire n3249;
wire n3250;
wire n3251;
wire n3252;
wire n3253;
wire n3254;
wire n3255;
wire n3256;
wire n3257;
wire n3258;
wire n3259;
wire n3260;
wire n3261;
wire n3262;
wire n3263;
wire n3264;
wire n3265;
wire n3266;
wire n3267;
wire n3268;
wire n3269;
wire n3270;
wire n3271;
wire n3272;
wire n3273;
wire n3274;
wire n3275;
wire n3276;
wire n3277;
wire n3278;
wire n3279;
wire n3280;
wire n3281;
wire n3282;
wire n3283;
wire n3284;
wire n3285;
wire n3286;
wire n3287;
wire n3288;
wire n3289;
wire n3290;
wire n3291;
wire n3292;
wire n3293;
wire n3294;
wire n3295;
wire n3296;
wire n3297;
wire n3298;
wire n3299;
wire n3300;
wire n3301;
wire n3302;
wire n3303;
wire n3304;
wire n3305;
wire n3306;
wire n3307;
wire n3308;
wire n3309;
wire n3310;
wire n3311;
wire n3312;
wire n3313;
wire n3314;
wire n3315;
wire n3316;
wire n3317;
wire n3318;
wire n3319;
wire n3320;
wire n3321;
wire n3322;
wire n3323;
wire n3324;
wire n3325;
wire n3326;
wire n3327;
wire n3328;
wire n3329;
wire n3330;
wire n3331;
wire n3332;
wire n3333;
wire n3334;
wire n3335;
wire n3336;
wire n3337;
wire n3338;
wire n3339;
wire n3340;
wire n3341;
wire n3342;
wire n3343;
wire n3344;
wire n3345;
wire n3346;
wire n3347;
wire n3348;
wire n3349;
wire n3350;
wire n3351;
wire n3352;
wire n3353;
wire n3354;
wire n3355;
wire n3356;
wire n3357;
wire n3358;
wire n3359;
wire n3360;
wire n3361;
wire n3362;
wire n3363;
wire n3364;
wire n3365;
wire n3366;
wire n3367;
wire n3368;
wire n3369;
wire n3370;
wire n3371;
wire n3372;
wire n3373;
wire n3374;
wire n3375;
wire n3376;
wire n3377;
wire n3378;
wire n3379;
wire n3380;
wire n3381;
wire n3382;
wire n3383;
wire n3384;
wire n3385;
wire n3386;
wire n3387;
wire n3388;
wire n3389;
wire n3390;
wire n3391;
wire n3392;
wire n3393;
wire n3394;
wire n3395;
wire n3396;
wire n3397;
wire n3398;
wire n3399;
wire n3400;
wire n3401;
wire n3402;
wire n3403;
wire n3404;
wire n3405;
wire n3406;
wire n3407;
wire n3408;
wire n3409;
wire n3410;
wire n3411;
wire n3412;
wire n3413;
wire n3414;
wire n3415;
wire n3416;
wire n3417;
wire n3418;
wire n3419;
wire n3420;
wire n3421;
wire n3422;
wire n3423;
wire n3424;
wire n3425;
wire n3426;
wire n3427;
wire n3428;
wire n3429;
wire n3430;
wire n3431;
wire n3432;
wire n3433;
wire n3434;
wire n3435;
wire n3436;
wire n3437;
wire n3438;
wire n3439;
wire n3440;
wire n3441;
wire n3442;
wire n3443;
wire n3444;
wire n3445;
wire n3446;
wire n3447;
wire n3448;
wire n3449;
wire n3450;
wire n3451;
wire n3452;
wire n3453;
wire n3454;
wire n3455;
wire n3456;
wire n3457;
wire n3458;
wire n3459;
wire n3460;
wire n3461;
wire n3462;
wire n3463;
wire n3464;
wire n3465;
wire n3466;
wire n3467;
wire n3468;
wire n3469;
wire n3470;
wire n3471;
wire n3472;
wire n3473;
wire n3474;
wire n3475;
wire n3476;
wire n3477;
wire n3478;
wire n3479;
wire n3480;
wire n3481;
wire n3482;
wire n3483;
wire n3484;
wire n3485;
wire n3486;
wire n3487;
wire n3488;
wire n3489;
wire n3490;
wire n3491;
wire n3492;
xor (out,n0,n1595);
nand (n0,n1,n1594);
or (n1,n2,n110);
not (n2,n3);
nand (n3,n4,n109);
or (n4,n5,n97);
or (n5,n6,n96);
and (n6,n7,n60);
xor (n7,n8,n35);
nand (n8,n9,n25);
or (n9,n10,n18);
not (n10,n11);
nand (n11,n12,n16);
or (n12,n13,n14);
not (n14,n15);
or (n16,n17,n15);
not (n17,n13);
nor (n18,n19,n23);
and (n19,n20,n21);
not (n21,n22);
and (n23,n24,n22);
not (n24,n20);
or (n25,n26,n30);
nand (n26,n27,n18);
or (n27,n28,n29);
and (n28,n21,n13);
and (n29,n22,n17);
nor (n30,n31,n33);
and (n31,n17,n32);
and (n33,n13,n34);
not (n34,n32);
not (n35,n36);
nand (n36,n37,n54);
or (n37,n38,n49);
nand (n38,n39,n44);
nor (n39,n40,n42);
and (n40,n17,n41);
and (n42,n13,n43);
not (n43,n41);
nand (n44,n45,n48);
or (n45,n46,n41);
not (n46,n47);
nand (n48,n46,n41);
nor (n49,n50,n52);
and (n50,n46,n51);
and (n52,n47,n53);
not (n53,n51);
or (n54,n39,n55);
nor (n55,n56,n58);
and (n56,n46,n57);
and (n58,n47,n59);
not (n59,n57);
or (n60,n61,n95);
and (n61,n62,n87);
xor (n62,n63,n81);
nand (n63,n64,n78);
or (n64,n65,n77);
not (n65,n66);
nand (n66,n67,n74);
nor (n67,n68,n72);
and (n68,n69,n71);
not (n69,n70);
and (n72,n70,n73);
not (n73,n71);
nand (n74,n75,n76);
nand (n75,n24,n71);
nand (n76,n20,n73);
not (n77,n67);
nand (n78,n79,n80);
or (n79,n20,n14);
or (n80,n24,n15);
nand (n81,n82,n86);
or (n82,n26,n83);
nor (n83,n84,n85);
and (n84,n17,n57);
and (n85,n13,n59);
or (n86,n18,n30);
nand (n87,n88,n94);
or (n88,n38,n89);
nor (n89,n90,n92);
and (n90,n46,n91);
and (n92,n47,n93);
not (n93,n91);
or (n94,n39,n49);
and (n95,n63,n81);
and (n96,n8,n35);
xor (n97,n98,n36);
xor (n98,n99,n103);
nand (n99,n100,n11);
or (n100,n101,n102);
not (n101,n26);
not (n102,n18);
nand (n103,n104,n105);
or (n104,n38,n55);
or (n105,n39,n106);
nor (n106,n107,n108);
and (n107,n46,n32);
and (n108,n47,n34);
nand (n109,n5,n97);
not (n110,n111);
nand (n111,n112,n1582);
or (n112,n113,n352);
not (n113,n114);
and (n114,n115,n332,n345);
and (n115,n116,n306);
nand (n116,n117,n270);
not (n117,n118);
or (n118,n119,n269);
and (n119,n120,n239);
xor (n120,n121,n167);
or (n121,n122,n166);
and (n122,n123,n146);
xor (n123,n124,n137);
nand (n124,n125,n131);
or (n125,n38,n126);
nor (n126,n127,n129);
and (n127,n46,n128);
and (n129,n47,n130);
not (n130,n128);
or (n131,n132,n39);
nor (n132,n133,n135);
and (n133,n46,n134);
and (n135,n47,n136);
not (n136,n134);
nand (n137,n138,n142);
or (n138,n66,n139);
nor (n139,n140,n141);
and (n140,n24,n91);
and (n141,n20,n93);
or (n142,n67,n143);
nor (n143,n144,n145);
and (n144,n24,n51);
and (n145,n20,n53);
nand (n146,n147,n162);
or (n147,n148,n159);
nand (n148,n149,n156);
nor (n149,n150,n154);
and (n150,n151,n153);
not (n151,n152);
and (n154,n152,n155);
not (n155,n153);
nand (n156,n157,n158);
or (n157,n69,n153);
nand (n158,n69,n153);
nor (n159,n160,n161);
and (n160,n69,n51);
and (n161,n70,n53);
or (n162,n149,n163);
nor (n163,n164,n165);
and (n164,n69,n57);
and (n165,n70,n59);
and (n166,n124,n137);
xor (n167,n168,n219);
xor (n168,n169,n179);
not (n169,n170);
nand (n170,n171,n175);
or (n171,n148,n172);
nor (n172,n173,n174);
and (n173,n69,n32);
and (n174,n70,n34);
or (n175,n149,n176);
nor (n176,n177,n178);
and (n177,n69,n15);
and (n178,n70,n14);
or (n179,n180,n218);
and (n180,n181,n204);
xor (n181,n182,n201);
nand (n182,n183,n197);
or (n183,n184,n192);
not (n184,n185);
nor (n185,n186,n190);
and (n186,n187,n189);
not (n187,n188);
and (n190,n188,n191);
not (n191,n189);
not (n192,n193);
nand (n193,n185,n194);
nand (n194,n195,n196);
or (n195,n189,n151);
nand (n196,n151,n189);
not (n197,n198);
nor (n198,n199,n200);
and (n199,n151,n15);
and (n200,n152,n14);
nand (n201,n202,n203);
or (n202,n148,n163);
or (n203,n149,n172);
nand (n204,n205,n212);
or (n205,n18,n206);
not (n206,n207);
nand (n207,n208,n211);
or (n208,n13,n209);
not (n209,n210);
or (n211,n17,n210);
or (n212,n26,n213);
nor (n213,n214,n216);
and (n214,n17,n215);
and (n216,n13,n217);
not (n217,n215);
and (n218,n182,n201);
xor (n219,n220,n233);
xor (n220,n221,n227);
nand (n221,n222,n223);
or (n222,n38,n132);
or (n223,n39,n224);
nor (n224,n225,n226);
and (n225,n46,n215);
and (n226,n47,n217);
nand (n227,n228,n229);
or (n228,n66,n143);
or (n229,n67,n230);
nor (n230,n231,n232);
and (n231,n24,n57);
and (n232,n20,n59);
nand (n233,n234,n235);
or (n234,n206,n26);
or (n235,n236,n18);
nor (n236,n237,n238);
and (n237,n17,n91);
and (n238,n13,n93);
or (n239,n240,n268);
and (n240,n241,n267);
xor (n241,n242,n266);
or (n242,n243,n265);
and (n243,n244,n259);
xor (n244,n245,n251);
nand (n245,n246,n250);
or (n246,n26,n247);
nor (n247,n248,n249);
and (n248,n134,n17);
and (n249,n13,n136);
or (n250,n213,n18);
nand (n251,n252,n258);
or (n252,n38,n253);
nor (n253,n254,n256);
and (n254,n255,n46);
and (n256,n47,n257);
not (n257,n255);
or (n258,n39,n126);
nand (n259,n260,n264);
or (n260,n193,n261);
nor (n261,n262,n263);
and (n262,n151,n32);
and (n263,n152,n34);
or (n264,n185,n198);
and (n265,n245,n251);
xor (n266,n181,n204);
xor (n267,n123,n146);
and (n268,n242,n266);
and (n269,n121,n167);
not (n270,n271);
xor (n271,n272,n303);
xor (n272,n273,n292);
xor (n273,n274,n286);
xor (n274,n275,n280);
nand (n275,n276,n279);
or (n276,n277,n278);
not (n277,n148);
not (n278,n149);
not (n279,n176);
nand (n280,n281,n282);
or (n281,n66,n230);
or (n282,n67,n283);
nor (n283,n284,n285);
and (n284,n24,n32);
and (n285,n20,n34);
nand (n286,n287,n288);
or (n287,n38,n224);
or (n288,n39,n289);
nor (n289,n290,n291);
and (n290,n46,n210);
and (n291,n47,n209);
xor (n292,n293,n300);
xor (n293,n294,n170);
nand (n294,n295,n296);
or (n295,n26,n236);
or (n296,n18,n297);
nor (n297,n298,n299);
and (n298,n17,n51);
and (n299,n13,n53);
or (n300,n301,n302);
and (n301,n220,n233);
and (n302,n221,n227);
or (n303,n304,n305);
and (n304,n168,n219);
and (n305,n169,n179);
nand (n306,n307,n311);
not (n307,n308);
or (n308,n309,n310);
and (n309,n272,n303);
and (n310,n273,n292);
not (n311,n312);
xor (n312,n313,n329);
xor (n313,n314,n317);
or (n314,n315,n316);
and (n315,n274,n286);
and (n316,n275,n280);
xor (n317,n318,n325);
xor (n318,n319,n322);
nand (n319,n320,n321);
or (n320,n26,n297);
or (n321,n83,n18);
nand (n322,n323,n324);
or (n323,n38,n289);
or (n324,n39,n89);
nor (n325,n326,n328);
and (n326,n65,n327);
not (n327,n283);
and (n328,n77,n78);
or (n329,n330,n331);
and (n330,n293,n300);
and (n331,n294,n170);
nand (n332,n333,n337);
not (n333,n334);
or (n334,n335,n336);
and (n335,n313,n329);
and (n336,n314,n317);
not (n337,n338);
xor (n338,n339,n342);
xor (n339,n340,n341);
not (n340,n325);
xor (n341,n62,n87);
or (n342,n343,n344);
and (n343,n318,n325);
and (n344,n319,n322);
nand (n345,n346,n350);
not (n346,n347);
or (n347,n348,n349);
and (n348,n339,n342);
and (n349,n340,n341);
not (n350,n351);
xor (n351,n7,n60);
not (n352,n353);
nand (n353,n354,n1077);
nor (n354,n355,n1065);
and (n355,n356,n968);
not (n356,n357);
nor (n357,n358,n967);
and (n358,n359,n900);
nand (n359,n360,n740);
not (n360,n361);
and (n361,n362,n672);
xor (n362,n363,n597);
xor (n363,n364,n478);
xor (n364,n365,n428);
xor (n365,n366,n405);
or (n366,n367,n404);
and (n367,n368,n391);
xor (n368,n369,n378);
nand (n369,n370,n374);
or (n370,n193,n371);
nor (n371,n372,n373);
and (n372,n151,n210);
and (n373,n152,n209);
or (n374,n185,n375);
nor (n375,n376,n377);
and (n376,n151,n91);
and (n377,n152,n93);
nand (n378,n379,n385);
or (n379,n26,n380);
nor (n380,n381,n383);
and (n381,n382,n17);
and (n383,n13,n384);
not (n384,n382);
or (n385,n386,n18);
nor (n386,n387,n389);
and (n387,n388,n17);
and (n389,n13,n390);
not (n390,n388);
nand (n391,n392,n398);
or (n392,n38,n393);
nor (n393,n394,n396);
and (n394,n395,n46);
and (n396,n47,n397);
not (n397,n395);
or (n398,n399,n39);
nor (n399,n400,n402);
and (n400,n401,n46);
and (n402,n47,n403);
not (n403,n401);
and (n404,n369,n378);
xor (n405,n406,n422);
xor (n406,n407,n416);
nand (n407,n408,n412);
or (n408,n66,n409);
nor (n409,n410,n411);
and (n410,n128,n24);
and (n411,n20,n130);
or (n412,n413,n67);
nor (n413,n414,n415);
and (n414,n134,n24);
and (n415,n20,n136);
nand (n416,n417,n418);
or (n417,n193,n375);
or (n418,n185,n419);
nor (n419,n420,n421);
and (n420,n151,n51);
and (n421,n152,n53);
nand (n422,n423,n424);
or (n423,n26,n386);
or (n424,n425,n18);
nor (n425,n426,n427);
and (n426,n255,n17);
and (n427,n13,n257);
xor (n428,n429,n468);
xor (n429,n430,n450);
nand (n430,n431,n445);
or (n431,n432,n438);
nand (n432,n433,n437);
or (n433,n434,n436);
not (n434,n435);
nand (n437,n434,n436);
not (n438,n439);
nand (n439,n440,n441);
not (n440,n432);
nand (n441,n442,n444);
or (n442,n434,n443);
nand (n444,n443,n434);
not (n445,n446);
nor (n446,n447,n449);
and (n447,n448,n15);
not (n448,n443);
and (n449,n443,n14);
nand (n450,n451,n464);
or (n451,n452,n461);
nand (n452,n453,n458);
nor (n453,n454,n457);
and (n454,n455,n443);
not (n455,n456);
and (n457,n456,n448);
nand (n458,n459,n460);
or (n459,n456,n187);
nand (n460,n187,n456);
nor (n461,n462,n463);
and (n462,n187,n57);
and (n463,n188,n59);
or (n464,n453,n465);
nor (n465,n466,n467);
and (n466,n187,n32);
and (n467,n188,n34);
nand (n468,n469,n474);
or (n469,n470,n149);
not (n470,n471);
nand (n471,n472,n473);
or (n472,n70,n209);
or (n473,n69,n210);
or (n474,n148,n475);
nor (n475,n476,n477);
and (n476,n69,n215);
and (n477,n70,n217);
xor (n478,n479,n567);
xor (n479,n480,n517);
xor (n480,n481,n494);
xor (n481,n482,n488);
nand (n482,n483,n484);
or (n483,n38,n399);
or (n484,n485,n39);
nor (n485,n486,n487);
and (n486,n46,n382);
and (n487,n47,n384);
nand (n488,n489,n493);
or (n489,n439,n490);
nor (n490,n491,n492);
and (n491,n448,n32);
and (n492,n443,n34);
or (n493,n440,n446);
or (n494,n495,n516);
and (n495,n496,n510);
xor (n496,n497,n504);
nand (n497,n498,n503);
or (n498,n499,n452);
not (n499,n500);
nand (n500,n501,n502);
or (n501,n188,n53);
or (n502,n187,n51);
or (n503,n453,n461);
nand (n504,n505,n509);
or (n505,n148,n506);
nor (n506,n507,n508);
and (n507,n69,n134);
and (n508,n70,n136);
or (n509,n149,n475);
nand (n510,n511,n515);
or (n511,n66,n512);
nor (n512,n513,n514);
and (n513,n255,n24);
and (n514,n20,n257);
or (n515,n67,n409);
and (n516,n497,n504);
or (n517,n518,n566);
and (n518,n519,n541);
xor (n519,n520,n521);
not (n520,n488);
nand (n521,n522,n534);
not (n522,n523);
nand (n523,n524,n529);
or (n524,n525,n528);
not (n525,n526);
nand (n526,n527,n436);
not (n527,n528);
not (n529,n530);
nor (n530,n531,n533);
and (n531,n532,n15);
not (n532,n436);
and (n533,n436,n14);
not (n534,n535);
nand (n535,n536,n540);
or (n536,n439,n537);
nor (n537,n538,n539);
and (n538,n448,n57);
and (n539,n443,n59);
or (n540,n440,n490);
or (n541,n542,n565);
and (n542,n543,n558);
xor (n543,n544,n552);
nand (n544,n545,n551);
or (n545,n38,n546);
nor (n546,n547,n549);
and (n547,n548,n46);
and (n549,n550,n47);
not (n550,n548);
or (n551,n393,n39);
nand (n552,n553,n557);
or (n553,n193,n554);
nor (n554,n555,n556);
and (n555,n151,n215);
and (n556,n152,n217);
or (n557,n185,n371);
nand (n558,n559,n564);
or (n559,n148,n560);
not (n560,n561);
nor (n561,n562,n563);
and (n562,n130,n69);
and (n563,n128,n70);
or (n564,n506,n149);
and (n565,n544,n552);
and (n566,n520,n521);
or (n567,n568,n596);
and (n568,n569,n595);
xor (n569,n570,n594);
or (n570,n571,n593);
and (n571,n572,n587);
xor (n572,n573,n581);
nand (n573,n574,n575);
or (n574,n453,n499);
nand (n575,n576,n580);
not (n576,n577);
nor (n577,n578,n579);
and (n578,n91,n187);
and (n579,n93,n188);
not (n580,n452);
nand (n581,n582,n586);
or (n582,n66,n583);
nor (n583,n584,n585);
and (n584,n388,n24);
and (n585,n20,n390);
or (n586,n512,n67);
nand (n587,n588,n592);
or (n588,n26,n589);
nor (n589,n590,n591);
and (n590,n401,n17);
and (n591,n13,n403);
or (n592,n380,n18);
and (n593,n573,n581);
xor (n594,n368,n391);
xor (n595,n496,n510);
and (n596,n570,n594);
or (n597,n598,n671);
and (n598,n599,n663);
xor (n599,n600,n662);
or (n600,n601,n661);
and (n601,n602,n639);
xor (n602,n603,n617);
and (n603,n604,n611);
nor (n604,n605,n46);
nor (n605,n606,n609);
and (n606,n607,n17);
nand (n607,n608,n41);
and (n609,n610,n43);
not (n610,n608);
nand (n611,n612,n616);
or (n612,n613,n526);
nor (n613,n614,n615);
and (n614,n32,n532);
and (n615,n34,n436);
or (n616,n530,n527);
or (n617,n618,n638);
and (n618,n619,n632);
xor (n619,n620,n626);
nand (n620,n621,n625);
or (n621,n439,n622);
nor (n622,n623,n624);
and (n623,n448,n51);
and (n624,n443,n53);
or (n625,n440,n537);
nand (n626,n627,n631);
or (n627,n38,n628);
nor (n628,n629,n630);
and (n629,n610,n47);
and (n630,n608,n46);
or (n631,n546,n39);
nand (n632,n633,n637);
or (n633,n193,n634);
nor (n634,n635,n636);
and (n635,n151,n134);
and (n636,n152,n136);
or (n637,n185,n554);
and (n638,n620,n626);
or (n639,n640,n660);
and (n640,n641,n654);
xor (n641,n642,n648);
nand (n642,n643,n644);
or (n643,n149,n560);
or (n644,n148,n645);
nor (n645,n646,n647);
and (n646,n69,n255);
and (n647,n70,n257);
nand (n648,n649,n653);
or (n649,n452,n650);
nor (n650,n651,n652);
and (n651,n187,n210);
and (n652,n188,n209);
or (n653,n453,n577);
nand (n654,n655,n659);
or (n655,n66,n656);
nor (n656,n657,n658);
and (n657,n24,n382);
and (n658,n20,n384);
or (n659,n67,n583);
and (n660,n642,n648);
and (n661,n603,n617);
xor (n662,n519,n541);
or (n663,n664,n670);
and (n664,n665,n669);
xor (n665,n666,n667);
xor (n666,n572,n587);
nand (n667,n668,n521);
or (n668,n522,n534);
xor (n669,n543,n558);
and (n670,n666,n667);
and (n671,n600,n662);
or (n672,n673,n739);
and (n673,n674,n738);
xor (n674,n675,n676);
xor (n675,n569,n595);
or (n676,n677,n737);
and (n677,n678,n709);
xor (n678,n679,n708);
or (n679,n680,n707);
and (n680,n681,n690);
xor (n681,n682,n689);
nand (n682,n683,n688);
or (n683,n26,n684);
not (n684,n685);
nand (n685,n686,n687);
or (n686,n397,n13);
or (n687,n17,n395);
or (n688,n589,n18);
xor (n689,n604,n611);
or (n690,n691,n706);
and (n691,n692,n700);
xor (n692,n693,n694);
nor (n693,n39,n610);
nand (n694,n695,n699);
or (n695,n696,n526);
nor (n696,n697,n698);
and (n697,n436,n59);
nor (n698,n436,n59);
or (n699,n613,n527);
nand (n700,n701,n705);
or (n701,n439,n702);
nor (n702,n703,n704);
and (n703,n448,n91);
and (n704,n443,n93);
or (n705,n440,n622);
and (n706,n693,n694);
and (n707,n682,n689);
xor (n708,n602,n639);
or (n709,n710,n736);
and (n710,n711,n735);
xor (n711,n712,n734);
or (n712,n713,n733);
and (n713,n714,n727);
xor (n714,n715,n721);
nand (n715,n716,n720);
or (n716,n193,n717);
nor (n717,n718,n719);
and (n718,n128,n151);
and (n719,n152,n130);
or (n720,n634,n185);
nand (n721,n722,n726);
or (n722,n148,n723);
nor (n723,n724,n725);
and (n724,n69,n388);
and (n725,n70,n390);
or (n726,n645,n149);
nand (n727,n728,n732);
or (n728,n452,n729);
nor (n729,n730,n731);
and (n730,n187,n215);
and (n731,n188,n217);
or (n732,n453,n650);
and (n733,n715,n721);
xor (n734,n641,n654);
xor (n735,n619,n632);
and (n736,n712,n734);
and (n737,n679,n708);
xor (n738,n599,n663);
and (n739,n675,n676);
nand (n740,n741,n899);
nand (n741,n742,n898);
or (n742,n743,n836);
nor (n743,n744,n745);
xor (n744,n674,n738);
or (n745,n746,n835);
and (n746,n747,n834);
xor (n747,n748,n749);
xor (n748,n665,n669);
or (n749,n750,n833);
and (n750,n751,n782);
xor (n751,n752,n781);
or (n752,n753,n780);
and (n753,n754,n768);
xor (n754,n755,n761);
nand (n755,n756,n760);
or (n756,n66,n757);
nor (n757,n758,n759);
and (n758,n401,n24);
and (n759,n20,n403);
or (n760,n67,n656);
nand (n761,n762,n763);
or (n762,n18,n684);
nand (n763,n764,n101);
not (n764,n765);
nor (n765,n766,n767);
and (n766,n17,n548);
and (n767,n550,n13);
and (n768,n769,n774);
nor (n769,n770,n17);
nor (n770,n771,n773);
and (n771,n772,n24);
nand (n772,n22,n608);
and (n773,n610,n21);
nand (n774,n775,n779);
or (n775,n776,n526);
nor (n776,n777,n778);
and (n777,n532,n51);
and (n778,n436,n53);
or (n779,n696,n527);
and (n780,n755,n761);
xor (n781,n681,n690);
or (n782,n783,n832);
and (n783,n784,n831);
xor (n784,n785,n809);
or (n785,n786,n808);
and (n786,n787,n801);
xor (n787,n788,n794);
nand (n788,n789,n793);
or (n789,n439,n790);
nor (n790,n791,n792);
and (n791,n210,n448);
and (n792,n209,n443);
or (n793,n440,n702);
nand (n794,n795,n800);
or (n795,n796,n193);
not (n796,n797);
nand (n797,n798,n799);
or (n798,n152,n257);
or (n799,n151,n255);
or (n800,n717,n185);
nand (n801,n802,n807);
or (n802,n148,n803);
not (n803,n804);
nor (n804,n805,n806);
and (n805,n384,n69);
and (n806,n382,n70);
or (n807,n723,n149);
and (n808,n788,n794);
or (n809,n810,n830);
and (n810,n811,n824);
xor (n811,n812,n818);
nand (n812,n813,n817);
or (n813,n452,n814);
nor (n814,n815,n816);
and (n815,n187,n134);
and (n816,n188,n136);
or (n817,n453,n729);
nand (n818,n819,n823);
or (n819,n66,n820);
nor (n820,n821,n822);
and (n821,n395,n24);
and (n822,n20,n397);
or (n823,n757,n67);
nand (n824,n825,n829);
or (n825,n26,n826);
nor (n826,n827,n828);
and (n827,n610,n13);
and (n828,n608,n17);
or (n829,n765,n18);
and (n830,n812,n818);
xor (n831,n692,n700);
and (n832,n785,n809);
and (n833,n752,n781);
xor (n834,n678,n709);
and (n835,n748,n749);
nand (n836,n837,n838);
xor (n837,n747,n834);
or (n838,n839,n897);
and (n839,n840,n896);
xor (n840,n841,n842);
xor (n841,n711,n735);
or (n842,n843,n895);
and (n843,n844,n847);
xor (n844,n845,n846);
xor (n845,n714,n727);
xor (n846,n754,n768);
or (n847,n848,n894);
and (n848,n849,n871);
xor (n849,n850,n851);
xor (n850,n769,n774);
or (n851,n852,n870);
and (n852,n853,n863);
xor (n853,n854,n855);
and (n854,n102,n608);
nand (n855,n856,n861);
or (n856,n857,n439);
not (n857,n858);
nand (n858,n859,n860);
or (n859,n443,n217);
or (n860,n448,n215);
nand (n861,n862,n432);
not (n862,n790);
nand (n863,n864,n869);
or (n864,n193,n865);
not (n865,n866);
nand (n866,n867,n868);
or (n867,n152,n390);
or (n868,n151,n388);
or (n869,n185,n796);
and (n870,n854,n855);
or (n871,n872,n893);
and (n872,n873,n887);
xor (n873,n874,n881);
nand (n874,n875,n880);
or (n875,n876,n148);
not (n876,n877);
nand (n877,n878,n879);
or (n878,n70,n403);
or (n879,n69,n401);
nand (n880,n804,n278);
nand (n881,n882,n883);
or (n882,n527,n776);
or (n883,n884,n526);
nor (n884,n885,n886);
and (n885,n532,n91);
and (n886,n436,n93);
nand (n887,n888,n892);
or (n888,n889,n66);
nor (n889,n890,n891);
and (n890,n548,n24);
and (n891,n20,n550);
or (n892,n820,n67);
and (n893,n874,n881);
and (n894,n850,n851);
and (n895,n845,n846);
xor (n896,n751,n782);
and (n897,n841,n842);
nand (n898,n744,n745);
or (n899,n362,n672);
or (n900,n901,n904);
or (n901,n902,n903);
and (n902,n363,n597);
and (n903,n364,n478);
xor (n904,n905,n964);
xor (n905,n906,n934);
xor (n906,n907,n914);
xor (n907,n908,n911);
or (n908,n909,n910);
and (n909,n406,n422);
and (n910,n407,n416);
or (n911,n912,n913);
and (n912,n429,n468);
and (n913,n430,n450);
xor (n914,n915,n928);
xor (n915,n916,n922);
nand (n916,n917,n918);
or (n917,n66,n413);
or (n918,n67,n919);
nor (n919,n920,n921);
and (n920,n24,n215);
and (n921,n20,n217);
nand (n922,n923,n924);
or (n923,n26,n425);
or (n924,n925,n18);
nor (n925,n926,n927);
and (n926,n17,n128);
and (n927,n13,n130);
nand (n928,n929,n930);
or (n929,n452,n465);
or (n930,n453,n931);
nor (n931,n932,n933);
and (n932,n187,n15);
and (n933,n188,n14);
xor (n934,n935,n961);
xor (n935,n936,n958);
xor (n936,n937,n951);
xor (n937,n938,n944);
nand (n938,n939,n940);
or (n939,n38,n485);
or (n940,n941,n39);
nor (n941,n942,n943);
and (n942,n388,n46);
and (n943,n47,n390);
nand (n944,n945,n946);
or (n945,n470,n148);
nand (n946,n947,n278);
not (n947,n948);
nor (n948,n949,n950);
and (n949,n69,n91);
and (n950,n70,n93);
not (n951,n952);
nand (n952,n953,n954);
or (n953,n193,n419);
or (n954,n185,n955);
nor (n955,n956,n957);
and (n956,n151,n57);
and (n957,n152,n59);
or (n958,n959,n960);
and (n959,n481,n494);
and (n960,n482,n488);
or (n961,n962,n963);
and (n962,n365,n428);
and (n963,n366,n405);
or (n964,n965,n966);
and (n965,n479,n567);
and (n966,n480,n517);
and (n967,n904,n901);
not (n968,n969);
nand (n969,n970,n1041,n1060);
not (n970,n971);
nor (n971,n972,n1019);
xor (n972,n973,n999);
xor (n973,n974,n998);
or (n974,n975,n997);
and (n975,n976,n984);
xor (n976,n977,n983);
nand (n977,n978,n982);
or (n978,n66,n979);
nor (n979,n980,n981);
and (n980,n24,n210);
and (n981,n20,n209);
or (n982,n67,n139);
not (n983,n146);
or (n984,n985,n996);
and (n985,n986,n993);
xor (n986,n987,n990);
nand (n987,n988,n989);
or (n988,n26,n925);
or (n989,n247,n18);
nand (n990,n991,n992);
or (n991,n148,n948);
or (n992,n149,n159);
nand (n993,n994,n995);
or (n994,n38,n941);
or (n995,n253,n39);
and (n996,n987,n990);
and (n997,n977,n983);
xor (n998,n241,n267);
or (n999,n1000,n1018);
and (n1000,n1001,n1017);
xor (n1001,n1002,n1016);
or (n1002,n1003,n1015);
and (n1003,n1004,n1012);
xor (n1004,n1005,n1009);
nand (n1005,n1006,n1008);
or (n1006,n580,n1007);
not (n1007,n453);
not (n1008,n931);
nand (n1009,n1010,n1011);
or (n1010,n193,n955);
or (n1011,n185,n261);
nand (n1012,n1013,n1014);
or (n1013,n66,n919);
or (n1014,n67,n979);
and (n1015,n1005,n1009);
xor (n1016,n244,n259);
xor (n1017,n976,n984);
and (n1018,n1002,n1016);
or (n1019,n1020,n1040);
and (n1020,n1021,n1031);
xor (n1021,n1022,n1030);
or (n1022,n1023,n1029);
and (n1023,n1024,n1028);
xor (n1024,n952,n1025);
or (n1025,n1026,n1027);
and (n1026,n915,n928);
and (n1027,n916,n922);
xor (n1028,n986,n993);
and (n1029,n952,n1025);
xor (n1030,n1001,n1017);
or (n1031,n1032,n1039);
and (n1032,n1033,n1038);
xor (n1033,n1034,n1035);
xor (n1034,n1004,n1012);
or (n1035,n1036,n1037);
and (n1036,n937,n951);
and (n1037,n938,n944);
xor (n1038,n1024,n1028);
and (n1039,n1034,n1035);
and (n1040,n1022,n1030);
nor (n1041,n1042,n1055);
nor (n1042,n1043,n1046);
or (n1043,n1044,n1045);
and (n1044,n905,n964);
and (n1045,n906,n934);
xor (n1046,n1047,n1052);
xor (n1047,n1048,n1051);
or (n1048,n1049,n1050);
and (n1049,n907,n914);
and (n1050,n908,n911);
xor (n1051,n1033,n1038);
or (n1052,n1053,n1054);
and (n1053,n935,n961);
and (n1054,n936,n958);
nor (n1055,n1056,n1059);
or (n1056,n1057,n1058);
and (n1057,n1047,n1052);
and (n1058,n1048,n1051);
xor (n1059,n1021,n1031);
or (n1060,n1061,n1064);
or (n1061,n1062,n1063);
and (n1062,n973,n999);
and (n1063,n974,n998);
xor (n1064,n120,n239);
nand (n1065,n1066,n1076);
or (n1066,n1067,n1068);
not (n1067,n1060);
not (n1068,n1069);
nand (n1069,n1070,n1075);
nand (n1070,n970,n1071);
nand (n1071,n1072,n1074);
or (n1072,n1073,n1055);
nand (n1073,n1043,n1046);
nand (n1074,n1056,n1059);
nand (n1075,n1019,n972);
nand (n1076,n1061,n1064);
nand (n1077,n1078,n1578);
or (n1078,n1079,n1577);
and (n1079,n1080,n1143);
xor (n1080,n1081,n1142);
or (n1081,n1082,n1141);
and (n1082,n1083,n1086);
xor (n1083,n1084,n1085);
xor (n1084,n784,n831);
xor (n1085,n844,n847);
or (n1086,n1087,n1140);
and (n1087,n1088,n1091);
xor (n1088,n1089,n1090);
xor (n1089,n811,n824);
xor (n1090,n787,n801);
or (n1091,n1092,n1139);
and (n1092,n1093,n1114);
xor (n1093,n1094,n1100);
nand (n1094,n1095,n1099);
or (n1095,n452,n1096);
nor (n1096,n1097,n1098);
and (n1097,n187,n128);
and (n1098,n188,n130);
or (n1099,n453,n814);
nor (n1100,n1101,n1108);
not (n1101,n1102);
nand (n1102,n1103,n1107);
or (n1103,n1104,n439);
nor (n1104,n1105,n1106);
and (n1105,n134,n448);
and (n1106,n136,n443);
nand (n1107,n432,n858);
nand (n1108,n1109,n20);
nand (n1109,n1110,n1111);
or (n1110,n608,n71);
nand (n1111,n1112,n69);
not (n1112,n1113);
and (n1113,n608,n71);
or (n1114,n1115,n1138);
and (n1115,n1116,n1131);
xor (n1116,n1117,n1124);
nand (n1117,n1118,n1119);
or (n1118,n185,n865);
nand (n1119,n1120,n192);
not (n1120,n1121);
nor (n1121,n1122,n1123);
and (n1122,n384,n152);
and (n1123,n382,n151);
nand (n1124,n1125,n1130);
or (n1125,n1126,n148);
not (n1126,n1127);
nor (n1127,n1128,n1129);
and (n1128,n69,n397);
and (n1129,n70,n395);
nand (n1130,n278,n877);
nand (n1131,n1132,n1137);
or (n1132,n1133,n526);
not (n1133,n1134);
or (n1134,n1135,n1136);
and (n1135,n209,n436);
and (n1136,n210,n532);
or (n1137,n884,n527);
and (n1138,n1117,n1124);
and (n1139,n1094,n1100);
and (n1140,n1089,n1090);
and (n1141,n1084,n1085);
xor (n1142,n840,n896);
or (n1143,n1144,n1576);
and (n1144,n1145,n1179);
xor (n1145,n1146,n1178);
or (n1146,n1147,n1177);
and (n1147,n1148,n1176);
xor (n1148,n1149,n1150);
xor (n1149,n849,n871);
or (n1150,n1151,n1175);
and (n1151,n1152,n1155);
xor (n1152,n1153,n1154);
xor (n1153,n873,n887);
xor (n1154,n853,n863);
or (n1155,n1156,n1174);
and (n1156,n1157,n1170);
xor (n1157,n1158,n1164);
nand (n1158,n1159,n1163);
or (n1159,n66,n1160);
nor (n1160,n1161,n1162);
and (n1161,n610,n20);
and (n1162,n608,n24);
or (n1163,n889,n67);
nand (n1164,n1165,n1169);
or (n1165,n452,n1166);
nor (n1166,n1167,n1168);
and (n1167,n187,n255);
and (n1168,n188,n257);
or (n1169,n453,n1096);
nand (n1170,n1171,n1173);
or (n1171,n1172,n1101);
not (n1172,n1108);
or (n1173,n1102,n1108);
and (n1174,n1158,n1164);
and (n1175,n1153,n1154);
xor (n1176,n1088,n1091);
and (n1177,n1149,n1150);
xor (n1178,n1083,n1086);
nand (n1179,n1180,n1572);
or (n1180,n1181,n1550);
nor (n1181,n1182,n1549);
and (n1182,n1183,n1530);
or (n1183,n1184,n1529);
and (n1184,n1185,n1327);
xor (n1185,n1186,n1296);
or (n1186,n1187,n1295);
and (n1187,n1188,n1258);
xor (n1188,n1189,n1219);
xor (n1189,n1190,n1209);
xor (n1190,n1191,n1200);
nand (n1191,n1192,n1196);
or (n1192,n193,n1193);
nor (n1193,n1194,n1195);
and (n1194,n395,n151);
and (n1195,n397,n152);
or (n1196,n1197,n185);
nor (n1197,n1198,n1199);
and (n1198,n151,n401);
and (n1199,n152,n403);
nand (n1200,n1201,n1205);
or (n1201,n148,n1202);
nor (n1202,n1203,n1204);
and (n1203,n610,n70);
and (n1204,n608,n69);
or (n1205,n1206,n149);
nor (n1206,n1207,n1208);
and (n1207,n548,n69);
and (n1208,n550,n70);
nand (n1209,n1210,n1215);
or (n1210,n526,n1211);
not (n1211,n1212);
nor (n1212,n1213,n1214);
and (n1213,n134,n436);
and (n1214,n136,n532);
or (n1215,n1216,n527);
nor (n1216,n1217,n1218);
and (n1217,n215,n532);
and (n1218,n217,n436);
or (n1219,n1220,n1257);
and (n1220,n1221,n1240);
xor (n1221,n1222,n1231);
nand (n1222,n1223,n1227);
or (n1223,n439,n1224);
nor (n1224,n1225,n1226);
and (n1225,n448,n388);
and (n1226,n443,n390);
or (n1227,n440,n1228);
nor (n1228,n1229,n1230);
and (n1229,n257,n443);
and (n1230,n255,n448);
nand (n1231,n1232,n1236);
or (n1232,n452,n1233);
nor (n1233,n1234,n1235);
and (n1234,n401,n187);
and (n1235,n188,n403);
or (n1236,n453,n1237);
nor (n1237,n1238,n1239);
and (n1238,n187,n382);
and (n1239,n188,n384);
and (n1240,n1241,n1247);
nor (n1241,n1242,n151);
nor (n1242,n1243,n1246);
and (n1243,n1244,n187);
not (n1244,n1245);
and (n1245,n608,n189);
and (n1246,n610,n191);
nand (n1247,n1248,n1253);
or (n1248,n1249,n526);
not (n1249,n1250);
nor (n1250,n1251,n1252);
and (n1251,n257,n532);
and (n1252,n255,n436);
or (n1253,n1254,n527);
nor (n1254,n1255,n1256);
and (n1255,n128,n532);
and (n1256,n130,n436);
and (n1257,n1222,n1231);
xor (n1258,n1259,n1280);
xor (n1259,n1260,n1266);
nand (n1260,n1261,n1262);
or (n1261,n452,n1237);
or (n1262,n453,n1263);
nor (n1263,n1264,n1265);
and (n1264,n187,n388);
and (n1265,n188,n390);
xor (n1266,n1267,n1272);
nor (n1267,n1268,n69);
nor (n1268,n1269,n1271);
and (n1269,n1270,n151);
nand (n1270,n608,n153);
and (n1271,n610,n155);
nand (n1272,n1273,n1278);
or (n1273,n440,n1274);
not (n1274,n1275);
nand (n1275,n1276,n1277);
or (n1276,n443,n130);
or (n1277,n448,n128);
nand (n1278,n1279,n438);
not (n1279,n1228);
or (n1280,n1281,n1294);
and (n1281,n1282,n1287);
xor (n1282,n1283,n1284);
nor (n1283,n149,n610);
nand (n1284,n1285,n1286);
or (n1285,n527,n1211);
or (n1286,n1254,n526);
nand (n1287,n1288,n1289);
or (n1288,n185,n1193);
nand (n1289,n1290,n192);
not (n1290,n1291);
or (n1291,n1292,n1293);
and (n1292,n550,n151);
and (n1293,n548,n152);
and (n1294,n1283,n1284);
and (n1295,n1189,n1219);
xor (n1296,n1297,n1312);
xor (n1297,n1298,n1309);
xor (n1298,n1299,n1306);
xor (n1299,n1300,n1303);
nand (n1300,n1301,n1302);
or (n1301,n149,n1126);
or (n1302,n148,n1206);
nand (n1303,n1304,n1305);
or (n1304,n1216,n526);
nand (n1305,n1134,n528);
nand (n1306,n1307,n1308);
or (n1307,n452,n1263);
or (n1308,n453,n1166);
or (n1309,n1310,n1311);
and (n1310,n1259,n1280);
and (n1311,n1260,n1266);
xor (n1312,n1313,n1318);
xor (n1313,n1314,n1315);
and (n1314,n1267,n1272);
or (n1315,n1316,n1317);
and (n1316,n1190,n1209);
and (n1317,n1191,n1200);
xor (n1318,n1319,n1324);
xor (n1319,n1320,n1321);
nor (n1320,n67,n610);
nand (n1321,n1322,n1323);
or (n1322,n1274,n439);
or (n1323,n440,n1104);
nand (n1324,n1325,n1326);
or (n1325,n193,n1197);
or (n1326,n185,n1121);
nand (n1327,n1328,n1525,n1528);
nand (n1328,n1329,n1383,n1518);
not (n1329,n1330);
nor (n1330,n1331,n1358);
xor (n1331,n1332,n1357);
xor (n1332,n1333,n1356);
or (n1333,n1334,n1355);
and (n1334,n1335,n1349);
xor (n1335,n1336,n1342);
nand (n1336,n1337,n1341);
or (n1337,n193,n1338);
nor (n1338,n1339,n1340);
and (n1339,n610,n152);
and (n1340,n608,n151);
or (n1341,n1291,n185);
nand (n1342,n1343,n1348);
or (n1343,n1344,n439);
not (n1344,n1345);
nor (n1345,n1346,n1347);
and (n1346,n382,n443);
and (n1347,n384,n448);
or (n1348,n440,n1224);
nand (n1349,n1350,n1354);
or (n1350,n452,n1351);
nor (n1351,n1352,n1353);
and (n1352,n395,n187);
and (n1353,n188,n397);
or (n1354,n453,n1233);
and (n1355,n1336,n1342);
xor (n1356,n1282,n1287);
xor (n1357,n1221,n1240);
or (n1358,n1359,n1382);
and (n1359,n1360,n1381);
xor (n1360,n1361,n1362);
xor (n1361,n1241,n1247);
or (n1362,n1363,n1380);
and (n1363,n1364,n1373);
xor (n1364,n1365,n1366);
and (n1365,n184,n608);
nand (n1366,n1367,n1372);
or (n1367,n526,n1368);
not (n1368,n1369);
nor (n1369,n1370,n1371);
and (n1370,n390,n532);
and (n1371,n388,n436);
nand (n1372,n1250,n528);
nand (n1373,n1374,n1379);
or (n1374,n1375,n439);
not (n1375,n1376);
nor (n1376,n1377,n1378);
and (n1377,n403,n448);
and (n1378,n401,n443);
nand (n1379,n1345,n432);
and (n1380,n1365,n1366);
xor (n1381,n1335,n1349);
and (n1382,n1361,n1362);
or (n1383,n1384,n1517);
and (n1384,n1385,n1411);
xor (n1385,n1386,n1410);
or (n1386,n1387,n1409);
and (n1387,n1388,n1408);
xor (n1388,n1389,n1395);
nand (n1389,n1390,n1394);
or (n1390,n452,n1391);
nor (n1391,n1392,n1393);
and (n1392,n187,n548);
and (n1393,n188,n550);
or (n1394,n1351,n453);
and (n1395,n1396,n1402);
and (n1396,n1397,n188);
nand (n1397,n1398,n1399);
or (n1398,n608,n456);
nand (n1399,n1400,n448);
not (n1400,n1401);
and (n1401,n608,n456);
nand (n1402,n1403,n1404);
or (n1403,n527,n1368);
or (n1404,n1405,n526);
nor (n1405,n1406,n1407);
and (n1406,n532,n382);
and (n1407,n436,n384);
xor (n1408,n1364,n1373);
and (n1409,n1389,n1395);
xor (n1410,n1360,n1381);
nand (n1411,n1412,n1516);
or (n1412,n1413,n1511);
nor (n1413,n1414,n1510);
and (n1414,n1415,n1489);
nand (n1415,n1416,n1487);
or (n1416,n1417,n1471);
not (n1417,n1418);
or (n1418,n1419,n1470);
and (n1419,n1420,n1449);
xor (n1420,n1421,n1430);
nand (n1421,n1422,n1426);
or (n1422,n439,n1423);
nor (n1423,n1424,n1425);
and (n1424,n443,n610);
and (n1425,n608,n448);
or (n1426,n440,n1427);
nor (n1427,n1428,n1429);
and (n1428,n550,n443);
and (n1429,n548,n448);
nand (n1430,n1431,n1448);
or (n1431,n1432,n1438);
not (n1432,n1433);
nand (n1433,n1434,n443);
nand (n1434,n1435,n1437);
or (n1435,n1436,n436);
and (n1436,n608,n435);
nand (n1437,n610,n434);
not (n1438,n1439);
nand (n1439,n1440,n1444);
or (n1440,n1441,n526);
or (n1441,n1442,n1443);
and (n1442,n395,n436);
and (n1443,n397,n532);
or (n1444,n1445,n527);
nor (n1445,n1446,n1447);
and (n1446,n403,n436);
and (n1447,n401,n532);
or (n1448,n1439,n1433);
or (n1449,n1450,n1469);
and (n1450,n1451,n1459);
xor (n1451,n1452,n1453);
nor (n1452,n440,n610);
nand (n1453,n1454,n1458);
or (n1454,n1455,n526);
nor (n1455,n1456,n1457);
and (n1456,n550,n436);
and (n1457,n548,n532);
or (n1458,n1441,n527);
nor (n1459,n1460,n1467);
nor (n1460,n1461,n1463);
and (n1461,n1462,n528);
not (n1462,n1455);
and (n1463,n1464,n525);
nand (n1464,n1465,n1466);
or (n1465,n610,n436);
nand (n1466,n436,n610);
or (n1467,n1468,n532);
and (n1468,n608,n528);
and (n1469,n1452,n1453);
and (n1470,n1421,n1430);
not (n1471,n1472);
nand (n1472,n1473,n1486);
not (n1473,n1474);
xor (n1474,n1475,n1483);
xor (n1475,n1476,n1477);
and (n1476,n1007,n608);
nand (n1477,n1478,n1479);
or (n1478,n1427,n439);
nand (n1479,n1480,n432);
nor (n1480,n1481,n1482);
and (n1481,n397,n448);
and (n1482,n395,n443);
nand (n1483,n1484,n1485);
or (n1484,n1445,n526);
or (n1485,n1405,n527);
nand (n1486,n1432,n1439);
nand (n1487,n1488,n1474);
not (n1488,n1486);
nand (n1489,n1490,n1506);
not (n1490,n1491);
xor (n1491,n1492,n1505);
xor (n1492,n1493,n1497);
nand (n1493,n1494,n1496);
or (n1494,n1495,n439);
not (n1495,n1480);
nand (n1496,n1376,n432);
nand (n1497,n1498,n1503);
or (n1498,n1499,n452);
not (n1499,n1500);
nand (n1500,n1501,n1502);
or (n1501,n608,n187);
or (n1502,n610,n188);
nand (n1503,n1504,n1007);
not (n1504,n1391);
xor (n1505,n1396,n1402);
not (n1506,n1507);
or (n1507,n1508,n1509);
and (n1508,n1475,n1483);
and (n1509,n1476,n1477);
nor (n1510,n1490,n1506);
nor (n1511,n1512,n1513);
xor (n1512,n1388,n1408);
or (n1513,n1514,n1515);
and (n1514,n1492,n1505);
and (n1515,n1493,n1497);
nand (n1516,n1512,n1513);
and (n1517,n1386,n1410);
nand (n1518,n1519,n1523);
not (n1519,n1520);
or (n1520,n1521,n1522);
and (n1521,n1332,n1357);
and (n1522,n1333,n1356);
not (n1523,n1524);
xor (n1524,n1188,n1258);
nand (n1525,n1526,n1518);
not (n1526,n1527);
nand (n1527,n1331,n1358);
nand (n1528,n1524,n1520);
and (n1529,n1186,n1296);
or (n1530,n1531,n1546);
xor (n1531,n1532,n1543);
xor (n1532,n1533,n1534);
xor (n1533,n1157,n1170);
xor (n1534,n1535,n1542);
xor (n1535,n1536,n1539);
or (n1536,n1537,n1538);
and (n1537,n1319,n1324);
and (n1538,n1320,n1321);
or (n1539,n1540,n1541);
and (n1540,n1299,n1306);
and (n1541,n1300,n1303);
xor (n1542,n1116,n1131);
or (n1543,n1544,n1545);
and (n1544,n1313,n1318);
and (n1545,n1314,n1315);
or (n1546,n1547,n1548);
and (n1547,n1297,n1312);
and (n1548,n1298,n1309);
and (n1549,n1531,n1546);
nand (n1550,n1551,n1565);
not (n1551,n1552);
and (n1552,n1553,n1561);
not (n1553,n1554);
xor (n1554,n1555,n1560);
xor (n1555,n1556,n1557);
xor (n1556,n1093,n1114);
or (n1557,n1558,n1559);
and (n1558,n1535,n1542);
and (n1559,n1536,n1539);
xor (n1560,n1152,n1155);
not (n1561,n1562);
or (n1562,n1563,n1564);
and (n1563,n1532,n1543);
and (n1564,n1533,n1534);
nand (n1565,n1566,n1568);
not (n1566,n1567);
xor (n1567,n1148,n1176);
not (n1568,n1569);
or (n1569,n1570,n1571);
and (n1570,n1555,n1560);
and (n1571,n1556,n1557);
nor (n1572,n1573,n1575);
and (n1573,n1565,n1574);
nor (n1574,n1553,n1561);
nor (n1575,n1566,n1568);
and (n1576,n1146,n1178);
and (n1577,n1081,n1142);
nor (n1578,n1579,n969);
nand (n1579,n1580,n900,n899);
nor (n1580,n743,n1581);
nor (n1581,n838,n837);
nor (n1582,n1583,n1593);
and (n1583,n1584,n345);
nand (n1584,n1585,n1587);
not (n1585,n1586);
nor (n1586,n333,n337);
nand (n1587,n1588,n332);
not (n1588,n1589);
nor (n1589,n1590,n1592);
and (n1590,n1591,n306);
nor (n1591,n117,n270);
nor (n1592,n307,n311);
nor (n1593,n346,n350);
or (n1594,n111,n3);
xor (n1595,n1596,n3138);
xor (n1596,n1597,n3491);
xor (n1597,n1598,n3133);
xor (n1598,n1599,n3484);
xor (n1599,n1600,n3127);
xor (n1600,n1601,n3472);
xor (n1601,n1602,n3121);
xor (n1602,n1603,n3455);
xor (n1603,n1604,n3115);
xor (n1604,n1605,n3433);
xor (n1605,n1606,n3109);
xor (n1606,n1607,n3406);
xor (n1607,n1608,n3103);
xor (n1608,n1609,n3374);
xor (n1609,n1610,n3097);
xor (n1610,n1611,n3337);
xor (n1611,n1612,n3091);
xor (n1612,n1613,n3295);
xor (n1613,n1614,n3085);
xor (n1614,n1615,n3248);
xor (n1615,n1616,n3079);
xor (n1616,n1617,n3196);
xor (n1617,n1618,n3073);
xor (n1618,n1619,n3139);
xor (n1619,n1620,n3067);
xor (n1620,n1621,n3064);
xor (n1621,n1622,n3063);
xor (n1622,n1623,n2982);
xor (n1623,n1624,n2981);
xor (n1624,n1625,n2894);
xor (n1625,n1626,n2893);
xor (n1626,n1627,n2801);
xor (n1627,n1628,n2800);
xor (n1628,n1629,n2703);
xor (n1629,n1630,n2702);
xor (n1630,n1631,n2601);
xor (n1631,n1632,n2600);
xor (n1632,n1633,n2496);
xor (n1633,n1634,n2495);
xor (n1634,n1635,n2383);
xor (n1635,n1636,n2382);
xor (n1636,n1637,n2266);
xor (n1637,n1638,n2265);
xor (n1638,n1639,n2144);
xor (n1639,n1640,n2143);
xor (n1640,n1641,n2016);
xor (n1641,n1642,n2015);
xor (n1642,n1643,n1658);
xor (n1643,n1644,n1657);
xor (n1644,n1645,n1656);
xor (n1645,n1646,n1655);
xor (n1646,n1647,n1654);
xor (n1647,n1648,n1653);
xor (n1648,n1649,n1652);
xor (n1649,n1650,n1651);
and (n1650,n15,n528);
and (n1651,n15,n436);
and (n1652,n1650,n1651);
and (n1653,n15,n435);
and (n1654,n1648,n1653);
and (n1655,n15,n443);
and (n1656,n1646,n1655);
and (n1657,n15,n456);
or (n1658,n1659,n1660);
and (n1659,n1644,n1657);
and (n1660,n1643,n1661);
or (n1661,n1659,n1662);
and (n1662,n1643,n1663);
or (n1663,n1659,n1664);
and (n1664,n1643,n1665);
or (n1665,n1659,n1666);
and (n1666,n1643,n1667);
or (n1667,n1659,n1668);
and (n1668,n1643,n1669);
or (n1669,n1659,n1670);
and (n1670,n1643,n1671);
or (n1671,n1659,n1672);
and (n1672,n1643,n1673);
or (n1673,n1659,n1674);
and (n1674,n1643,n1675);
or (n1675,n1659,n1676);
and (n1676,n1643,n1677);
or (n1677,n1678,n1933);
and (n1678,n1679,n1932);
xor (n1679,n1645,n1680);
or (n1680,n1681,n1852);
and (n1681,n1682,n1851);
xor (n1682,n1647,n1683);
or (n1683,n1684,n1769);
and (n1684,n1685,n1768);
xor (n1685,n1649,n1686);
or (n1686,n1687,n1689);
and (n1687,n1650,n1688);
and (n1688,n32,n436);
and (n1689,n1690,n1691);
xor (n1690,n1650,n1688);
or (n1691,n1692,n1695);
and (n1692,n1693,n1694);
and (n1693,n32,n528);
and (n1694,n57,n436);
and (n1695,n1696,n1697);
xor (n1696,n1693,n1694);
or (n1697,n1698,n1701);
and (n1698,n1699,n1700);
and (n1699,n57,n528);
and (n1700,n51,n436);
and (n1701,n1702,n1703);
xor (n1702,n1699,n1700);
or (n1703,n1704,n1707);
and (n1704,n1705,n1706);
and (n1705,n51,n528);
and (n1706,n91,n436);
and (n1707,n1708,n1709);
xor (n1708,n1705,n1706);
or (n1709,n1710,n1713);
and (n1710,n1711,n1712);
and (n1711,n91,n528);
and (n1712,n210,n436);
and (n1713,n1714,n1715);
xor (n1714,n1711,n1712);
or (n1715,n1716,n1719);
and (n1716,n1717,n1718);
and (n1717,n210,n528);
and (n1718,n215,n436);
and (n1719,n1720,n1721);
xor (n1720,n1717,n1718);
or (n1721,n1722,n1724);
and (n1722,n1723,n1213);
and (n1723,n215,n528);
and (n1724,n1725,n1726);
xor (n1725,n1723,n1213);
or (n1726,n1727,n1730);
and (n1727,n1728,n1729);
and (n1728,n134,n528);
and (n1729,n128,n436);
and (n1730,n1731,n1732);
xor (n1731,n1728,n1729);
or (n1732,n1733,n1735);
and (n1733,n1734,n1252);
and (n1734,n128,n528);
and (n1735,n1736,n1737);
xor (n1736,n1734,n1252);
or (n1737,n1738,n1740);
and (n1738,n1739,n1371);
and (n1739,n255,n528);
and (n1740,n1741,n1742);
xor (n1741,n1739,n1371);
or (n1742,n1743,n1746);
and (n1743,n1744,n1745);
and (n1744,n388,n528);
and (n1745,n382,n436);
and (n1746,n1747,n1748);
xor (n1747,n1744,n1745);
or (n1748,n1749,n1752);
and (n1749,n1750,n1751);
and (n1750,n382,n528);
and (n1751,n401,n436);
and (n1752,n1753,n1754);
xor (n1753,n1750,n1751);
or (n1754,n1755,n1757);
and (n1755,n1756,n1442);
and (n1756,n401,n528);
and (n1757,n1758,n1759);
xor (n1758,n1756,n1442);
or (n1759,n1760,n1763);
and (n1760,n1761,n1762);
and (n1761,n395,n528);
and (n1762,n548,n436);
and (n1763,n1764,n1765);
xor (n1764,n1761,n1762);
and (n1765,n1766,n1767);
and (n1766,n548,n528);
and (n1767,n608,n436);
and (n1768,n32,n435);
and (n1769,n1770,n1771);
xor (n1770,n1685,n1768);
or (n1771,n1772,n1775);
and (n1772,n1773,n1774);
xor (n1773,n1690,n1691);
and (n1774,n57,n435);
and (n1775,n1776,n1777);
xor (n1776,n1773,n1774);
or (n1777,n1778,n1781);
and (n1778,n1779,n1780);
xor (n1779,n1696,n1697);
and (n1780,n51,n435);
and (n1781,n1782,n1783);
xor (n1782,n1779,n1780);
or (n1783,n1784,n1787);
and (n1784,n1785,n1786);
xor (n1785,n1702,n1703);
and (n1786,n91,n435);
and (n1787,n1788,n1789);
xor (n1788,n1785,n1786);
or (n1789,n1790,n1793);
and (n1790,n1791,n1792);
xor (n1791,n1708,n1709);
and (n1792,n210,n435);
and (n1793,n1794,n1795);
xor (n1794,n1791,n1792);
or (n1795,n1796,n1799);
and (n1796,n1797,n1798);
xor (n1797,n1714,n1715);
and (n1798,n215,n435);
and (n1799,n1800,n1801);
xor (n1800,n1797,n1798);
or (n1801,n1802,n1805);
and (n1802,n1803,n1804);
xor (n1803,n1720,n1721);
and (n1804,n134,n435);
and (n1805,n1806,n1807);
xor (n1806,n1803,n1804);
or (n1807,n1808,n1811);
and (n1808,n1809,n1810);
xor (n1809,n1725,n1726);
and (n1810,n128,n435);
and (n1811,n1812,n1813);
xor (n1812,n1809,n1810);
or (n1813,n1814,n1817);
and (n1814,n1815,n1816);
xor (n1815,n1731,n1732);
and (n1816,n255,n435);
and (n1817,n1818,n1819);
xor (n1818,n1815,n1816);
or (n1819,n1820,n1823);
and (n1820,n1821,n1822);
xor (n1821,n1736,n1737);
and (n1822,n388,n435);
and (n1823,n1824,n1825);
xor (n1824,n1821,n1822);
or (n1825,n1826,n1829);
and (n1826,n1827,n1828);
xor (n1827,n1741,n1742);
and (n1828,n382,n435);
and (n1829,n1830,n1831);
xor (n1830,n1827,n1828);
or (n1831,n1832,n1835);
and (n1832,n1833,n1834);
xor (n1833,n1747,n1748);
and (n1834,n401,n435);
and (n1835,n1836,n1837);
xor (n1836,n1833,n1834);
or (n1837,n1838,n1841);
and (n1838,n1839,n1840);
xor (n1839,n1753,n1754);
and (n1840,n395,n435);
and (n1841,n1842,n1843);
xor (n1842,n1839,n1840);
or (n1843,n1844,n1847);
and (n1844,n1845,n1846);
xor (n1845,n1758,n1759);
and (n1846,n548,n435);
and (n1847,n1848,n1849);
xor (n1848,n1845,n1846);
and (n1849,n1850,n1436);
xor (n1850,n1764,n1765);
and (n1851,n32,n443);
and (n1852,n1853,n1854);
xor (n1853,n1682,n1851);
or (n1854,n1855,n1858);
and (n1855,n1856,n1857);
xor (n1856,n1770,n1771);
and (n1857,n57,n443);
and (n1858,n1859,n1860);
xor (n1859,n1856,n1857);
or (n1860,n1861,n1864);
and (n1861,n1862,n1863);
xor (n1862,n1776,n1777);
and (n1863,n51,n443);
and (n1864,n1865,n1866);
xor (n1865,n1862,n1863);
or (n1866,n1867,n1870);
and (n1867,n1868,n1869);
xor (n1868,n1782,n1783);
and (n1869,n91,n443);
and (n1870,n1871,n1872);
xor (n1871,n1868,n1869);
or (n1872,n1873,n1876);
and (n1873,n1874,n1875);
xor (n1874,n1788,n1789);
and (n1875,n210,n443);
and (n1876,n1877,n1878);
xor (n1877,n1874,n1875);
or (n1878,n1879,n1882);
and (n1879,n1880,n1881);
xor (n1880,n1794,n1795);
and (n1881,n215,n443);
and (n1882,n1883,n1884);
xor (n1883,n1880,n1881);
or (n1884,n1885,n1888);
and (n1885,n1886,n1887);
xor (n1886,n1800,n1801);
and (n1887,n134,n443);
and (n1888,n1889,n1890);
xor (n1889,n1886,n1887);
or (n1890,n1891,n1894);
and (n1891,n1892,n1893);
xor (n1892,n1806,n1807);
and (n1893,n128,n443);
and (n1894,n1895,n1896);
xor (n1895,n1892,n1893);
or (n1896,n1897,n1900);
and (n1897,n1898,n1899);
xor (n1898,n1812,n1813);
and (n1899,n255,n443);
and (n1900,n1901,n1902);
xor (n1901,n1898,n1899);
or (n1902,n1903,n1906);
and (n1903,n1904,n1905);
xor (n1904,n1818,n1819);
and (n1905,n388,n443);
and (n1906,n1907,n1908);
xor (n1907,n1904,n1905);
or (n1908,n1909,n1911);
and (n1909,n1910,n1346);
xor (n1910,n1824,n1825);
and (n1911,n1912,n1913);
xor (n1912,n1910,n1346);
or (n1913,n1914,n1916);
and (n1914,n1915,n1378);
xor (n1915,n1830,n1831);
and (n1916,n1917,n1918);
xor (n1917,n1915,n1378);
or (n1918,n1919,n1921);
and (n1919,n1920,n1482);
xor (n1920,n1836,n1837);
and (n1921,n1922,n1923);
xor (n1922,n1920,n1482);
or (n1923,n1924,n1927);
and (n1924,n1925,n1926);
xor (n1925,n1842,n1843);
and (n1926,n548,n443);
and (n1927,n1928,n1929);
xor (n1928,n1925,n1926);
and (n1929,n1930,n1931);
xor (n1930,n1848,n1849);
and (n1931,n608,n443);
and (n1932,n32,n456);
and (n1933,n1934,n1935);
xor (n1934,n1679,n1932);
or (n1935,n1936,n1939);
and (n1936,n1937,n1938);
xor (n1937,n1853,n1854);
and (n1938,n57,n456);
and (n1939,n1940,n1941);
xor (n1940,n1937,n1938);
or (n1941,n1942,n1945);
and (n1942,n1943,n1944);
xor (n1943,n1859,n1860);
and (n1944,n51,n456);
and (n1945,n1946,n1947);
xor (n1946,n1943,n1944);
or (n1947,n1948,n1951);
and (n1948,n1949,n1950);
xor (n1949,n1865,n1866);
and (n1950,n91,n456);
and (n1951,n1952,n1953);
xor (n1952,n1949,n1950);
or (n1953,n1954,n1957);
and (n1954,n1955,n1956);
xor (n1955,n1871,n1872);
and (n1956,n210,n456);
and (n1957,n1958,n1959);
xor (n1958,n1955,n1956);
or (n1959,n1960,n1963);
and (n1960,n1961,n1962);
xor (n1961,n1877,n1878);
and (n1962,n215,n456);
and (n1963,n1964,n1965);
xor (n1964,n1961,n1962);
or (n1965,n1966,n1969);
and (n1966,n1967,n1968);
xor (n1967,n1883,n1884);
and (n1968,n134,n456);
and (n1969,n1970,n1971);
xor (n1970,n1967,n1968);
or (n1971,n1972,n1975);
and (n1972,n1973,n1974);
xor (n1973,n1889,n1890);
and (n1974,n128,n456);
and (n1975,n1976,n1977);
xor (n1976,n1973,n1974);
or (n1977,n1978,n1981);
and (n1978,n1979,n1980);
xor (n1979,n1895,n1896);
and (n1980,n255,n456);
and (n1981,n1982,n1983);
xor (n1982,n1979,n1980);
or (n1983,n1984,n1987);
and (n1984,n1985,n1986);
xor (n1985,n1901,n1902);
and (n1986,n388,n456);
and (n1987,n1988,n1989);
xor (n1988,n1985,n1986);
or (n1989,n1990,n1993);
and (n1990,n1991,n1992);
xor (n1991,n1907,n1908);
and (n1992,n382,n456);
and (n1993,n1994,n1995);
xor (n1994,n1991,n1992);
or (n1995,n1996,n1999);
and (n1996,n1997,n1998);
xor (n1997,n1912,n1913);
and (n1998,n401,n456);
and (n1999,n2000,n2001);
xor (n2000,n1997,n1998);
or (n2001,n2002,n2005);
and (n2002,n2003,n2004);
xor (n2003,n1917,n1918);
and (n2004,n395,n456);
and (n2005,n2006,n2007);
xor (n2006,n2003,n2004);
or (n2007,n2008,n2011);
and (n2008,n2009,n2010);
xor (n2009,n1922,n1923);
and (n2010,n548,n456);
and (n2011,n2012,n2013);
xor (n2012,n2009,n2010);
and (n2013,n2014,n1401);
xor (n2014,n1928,n1929);
and (n2015,n15,n188);
or (n2016,n2017,n2019);
and (n2017,n2018,n2015);
xor (n2018,n1643,n1661);
and (n2019,n2020,n2021);
xor (n2020,n2018,n2015);
or (n2021,n2022,n2024);
and (n2022,n2023,n2015);
xor (n2023,n1643,n1663);
and (n2024,n2025,n2026);
xor (n2025,n2023,n2015);
or (n2026,n2027,n2029);
and (n2027,n2028,n2015);
xor (n2028,n1643,n1665);
and (n2029,n2030,n2031);
xor (n2030,n2028,n2015);
or (n2031,n2032,n2034);
and (n2032,n2033,n2015);
xor (n2033,n1643,n1667);
and (n2034,n2035,n2036);
xor (n2035,n2033,n2015);
or (n2036,n2037,n2039);
and (n2037,n2038,n2015);
xor (n2038,n1643,n1669);
and (n2039,n2040,n2041);
xor (n2040,n2038,n2015);
or (n2041,n2042,n2044);
and (n2042,n2043,n2015);
xor (n2043,n1643,n1671);
and (n2044,n2045,n2046);
xor (n2045,n2043,n2015);
or (n2046,n2047,n2049);
and (n2047,n2048,n2015);
xor (n2048,n1643,n1673);
and (n2049,n2050,n2051);
xor (n2050,n2048,n2015);
or (n2051,n2052,n2054);
and (n2052,n2053,n2015);
xor (n2053,n1643,n1675);
and (n2054,n2055,n2056);
xor (n2055,n2053,n2015);
or (n2056,n2057,n2060);
and (n2057,n2058,n2059);
xor (n2058,n1643,n1677);
and (n2059,n32,n188);
and (n2060,n2061,n2062);
xor (n2061,n2058,n2059);
or (n2062,n2063,n2066);
and (n2063,n2064,n2065);
xor (n2064,n1934,n1935);
and (n2065,n57,n188);
and (n2066,n2067,n2068);
xor (n2067,n2064,n2065);
or (n2068,n2069,n2072);
and (n2069,n2070,n2071);
xor (n2070,n1940,n1941);
and (n2071,n51,n188);
and (n2072,n2073,n2074);
xor (n2073,n2070,n2071);
or (n2074,n2075,n2078);
and (n2075,n2076,n2077);
xor (n2076,n1946,n1947);
and (n2077,n91,n188);
and (n2078,n2079,n2080);
xor (n2079,n2076,n2077);
or (n2080,n2081,n2084);
and (n2081,n2082,n2083);
xor (n2082,n1952,n1953);
and (n2083,n210,n188);
and (n2084,n2085,n2086);
xor (n2085,n2082,n2083);
or (n2086,n2087,n2090);
and (n2087,n2088,n2089);
xor (n2088,n1958,n1959);
and (n2089,n215,n188);
and (n2090,n2091,n2092);
xor (n2091,n2088,n2089);
or (n2092,n2093,n2096);
and (n2093,n2094,n2095);
xor (n2094,n1964,n1965);
and (n2095,n134,n188);
and (n2096,n2097,n2098);
xor (n2097,n2094,n2095);
or (n2098,n2099,n2102);
and (n2099,n2100,n2101);
xor (n2100,n1970,n1971);
and (n2101,n128,n188);
and (n2102,n2103,n2104);
xor (n2103,n2100,n2101);
or (n2104,n2105,n2108);
and (n2105,n2106,n2107);
xor (n2106,n1976,n1977);
and (n2107,n255,n188);
and (n2108,n2109,n2110);
xor (n2109,n2106,n2107);
or (n2110,n2111,n2114);
and (n2111,n2112,n2113);
xor (n2112,n1982,n1983);
and (n2113,n388,n188);
and (n2114,n2115,n2116);
xor (n2115,n2112,n2113);
or (n2116,n2117,n2120);
and (n2117,n2118,n2119);
xor (n2118,n1988,n1989);
and (n2119,n382,n188);
and (n2120,n2121,n2122);
xor (n2121,n2118,n2119);
or (n2122,n2123,n2126);
and (n2123,n2124,n2125);
xor (n2124,n1994,n1995);
and (n2125,n401,n188);
and (n2126,n2127,n2128);
xor (n2127,n2124,n2125);
or (n2128,n2129,n2132);
and (n2129,n2130,n2131);
xor (n2130,n2000,n2001);
and (n2131,n395,n188);
and (n2132,n2133,n2134);
xor (n2133,n2130,n2131);
or (n2134,n2135,n2138);
and (n2135,n2136,n2137);
xor (n2136,n2006,n2007);
and (n2137,n548,n188);
and (n2138,n2139,n2140);
xor (n2139,n2136,n2137);
and (n2140,n2141,n2142);
xor (n2141,n2012,n2013);
and (n2142,n608,n188);
and (n2143,n15,n189);
or (n2144,n2145,n2147);
and (n2145,n2146,n2143);
xor (n2146,n2020,n2021);
and (n2147,n2148,n2149);
xor (n2148,n2146,n2143);
or (n2149,n2150,n2152);
and (n2150,n2151,n2143);
xor (n2151,n2025,n2026);
and (n2152,n2153,n2154);
xor (n2153,n2151,n2143);
or (n2154,n2155,n2157);
and (n2155,n2156,n2143);
xor (n2156,n2030,n2031);
and (n2157,n2158,n2159);
xor (n2158,n2156,n2143);
or (n2159,n2160,n2162);
and (n2160,n2161,n2143);
xor (n2161,n2035,n2036);
and (n2162,n2163,n2164);
xor (n2163,n2161,n2143);
or (n2164,n2165,n2167);
and (n2165,n2166,n2143);
xor (n2166,n2040,n2041);
and (n2167,n2168,n2169);
xor (n2168,n2166,n2143);
or (n2169,n2170,n2172);
and (n2170,n2171,n2143);
xor (n2171,n2045,n2046);
and (n2172,n2173,n2174);
xor (n2173,n2171,n2143);
or (n2174,n2175,n2177);
and (n2175,n2176,n2143);
xor (n2176,n2050,n2051);
and (n2177,n2178,n2179);
xor (n2178,n2176,n2143);
or (n2179,n2180,n2183);
and (n2180,n2181,n2182);
xor (n2181,n2055,n2056);
and (n2182,n32,n189);
and (n2183,n2184,n2185);
xor (n2184,n2181,n2182);
or (n2185,n2186,n2189);
and (n2186,n2187,n2188);
xor (n2187,n2061,n2062);
and (n2188,n57,n189);
and (n2189,n2190,n2191);
xor (n2190,n2187,n2188);
or (n2191,n2192,n2195);
and (n2192,n2193,n2194);
xor (n2193,n2067,n2068);
and (n2194,n51,n189);
and (n2195,n2196,n2197);
xor (n2196,n2193,n2194);
or (n2197,n2198,n2201);
and (n2198,n2199,n2200);
xor (n2199,n2073,n2074);
and (n2200,n91,n189);
and (n2201,n2202,n2203);
xor (n2202,n2199,n2200);
or (n2203,n2204,n2207);
and (n2204,n2205,n2206);
xor (n2205,n2079,n2080);
and (n2206,n210,n189);
and (n2207,n2208,n2209);
xor (n2208,n2205,n2206);
or (n2209,n2210,n2213);
and (n2210,n2211,n2212);
xor (n2211,n2085,n2086);
and (n2212,n215,n189);
and (n2213,n2214,n2215);
xor (n2214,n2211,n2212);
or (n2215,n2216,n2219);
and (n2216,n2217,n2218);
xor (n2217,n2091,n2092);
and (n2218,n134,n189);
and (n2219,n2220,n2221);
xor (n2220,n2217,n2218);
or (n2221,n2222,n2225);
and (n2222,n2223,n2224);
xor (n2223,n2097,n2098);
and (n2224,n128,n189);
and (n2225,n2226,n2227);
xor (n2226,n2223,n2224);
or (n2227,n2228,n2231);
and (n2228,n2229,n2230);
xor (n2229,n2103,n2104);
and (n2230,n255,n189);
and (n2231,n2232,n2233);
xor (n2232,n2229,n2230);
or (n2233,n2234,n2237);
and (n2234,n2235,n2236);
xor (n2235,n2109,n2110);
and (n2236,n388,n189);
and (n2237,n2238,n2239);
xor (n2238,n2235,n2236);
or (n2239,n2240,n2243);
and (n2240,n2241,n2242);
xor (n2241,n2115,n2116);
and (n2242,n382,n189);
and (n2243,n2244,n2245);
xor (n2244,n2241,n2242);
or (n2245,n2246,n2249);
and (n2246,n2247,n2248);
xor (n2247,n2121,n2122);
and (n2248,n401,n189);
and (n2249,n2250,n2251);
xor (n2250,n2247,n2248);
or (n2251,n2252,n2255);
and (n2252,n2253,n2254);
xor (n2253,n2127,n2128);
and (n2254,n395,n189);
and (n2255,n2256,n2257);
xor (n2256,n2253,n2254);
or (n2257,n2258,n2261);
and (n2258,n2259,n2260);
xor (n2259,n2133,n2134);
and (n2260,n548,n189);
and (n2261,n2262,n2263);
xor (n2262,n2259,n2260);
and (n2263,n2264,n1245);
xor (n2264,n2139,n2140);
and (n2265,n15,n152);
or (n2266,n2267,n2269);
and (n2267,n2268,n2265);
xor (n2268,n2148,n2149);
and (n2269,n2270,n2271);
xor (n2270,n2268,n2265);
or (n2271,n2272,n2274);
and (n2272,n2273,n2265);
xor (n2273,n2153,n2154);
and (n2274,n2275,n2276);
xor (n2275,n2273,n2265);
or (n2276,n2277,n2279);
and (n2277,n2278,n2265);
xor (n2278,n2158,n2159);
and (n2279,n2280,n2281);
xor (n2280,n2278,n2265);
or (n2281,n2282,n2284);
and (n2282,n2283,n2265);
xor (n2283,n2163,n2164);
and (n2284,n2285,n2286);
xor (n2285,n2283,n2265);
or (n2286,n2287,n2289);
and (n2287,n2288,n2265);
xor (n2288,n2168,n2169);
and (n2289,n2290,n2291);
xor (n2290,n2288,n2265);
or (n2291,n2292,n2294);
and (n2292,n2293,n2265);
xor (n2293,n2173,n2174);
and (n2294,n2295,n2296);
xor (n2295,n2293,n2265);
or (n2296,n2297,n2300);
and (n2297,n2298,n2299);
xor (n2298,n2178,n2179);
and (n2299,n32,n152);
and (n2300,n2301,n2302);
xor (n2301,n2298,n2299);
or (n2302,n2303,n2306);
and (n2303,n2304,n2305);
xor (n2304,n2184,n2185);
and (n2305,n57,n152);
and (n2306,n2307,n2308);
xor (n2307,n2304,n2305);
or (n2308,n2309,n2312);
and (n2309,n2310,n2311);
xor (n2310,n2190,n2191);
and (n2311,n51,n152);
and (n2312,n2313,n2314);
xor (n2313,n2310,n2311);
or (n2314,n2315,n2318);
and (n2315,n2316,n2317);
xor (n2316,n2196,n2197);
and (n2317,n91,n152);
and (n2318,n2319,n2320);
xor (n2319,n2316,n2317);
or (n2320,n2321,n2324);
and (n2321,n2322,n2323);
xor (n2322,n2202,n2203);
and (n2323,n210,n152);
and (n2324,n2325,n2326);
xor (n2325,n2322,n2323);
or (n2326,n2327,n2330);
and (n2327,n2328,n2329);
xor (n2328,n2208,n2209);
and (n2329,n215,n152);
and (n2330,n2331,n2332);
xor (n2331,n2328,n2329);
or (n2332,n2333,n2336);
and (n2333,n2334,n2335);
xor (n2334,n2214,n2215);
and (n2335,n134,n152);
and (n2336,n2337,n2338);
xor (n2337,n2334,n2335);
or (n2338,n2339,n2342);
and (n2339,n2340,n2341);
xor (n2340,n2220,n2221);
and (n2341,n128,n152);
and (n2342,n2343,n2344);
xor (n2343,n2340,n2341);
or (n2344,n2345,n2348);
and (n2345,n2346,n2347);
xor (n2346,n2226,n2227);
and (n2347,n255,n152);
and (n2348,n2349,n2350);
xor (n2349,n2346,n2347);
or (n2350,n2351,n2354);
and (n2351,n2352,n2353);
xor (n2352,n2232,n2233);
and (n2353,n388,n152);
and (n2354,n2355,n2356);
xor (n2355,n2352,n2353);
or (n2356,n2357,n2360);
and (n2357,n2358,n2359);
xor (n2358,n2238,n2239);
and (n2359,n382,n152);
and (n2360,n2361,n2362);
xor (n2361,n2358,n2359);
or (n2362,n2363,n2366);
and (n2363,n2364,n2365);
xor (n2364,n2244,n2245);
and (n2365,n401,n152);
and (n2366,n2367,n2368);
xor (n2367,n2364,n2365);
or (n2368,n2369,n2372);
and (n2369,n2370,n2371);
xor (n2370,n2250,n2251);
and (n2371,n395,n152);
and (n2372,n2373,n2374);
xor (n2373,n2370,n2371);
or (n2374,n2375,n2377);
and (n2375,n2376,n1293);
xor (n2376,n2256,n2257);
and (n2377,n2378,n2379);
xor (n2378,n2376,n1293);
and (n2379,n2380,n2381);
xor (n2380,n2262,n2263);
and (n2381,n608,n152);
and (n2382,n15,n153);
or (n2383,n2384,n2386);
and (n2384,n2385,n2382);
xor (n2385,n2270,n2271);
and (n2386,n2387,n2388);
xor (n2387,n2385,n2382);
or (n2388,n2389,n2391);
and (n2389,n2390,n2382);
xor (n2390,n2275,n2276);
and (n2391,n2392,n2393);
xor (n2392,n2390,n2382);
or (n2393,n2394,n2396);
and (n2394,n2395,n2382);
xor (n2395,n2280,n2281);
and (n2396,n2397,n2398);
xor (n2397,n2395,n2382);
or (n2398,n2399,n2401);
and (n2399,n2400,n2382);
xor (n2400,n2285,n2286);
and (n2401,n2402,n2403);
xor (n2402,n2400,n2382);
or (n2403,n2404,n2406);
and (n2404,n2405,n2382);
xor (n2405,n2290,n2291);
and (n2406,n2407,n2408);
xor (n2407,n2405,n2382);
or (n2408,n2409,n2412);
and (n2409,n2410,n2411);
xor (n2410,n2295,n2296);
and (n2411,n32,n153);
and (n2412,n2413,n2414);
xor (n2413,n2410,n2411);
or (n2414,n2415,n2418);
and (n2415,n2416,n2417);
xor (n2416,n2301,n2302);
and (n2417,n57,n153);
and (n2418,n2419,n2420);
xor (n2419,n2416,n2417);
or (n2420,n2421,n2424);
and (n2421,n2422,n2423);
xor (n2422,n2307,n2308);
and (n2423,n51,n153);
and (n2424,n2425,n2426);
xor (n2425,n2422,n2423);
or (n2426,n2427,n2430);
and (n2427,n2428,n2429);
xor (n2428,n2313,n2314);
and (n2429,n91,n153);
and (n2430,n2431,n2432);
xor (n2431,n2428,n2429);
or (n2432,n2433,n2436);
and (n2433,n2434,n2435);
xor (n2434,n2319,n2320);
and (n2435,n210,n153);
and (n2436,n2437,n2438);
xor (n2437,n2434,n2435);
or (n2438,n2439,n2442);
and (n2439,n2440,n2441);
xor (n2440,n2325,n2326);
and (n2441,n215,n153);
and (n2442,n2443,n2444);
xor (n2443,n2440,n2441);
or (n2444,n2445,n2448);
and (n2445,n2446,n2447);
xor (n2446,n2331,n2332);
and (n2447,n134,n153);
and (n2448,n2449,n2450);
xor (n2449,n2446,n2447);
or (n2450,n2451,n2454);
and (n2451,n2452,n2453);
xor (n2452,n2337,n2338);
and (n2453,n128,n153);
and (n2454,n2455,n2456);
xor (n2455,n2452,n2453);
or (n2456,n2457,n2460);
and (n2457,n2458,n2459);
xor (n2458,n2343,n2344);
and (n2459,n255,n153);
and (n2460,n2461,n2462);
xor (n2461,n2458,n2459);
or (n2462,n2463,n2466);
and (n2463,n2464,n2465);
xor (n2464,n2349,n2350);
and (n2465,n388,n153);
and (n2466,n2467,n2468);
xor (n2467,n2464,n2465);
or (n2468,n2469,n2472);
and (n2469,n2470,n2471);
xor (n2470,n2355,n2356);
and (n2471,n382,n153);
and (n2472,n2473,n2474);
xor (n2473,n2470,n2471);
or (n2474,n2475,n2478);
and (n2475,n2476,n2477);
xor (n2476,n2361,n2362);
and (n2477,n401,n153);
and (n2478,n2479,n2480);
xor (n2479,n2476,n2477);
or (n2480,n2481,n2484);
and (n2481,n2482,n2483);
xor (n2482,n2367,n2368);
and (n2483,n395,n153);
and (n2484,n2485,n2486);
xor (n2485,n2482,n2483);
or (n2486,n2487,n2490);
and (n2487,n2488,n2489);
xor (n2488,n2373,n2374);
and (n2489,n548,n153);
and (n2490,n2491,n2492);
xor (n2491,n2488,n2489);
and (n2492,n2493,n2494);
xor (n2493,n2378,n2379);
not (n2494,n1270);
and (n2495,n15,n70);
or (n2496,n2497,n2499);
and (n2497,n2498,n2495);
xor (n2498,n2387,n2388);
and (n2499,n2500,n2501);
xor (n2500,n2498,n2495);
or (n2501,n2502,n2504);
and (n2502,n2503,n2495);
xor (n2503,n2392,n2393);
and (n2504,n2505,n2506);
xor (n2505,n2503,n2495);
or (n2506,n2507,n2509);
and (n2507,n2508,n2495);
xor (n2508,n2397,n2398);
and (n2509,n2510,n2511);
xor (n2510,n2508,n2495);
or (n2511,n2512,n2514);
and (n2512,n2513,n2495);
xor (n2513,n2402,n2403);
and (n2514,n2515,n2516);
xor (n2515,n2513,n2495);
or (n2516,n2517,n2520);
and (n2517,n2518,n2519);
xor (n2518,n2407,n2408);
and (n2519,n32,n70);
and (n2520,n2521,n2522);
xor (n2521,n2518,n2519);
or (n2522,n2523,n2526);
and (n2523,n2524,n2525);
xor (n2524,n2413,n2414);
and (n2525,n57,n70);
and (n2526,n2527,n2528);
xor (n2527,n2524,n2525);
or (n2528,n2529,n2532);
and (n2529,n2530,n2531);
xor (n2530,n2419,n2420);
and (n2531,n51,n70);
and (n2532,n2533,n2534);
xor (n2533,n2530,n2531);
or (n2534,n2535,n2538);
and (n2535,n2536,n2537);
xor (n2536,n2425,n2426);
and (n2537,n91,n70);
and (n2538,n2539,n2540);
xor (n2539,n2536,n2537);
or (n2540,n2541,n2544);
and (n2541,n2542,n2543);
xor (n2542,n2431,n2432);
and (n2543,n210,n70);
and (n2544,n2545,n2546);
xor (n2545,n2542,n2543);
or (n2546,n2547,n2550);
and (n2547,n2548,n2549);
xor (n2548,n2437,n2438);
and (n2549,n215,n70);
and (n2550,n2551,n2552);
xor (n2551,n2548,n2549);
or (n2552,n2553,n2556);
and (n2553,n2554,n2555);
xor (n2554,n2443,n2444);
and (n2555,n134,n70);
and (n2556,n2557,n2558);
xor (n2557,n2554,n2555);
or (n2558,n2559,n2561);
and (n2559,n2560,n563);
xor (n2560,n2449,n2450);
and (n2561,n2562,n2563);
xor (n2562,n2560,n563);
or (n2563,n2564,n2567);
and (n2564,n2565,n2566);
xor (n2565,n2455,n2456);
and (n2566,n255,n70);
and (n2567,n2568,n2569);
xor (n2568,n2565,n2566);
or (n2569,n2570,n2573);
and (n2570,n2571,n2572);
xor (n2571,n2461,n2462);
and (n2572,n388,n70);
and (n2573,n2574,n2575);
xor (n2574,n2571,n2572);
or (n2575,n2576,n2578);
and (n2576,n2577,n806);
xor (n2577,n2467,n2468);
and (n2578,n2579,n2580);
xor (n2579,n2577,n806);
or (n2580,n2581,n2584);
and (n2581,n2582,n2583);
xor (n2582,n2473,n2474);
and (n2583,n401,n70);
and (n2584,n2585,n2586);
xor (n2585,n2582,n2583);
or (n2586,n2587,n2589);
and (n2587,n2588,n1129);
xor (n2588,n2479,n2480);
and (n2589,n2590,n2591);
xor (n2590,n2588,n1129);
or (n2591,n2592,n2595);
and (n2592,n2593,n2594);
xor (n2593,n2485,n2486);
and (n2594,n548,n70);
and (n2595,n2596,n2597);
xor (n2596,n2593,n2594);
and (n2597,n2598,n2599);
xor (n2598,n2491,n2492);
and (n2599,n608,n70);
and (n2600,n15,n71);
or (n2601,n2602,n2604);
and (n2602,n2603,n2600);
xor (n2603,n2500,n2501);
and (n2604,n2605,n2606);
xor (n2605,n2603,n2600);
or (n2606,n2607,n2609);
and (n2607,n2608,n2600);
xor (n2608,n2505,n2506);
and (n2609,n2610,n2611);
xor (n2610,n2608,n2600);
or (n2611,n2612,n2614);
and (n2612,n2613,n2600);
xor (n2613,n2510,n2511);
and (n2614,n2615,n2616);
xor (n2615,n2613,n2600);
or (n2616,n2617,n2620);
and (n2617,n2618,n2619);
xor (n2618,n2515,n2516);
and (n2619,n32,n71);
and (n2620,n2621,n2622);
xor (n2621,n2618,n2619);
or (n2622,n2623,n2626);
and (n2623,n2624,n2625);
xor (n2624,n2521,n2522);
and (n2625,n57,n71);
and (n2626,n2627,n2628);
xor (n2627,n2624,n2625);
or (n2628,n2629,n2632);
and (n2629,n2630,n2631);
xor (n2630,n2527,n2528);
and (n2631,n51,n71);
and (n2632,n2633,n2634);
xor (n2633,n2630,n2631);
or (n2634,n2635,n2638);
and (n2635,n2636,n2637);
xor (n2636,n2533,n2534);
and (n2637,n91,n71);
and (n2638,n2639,n2640);
xor (n2639,n2636,n2637);
or (n2640,n2641,n2644);
and (n2641,n2642,n2643);
xor (n2642,n2539,n2540);
and (n2643,n210,n71);
and (n2644,n2645,n2646);
xor (n2645,n2642,n2643);
or (n2646,n2647,n2650);
and (n2647,n2648,n2649);
xor (n2648,n2545,n2546);
and (n2649,n215,n71);
and (n2650,n2651,n2652);
xor (n2651,n2648,n2649);
or (n2652,n2653,n2656);
and (n2653,n2654,n2655);
xor (n2654,n2551,n2552);
and (n2655,n134,n71);
and (n2656,n2657,n2658);
xor (n2657,n2654,n2655);
or (n2658,n2659,n2662);
and (n2659,n2660,n2661);
xor (n2660,n2557,n2558);
and (n2661,n128,n71);
and (n2662,n2663,n2664);
xor (n2663,n2660,n2661);
or (n2664,n2665,n2668);
and (n2665,n2666,n2667);
xor (n2666,n2562,n2563);
and (n2667,n255,n71);
and (n2668,n2669,n2670);
xor (n2669,n2666,n2667);
or (n2670,n2671,n2674);
and (n2671,n2672,n2673);
xor (n2672,n2568,n2569);
and (n2673,n388,n71);
and (n2674,n2675,n2676);
xor (n2675,n2672,n2673);
or (n2676,n2677,n2680);
and (n2677,n2678,n2679);
xor (n2678,n2574,n2575);
and (n2679,n382,n71);
and (n2680,n2681,n2682);
xor (n2681,n2678,n2679);
or (n2682,n2683,n2686);
and (n2683,n2684,n2685);
xor (n2684,n2579,n2580);
and (n2685,n401,n71);
and (n2686,n2687,n2688);
xor (n2687,n2684,n2685);
or (n2688,n2689,n2692);
and (n2689,n2690,n2691);
xor (n2690,n2585,n2586);
and (n2691,n395,n71);
and (n2692,n2693,n2694);
xor (n2693,n2690,n2691);
or (n2694,n2695,n2698);
and (n2695,n2696,n2697);
xor (n2696,n2590,n2591);
and (n2697,n548,n71);
and (n2698,n2699,n2700);
xor (n2699,n2696,n2697);
and (n2700,n2701,n1113);
xor (n2701,n2596,n2597);
and (n2702,n15,n20);
or (n2703,n2704,n2706);
and (n2704,n2705,n2702);
xor (n2705,n2605,n2606);
and (n2706,n2707,n2708);
xor (n2707,n2705,n2702);
or (n2708,n2709,n2711);
and (n2709,n2710,n2702);
xor (n2710,n2610,n2611);
and (n2711,n2712,n2713);
xor (n2712,n2710,n2702);
or (n2713,n2714,n2717);
and (n2714,n2715,n2716);
xor (n2715,n2615,n2616);
and (n2716,n32,n20);
and (n2717,n2718,n2719);
xor (n2718,n2715,n2716);
or (n2719,n2720,n2723);
and (n2720,n2721,n2722);
xor (n2721,n2621,n2622);
and (n2722,n57,n20);
and (n2723,n2724,n2725);
xor (n2724,n2721,n2722);
or (n2725,n2726,n2729);
and (n2726,n2727,n2728);
xor (n2727,n2627,n2628);
and (n2728,n51,n20);
and (n2729,n2730,n2731);
xor (n2730,n2727,n2728);
or (n2731,n2732,n2735);
and (n2732,n2733,n2734);
xor (n2733,n2633,n2634);
and (n2734,n91,n20);
and (n2735,n2736,n2737);
xor (n2736,n2733,n2734);
or (n2737,n2738,n2741);
and (n2738,n2739,n2740);
xor (n2739,n2639,n2640);
and (n2740,n210,n20);
and (n2741,n2742,n2743);
xor (n2742,n2739,n2740);
or (n2743,n2744,n2747);
and (n2744,n2745,n2746);
xor (n2745,n2645,n2646);
and (n2746,n215,n20);
and (n2747,n2748,n2749);
xor (n2748,n2745,n2746);
or (n2749,n2750,n2753);
and (n2750,n2751,n2752);
xor (n2751,n2651,n2652);
and (n2752,n134,n20);
and (n2753,n2754,n2755);
xor (n2754,n2751,n2752);
or (n2755,n2756,n2759);
and (n2756,n2757,n2758);
xor (n2757,n2657,n2658);
and (n2758,n128,n20);
and (n2759,n2760,n2761);
xor (n2760,n2757,n2758);
or (n2761,n2762,n2765);
and (n2762,n2763,n2764);
xor (n2763,n2663,n2664);
and (n2764,n255,n20);
and (n2765,n2766,n2767);
xor (n2766,n2763,n2764);
or (n2767,n2768,n2771);
and (n2768,n2769,n2770);
xor (n2769,n2669,n2670);
and (n2770,n388,n20);
and (n2771,n2772,n2773);
xor (n2772,n2769,n2770);
or (n2773,n2774,n2777);
and (n2774,n2775,n2776);
xor (n2775,n2675,n2676);
and (n2776,n382,n20);
and (n2777,n2778,n2779);
xor (n2778,n2775,n2776);
or (n2779,n2780,n2783);
and (n2780,n2781,n2782);
xor (n2781,n2681,n2682);
and (n2782,n401,n20);
and (n2783,n2784,n2785);
xor (n2784,n2781,n2782);
or (n2785,n2786,n2789);
and (n2786,n2787,n2788);
xor (n2787,n2687,n2688);
and (n2788,n395,n20);
and (n2789,n2790,n2791);
xor (n2790,n2787,n2788);
or (n2791,n2792,n2795);
and (n2792,n2793,n2794);
xor (n2793,n2693,n2694);
and (n2794,n548,n20);
and (n2795,n2796,n2797);
xor (n2796,n2793,n2794);
and (n2797,n2798,n2799);
xor (n2798,n2699,n2700);
and (n2799,n608,n20);
and (n2800,n15,n22);
or (n2801,n2802,n2804);
and (n2802,n2803,n2800);
xor (n2803,n2707,n2708);
and (n2804,n2805,n2806);
xor (n2805,n2803,n2800);
or (n2806,n2807,n2810);
and (n2807,n2808,n2809);
xor (n2808,n2712,n2713);
and (n2809,n32,n22);
and (n2810,n2811,n2812);
xor (n2811,n2808,n2809);
or (n2812,n2813,n2816);
and (n2813,n2814,n2815);
xor (n2814,n2718,n2719);
and (n2815,n57,n22);
and (n2816,n2817,n2818);
xor (n2817,n2814,n2815);
or (n2818,n2819,n2822);
and (n2819,n2820,n2821);
xor (n2820,n2724,n2725);
and (n2821,n51,n22);
and (n2822,n2823,n2824);
xor (n2823,n2820,n2821);
or (n2824,n2825,n2828);
and (n2825,n2826,n2827);
xor (n2826,n2730,n2731);
and (n2827,n91,n22);
and (n2828,n2829,n2830);
xor (n2829,n2826,n2827);
or (n2830,n2831,n2834);
and (n2831,n2832,n2833);
xor (n2832,n2736,n2737);
and (n2833,n210,n22);
and (n2834,n2835,n2836);
xor (n2835,n2832,n2833);
or (n2836,n2837,n2840);
and (n2837,n2838,n2839);
xor (n2838,n2742,n2743);
and (n2839,n215,n22);
and (n2840,n2841,n2842);
xor (n2841,n2838,n2839);
or (n2842,n2843,n2846);
and (n2843,n2844,n2845);
xor (n2844,n2748,n2749);
and (n2845,n134,n22);
and (n2846,n2847,n2848);
xor (n2847,n2844,n2845);
or (n2848,n2849,n2852);
and (n2849,n2850,n2851);
xor (n2850,n2754,n2755);
and (n2851,n128,n22);
and (n2852,n2853,n2854);
xor (n2853,n2850,n2851);
or (n2854,n2855,n2858);
and (n2855,n2856,n2857);
xor (n2856,n2760,n2761);
and (n2857,n255,n22);
and (n2858,n2859,n2860);
xor (n2859,n2856,n2857);
or (n2860,n2861,n2864);
and (n2861,n2862,n2863);
xor (n2862,n2766,n2767);
and (n2863,n388,n22);
and (n2864,n2865,n2866);
xor (n2865,n2862,n2863);
or (n2866,n2867,n2870);
and (n2867,n2868,n2869);
xor (n2868,n2772,n2773);
and (n2869,n382,n22);
and (n2870,n2871,n2872);
xor (n2871,n2868,n2869);
or (n2872,n2873,n2876);
and (n2873,n2874,n2875);
xor (n2874,n2778,n2779);
and (n2875,n401,n22);
and (n2876,n2877,n2878);
xor (n2877,n2874,n2875);
or (n2878,n2879,n2882);
and (n2879,n2880,n2881);
xor (n2880,n2784,n2785);
and (n2881,n395,n22);
and (n2882,n2883,n2884);
xor (n2883,n2880,n2881);
or (n2884,n2885,n2888);
and (n2885,n2886,n2887);
xor (n2886,n2790,n2791);
and (n2887,n548,n22);
and (n2888,n2889,n2890);
xor (n2889,n2886,n2887);
and (n2890,n2891,n2892);
xor (n2891,n2796,n2797);
not (n2892,n772);
and (n2893,n15,n13);
or (n2894,n2895,n2898);
and (n2895,n2896,n2897);
xor (n2896,n2805,n2806);
and (n2897,n32,n13);
and (n2898,n2899,n2900);
xor (n2899,n2896,n2897);
or (n2900,n2901,n2904);
and (n2901,n2902,n2903);
xor (n2902,n2811,n2812);
and (n2903,n57,n13);
and (n2904,n2905,n2906);
xor (n2905,n2902,n2903);
or (n2906,n2907,n2910);
and (n2907,n2908,n2909);
xor (n2908,n2817,n2818);
and (n2909,n51,n13);
and (n2910,n2911,n2912);
xor (n2911,n2908,n2909);
or (n2912,n2913,n2916);
and (n2913,n2914,n2915);
xor (n2914,n2823,n2824);
and (n2915,n91,n13);
and (n2916,n2917,n2918);
xor (n2917,n2914,n2915);
or (n2918,n2919,n2922);
and (n2919,n2920,n2921);
xor (n2920,n2829,n2830);
and (n2921,n210,n13);
and (n2922,n2923,n2924);
xor (n2923,n2920,n2921);
or (n2924,n2925,n2928);
and (n2925,n2926,n2927);
xor (n2926,n2835,n2836);
and (n2927,n215,n13);
and (n2928,n2929,n2930);
xor (n2929,n2926,n2927);
or (n2930,n2931,n2934);
and (n2931,n2932,n2933);
xor (n2932,n2841,n2842);
and (n2933,n134,n13);
and (n2934,n2935,n2936);
xor (n2935,n2932,n2933);
or (n2936,n2937,n2940);
and (n2937,n2938,n2939);
xor (n2938,n2847,n2848);
and (n2939,n128,n13);
and (n2940,n2941,n2942);
xor (n2941,n2938,n2939);
or (n2942,n2943,n2946);
and (n2943,n2944,n2945);
xor (n2944,n2853,n2854);
and (n2945,n255,n13);
and (n2946,n2947,n2948);
xor (n2947,n2944,n2945);
or (n2948,n2949,n2952);
and (n2949,n2950,n2951);
xor (n2950,n2859,n2860);
and (n2951,n388,n13);
and (n2952,n2953,n2954);
xor (n2953,n2950,n2951);
or (n2954,n2955,n2958);
and (n2955,n2956,n2957);
xor (n2956,n2865,n2866);
and (n2957,n382,n13);
and (n2958,n2959,n2960);
xor (n2959,n2956,n2957);
or (n2960,n2961,n2964);
and (n2961,n2962,n2963);
xor (n2962,n2871,n2872);
and (n2963,n401,n13);
and (n2964,n2965,n2966);
xor (n2965,n2962,n2963);
or (n2966,n2967,n2970);
and (n2967,n2968,n2969);
xor (n2968,n2877,n2878);
and (n2969,n395,n13);
and (n2970,n2971,n2972);
xor (n2971,n2968,n2969);
or (n2972,n2973,n2976);
and (n2973,n2974,n2975);
xor (n2974,n2883,n2884);
and (n2975,n548,n13);
and (n2976,n2977,n2978);
xor (n2977,n2974,n2975);
and (n2978,n2979,n2980);
xor (n2979,n2889,n2890);
and (n2980,n608,n13);
and (n2981,n32,n41);
or (n2982,n2983,n2986);
and (n2983,n2984,n2985);
xor (n2984,n2899,n2900);
and (n2985,n57,n41);
and (n2986,n2987,n2988);
xor (n2987,n2984,n2985);
or (n2988,n2989,n2992);
and (n2989,n2990,n2991);
xor (n2990,n2905,n2906);
and (n2991,n51,n41);
and (n2992,n2993,n2994);
xor (n2993,n2990,n2991);
or (n2994,n2995,n2998);
and (n2995,n2996,n2997);
xor (n2996,n2911,n2912);
and (n2997,n91,n41);
and (n2998,n2999,n3000);
xor (n2999,n2996,n2997);
or (n3000,n3001,n3004);
and (n3001,n3002,n3003);
xor (n3002,n2917,n2918);
and (n3003,n210,n41);
and (n3004,n3005,n3006);
xor (n3005,n3002,n3003);
or (n3006,n3007,n3010);
and (n3007,n3008,n3009);
xor (n3008,n2923,n2924);
and (n3009,n215,n41);
and (n3010,n3011,n3012);
xor (n3011,n3008,n3009);
or (n3012,n3013,n3016);
and (n3013,n3014,n3015);
xor (n3014,n2929,n2930);
and (n3015,n134,n41);
and (n3016,n3017,n3018);
xor (n3017,n3014,n3015);
or (n3018,n3019,n3022);
and (n3019,n3020,n3021);
xor (n3020,n2935,n2936);
and (n3021,n128,n41);
and (n3022,n3023,n3024);
xor (n3023,n3020,n3021);
or (n3024,n3025,n3028);
and (n3025,n3026,n3027);
xor (n3026,n2941,n2942);
and (n3027,n255,n41);
and (n3028,n3029,n3030);
xor (n3029,n3026,n3027);
or (n3030,n3031,n3034);
and (n3031,n3032,n3033);
xor (n3032,n2947,n2948);
and (n3033,n388,n41);
and (n3034,n3035,n3036);
xor (n3035,n3032,n3033);
or (n3036,n3037,n3040);
and (n3037,n3038,n3039);
xor (n3038,n2953,n2954);
and (n3039,n382,n41);
and (n3040,n3041,n3042);
xor (n3041,n3038,n3039);
or (n3042,n3043,n3046);
and (n3043,n3044,n3045);
xor (n3044,n2959,n2960);
and (n3045,n401,n41);
and (n3046,n3047,n3048);
xor (n3047,n3044,n3045);
or (n3048,n3049,n3052);
and (n3049,n3050,n3051);
xor (n3050,n2965,n2966);
and (n3051,n395,n41);
and (n3052,n3053,n3054);
xor (n3053,n3050,n3051);
or (n3054,n3055,n3058);
and (n3055,n3056,n3057);
xor (n3056,n2971,n2972);
and (n3057,n548,n41);
and (n3058,n3059,n3060);
xor (n3059,n3056,n3057);
and (n3060,n3061,n3062);
xor (n3061,n2977,n2978);
not (n3062,n607);
and (n3063,n57,n47);
or (n3064,n3065,n3068);
and (n3065,n3066,n3067);
xor (n3066,n2987,n2988);
and (n3067,n51,n47);
and (n3068,n3069,n3070);
xor (n3069,n3066,n3067);
or (n3070,n3071,n3074);
and (n3071,n3072,n3073);
xor (n3072,n2993,n2994);
and (n3073,n91,n47);
and (n3074,n3075,n3076);
xor (n3075,n3072,n3073);
or (n3076,n3077,n3080);
and (n3077,n3078,n3079);
xor (n3078,n2999,n3000);
and (n3079,n210,n47);
and (n3080,n3081,n3082);
xor (n3081,n3078,n3079);
or (n3082,n3083,n3086);
and (n3083,n3084,n3085);
xor (n3084,n3005,n3006);
and (n3085,n215,n47);
and (n3086,n3087,n3088);
xor (n3087,n3084,n3085);
or (n3088,n3089,n3092);
and (n3089,n3090,n3091);
xor (n3090,n3011,n3012);
and (n3091,n134,n47);
and (n3092,n3093,n3094);
xor (n3093,n3090,n3091);
or (n3094,n3095,n3098);
and (n3095,n3096,n3097);
xor (n3096,n3017,n3018);
and (n3097,n128,n47);
and (n3098,n3099,n3100);
xor (n3099,n3096,n3097);
or (n3100,n3101,n3104);
and (n3101,n3102,n3103);
xor (n3102,n3023,n3024);
and (n3103,n255,n47);
and (n3104,n3105,n3106);
xor (n3105,n3102,n3103);
or (n3106,n3107,n3110);
and (n3107,n3108,n3109);
xor (n3108,n3029,n3030);
and (n3109,n388,n47);
and (n3110,n3111,n3112);
xor (n3111,n3108,n3109);
or (n3112,n3113,n3116);
and (n3113,n3114,n3115);
xor (n3114,n3035,n3036);
and (n3115,n382,n47);
and (n3116,n3117,n3118);
xor (n3117,n3114,n3115);
or (n3118,n3119,n3122);
and (n3119,n3120,n3121);
xor (n3120,n3041,n3042);
and (n3121,n401,n47);
and (n3122,n3123,n3124);
xor (n3123,n3120,n3121);
or (n3124,n3125,n3128);
and (n3125,n3126,n3127);
xor (n3126,n3047,n3048);
and (n3127,n395,n47);
and (n3128,n3129,n3130);
xor (n3129,n3126,n3127);
or (n3130,n3131,n3134);
and (n3131,n3132,n3133);
xor (n3132,n3053,n3054);
and (n3133,n548,n47);
and (n3134,n3135,n3136);
xor (n3135,n3132,n3133);
and (n3136,n3137,n3138);
xor (n3137,n3059,n3060);
and (n3138,n608,n47);
or (n3139,n3140,n3142);
and (n3140,n3141,n3073);
xor (n3141,n3069,n3070);
and (n3142,n3143,n3144);
xor (n3143,n3141,n3073);
or (n3144,n3145,n3147);
and (n3145,n3146,n3079);
xor (n3146,n3075,n3076);
and (n3147,n3148,n3149);
xor (n3148,n3146,n3079);
or (n3149,n3150,n3152);
and (n3150,n3151,n3085);
xor (n3151,n3081,n3082);
and (n3152,n3153,n3154);
xor (n3153,n3151,n3085);
or (n3154,n3155,n3157);
and (n3155,n3156,n3091);
xor (n3156,n3087,n3088);
and (n3157,n3158,n3159);
xor (n3158,n3156,n3091);
or (n3159,n3160,n3162);
and (n3160,n3161,n3097);
xor (n3161,n3093,n3094);
and (n3162,n3163,n3164);
xor (n3163,n3161,n3097);
or (n3164,n3165,n3167);
and (n3165,n3166,n3103);
xor (n3166,n3099,n3100);
and (n3167,n3168,n3169);
xor (n3168,n3166,n3103);
or (n3169,n3170,n3172);
and (n3170,n3171,n3109);
xor (n3171,n3105,n3106);
and (n3172,n3173,n3174);
xor (n3173,n3171,n3109);
or (n3174,n3175,n3177);
and (n3175,n3176,n3115);
xor (n3176,n3111,n3112);
and (n3177,n3178,n3179);
xor (n3178,n3176,n3115);
or (n3179,n3180,n3182);
and (n3180,n3181,n3121);
xor (n3181,n3117,n3118);
and (n3182,n3183,n3184);
xor (n3183,n3181,n3121);
or (n3184,n3185,n3187);
and (n3185,n3186,n3127);
xor (n3186,n3123,n3124);
and (n3187,n3188,n3189);
xor (n3188,n3186,n3127);
or (n3189,n3190,n3192);
and (n3190,n3191,n3133);
xor (n3191,n3129,n3130);
and (n3192,n3193,n3194);
xor (n3193,n3191,n3133);
and (n3194,n3195,n3138);
xor (n3195,n3135,n3136);
or (n3196,n3197,n3199);
and (n3197,n3198,n3079);
xor (n3198,n3143,n3144);
and (n3199,n3200,n3201);
xor (n3200,n3198,n3079);
or (n3201,n3202,n3204);
and (n3202,n3203,n3085);
xor (n3203,n3148,n3149);
and (n3204,n3205,n3206);
xor (n3205,n3203,n3085);
or (n3206,n3207,n3209);
and (n3207,n3208,n3091);
xor (n3208,n3153,n3154);
and (n3209,n3210,n3211);
xor (n3210,n3208,n3091);
or (n3211,n3212,n3214);
and (n3212,n3213,n3097);
xor (n3213,n3158,n3159);
and (n3214,n3215,n3216);
xor (n3215,n3213,n3097);
or (n3216,n3217,n3219);
and (n3217,n3218,n3103);
xor (n3218,n3163,n3164);
and (n3219,n3220,n3221);
xor (n3220,n3218,n3103);
or (n3221,n3222,n3224);
and (n3222,n3223,n3109);
xor (n3223,n3168,n3169);
and (n3224,n3225,n3226);
xor (n3225,n3223,n3109);
or (n3226,n3227,n3229);
and (n3227,n3228,n3115);
xor (n3228,n3173,n3174);
and (n3229,n3230,n3231);
xor (n3230,n3228,n3115);
or (n3231,n3232,n3234);
and (n3232,n3233,n3121);
xor (n3233,n3178,n3179);
and (n3234,n3235,n3236);
xor (n3235,n3233,n3121);
or (n3236,n3237,n3239);
and (n3237,n3238,n3127);
xor (n3238,n3183,n3184);
and (n3239,n3240,n3241);
xor (n3240,n3238,n3127);
or (n3241,n3242,n3244);
and (n3242,n3243,n3133);
xor (n3243,n3188,n3189);
and (n3244,n3245,n3246);
xor (n3245,n3243,n3133);
and (n3246,n3247,n3138);
xor (n3247,n3193,n3194);
or (n3248,n3249,n3251);
and (n3249,n3250,n3085);
xor (n3250,n3200,n3201);
and (n3251,n3252,n3253);
xor (n3252,n3250,n3085);
or (n3253,n3254,n3256);
and (n3254,n3255,n3091);
xor (n3255,n3205,n3206);
and (n3256,n3257,n3258);
xor (n3257,n3255,n3091);
or (n3258,n3259,n3261);
and (n3259,n3260,n3097);
xor (n3260,n3210,n3211);
and (n3261,n3262,n3263);
xor (n3262,n3260,n3097);
or (n3263,n3264,n3266);
and (n3264,n3265,n3103);
xor (n3265,n3215,n3216);
and (n3266,n3267,n3268);
xor (n3267,n3265,n3103);
or (n3268,n3269,n3271);
and (n3269,n3270,n3109);
xor (n3270,n3220,n3221);
and (n3271,n3272,n3273);
xor (n3272,n3270,n3109);
or (n3273,n3274,n3276);
and (n3274,n3275,n3115);
xor (n3275,n3225,n3226);
and (n3276,n3277,n3278);
xor (n3277,n3275,n3115);
or (n3278,n3279,n3281);
and (n3279,n3280,n3121);
xor (n3280,n3230,n3231);
and (n3281,n3282,n3283);
xor (n3282,n3280,n3121);
or (n3283,n3284,n3286);
and (n3284,n3285,n3127);
xor (n3285,n3235,n3236);
and (n3286,n3287,n3288);
xor (n3287,n3285,n3127);
or (n3288,n3289,n3291);
and (n3289,n3290,n3133);
xor (n3290,n3240,n3241);
and (n3291,n3292,n3293);
xor (n3292,n3290,n3133);
and (n3293,n3294,n3138);
xor (n3294,n3245,n3246);
or (n3295,n3296,n3298);
and (n3296,n3297,n3091);
xor (n3297,n3252,n3253);
and (n3298,n3299,n3300);
xor (n3299,n3297,n3091);
or (n3300,n3301,n3303);
and (n3301,n3302,n3097);
xor (n3302,n3257,n3258);
and (n3303,n3304,n3305);
xor (n3304,n3302,n3097);
or (n3305,n3306,n3308);
and (n3306,n3307,n3103);
xor (n3307,n3262,n3263);
and (n3308,n3309,n3310);
xor (n3309,n3307,n3103);
or (n3310,n3311,n3313);
and (n3311,n3312,n3109);
xor (n3312,n3267,n3268);
and (n3313,n3314,n3315);
xor (n3314,n3312,n3109);
or (n3315,n3316,n3318);
and (n3316,n3317,n3115);
xor (n3317,n3272,n3273);
and (n3318,n3319,n3320);
xor (n3319,n3317,n3115);
or (n3320,n3321,n3323);
and (n3321,n3322,n3121);
xor (n3322,n3277,n3278);
and (n3323,n3324,n3325);
xor (n3324,n3322,n3121);
or (n3325,n3326,n3328);
and (n3326,n3327,n3127);
xor (n3327,n3282,n3283);
and (n3328,n3329,n3330);
xor (n3329,n3327,n3127);
or (n3330,n3331,n3333);
and (n3331,n3332,n3133);
xor (n3332,n3287,n3288);
and (n3333,n3334,n3335);
xor (n3334,n3332,n3133);
and (n3335,n3336,n3138);
xor (n3336,n3292,n3293);
or (n3337,n3338,n3340);
and (n3338,n3339,n3097);
xor (n3339,n3299,n3300);
and (n3340,n3341,n3342);
xor (n3341,n3339,n3097);
or (n3342,n3343,n3345);
and (n3343,n3344,n3103);
xor (n3344,n3304,n3305);
and (n3345,n3346,n3347);
xor (n3346,n3344,n3103);
or (n3347,n3348,n3350);
and (n3348,n3349,n3109);
xor (n3349,n3309,n3310);
and (n3350,n3351,n3352);
xor (n3351,n3349,n3109);
or (n3352,n3353,n3355);
and (n3353,n3354,n3115);
xor (n3354,n3314,n3315);
and (n3355,n3356,n3357);
xor (n3356,n3354,n3115);
or (n3357,n3358,n3360);
and (n3358,n3359,n3121);
xor (n3359,n3319,n3320);
and (n3360,n3361,n3362);
xor (n3361,n3359,n3121);
or (n3362,n3363,n3365);
and (n3363,n3364,n3127);
xor (n3364,n3324,n3325);
and (n3365,n3366,n3367);
xor (n3366,n3364,n3127);
or (n3367,n3368,n3370);
and (n3368,n3369,n3133);
xor (n3369,n3329,n3330);
and (n3370,n3371,n3372);
xor (n3371,n3369,n3133);
and (n3372,n3373,n3138);
xor (n3373,n3334,n3335);
or (n3374,n3375,n3377);
and (n3375,n3376,n3103);
xor (n3376,n3341,n3342);
and (n3377,n3378,n3379);
xor (n3378,n3376,n3103);
or (n3379,n3380,n3382);
and (n3380,n3381,n3109);
xor (n3381,n3346,n3347);
and (n3382,n3383,n3384);
xor (n3383,n3381,n3109);
or (n3384,n3385,n3387);
and (n3385,n3386,n3115);
xor (n3386,n3351,n3352);
and (n3387,n3388,n3389);
xor (n3388,n3386,n3115);
or (n3389,n3390,n3392);
and (n3390,n3391,n3121);
xor (n3391,n3356,n3357);
and (n3392,n3393,n3394);
xor (n3393,n3391,n3121);
or (n3394,n3395,n3397);
and (n3395,n3396,n3127);
xor (n3396,n3361,n3362);
and (n3397,n3398,n3399);
xor (n3398,n3396,n3127);
or (n3399,n3400,n3402);
and (n3400,n3401,n3133);
xor (n3401,n3366,n3367);
and (n3402,n3403,n3404);
xor (n3403,n3401,n3133);
and (n3404,n3405,n3138);
xor (n3405,n3371,n3372);
or (n3406,n3407,n3409);
and (n3407,n3408,n3109);
xor (n3408,n3378,n3379);
and (n3409,n3410,n3411);
xor (n3410,n3408,n3109);
or (n3411,n3412,n3414);
and (n3412,n3413,n3115);
xor (n3413,n3383,n3384);
and (n3414,n3415,n3416);
xor (n3415,n3413,n3115);
or (n3416,n3417,n3419);
and (n3417,n3418,n3121);
xor (n3418,n3388,n3389);
and (n3419,n3420,n3421);
xor (n3420,n3418,n3121);
or (n3421,n3422,n3424);
and (n3422,n3423,n3127);
xor (n3423,n3393,n3394);
and (n3424,n3425,n3426);
xor (n3425,n3423,n3127);
or (n3426,n3427,n3429);
and (n3427,n3428,n3133);
xor (n3428,n3398,n3399);
and (n3429,n3430,n3431);
xor (n3430,n3428,n3133);
and (n3431,n3432,n3138);
xor (n3432,n3403,n3404);
or (n3433,n3434,n3436);
and (n3434,n3435,n3115);
xor (n3435,n3410,n3411);
and (n3436,n3437,n3438);
xor (n3437,n3435,n3115);
or (n3438,n3439,n3441);
and (n3439,n3440,n3121);
xor (n3440,n3415,n3416);
and (n3441,n3442,n3443);
xor (n3442,n3440,n3121);
or (n3443,n3444,n3446);
and (n3444,n3445,n3127);
xor (n3445,n3420,n3421);
and (n3446,n3447,n3448);
xor (n3447,n3445,n3127);
or (n3448,n3449,n3451);
and (n3449,n3450,n3133);
xor (n3450,n3425,n3426);
and (n3451,n3452,n3453);
xor (n3452,n3450,n3133);
and (n3453,n3454,n3138);
xor (n3454,n3430,n3431);
or (n3455,n3456,n3458);
and (n3456,n3457,n3121);
xor (n3457,n3437,n3438);
and (n3458,n3459,n3460);
xor (n3459,n3457,n3121);
or (n3460,n3461,n3463);
and (n3461,n3462,n3127);
xor (n3462,n3442,n3443);
and (n3463,n3464,n3465);
xor (n3464,n3462,n3127);
or (n3465,n3466,n3468);
and (n3466,n3467,n3133);
xor (n3467,n3447,n3448);
and (n3468,n3469,n3470);
xor (n3469,n3467,n3133);
and (n3470,n3471,n3138);
xor (n3471,n3452,n3453);
or (n3472,n3473,n3475);
and (n3473,n3474,n3127);
xor (n3474,n3459,n3460);
and (n3475,n3476,n3477);
xor (n3476,n3474,n3127);
or (n3477,n3478,n3480);
and (n3478,n3479,n3133);
xor (n3479,n3464,n3465);
and (n3480,n3481,n3482);
xor (n3481,n3479,n3133);
and (n3482,n3483,n3138);
xor (n3483,n3469,n3470);
or (n3484,n3485,n3487);
and (n3485,n3486,n3133);
xor (n3486,n3476,n3477);
and (n3487,n3488,n3489);
xor (n3488,n3486,n3133);
and (n3489,n3490,n3138);
xor (n3490,n3481,n3482);
and (n3491,n3492,n3138);
xor (n3492,n3488,n3489);
endmodule
