module top (out,n5,n6,n15,n19,n20,n23,n24,n55,n61
        ,n70,n107,n111,n159,n189,n242,n344,n353,n356,n359
        ,n389,n440,n515,n567);
output out;
input n5;
input n6;
input n15;
input n19;
input n20;
input n23;
input n24;
input n55;
input n61;
input n70;
input n107;
input n111;
input n159;
input n189;
input n242;
input n344;
input n353;
input n356;
input n359;
input n389;
input n440;
input n515;
input n567;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n16;
wire n17;
wire n18;
wire n21;
wire n22;
wire n25;
wire n26;
wire n27;
wire n28;
wire n29;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n108;
wire n109;
wire n110;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n354;
wire n355;
wire n357;
wire n358;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
xor (out,n0,n751);
xor (n0,n1,n666);
xor (n1,n2,n341);
or (n2,n3,n41);
and (n3,n4,n7);
and (n4,n5,n6);
or (n7,n8,n35,n40);
and (n8,n9,n32);
or (n9,n10,n29,n31);
and (n10,n11,n26);
or (n11,n12,n21,n25);
and (n12,n13,n18);
nor (n13,n14,n16);
not (n14,n15);
and (n16,n17,n15);
not (n17,n6);
and (n18,n19,n20);
and (n21,n18,n22);
and (n22,n23,n24);
and (n25,n13,n22);
nor (n26,n27,n28);
not (n27,n19);
and (n28,n17,n19);
and (n29,n26,n30);
and (n30,n23,n20);
and (n31,n11,n30);
nor (n32,n33,n34);
not (n33,n23);
and (n34,n17,n23);
and (n35,n32,n36);
nor (n36,n37,n39);
and (n37,n38,n20);
not (n38,n5);
not (n39,n20);
and (n40,n9,n36);
and (n41,n42,n43);
xor (n42,n4,n7);
or (n43,n44,n89);
and (n44,n45,n47);
xor (n45,n46,n36);
xor (n46,n9,n32);
or (n47,n48,n85,n88);
and (n48,n49,n82);
or (n49,n50,n78,n81);
and (n50,n51,n64);
or (n51,n52,n58,n63);
and (n52,n53,n57);
nor (n53,n54,n56);
not (n54,n55);
and (n56,n17,n55);
and (n57,n15,n20);
and (n58,n57,n59);
nor (n59,n60,n62);
and (n60,n38,n61);
not (n62,n61);
and (n63,n53,n59);
or (n64,n65,n75,n77);
and (n65,n66,n74);
or (n66,n67,n71,n73);
and (n67,n68,n69);
and (n68,n15,n24);
and (n69,n19,n70);
and (n71,n69,n72);
and (n72,n23,n61);
and (n73,n68,n72);
and (n74,n19,n24);
and (n75,n74,n76);
and (n76,n23,n70);
and (n77,n66,n76);
and (n78,n64,n79);
xor (n79,n80,n22);
xor (n80,n13,n18);
and (n81,n51,n79);
nor (n82,n83,n84);
and (n83,n38,n24);
not (n84,n24);
and (n85,n82,n86);
xor (n86,n87,n30);
xor (n87,n11,n26);
and (n88,n49,n86);
and (n89,n90,n91);
xor (n90,n45,n47);
or (n91,n92,n130);
and (n92,n93,n95);
xor (n93,n94,n86);
xor (n94,n49,n82);
or (n95,n96,n126,n129);
and (n96,n97,n123);
or (n97,n98,n119,n122);
and (n98,n99,n117);
or (n99,n100,n113,n116);
and (n100,n101,n109);
or (n101,n102,n105,n108);
and (n102,n103,n104);
and (n103,n15,n70);
and (n104,n19,n61);
and (n105,n104,n106);
and (n106,n23,n107);
and (n108,n103,n106);
and (n109,n110,n112);
and (n110,n111,n20);
and (n112,n55,n24);
and (n113,n109,n114);
xor (n114,n115,n72);
xor (n115,n68,n69);
and (n116,n101,n114);
xor (n117,n118,n59);
xor (n118,n53,n57);
and (n119,n117,n120);
xor (n120,n121,n76);
xor (n121,n66,n74);
and (n122,n99,n120);
nor (n123,n124,n125);
and (n124,n38,n70);
not (n125,n70);
and (n126,n123,n127);
xor (n127,n128,n79);
xor (n128,n51,n64);
and (n129,n97,n127);
and (n130,n131,n132);
xor (n131,n93,n95);
or (n132,n133,n176);
and (n133,n134,n136);
xor (n134,n135,n127);
xor (n135,n97,n123);
or (n136,n137,n172,n175);
and (n137,n138,n149);
or (n138,n139,n144,n148);
and (n139,n140,n143);
nor (n140,n141,n142);
not (n141,n111);
and (n142,n17,n111);
and (n143,n55,n20);
and (n144,n143,n145);
nor (n145,n146,n147);
and (n146,n38,n107);
not (n147,n107);
and (n148,n140,n145);
or (n149,n150,n168,n171);
and (n150,n151,n166);
or (n151,n152,n163,n165);
and (n152,n153,n161);
or (n153,n154,n157,n160);
and (n154,n155,n156);
and (n155,n15,n61);
and (n156,n19,n107);
and (n157,n156,n158);
and (n158,n23,n159);
and (n160,n155,n158);
xor (n161,n162,n106);
xor (n162,n103,n104);
and (n163,n161,n164);
xor (n164,n110,n112);
and (n165,n153,n164);
xor (n166,n167,n145);
xor (n167,n140,n143);
and (n168,n166,n169);
xor (n169,n170,n114);
xor (n170,n101,n109);
and (n171,n151,n169);
and (n172,n149,n173);
xor (n173,n174,n120);
xor (n174,n99,n117);
and (n175,n138,n173);
and (n176,n177,n178);
xor (n177,n134,n136);
or (n178,n179,n225);
and (n179,n180,n182);
xor (n180,n181,n173);
xor (n181,n138,n149);
or (n182,n183,n221,n224);
and (n183,n184,n202);
or (n184,n185,n197,n201);
and (n185,n186,n194);
or (n186,n187,n191,n193);
and (n187,n188,n190);
and (n188,n189,n20);
and (n190,n111,n24);
and (n191,n190,n192);
and (n192,n55,n70);
and (n193,n188,n192);
nor (n194,n195,n196);
not (n195,n189);
and (n196,n17,n189);
and (n197,n194,n198);
nor (n198,n199,n200);
and (n199,n38,n159);
not (n200,n159);
and (n201,n186,n198);
or (n202,n203,n217,n220);
and (n203,n204,n215);
or (n204,n205,n211,n214);
and (n205,n206,n209);
and (n206,n207,n208);
and (n207,n15,n107);
and (n208,n19,n159);
xor (n209,n210,n192);
xor (n210,n188,n190);
and (n211,n209,n212);
xor (n212,n213,n158);
xor (n213,n155,n156);
and (n214,n206,n212);
xor (n215,n216,n198);
xor (n216,n186,n194);
and (n217,n215,n218);
xor (n218,n219,n164);
xor (n219,n153,n161);
and (n220,n204,n218);
and (n221,n202,n222);
xor (n222,n223,n169);
xor (n223,n151,n166);
and (n224,n184,n222);
and (n225,n226,n227);
xor (n226,n180,n182);
or (n227,n228,n247);
and (n228,n229,n231);
xor (n229,n230,n222);
xor (n230,n184,n202);
and (n231,n232,n245);
or (n232,n233,n239,n244);
and (n233,n234,n237);
and (n234,n235,n236);
and (n235,n55,n61);
xor (n236,n207,n208);
xor (n237,n238,n212);
xor (n238,n206,n209);
and (n239,n237,n240);
nor (n240,n241,n243);
not (n241,n242);
and (n243,n17,n242);
and (n244,n234,n240);
xor (n245,n246,n218);
xor (n246,n204,n215);
and (n247,n248,n249);
xor (n248,n229,n231);
or (n249,n250,n280);
and (n250,n251,n252);
xor (n251,n232,n245);
or (n252,n253,n276,n279);
and (n253,n254,n261);
or (n254,n255,n258,n260);
and (n255,n256,n257);
and (n256,n242,n20);
and (n257,n189,n24);
and (n258,n257,n259);
and (n259,n111,n70);
and (n260,n256,n259);
or (n261,n262,n273,n275);
and (n262,n263,n271);
or (n263,n264,n267,n270);
and (n264,n265,n266);
and (n265,n111,n107);
and (n266,n55,n159);
and (n267,n268,n269);
and (n268,n55,n107);
and (n269,n15,n159);
and (n270,n264,n269);
xor (n271,n272,n259);
xor (n272,n256,n257);
and (n273,n271,n274);
xor (n274,n235,n236);
and (n275,n263,n274);
and (n276,n261,n277);
xor (n277,n278,n240);
xor (n278,n234,n237);
and (n279,n254,n277);
and (n280,n281,n282);
xor (n281,n251,n252);
or (n282,n283,n311);
and (n283,n284,n286);
xor (n284,n285,n277);
xor (n285,n254,n261);
or (n286,n287,n307,n310);
and (n287,n288,n291);
and (n288,n289,n290);
and (n289,n189,n70);
and (n290,n111,n61);
or (n291,n292,n303,n306);
and (n292,n293,n302);
or (n293,n294,n299,n301);
and (n294,n295,n298);
and (n295,n296,n297);
and (n296,n189,n107);
and (n297,n111,n159);
and (n298,n189,n61);
and (n299,n298,n300);
xor (n300,n265,n266);
and (n301,n295,n300);
xor (n302,n289,n290);
and (n303,n302,n304);
xor (n304,n305,n269);
xor (n305,n264,n268);
and (n306,n293,n304);
and (n307,n291,n308);
xor (n308,n309,n274);
xor (n309,n263,n271);
and (n310,n288,n308);
and (n311,n312,n313);
xor (n312,n284,n286);
or (n313,n314,n336);
and (n314,n315,n317);
xor (n315,n316,n308);
xor (n316,n288,n291);
and (n317,n318,n334);
or (n318,n319,n330,n333);
and (n319,n320,n329);
or (n320,n321,n326,n328);
and (n321,n322,n325);
and (n322,n323,n324);
and (n323,n242,n107);
and (n324,n189,n159);
and (n325,n242,n61);
and (n326,n325,n327);
xor (n327,n296,n297);
and (n328,n322,n327);
and (n329,n242,n70);
and (n330,n329,n331);
xor (n331,n332,n300);
xor (n332,n295,n298);
and (n333,n320,n331);
xor (n334,n335,n304);
xor (n335,n293,n302);
and (n336,n337,n338);
xor (n337,n315,n317);
and (n338,n339,n340);
and (n339,n242,n24);
xor (n340,n318,n334);
or (n341,n342,n375);
and (n342,n343,n345);
and (n343,n344,n6);
or (n345,n346,n370,n374);
and (n346,n347,n367);
or (n347,n348,n364,n366);
and (n348,n349,n361);
or (n349,n350,n357,n360);
and (n350,n351,n355);
nor (n351,n352,n354);
not (n352,n353);
and (n354,n17,n353);
and (n355,n356,n20);
and (n357,n355,n358);
and (n358,n359,n24);
and (n360,n351,n358);
nor (n361,n362,n363);
not (n362,n356);
and (n363,n17,n356);
and (n364,n361,n365);
and (n365,n359,n20);
and (n366,n349,n365);
nor (n367,n368,n369);
not (n368,n359);
and (n369,n17,n359);
and (n370,n367,n371);
nor (n371,n372,n39);
and (n372,n373,n20);
not (n373,n344);
and (n374,n347,n371);
and (n375,n376,n377);
xor (n376,n343,n345);
or (n377,n378,n419);
and (n378,n379,n381);
xor (n379,n380,n371);
xor (n380,n347,n367);
or (n381,n382,n415,n418);
and (n382,n383,n413);
or (n383,n384,n409,n412);
and (n384,n385,n396);
or (n385,n386,n392,n395);
and (n386,n387,n391);
nor (n387,n388,n390);
not (n388,n389);
and (n390,n17,n389);
and (n391,n353,n20);
and (n392,n391,n393);
nor (n393,n394,n62);
and (n394,n373,n61);
and (n395,n387,n393);
or (n396,n397,n406,n408);
and (n397,n398,n405);
or (n398,n399,n402,n404);
and (n399,n400,n401);
and (n400,n353,n24);
and (n401,n356,n70);
and (n402,n401,n403);
and (n403,n359,n61);
and (n404,n400,n403);
and (n405,n356,n24);
and (n406,n405,n407);
and (n407,n359,n70);
and (n408,n398,n407);
and (n409,n396,n410);
xor (n410,n411,n358);
xor (n411,n351,n355);
and (n412,n385,n410);
nor (n413,n414,n84);
and (n414,n373,n24);
and (n415,n413,n416);
xor (n416,n417,n365);
xor (n417,n349,n361);
and (n418,n383,n416);
and (n419,n420,n421);
xor (n420,n379,n381);
or (n421,n422,n458);
and (n422,n423,n425);
xor (n423,n424,n416);
xor (n424,n383,n413);
or (n425,n426,n454,n457);
and (n426,n427,n452);
or (n427,n428,n448,n451);
and (n428,n429,n446);
or (n429,n430,n442,n445);
and (n430,n431,n438);
or (n431,n432,n435,n437);
and (n432,n433,n434);
and (n433,n353,n70);
and (n434,n356,n61);
and (n435,n434,n436);
and (n436,n359,n107);
and (n437,n433,n436);
and (n438,n439,n441);
and (n439,n440,n20);
and (n441,n389,n24);
and (n442,n438,n443);
xor (n443,n444,n403);
xor (n444,n400,n401);
and (n445,n431,n443);
xor (n446,n447,n393);
xor (n447,n387,n391);
and (n448,n446,n449);
xor (n449,n450,n407);
xor (n450,n398,n405);
and (n451,n429,n449);
nor (n452,n453,n125);
and (n453,n373,n70);
and (n454,n452,n455);
xor (n455,n456,n410);
xor (n456,n385,n396);
and (n457,n427,n455);
and (n458,n459,n460);
xor (n459,n423,n425);
or (n460,n461,n502);
and (n461,n462,n464);
xor (n462,n463,n455);
xor (n463,n427,n452);
or (n464,n465,n498,n501);
and (n465,n466,n476);
or (n466,n467,n472,n475);
and (n467,n468,n471);
nor (n468,n469,n470);
not (n469,n440);
and (n470,n17,n440);
and (n471,n389,n20);
and (n472,n471,n473);
nor (n473,n474,n147);
and (n474,n373,n107);
and (n475,n468,n473);
or (n476,n477,n494,n497);
and (n477,n478,n492);
or (n478,n479,n489,n491);
and (n479,n480,n487);
or (n480,n481,n484,n486);
and (n481,n482,n483);
and (n482,n353,n61);
and (n483,n356,n107);
and (n484,n483,n485);
and (n485,n359,n159);
and (n486,n482,n485);
xor (n487,n488,n436);
xor (n488,n433,n434);
and (n489,n487,n490);
xor (n490,n439,n441);
and (n491,n480,n490);
xor (n492,n493,n473);
xor (n493,n468,n471);
and (n494,n492,n495);
xor (n495,n496,n443);
xor (n496,n431,n438);
and (n497,n478,n495);
and (n498,n476,n499);
xor (n499,n500,n449);
xor (n500,n429,n446);
and (n501,n466,n499);
and (n502,n503,n504);
xor (n503,n462,n464);
or (n504,n505,n550);
and (n505,n506,n508);
xor (n506,n507,n499);
xor (n507,n466,n476);
or (n508,n509,n546,n549);
and (n509,n510,n527);
or (n510,n511,n523,n526);
and (n511,n512,n520);
or (n512,n513,n517,n519);
and (n513,n514,n516);
and (n514,n515,n20);
and (n516,n440,n24);
and (n517,n516,n518);
and (n518,n389,n70);
and (n519,n514,n518);
nor (n520,n521,n522);
not (n521,n515);
and (n522,n17,n515);
and (n523,n520,n524);
nor (n524,n525,n200);
and (n525,n373,n159);
and (n526,n512,n524);
or (n527,n528,n542,n545);
and (n528,n529,n540);
or (n529,n530,n536,n539);
and (n530,n531,n534);
and (n531,n532,n533);
and (n532,n353,n107);
and (n533,n356,n159);
xor (n534,n535,n518);
xor (n535,n514,n516);
and (n536,n534,n537);
xor (n537,n538,n485);
xor (n538,n482,n483);
and (n539,n531,n537);
xor (n540,n541,n524);
xor (n541,n512,n520);
and (n542,n540,n543);
xor (n543,n544,n490);
xor (n544,n480,n487);
and (n545,n529,n543);
and (n546,n527,n547);
xor (n547,n548,n495);
xor (n548,n478,n492);
and (n549,n510,n547);
and (n550,n551,n552);
xor (n551,n506,n508);
or (n552,n553,n572);
and (n553,n554,n556);
xor (n554,n555,n547);
xor (n555,n510,n527);
and (n556,n557,n570);
or (n557,n558,n564,n569);
and (n558,n559,n562);
and (n559,n560,n561);
and (n560,n389,n61);
xor (n561,n532,n533);
xor (n562,n563,n537);
xor (n563,n531,n534);
and (n564,n562,n565);
nor (n565,n566,n568);
not (n566,n567);
and (n568,n17,n567);
and (n569,n559,n565);
xor (n570,n571,n543);
xor (n571,n529,n540);
and (n572,n573,n574);
xor (n573,n554,n556);
or (n574,n575,n605);
and (n575,n576,n577);
xor (n576,n557,n570);
or (n577,n578,n601,n604);
and (n578,n579,n586);
or (n579,n580,n583,n585);
and (n580,n581,n582);
and (n581,n567,n20);
and (n582,n515,n24);
and (n583,n582,n584);
and (n584,n440,n70);
and (n585,n581,n584);
or (n586,n587,n598,n600);
and (n587,n588,n596);
or (n588,n589,n592,n595);
and (n589,n590,n591);
and (n590,n440,n107);
and (n591,n389,n159);
and (n592,n593,n594);
and (n593,n389,n107);
and (n594,n353,n159);
and (n595,n589,n594);
xor (n596,n597,n584);
xor (n597,n581,n582);
and (n598,n596,n599);
xor (n599,n560,n561);
and (n600,n588,n599);
and (n601,n586,n602);
xor (n602,n603,n565);
xor (n603,n559,n562);
and (n604,n579,n602);
and (n605,n606,n607);
xor (n606,n576,n577);
or (n607,n608,n636);
and (n608,n609,n611);
xor (n609,n610,n602);
xor (n610,n579,n586);
or (n611,n612,n632,n635);
and (n612,n613,n616);
and (n613,n614,n615);
and (n614,n515,n70);
and (n615,n440,n61);
or (n616,n617,n628,n631);
and (n617,n618,n627);
or (n618,n619,n624,n626);
and (n619,n620,n623);
and (n620,n621,n622);
and (n621,n515,n107);
and (n622,n440,n159);
and (n623,n515,n61);
and (n624,n623,n625);
xor (n625,n590,n591);
and (n626,n620,n625);
xor (n627,n614,n615);
and (n628,n627,n629);
xor (n629,n630,n594);
xor (n630,n589,n593);
and (n631,n618,n629);
and (n632,n616,n633);
xor (n633,n634,n599);
xor (n634,n588,n596);
and (n635,n613,n633);
and (n636,n637,n638);
xor (n637,n609,n611);
or (n638,n639,n661);
and (n639,n640,n642);
xor (n640,n641,n633);
xor (n641,n613,n616);
and (n642,n643,n659);
or (n643,n644,n655,n658);
and (n644,n645,n654);
or (n645,n646,n651,n653);
and (n646,n647,n650);
and (n647,n648,n649);
and (n648,n567,n107);
and (n649,n515,n159);
and (n650,n567,n61);
and (n651,n650,n652);
xor (n652,n621,n622);
and (n653,n647,n652);
and (n654,n567,n70);
and (n655,n654,n656);
xor (n656,n657,n625);
xor (n657,n620,n623);
and (n658,n645,n656);
xor (n659,n660,n629);
xor (n660,n618,n627);
and (n661,n662,n663);
xor (n662,n640,n642);
and (n663,n664,n665);
and (n664,n567,n24);
xor (n665,n643,n659);
or (n666,n667,n670,n750);
and (n667,n668,n669);
xor (n668,n42,n43);
xor (n669,n376,n377);
and (n670,n669,n671);
or (n671,n672,n675,n749);
and (n672,n673,n674);
xor (n673,n90,n91);
xor (n674,n420,n421);
and (n675,n674,n676);
or (n676,n677,n680,n748);
and (n677,n678,n679);
xor (n678,n131,n132);
xor (n679,n459,n460);
and (n680,n679,n681);
or (n681,n682,n685,n747);
and (n682,n683,n684);
xor (n683,n177,n178);
xor (n684,n503,n504);
and (n685,n684,n686);
or (n686,n687,n690,n746);
and (n687,n688,n689);
xor (n688,n226,n227);
xor (n689,n551,n552);
and (n690,n689,n691);
or (n691,n692,n695,n745);
and (n692,n693,n694);
xor (n693,n248,n249);
xor (n694,n573,n574);
and (n695,n694,n696);
or (n696,n697,n700,n744);
and (n697,n698,n699);
xor (n698,n281,n282);
xor (n699,n606,n607);
and (n700,n699,n701);
or (n701,n702,n705,n743);
and (n702,n703,n704);
xor (n703,n312,n313);
xor (n704,n637,n638);
and (n705,n704,n706);
or (n706,n707,n710,n742);
and (n707,n708,n709);
xor (n708,n337,n338);
xor (n709,n662,n663);
and (n710,n709,n711);
or (n711,n712,n715,n741);
and (n712,n713,n714);
xor (n713,n339,n340);
xor (n714,n664,n665);
and (n715,n714,n716);
or (n716,n717,n722,n740);
and (n717,n718,n720);
xor (n718,n719,n331);
xor (n719,n320,n329);
xor (n720,n721,n656);
xor (n721,n645,n654);
and (n722,n720,n723);
or (n723,n724,n729,n739);
and (n724,n725,n727);
xor (n725,n726,n327);
xor (n726,n322,n325);
xor (n727,n728,n652);
xor (n728,n647,n650);
and (n729,n727,n730);
or (n730,n731,n734,n738);
and (n731,n732,n733);
xor (n732,n323,n324);
xor (n733,n648,n649);
and (n734,n733,n735);
and (n735,n736,n737);
and (n736,n242,n159);
and (n737,n567,n159);
and (n738,n732,n735);
and (n739,n725,n730);
and (n740,n718,n723);
and (n741,n713,n716);
and (n742,n708,n711);
and (n743,n703,n706);
and (n744,n698,n701);
and (n745,n693,n696);
and (n746,n688,n691);
and (n747,n683,n686);
and (n748,n678,n681);
and (n749,n673,n676);
and (n750,n668,n671);
xor (n751,n752,n816);
xor (n752,n753,n783);
and (n753,n754,n6);
or (n754,n755,n756,n782);
and (n755,n5,n344);
and (n756,n344,n757);
or (n757,n758,n759,n781);
and (n758,n23,n359);
and (n759,n359,n760);
or (n760,n761,n762,n780);
and (n761,n19,n356);
and (n762,n356,n763);
or (n763,n764,n765,n779);
and (n764,n15,n353);
and (n765,n353,n766);
or (n766,n767,n768,n778);
and (n767,n55,n389);
and (n768,n389,n769);
or (n769,n770,n771,n777);
and (n770,n111,n440);
and (n771,n440,n772);
or (n772,n773,n774,n776);
and (n773,n189,n515);
and (n774,n515,n775);
and (n775,n242,n567);
and (n776,n189,n775);
and (n777,n111,n772);
and (n778,n55,n769);
and (n779,n15,n766);
and (n780,n19,n763);
and (n781,n23,n760);
and (n782,n5,n757);
or (n783,n784,n811,n815);
and (n784,n785,n808);
or (n785,n786,n805,n807);
and (n786,n787,n802);
or (n787,n788,n797,n801);
and (n788,n789,n794);
nor (n789,n790,n793);
not (n790,n791);
xor (n791,n792,n763);
xor (n792,n19,n356);
and (n793,n17,n791);
and (n794,n795,n20);
xor (n795,n796,n760);
xor (n796,n23,n359);
and (n797,n794,n798);
and (n798,n799,n24);
xor (n799,n800,n757);
xor (n800,n5,n344);
and (n801,n789,n798);
nor (n802,n803,n804);
not (n803,n795);
and (n804,n17,n795);
and (n805,n802,n806);
and (n806,n799,n20);
and (n807,n787,n806);
nor (n808,n809,n810);
not (n809,n799);
and (n810,n17,n799);
and (n811,n808,n812);
nor (n812,n813,n39);
and (n813,n814,n20);
not (n814,n754);
and (n815,n785,n812);
or (n816,n817,n859);
and (n817,n818,n820);
xor (n818,n819,n812);
xor (n819,n785,n808);
or (n820,n821,n855,n858);
and (n821,n822,n853);
or (n822,n823,n849,n852);
and (n823,n824,n836);
or (n824,n825,n832,n835);
and (n825,n826,n831);
nor (n826,n827,n830);
not (n827,n828);
xor (n828,n829,n766);
xor (n829,n15,n353);
and (n830,n17,n828);
and (n831,n791,n20);
and (n832,n831,n833);
nor (n833,n834,n62);
and (n834,n814,n61);
and (n835,n826,n833);
or (n836,n837,n846,n848);
and (n837,n838,n845);
or (n838,n839,n842,n844);
and (n839,n840,n841);
and (n840,n791,n24);
and (n841,n795,n70);
and (n842,n841,n843);
and (n843,n799,n61);
and (n844,n840,n843);
and (n845,n795,n24);
and (n846,n845,n847);
and (n847,n799,n70);
and (n848,n838,n847);
and (n849,n836,n850);
xor (n850,n851,n798);
xor (n851,n789,n794);
and (n852,n824,n850);
nor (n853,n854,n84);
and (n854,n814,n24);
and (n855,n853,n856);
xor (n856,n857,n806);
xor (n857,n787,n802);
and (n858,n822,n856);
and (n859,n860,n861);
xor (n860,n818,n820);
or (n861,n862,n907);
and (n862,n863,n865);
xor (n863,n864,n856);
xor (n864,n822,n853);
or (n865,n866,n903,n906);
and (n866,n867,n901);
or (n867,n868,n897,n900);
and (n868,n869,n895);
or (n869,n870,n891,n894);
and (n870,n871,n878);
or (n871,n872,n875,n877);
and (n872,n873,n874);
and (n873,n791,n70);
and (n874,n795,n61);
and (n875,n874,n876);
and (n876,n799,n107);
and (n877,n873,n876);
or (n878,n879,n888,n890);
and (n879,n880,n885);
nor (n880,n881,n884);
not (n881,n882);
xor (n882,n883,n772);
xor (n883,n111,n440);
and (n884,n17,n882);
and (n885,n886,n20);
xor (n886,n887,n769);
xor (n887,n55,n389);
and (n888,n885,n889);
and (n889,n828,n24);
and (n890,n880,n889);
and (n891,n878,n892);
xor (n892,n893,n843);
xor (n893,n840,n841);
and (n894,n871,n892);
xor (n895,n896,n833);
xor (n896,n826,n831);
and (n897,n895,n898);
xor (n898,n899,n847);
xor (n899,n838,n845);
and (n900,n869,n898);
nor (n901,n902,n125);
and (n902,n814,n70);
and (n903,n901,n904);
xor (n904,n905,n850);
xor (n905,n824,n836);
and (n906,n867,n904);
and (n907,n908,n909);
xor (n908,n863,n865);
or (n909,n910,n952);
and (n910,n911,n913);
xor (n911,n912,n904);
xor (n912,n867,n901);
or (n913,n914,n948,n951);
and (n914,n915,n925);
or (n915,n916,n921,n924);
and (n916,n917,n920);
nor (n917,n918,n919);
not (n918,n886);
and (n919,n17,n886);
and (n920,n828,n20);
and (n921,n920,n922);
nor (n922,n923,n147);
and (n923,n814,n107);
and (n924,n917,n922);
or (n925,n926,n944,n947);
and (n926,n927,n942);
or (n927,n928,n938,n941);
and (n928,n929,n936);
or (n929,n930,n933,n935);
and (n930,n931,n932);
and (n931,n791,n61);
and (n932,n795,n107);
and (n933,n932,n934);
and (n934,n799,n159);
and (n935,n931,n934);
xor (n936,n937,n876);
xor (n937,n873,n874);
and (n938,n936,n939);
xor (n939,n940,n889);
xor (n940,n880,n885);
and (n941,n929,n939);
xor (n942,n943,n922);
xor (n943,n917,n920);
and (n944,n942,n945);
xor (n945,n946,n892);
xor (n946,n871,n878);
and (n947,n927,n945);
and (n948,n925,n949);
xor (n949,n950,n898);
xor (n950,n869,n895);
and (n951,n915,n949);
and (n952,n953,n954);
xor (n953,n911,n913);
or (n954,n955,n994);
and (n955,n956,n958);
xor (n956,n957,n949);
xor (n957,n915,n925);
or (n958,n959,n990,n993);
and (n959,n960,n970);
and (n960,n961,n968);
or (n961,n962,n965,n967);
and (n962,n963,n964);
and (n963,n882,n20);
and (n964,n886,n24);
and (n965,n964,n966);
and (n966,n828,n70);
and (n967,n963,n966);
nor (n968,n969,n200);
and (n969,n814,n159);
or (n970,n971,n987,n989);
and (n971,n972,n985);
or (n972,n973,n981,n984);
and (n973,n974,n979);
nor (n974,n975,n978);
not (n975,n976);
xor (n976,n977,n775);
xor (n977,n189,n515);
and (n978,n17,n976);
xor (n979,n980,n934);
xor (n980,n931,n932);
and (n981,n979,n982);
xor (n982,n983,n966);
xor (n983,n963,n964);
and (n984,n974,n982);
xor (n985,n986,n939);
xor (n986,n929,n936);
and (n987,n985,n988);
xor (n988,n961,n968);
and (n989,n972,n988);
and (n990,n970,n991);
xor (n991,n992,n945);
xor (n992,n927,n942);
and (n993,n960,n991);
and (n994,n995,n996);
xor (n995,n956,n958);
or (n996,n997,n1034);
and (n997,n998,n1000);
xor (n998,n999,n991);
xor (n999,n960,n970);
or (n1000,n1001,n1030,n1033);
and (n1001,n1002,n1013);
and (n1002,n1003,n1010);
or (n1003,n1004,n1007,n1009);
and (n1004,n1005,n1006);
and (n1005,n882,n24);
and (n1006,n886,n70);
and (n1007,n1006,n1008);
and (n1008,n828,n61);
and (n1009,n1005,n1008);
and (n1010,n1011,n1012);
and (n1011,n791,n107);
and (n1012,n795,n159);
or (n1013,n1014,n1026,n1029);
and (n1014,n1015,n1025);
or (n1015,n1016,n1022,n1024);
and (n1016,n1017,n1020);
and (n1017,n1018,n1019);
and (n1018,n828,n107);
and (n1019,n791,n159);
xor (n1020,n1021,n1008);
xor (n1021,n1005,n1006);
and (n1022,n1020,n1023);
xor (n1023,n1011,n1012);
and (n1024,n1017,n1023);
xor (n1025,n1003,n1010);
and (n1026,n1025,n1027);
xor (n1027,n1028,n982);
xor (n1028,n974,n979);
and (n1029,n1015,n1027);
and (n1030,n1013,n1031);
xor (n1031,n1032,n988);
xor (n1032,n972,n985);
and (n1033,n1002,n1031);
and (n1034,n1035,n1036);
xor (n1035,n998,n1000);
or (n1036,n1037,n1062);
and (n1037,n1038,n1040);
xor (n1038,n1039,n1031);
xor (n1039,n1002,n1013);
or (n1040,n1041,n1058,n1061);
and (n1041,n1042,n1048);
and (n1042,n1043,n1047);
nor (n1043,n1044,n1046);
not (n1044,n1045);
xor (n1045,n242,n567);
and (n1046,n17,n1045);
and (n1047,n976,n20);
or (n1048,n1049,n1055,n1057);
and (n1049,n1050,n1053);
and (n1050,n1051,n1052);
and (n1051,n886,n61);
xor (n1052,n1018,n1019);
xor (n1053,n1054,n1023);
xor (n1054,n1017,n1020);
and (n1055,n1053,n1056);
xor (n1056,n1043,n1047);
and (n1057,n1050,n1056);
and (n1058,n1048,n1059);
xor (n1059,n1060,n1027);
xor (n1060,n1015,n1025);
and (n1061,n1042,n1059);
and (n1062,n1063,n1064);
xor (n1063,n1038,n1040);
or (n1064,n1065,n1096);
and (n1065,n1066,n1068);
xor (n1066,n1067,n1059);
xor (n1067,n1042,n1048);
or (n1068,n1069,n1092,n1095);
and (n1069,n1070,n1077);
or (n1070,n1071,n1074,n1076);
and (n1071,n1072,n1073);
and (n1072,n1045,n20);
and (n1073,n976,n24);
and (n1074,n1073,n1075);
and (n1075,n882,n70);
and (n1076,n1072,n1075);
or (n1077,n1078,n1089,n1091);
and (n1078,n1079,n1087);
or (n1079,n1080,n1083,n1086);
and (n1080,n1081,n1082);
and (n1081,n882,n107);
and (n1082,n886,n159);
and (n1083,n1084,n1085);
and (n1084,n886,n107);
and (n1085,n828,n159);
and (n1086,n1080,n1085);
xor (n1087,n1088,n1075);
xor (n1088,n1072,n1073);
and (n1089,n1087,n1090);
xor (n1090,n1051,n1052);
and (n1091,n1079,n1090);
and (n1092,n1077,n1093);
xor (n1093,n1094,n1056);
xor (n1094,n1050,n1053);
and (n1095,n1070,n1093);
and (n1096,n1097,n1098);
xor (n1097,n1066,n1068);
or (n1098,n1099,n1127);
and (n1099,n1100,n1102);
xor (n1100,n1101,n1093);
xor (n1101,n1070,n1077);
or (n1102,n1103,n1123,n1126);
and (n1103,n1104,n1107);
and (n1104,n1105,n1106);
and (n1105,n976,n70);
and (n1106,n882,n61);
or (n1107,n1108,n1119,n1122);
and (n1108,n1109,n1118);
or (n1109,n1110,n1115,n1117);
and (n1110,n1111,n1114);
and (n1111,n1112,n1113);
and (n1112,n976,n107);
and (n1113,n882,n159);
and (n1114,n976,n61);
and (n1115,n1114,n1116);
xor (n1116,n1081,n1082);
and (n1117,n1111,n1116);
xor (n1118,n1105,n1106);
and (n1119,n1118,n1120);
xor (n1120,n1121,n1085);
xor (n1121,n1080,n1084);
and (n1122,n1109,n1120);
and (n1123,n1107,n1124);
xor (n1124,n1125,n1090);
xor (n1125,n1079,n1087);
and (n1126,n1104,n1124);
and (n1127,n1128,n1129);
xor (n1128,n1100,n1102);
or (n1129,n1130,n1152);
and (n1130,n1131,n1133);
xor (n1131,n1132,n1124);
xor (n1132,n1104,n1107);
and (n1133,n1134,n1150);
or (n1134,n1135,n1146,n1149);
and (n1135,n1136,n1145);
or (n1136,n1137,n1142,n1144);
and (n1137,n1138,n1141);
and (n1138,n1139,n1140);
and (n1139,n1045,n107);
and (n1140,n976,n159);
and (n1141,n1045,n61);
and (n1142,n1141,n1143);
xor (n1143,n1112,n1113);
and (n1144,n1138,n1143);
and (n1145,n1045,n70);
and (n1146,n1145,n1147);
xor (n1147,n1148,n1116);
xor (n1148,n1111,n1114);
and (n1149,n1136,n1147);
xor (n1150,n1151,n1120);
xor (n1151,n1109,n1118);
and (n1152,n1153,n1154);
xor (n1153,n1131,n1133);
and (n1154,n1155,n1156);
and (n1155,n1045,n24);
xor (n1156,n1134,n1150);
endmodule
