module top (out,n3,n7,n9,n10,n30,n32,n37,n43,n52
        ,n56,n61,n67,n76,n78,n83,n88,n95,n106,n108
        ,n114,n118,n124,n134,n140,n144,n150,n159,n166,n172
        ,n184,n185,n190,n195,n201,n209,n217,n223,n232,n238
        ,n243,n249,n265,n266,n274,n281,n290,n292,n298,n302
        ,n308,n348,n377,n398,n414,n415,n436,n443,n449,n533
        ,n551,n670,n781,n783,n889,n1064,n1086,n1103,n1266);
output out;
input n3;
input n7;
input n9;
input n10;
input n30;
input n32;
input n37;
input n43;
input n52;
input n56;
input n61;
input n67;
input n76;
input n78;
input n83;
input n88;
input n95;
input n106;
input n108;
input n114;
input n118;
input n124;
input n134;
input n140;
input n144;
input n150;
input n159;
input n166;
input n172;
input n184;
input n185;
input n190;
input n195;
input n201;
input n209;
input n217;
input n223;
input n232;
input n238;
input n243;
input n249;
input n265;
input n266;
input n274;
input n281;
input n290;
input n292;
input n298;
input n302;
input n308;
input n348;
input n377;
input n398;
input n414;
input n415;
input n436;
input n443;
input n449;
input n533;
input n551;
input n670;
input n781;
input n783;
input n889;
input n1064;
input n1086;
input n1103;
input n1266;
wire n0;
wire n1;
wire n2;
wire n4;
wire n5;
wire n6;
wire n8;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n24;
wire n25;
wire n26;
wire n27;
wire n28;
wire n29;
wire n31;
wire n33;
wire n34;
wire n35;
wire n36;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n53;
wire n54;
wire n55;
wire n57;
wire n58;
wire n59;
wire n60;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n77;
wire n79;
wire n80;
wire n81;
wire n82;
wire n84;
wire n85;
wire n86;
wire n87;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n107;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n115;
wire n116;
wire n117;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n141;
wire n142;
wire n143;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n186;
wire n187;
wire n188;
wire n189;
wire n191;
wire n192;
wire n193;
wire n194;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n239;
wire n240;
wire n241;
wire n242;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n291;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n299;
wire n300;
wire n301;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n782;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2988;
wire n2989;
wire n2990;
wire n2991;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2996;
wire n2997;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3003;
wire n3004;
wire n3005;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3010;
wire n3011;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3038;
wire n3039;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
wire n3056;
wire n3057;
wire n3058;
wire n3059;
wire n3060;
wire n3061;
wire n3062;
wire n3063;
wire n3064;
wire n3065;
wire n3066;
wire n3067;
wire n3068;
wire n3069;
wire n3070;
wire n3071;
wire n3072;
wire n3073;
wire n3074;
wire n3075;
wire n3076;
wire n3077;
wire n3078;
wire n3079;
wire n3080;
wire n3081;
wire n3082;
wire n3083;
wire n3084;
wire n3085;
wire n3086;
wire n3087;
wire n3088;
wire n3089;
wire n3090;
wire n3091;
wire n3092;
wire n3093;
wire n3094;
wire n3095;
wire n3096;
wire n3097;
wire n3098;
wire n3099;
wire n3100;
wire n3101;
wire n3102;
wire n3103;
wire n3104;
wire n3105;
wire n3106;
wire n3107;
wire n3108;
wire n3109;
wire n3110;
wire n3111;
wire n3112;
wire n3113;
wire n3114;
wire n3115;
wire n3116;
wire n3117;
wire n3118;
wire n3119;
wire n3120;
wire n3121;
wire n3122;
wire n3123;
wire n3124;
wire n3125;
wire n3126;
wire n3127;
wire n3128;
wire n3129;
wire n3130;
wire n3131;
wire n3132;
wire n3133;
wire n3134;
wire n3135;
wire n3136;
wire n3137;
wire n3138;
wire n3139;
wire n3140;
wire n3141;
wire n3142;
wire n3143;
wire n3144;
wire n3145;
wire n3146;
wire n3147;
wire n3148;
wire n3149;
wire n3150;
wire n3151;
wire n3152;
wire n3153;
wire n3154;
wire n3155;
wire n3156;
wire n3157;
wire n3158;
wire n3159;
wire n3160;
wire n3161;
wire n3162;
wire n3163;
wire n3164;
wire n3165;
wire n3166;
wire n3167;
wire n3168;
wire n3169;
wire n3170;
wire n3171;
wire n3172;
wire n3173;
wire n3174;
wire n3175;
wire n3176;
wire n3177;
wire n3178;
wire n3179;
wire n3180;
wire n3181;
wire n3182;
wire n3183;
wire n3184;
wire n3185;
wire n3186;
wire n3187;
wire n3188;
wire n3189;
wire n3190;
wire n3191;
wire n3192;
wire n3193;
wire n3194;
wire n3195;
wire n3196;
wire n3197;
wire n3198;
wire n3199;
wire n3200;
wire n3201;
wire n3202;
wire n3203;
wire n3204;
wire n3205;
wire n3206;
wire n3207;
wire n3208;
wire n3209;
wire n3210;
wire n3211;
wire n3212;
wire n3213;
wire n3214;
wire n3215;
wire n3216;
wire n3217;
wire n3218;
wire n3219;
wire n3220;
wire n3221;
wire n3222;
wire n3223;
wire n3224;
wire n3225;
wire n3226;
wire n3227;
wire n3228;
wire n3229;
wire n3230;
wire n3231;
wire n3232;
wire n3233;
wire n3234;
wire n3235;
wire n3236;
wire n3237;
wire n3238;
wire n3239;
wire n3240;
wire n3241;
wire n3242;
wire n3243;
wire n3244;
wire n3245;
wire n3246;
wire n3247;
wire n3248;
wire n3249;
wire n3250;
wire n3251;
wire n3252;
wire n3253;
wire n3254;
wire n3255;
wire n3256;
wire n3257;
wire n3258;
wire n3259;
wire n3260;
wire n3261;
wire n3262;
wire n3263;
wire n3264;
wire n3265;
wire n3266;
wire n3267;
wire n3268;
wire n3269;
wire n3270;
wire n3271;
wire n3272;
wire n3273;
wire n3274;
wire n3275;
wire n3276;
wire n3277;
wire n3278;
wire n3279;
wire n3280;
wire n3281;
wire n3282;
wire n3283;
wire n3284;
wire n3285;
wire n3286;
wire n3287;
wire n3288;
wire n3289;
wire n3290;
wire n3291;
wire n3292;
wire n3293;
wire n3294;
wire n3295;
wire n3296;
wire n3297;
wire n3298;
wire n3299;
wire n3300;
wire n3301;
wire n3302;
wire n3303;
wire n3304;
wire n3305;
wire n3306;
wire n3307;
wire n3308;
wire n3309;
wire n3310;
wire n3311;
wire n3312;
wire n3313;
wire n3314;
wire n3315;
wire n3316;
wire n3317;
wire n3318;
wire n3319;
wire n3320;
wire n3321;
wire n3322;
wire n3323;
wire n3324;
wire n3325;
wire n3326;
wire n3327;
wire n3328;
wire n3329;
wire n3330;
wire n3331;
wire n3332;
wire n3333;
wire n3334;
wire n3335;
wire n3336;
wire n3337;
wire n3338;
wire n3339;
wire n3340;
wire n3341;
wire n3342;
wire n3343;
wire n3344;
wire n3345;
wire n3346;
wire n3347;
wire n3348;
wire n3349;
wire n3350;
wire n3351;
wire n3352;
wire n3353;
wire n3354;
wire n3355;
wire n3356;
wire n3357;
wire n3358;
wire n3359;
wire n3360;
wire n3361;
wire n3362;
wire n3363;
wire n3364;
wire n3365;
wire n3366;
wire n3367;
wire n3368;
wire n3369;
wire n3370;
wire n3371;
wire n3372;
wire n3373;
wire n3374;
wire n3375;
wire n3376;
wire n3377;
wire n3378;
wire n3379;
wire n3380;
wire n3381;
wire n3382;
wire n3383;
wire n3384;
wire n3385;
wire n3386;
wire n3387;
wire n3388;
wire n3389;
wire n3390;
wire n3391;
wire n3392;
wire n3393;
wire n3394;
wire n3395;
wire n3396;
wire n3397;
wire n3398;
wire n3399;
wire n3400;
wire n3401;
wire n3402;
wire n3403;
wire n3404;
wire n3405;
wire n3406;
wire n3407;
wire n3408;
wire n3409;
wire n3410;
wire n3411;
wire n3412;
wire n3413;
wire n3414;
wire n3415;
wire n3416;
wire n3417;
wire n3418;
wire n3419;
wire n3420;
wire n3421;
wire n3422;
wire n3423;
wire n3424;
wire n3425;
wire n3426;
wire n3427;
wire n3428;
wire n3429;
wire n3430;
wire n3431;
wire n3432;
wire n3433;
wire n3434;
wire n3435;
wire n3436;
wire n3437;
wire n3438;
wire n3439;
wire n3440;
wire n3441;
wire n3442;
wire n3443;
wire n3444;
wire n3445;
wire n3446;
wire n3447;
wire n3448;
wire n3449;
wire n3450;
wire n3451;
wire n3452;
wire n3453;
wire n3454;
wire n3455;
wire n3456;
wire n3457;
wire n3458;
wire n3459;
wire n3460;
wire n3461;
wire n3462;
wire n3463;
wire n3464;
wire n3465;
wire n3466;
wire n3467;
wire n3468;
wire n3469;
wire n3470;
wire n3471;
wire n3472;
wire n3473;
wire n3474;
wire n3475;
wire n3476;
wire n3477;
wire n3478;
wire n3479;
wire n3480;
wire n3481;
wire n3482;
wire n3483;
wire n3484;
wire n3485;
wire n3486;
wire n3487;
wire n3488;
wire n3489;
wire n3490;
wire n3491;
wire n3492;
wire n3493;
wire n3494;
wire n3495;
wire n3496;
wire n3497;
wire n3498;
wire n3499;
wire n3500;
wire n3501;
wire n3502;
wire n3503;
wire n3504;
wire n3505;
wire n3506;
wire n3507;
wire n3508;
wire n3509;
wire n3510;
wire n3511;
wire n3512;
wire n3513;
wire n3514;
wire n3515;
wire n3516;
wire n3517;
wire n3518;
wire n3519;
wire n3520;
wire n3521;
wire n3522;
wire n3523;
wire n3524;
wire n3525;
wire n3526;
wire n3527;
wire n3528;
wire n3529;
wire n3530;
wire n3531;
wire n3532;
wire n3533;
wire n3534;
wire n3535;
wire n3536;
wire n3537;
wire n3538;
wire n3539;
wire n3540;
wire n3541;
wire n3542;
wire n3543;
wire n3544;
wire n3545;
wire n3546;
wire n3547;
wire n3548;
wire n3549;
wire n3550;
wire n3551;
wire n3552;
wire n3553;
wire n3554;
wire n3555;
wire n3556;
wire n3557;
wire n3558;
wire n3559;
wire n3560;
wire n3561;
wire n3562;
wire n3563;
wire n3564;
wire n3565;
wire n3566;
wire n3567;
wire n3568;
wire n3569;
wire n3570;
wire n3571;
wire n3572;
wire n3573;
wire n3574;
wire n3575;
wire n3576;
wire n3577;
wire n3578;
wire n3579;
wire n3580;
wire n3581;
wire n3582;
wire n3583;
wire n3584;
wire n3585;
wire n3586;
wire n3587;
wire n3588;
wire n3589;
wire n3590;
wire n3591;
wire n3592;
wire n3593;
wire n3594;
wire n3595;
wire n3596;
wire n3597;
wire n3598;
wire n3599;
wire n3600;
wire n3601;
wire n3602;
wire n3603;
wire n3604;
wire n3605;
wire n3606;
wire n3607;
wire n3608;
wire n3609;
wire n3610;
wire n3611;
wire n3612;
wire n3613;
wire n3614;
wire n3615;
wire n3616;
wire n3617;
wire n3618;
wire n3619;
wire n3620;
wire n3621;
wire n3622;
wire n3623;
wire n3624;
wire n3625;
wire n3626;
wire n3627;
wire n3628;
wire n3629;
wire n3630;
wire n3631;
wire n3632;
wire n3633;
wire n3634;
wire n3635;
wire n3636;
wire n3637;
wire n3638;
wire n3639;
wire n3640;
wire n3641;
wire n3642;
wire n3643;
wire n3644;
wire n3645;
wire n3646;
wire n3647;
wire n3648;
wire n3649;
wire n3650;
wire n3651;
wire n3652;
wire n3653;
wire n3654;
wire n3655;
wire n3656;
wire n3657;
wire n3658;
wire n3659;
wire n3660;
wire n3661;
wire n3662;
wire n3663;
wire n3664;
wire n3665;
wire n3666;
wire n3667;
wire n3668;
wire n3669;
wire n3670;
wire n3671;
wire n3672;
wire n3673;
wire n3674;
wire n3675;
wire n3676;
wire n3677;
wire n3678;
wire n3679;
wire n3680;
wire n3681;
wire n3682;
wire n3683;
wire n3684;
wire n3685;
wire n3686;
wire n3687;
wire n3688;
wire n3689;
wire n3690;
wire n3691;
wire n3692;
wire n3693;
wire n3694;
wire n3695;
wire n3696;
wire n3697;
wire n3698;
wire n3699;
wire n3700;
wire n3701;
wire n3702;
wire n3703;
wire n3704;
wire n3705;
wire n3706;
wire n3707;
wire n3708;
wire n3709;
wire n3710;
wire n3711;
wire n3712;
wire n3713;
wire n3714;
wire n3715;
wire n3716;
wire n3717;
wire n3718;
wire n3719;
wire n3720;
wire n3721;
wire n3722;
wire n3723;
wire n3724;
wire n3725;
wire n3726;
wire n3727;
wire n3728;
wire n3729;
wire n3730;
wire n3731;
wire n3732;
wire n3733;
wire n3734;
wire n3735;
wire n3736;
wire n3737;
wire n3738;
wire n3739;
wire n3740;
wire n3741;
wire n3742;
wire n3743;
wire n3744;
wire n3745;
wire n3746;
wire n3747;
wire n3748;
wire n3749;
wire n3750;
wire n3751;
wire n3752;
wire n3753;
wire n3754;
wire n3755;
wire n3756;
wire n3757;
wire n3758;
wire n3759;
wire n3760;
wire n3761;
wire n3762;
wire n3763;
wire n3764;
wire n3765;
wire n3766;
wire n3767;
wire n3768;
wire n3769;
wire n3770;
wire n3771;
wire n3772;
wire n3773;
wire n3774;
wire n3775;
wire n3776;
wire n3777;
wire n3778;
wire n3779;
wire n3780;
wire n3781;
wire n3782;
wire n3783;
wire n3784;
wire n3785;
wire n3786;
wire n3787;
wire n3788;
wire n3789;
wire n3790;
wire n3791;
wire n3792;
wire n3793;
wire n3794;
wire n3795;
wire n3796;
wire n3797;
wire n3798;
wire n3799;
wire n3800;
wire n3801;
wire n3802;
wire n3803;
wire n3804;
wire n3805;
wire n3806;
wire n3807;
wire n3808;
wire n3809;
wire n3810;
wire n3811;
wire n3812;
wire n3813;
wire n3814;
wire n3815;
wire n3816;
wire n3817;
wire n3818;
wire n3819;
wire n3820;
wire n3821;
wire n3822;
wire n3823;
wire n3824;
wire n3825;
wire n3826;
wire n3827;
wire n3828;
wire n3829;
wire n3830;
wire n3831;
wire n3832;
wire n3833;
wire n3834;
wire n3835;
wire n3836;
wire n3837;
wire n3838;
wire n3839;
wire n3840;
wire n3841;
wire n3842;
wire n3843;
wire n3844;
wire n3845;
wire n3846;
wire n3847;
wire n3848;
wire n3849;
wire n3850;
wire n3851;
wire n3852;
wire n3853;
wire n3854;
wire n3855;
wire n3856;
wire n3857;
wire n3858;
wire n3859;
wire n3860;
wire n3861;
wire n3862;
wire n3863;
wire n3864;
wire n3865;
wire n3866;
wire n3867;
wire n3868;
wire n3869;
wire n3870;
wire n3871;
wire n3872;
wire n3873;
wire n3874;
wire n3875;
wire n3876;
wire n3877;
wire n3878;
wire n3879;
wire n3880;
wire n3881;
wire n3882;
wire n3883;
wire n3884;
wire n3885;
wire n3886;
wire n3887;
wire n3888;
wire n3889;
wire n3890;
wire n3891;
wire n3892;
wire n3893;
wire n3894;
wire n3895;
wire n3896;
wire n3897;
wire n3898;
wire n3899;
wire n3900;
wire n3901;
wire n3902;
wire n3903;
wire n3904;
wire n3905;
wire n3906;
wire n3907;
wire n3908;
wire n3909;
wire n3910;
wire n3911;
wire n3912;
wire n3913;
wire n3914;
wire n3915;
wire n3916;
wire n3917;
wire n3918;
wire n3919;
wire n3920;
wire n3921;
wire n3922;
wire n3923;
wire n3924;
wire n3925;
wire n3926;
wire n3927;
wire n3928;
wire n3929;
wire n3930;
wire n3931;
wire n3932;
wire n3933;
wire n3934;
wire n3935;
wire n3936;
wire n3937;
wire n3938;
wire n3939;
wire n3940;
wire n3941;
wire n3942;
wire n3943;
wire n3944;
wire n3945;
wire n3946;
wire n3947;
wire n3948;
wire n3949;
wire n3950;
wire n3951;
wire n3952;
wire n3953;
wire n3954;
wire n3955;
wire n3956;
wire n3957;
wire n3958;
wire n3959;
wire n3960;
wire n3961;
wire n3962;
wire n3963;
wire n3964;
wire n3965;
wire n3966;
wire n3967;
wire n3968;
wire n3969;
wire n3970;
wire n3971;
wire n3972;
wire n3973;
wire n3974;
wire n3975;
wire n3976;
wire n3977;
wire n3978;
wire n3979;
wire n3980;
wire n3981;
wire n3982;
wire n3983;
wire n3984;
wire n3985;
wire n3986;
wire n3987;
wire n3988;
wire n3989;
wire n3990;
wire n3991;
wire n3992;
wire n3993;
wire n3994;
wire n3995;
wire n3996;
wire n3997;
wire n3998;
wire n3999;
wire n4000;
wire n4001;
wire n4002;
wire n4003;
wire n4004;
wire n4005;
wire n4006;
wire n4007;
wire n4008;
wire n4009;
wire n4010;
wire n4011;
wire n4012;
wire n4013;
wire n4014;
wire n4015;
wire n4016;
wire n4017;
wire n4018;
wire n4019;
wire n4020;
wire n4021;
wire n4022;
wire n4023;
wire n4024;
wire n4025;
wire n4026;
wire n4027;
wire n4028;
wire n4029;
wire n4030;
wire n4031;
wire n4032;
wire n4033;
wire n4034;
wire n4035;
wire n4036;
wire n4037;
wire n4038;
wire n4039;
wire n4040;
wire n4041;
wire n4042;
wire n4043;
wire n4044;
wire n4045;
wire n4046;
wire n4047;
wire n4048;
wire n4049;
wire n4050;
wire n4051;
wire n4052;
wire n4053;
wire n4054;
wire n4055;
wire n4056;
wire n4057;
wire n4058;
wire n4059;
wire n4060;
wire n4061;
wire n4062;
wire n4063;
wire n4064;
wire n4065;
wire n4066;
wire n4067;
wire n4068;
wire n4069;
wire n4070;
wire n4071;
wire n4072;
wire n4073;
wire n4074;
wire n4075;
wire n4076;
wire n4077;
wire n4078;
wire n4079;
wire n4080;
wire n4081;
wire n4082;
wire n4083;
wire n4084;
wire n4085;
wire n4086;
wire n4087;
wire n4088;
wire n4089;
wire n4090;
wire n4091;
wire n4092;
wire n4093;
wire n4094;
wire n4095;
wire n4096;
wire n4097;
wire n4098;
wire n4099;
wire n4100;
wire n4101;
wire n4102;
wire n4103;
wire n4104;
wire n4105;
wire n4106;
wire n4107;
wire n4108;
wire n4109;
wire n4110;
wire n4111;
wire n4112;
wire n4113;
wire n4114;
wire n4115;
wire n4116;
wire n4117;
wire n4118;
wire n4119;
wire n4120;
wire n4121;
wire n4122;
wire n4123;
wire n4124;
wire n4125;
wire n4126;
wire n4127;
wire n4128;
wire n4129;
wire n4130;
wire n4131;
wire n4132;
wire n4133;
wire n4134;
wire n4135;
wire n4136;
wire n4137;
wire n4138;
wire n4139;
wire n4140;
wire n4141;
wire n4142;
wire n4143;
wire n4144;
wire n4145;
wire n4146;
wire n4147;
wire n4148;
wire n4149;
wire n4150;
wire n4151;
wire n4152;
wire n4153;
wire n4154;
wire n4155;
wire n4156;
wire n4157;
wire n4158;
wire n4159;
wire n4160;
wire n4161;
wire n4162;
wire n4163;
wire n4164;
wire n4165;
wire n4166;
wire n4167;
wire n4168;
wire n4169;
wire n4170;
wire n4171;
wire n4172;
wire n4173;
wire n4174;
wire n4175;
wire n4176;
wire n4177;
wire n4178;
wire n4179;
wire n4180;
wire n4181;
wire n4182;
wire n4183;
wire n4184;
wire n4185;
wire n4186;
wire n4187;
wire n4188;
wire n4189;
wire n4190;
wire n4191;
wire n4192;
wire n4193;
wire n4194;
wire n4195;
wire n4196;
wire n4197;
wire n4198;
wire n4199;
wire n4200;
wire n4201;
wire n4202;
wire n4203;
wire n4204;
wire n4205;
wire n4206;
wire n4207;
wire n4208;
wire n4209;
wire n4210;
wire n4211;
wire n4212;
wire n4213;
wire n4214;
wire n4215;
wire n4216;
wire n4217;
wire n4218;
wire n4219;
wire n4220;
wire n4221;
wire n4222;
wire n4223;
wire n4224;
wire n4225;
wire n4226;
wire n4227;
wire n4228;
wire n4229;
wire n4230;
wire n4231;
wire n4232;
wire n4233;
wire n4234;
wire n4235;
wire n4236;
wire n4237;
wire n4238;
wire n4239;
wire n4240;
wire n4241;
wire n4242;
wire n4243;
wire n4244;
wire n4245;
wire n4246;
wire n4247;
wire n4248;
wire n4249;
wire n4250;
wire n4251;
wire n4252;
wire n4253;
wire n4254;
wire n4255;
wire n4256;
wire n4257;
wire n4258;
wire n4259;
wire n4260;
wire n4261;
wire n4262;
wire n4263;
wire n4264;
wire n4265;
wire n4266;
wire n4267;
wire n4268;
wire n4269;
wire n4270;
wire n4271;
wire n4272;
wire n4273;
wire n4274;
wire n4275;
wire n4276;
wire n4277;
wire n4278;
wire n4279;
wire n4280;
wire n4281;
wire n4282;
wire n4283;
wire n4284;
wire n4285;
wire n4286;
wire n4287;
wire n4288;
wire n4289;
wire n4290;
wire n4291;
wire n4292;
wire n4293;
wire n4294;
wire n4295;
wire n4296;
wire n4297;
wire n4298;
wire n4299;
wire n4300;
wire n4301;
wire n4302;
wire n4303;
wire n4304;
wire n4305;
wire n4306;
wire n4307;
wire n4308;
wire n4309;
wire n4310;
wire n4311;
wire n4312;
wire n4313;
wire n4314;
wire n4315;
wire n4316;
wire n4317;
wire n4318;
wire n4319;
wire n4320;
wire n4321;
wire n4322;
wire n4323;
wire n4324;
wire n4325;
wire n4326;
wire n4327;
wire n4328;
wire n4329;
wire n4330;
wire n4331;
wire n4332;
wire n4333;
wire n4334;
wire n4335;
wire n4336;
wire n4337;
wire n4338;
wire n4339;
wire n4340;
wire n4341;
wire n4342;
wire n4343;
wire n4344;
wire n4345;
wire n4346;
wire n4347;
wire n4348;
wire n4349;
wire n4350;
wire n4351;
wire n4352;
wire n4353;
wire n4354;
wire n4355;
wire n4356;
wire n4357;
wire n4358;
wire n4359;
wire n4360;
wire n4361;
wire n4362;
wire n4363;
wire n4364;
wire n4365;
wire n4366;
wire n4367;
wire n4368;
wire n4369;
wire n4370;
wire n4371;
wire n4372;
wire n4373;
wire n4374;
wire n4375;
wire n4376;
wire n4377;
wire n4378;
wire n4379;
wire n4380;
wire n4381;
wire n4382;
wire n4383;
wire n4384;
wire n4385;
wire n4386;
wire n4387;
wire n4388;
wire n4389;
wire n4390;
wire n4391;
wire n4392;
wire n4393;
wire n4394;
wire n4395;
wire n4396;
wire n4397;
wire n4398;
wire n4399;
wire n4400;
wire n4401;
wire n4402;
wire n4403;
wire n4404;
wire n4405;
wire n4406;
wire n4407;
wire n4408;
wire n4409;
wire n4410;
wire n4411;
wire n4412;
wire n4413;
wire n4414;
wire n4415;
wire n4416;
wire n4417;
wire n4418;
wire n4419;
wire n4420;
wire n4421;
wire n4422;
wire n4423;
wire n4424;
wire n4425;
wire n4426;
wire n4427;
wire n4428;
wire n4429;
wire n4430;
wire n4431;
wire n4432;
wire n4433;
wire n4434;
wire n4435;
wire n4436;
wire n4437;
wire n4438;
wire n4439;
wire n4440;
wire n4441;
wire n4442;
wire n4443;
wire n4444;
wire n4445;
wire n4446;
wire n4447;
wire n4448;
wire n4449;
wire n4450;
wire n4451;
wire n4452;
wire n4453;
wire n4454;
wire n4455;
wire n4456;
wire n4457;
wire n4458;
wire n4459;
wire n4460;
wire n4461;
wire n4462;
wire n4463;
wire n4464;
wire n4465;
wire n4466;
wire n4467;
wire n4468;
wire n4469;
wire n4470;
wire n4471;
wire n4472;
wire n4473;
wire n4474;
wire n4475;
wire n4476;
wire n4477;
wire n4478;
wire n4479;
wire n4480;
wire n4481;
wire n4482;
wire n4483;
wire n4484;
wire n4485;
wire n4486;
wire n4487;
wire n4488;
wire n4489;
wire n4490;
wire n4491;
wire n4492;
wire n4493;
wire n4494;
wire n4495;
wire n4496;
wire n4497;
wire n4498;
wire n4499;
wire n4500;
wire n4501;
wire n4502;
wire n4503;
wire n4504;
wire n4505;
wire n4506;
wire n4507;
wire n4508;
wire n4509;
wire n4510;
wire n4511;
wire n4512;
wire n4513;
wire n4514;
wire n4515;
wire n4516;
wire n4517;
wire n4518;
wire n4519;
wire n4520;
wire n4521;
wire n4522;
wire n4523;
wire n4524;
wire n4525;
wire n4526;
wire n4527;
wire n4528;
wire n4529;
wire n4530;
wire n4531;
wire n4532;
wire n4533;
wire n4534;
wire n4535;
wire n4536;
wire n4537;
wire n4538;
wire n4539;
wire n4540;
wire n4541;
wire n4542;
wire n4543;
wire n4544;
wire n4545;
wire n4546;
wire n4547;
wire n4548;
wire n4549;
wire n4550;
wire n4551;
wire n4552;
wire n4553;
wire n4554;
wire n4555;
wire n4556;
wire n4557;
wire n4558;
wire n4559;
wire n4560;
wire n4561;
wire n4562;
wire n4563;
wire n4564;
wire n4565;
wire n4566;
wire n4567;
wire n4568;
wire n4569;
wire n4570;
wire n4571;
wire n4572;
wire n4573;
wire n4574;
wire n4575;
wire n4576;
wire n4577;
wire n4578;
wire n4579;
wire n4580;
wire n4581;
wire n4582;
wire n4583;
wire n4584;
wire n4585;
wire n4586;
wire n4587;
wire n4588;
wire n4589;
wire n4590;
wire n4591;
wire n4592;
wire n4593;
wire n4594;
wire n4595;
wire n4596;
wire n4597;
wire n4598;
wire n4599;
wire n4600;
wire n4601;
wire n4602;
wire n4603;
wire n4604;
wire n4605;
wire n4606;
wire n4607;
wire n4608;
wire n4609;
wire n4610;
wire n4611;
wire n4612;
wire n4613;
wire n4614;
wire n4615;
wire n4616;
wire n4617;
wire n4618;
wire n4619;
wire n4620;
wire n4621;
wire n4622;
wire n4623;
wire n4624;
wire n4625;
wire n4626;
wire n4627;
wire n4628;
wire n4629;
wire n4630;
wire n4631;
wire n4632;
wire n4633;
wire n4634;
wire n4635;
wire n4636;
wire n4637;
wire n4638;
wire n4639;
wire n4640;
wire n4641;
wire n4642;
wire n4643;
wire n4644;
wire n4645;
wire n4646;
wire n4647;
wire n4648;
wire n4649;
wire n4650;
wire n4651;
wire n4652;
wire n4653;
wire n4654;
wire n4655;
wire n4656;
wire n4657;
wire n4658;
wire n4659;
wire n4660;
wire n4661;
wire n4662;
wire n4663;
wire n4664;
wire n4665;
wire n4666;
wire n4667;
wire n4668;
wire n4669;
wire n4670;
wire n4671;
wire n4672;
wire n4673;
wire n4674;
wire n4675;
wire n4676;
wire n4677;
wire n4678;
wire n4679;
wire n4680;
wire n4681;
wire n4682;
wire n4683;
wire n4684;
wire n4685;
wire n4686;
wire n4687;
wire n4688;
wire n4689;
wire n4690;
wire n4691;
wire n4692;
wire n4693;
wire n4694;
wire n4695;
wire n4696;
wire n4697;
wire n4698;
wire n4699;
wire n4700;
wire n4701;
wire n4702;
wire n4703;
wire n4704;
wire n4705;
wire n4706;
wire n4707;
wire n4708;
wire n4709;
wire n4710;
wire n4711;
wire n4712;
wire n4713;
wire n4714;
wire n4715;
wire n4716;
wire n4717;
wire n4718;
wire n4719;
wire n4720;
wire n4721;
wire n4722;
wire n4723;
wire n4724;
wire n4725;
wire n4726;
wire n4727;
wire n4728;
wire n4729;
wire n4730;
wire n4731;
wire n4732;
wire n4733;
wire n4734;
wire n4735;
wire n4736;
wire n4737;
wire n4738;
wire n4739;
wire n4740;
wire n4741;
wire n4742;
wire n4743;
wire n4744;
wire n4745;
wire n4746;
wire n4747;
wire n4748;
wire n4749;
wire n4750;
wire n4751;
wire n4752;
wire n4753;
wire n4754;
wire n4755;
wire n4756;
wire n4757;
wire n4758;
wire n4759;
wire n4760;
wire n4761;
wire n4762;
wire n4763;
wire n4764;
wire n4765;
wire n4766;
wire n4767;
wire n4768;
wire n4769;
wire n4770;
wire n4771;
wire n4772;
wire n4773;
wire n4774;
wire n4775;
wire n4776;
wire n4777;
wire n4778;
wire n4779;
wire n4780;
wire n4781;
wire n4782;
wire n4783;
wire n4784;
wire n4785;
wire n4786;
wire n4787;
wire n4788;
wire n4789;
wire n4790;
wire n4791;
wire n4792;
wire n4793;
wire n4794;
wire n4795;
wire n4796;
wire n4797;
wire n4798;
wire n4799;
wire n4800;
wire n4801;
wire n4802;
wire n4803;
wire n4804;
wire n4805;
wire n4806;
wire n4807;
wire n4808;
wire n4809;
wire n4810;
wire n4811;
wire n4812;
wire n4813;
wire n4814;
wire n4815;
wire n4816;
wire n4817;
wire n4818;
wire n4819;
wire n4820;
wire n4821;
wire n4822;
wire n4823;
wire n4824;
wire n4825;
wire n4826;
wire n4827;
wire n4828;
wire n4829;
wire n4830;
wire n4831;
wire n4832;
wire n4833;
wire n4834;
wire n4835;
wire n4836;
wire n4837;
wire n4838;
wire n4839;
wire n4840;
wire n4841;
wire n4842;
wire n4843;
wire n4844;
wire n4845;
wire n4846;
wire n4847;
wire n4848;
wire n4849;
wire n4850;
wire n4851;
wire n4852;
wire n4853;
wire n4854;
wire n4855;
wire n4856;
wire n4857;
wire n4858;
wire n4859;
wire n4860;
wire n4861;
wire n4862;
wire n4863;
wire n4864;
wire n4865;
wire n4866;
wire n4867;
wire n4868;
wire n4869;
wire n4870;
wire n4871;
wire n4872;
wire n4873;
wire n4874;
wire n4875;
wire n4876;
wire n4877;
wire n4878;
wire n4879;
wire n4880;
wire n4881;
wire n4882;
wire n4883;
wire n4884;
wire n4885;
wire n4886;
wire n4887;
wire n4888;
wire n4889;
wire n4890;
wire n4891;
wire n4892;
wire n4893;
wire n4894;
wire n4895;
wire n4896;
wire n4897;
wire n4898;
wire n4899;
wire n4900;
wire n4901;
wire n4902;
wire n4903;
wire n4904;
wire n4905;
wire n4906;
wire n4907;
wire n4908;
wire n4909;
wire n4910;
wire n4911;
wire n4912;
wire n4913;
wire n4914;
wire n4915;
wire n4916;
wire n4917;
wire n4918;
wire n4919;
wire n4920;
wire n4921;
wire n4922;
wire n4923;
wire n4924;
wire n4925;
wire n4926;
wire n4927;
wire n4928;
wire n4929;
wire n4930;
wire n4931;
wire n4932;
wire n4933;
wire n4934;
wire n4935;
wire n4936;
wire n4937;
wire n4938;
wire n4939;
wire n4940;
wire n4941;
wire n4942;
wire n4943;
wire n4944;
wire n4945;
wire n4946;
wire n4947;
wire n4948;
wire n4949;
wire n4950;
wire n4951;
wire n4952;
wire n4953;
wire n4954;
wire n4955;
wire n4956;
wire n4957;
wire n4958;
wire n4959;
wire n4960;
wire n4961;
wire n4962;
wire n4963;
wire n4964;
wire n4965;
wire n4966;
wire n4967;
wire n4968;
wire n4969;
wire n4970;
wire n4971;
wire n4972;
wire n4973;
wire n4974;
wire n4975;
wire n4976;
wire n4977;
wire n4978;
wire n4979;
wire n4980;
wire n4981;
wire n4982;
wire n4983;
wire n4984;
wire n4985;
wire n4986;
wire n4987;
wire n4988;
wire n4989;
wire n4990;
wire n4991;
wire n4992;
wire n4993;
wire n4994;
wire n4995;
wire n4996;
wire n4997;
wire n4998;
wire n4999;
wire n5000;
wire n5001;
wire n5002;
wire n5003;
wire n5004;
wire n5005;
wire n5006;
wire n5007;
wire n5008;
wire n5009;
wire n5010;
wire n5011;
wire n5012;
wire n5013;
wire n5014;
wire n5015;
wire n5016;
wire n5017;
wire n5018;
wire n5019;
wire n5020;
wire n5021;
wire n5022;
wire n5023;
wire n5024;
wire n5025;
wire n5026;
wire n5027;
wire n5028;
wire n5029;
wire n5030;
wire n5031;
wire n5032;
wire n5033;
wire n5034;
wire n5035;
wire n5036;
wire n5037;
wire n5038;
wire n5039;
wire n5040;
wire n5041;
wire n5042;
wire n5043;
wire n5044;
wire n5045;
wire n5046;
wire n5047;
wire n5048;
wire n5049;
wire n5050;
wire n5051;
wire n5052;
wire n5053;
wire n5054;
wire n5055;
wire n5056;
wire n5057;
wire n5058;
wire n5059;
wire n5060;
wire n5061;
wire n5062;
wire n5063;
wire n5064;
wire n5065;
wire n5066;
wire n5067;
wire n5068;
wire n5069;
wire n5070;
wire n5071;
wire n5072;
wire n5073;
wire n5074;
wire n5075;
wire n5076;
wire n5077;
wire n5078;
wire n5079;
wire n5080;
wire n5081;
wire n5082;
wire n5083;
wire n5084;
wire n5085;
wire n5086;
wire n5087;
wire n5088;
wire n5089;
wire n5090;
wire n5091;
wire n5092;
wire n5093;
wire n5094;
wire n5095;
wire n5096;
wire n5097;
wire n5098;
wire n5099;
wire n5100;
wire n5101;
wire n5102;
wire n5103;
wire n5104;
wire n5105;
wire n5106;
wire n5107;
wire n5108;
wire n5109;
wire n5110;
wire n5111;
wire n5112;
wire n5113;
wire n5114;
wire n5115;
wire n5116;
wire n5117;
wire n5118;
wire n5119;
wire n5120;
wire n5121;
wire n5122;
wire n5123;
wire n5124;
wire n5125;
wire n5126;
wire n5127;
wire n5128;
wire n5129;
wire n5130;
wire n5131;
wire n5132;
wire n5133;
wire n5134;
wire n5135;
wire n5136;
wire n5137;
wire n5138;
wire n5139;
wire n5140;
wire n5141;
wire n5142;
wire n5143;
wire n5144;
wire n5145;
wire n5146;
wire n5147;
wire n5148;
wire n5149;
wire n5150;
wire n5151;
wire n5152;
wire n5153;
wire n5154;
wire n5155;
wire n5156;
wire n5157;
wire n5158;
wire n5159;
wire n5160;
wire n5161;
wire n5162;
wire n5163;
wire n5164;
wire n5165;
wire n5166;
wire n5167;
wire n5168;
wire n5169;
wire n5170;
wire n5171;
wire n5172;
wire n5173;
wire n5174;
wire n5175;
wire n5176;
wire n5177;
wire n5178;
wire n5179;
wire n5180;
wire n5181;
wire n5182;
wire n5183;
wire n5184;
wire n5185;
wire n5186;
wire n5187;
wire n5188;
wire n5189;
wire n5190;
wire n5191;
wire n5192;
wire n5193;
wire n5194;
wire n5195;
wire n5196;
wire n5197;
wire n5198;
wire n5199;
wire n5200;
wire n5201;
wire n5202;
wire n5203;
wire n5204;
wire n5205;
wire n5206;
wire n5207;
wire n5208;
wire n5209;
wire n5210;
wire n5211;
wire n5212;
wire n5213;
wire n5214;
wire n5215;
wire n5216;
wire n5217;
wire n5218;
wire n5219;
wire n5220;
wire n5221;
wire n5222;
wire n5223;
wire n5224;
wire n5225;
wire n5226;
wire n5227;
wire n5228;
wire n5229;
wire n5230;
wire n5231;
wire n5232;
wire n5233;
wire n5234;
wire n5235;
wire n5236;
wire n5237;
wire n5238;
wire n5239;
wire n5240;
wire n5241;
wire n5242;
wire n5243;
wire n5244;
wire n5245;
wire n5246;
wire n5247;
wire n5248;
wire n5249;
wire n5250;
wire n5251;
wire n5252;
wire n5253;
wire n5254;
wire n5255;
wire n5256;
wire n5257;
wire n5258;
wire n5259;
wire n5260;
wire n5261;
wire n5262;
wire n5263;
wire n5264;
wire n5265;
wire n5266;
wire n5267;
wire n5268;
wire n5269;
wire n5270;
wire n5271;
wire n5272;
wire n5273;
wire n5274;
wire n5275;
wire n5276;
wire n5277;
wire n5278;
wire n5279;
wire n5280;
wire n5281;
wire n5282;
wire n5283;
wire n5284;
wire n5285;
wire n5286;
wire n5287;
wire n5288;
wire n5289;
wire n5290;
wire n5291;
wire n5292;
wire n5293;
wire n5294;
wire n5295;
wire n5296;
wire n5297;
wire n5298;
wire n5299;
wire n5300;
wire n5301;
wire n5302;
wire n5303;
wire n5304;
wire n5305;
wire n5306;
wire n5307;
wire n5308;
wire n5309;
wire n5310;
wire n5311;
wire n5312;
wire n5313;
wire n5314;
wire n5315;
wire n5316;
wire n5317;
wire n5318;
wire n5319;
wire n5320;
wire n5321;
wire n5322;
wire n5323;
wire n5324;
wire n5325;
wire n5326;
wire n5327;
wire n5328;
wire n5329;
wire n5330;
wire n5331;
wire n5332;
wire n5333;
wire n5334;
wire n5335;
wire n5336;
wire n5337;
wire n5338;
wire n5339;
wire n5340;
wire n5341;
wire n5342;
wire n5343;
wire n5344;
wire n5345;
wire n5346;
wire n5347;
wire n5348;
wire n5349;
wire n5350;
wire n5351;
wire n5352;
wire n5353;
wire n5354;
wire n5355;
wire n5356;
wire n5357;
wire n5358;
wire n5359;
wire n5360;
wire n5361;
wire n5362;
wire n5363;
wire n5364;
wire n5365;
wire n5366;
wire n5367;
wire n5368;
wire n5369;
wire n5370;
wire n5371;
wire n5372;
wire n5373;
wire n5374;
wire n5375;
wire n5376;
wire n5377;
wire n5378;
wire n5379;
wire n5380;
wire n5381;
wire n5382;
wire n5383;
wire n5384;
wire n5385;
wire n5386;
wire n5387;
wire n5388;
wire n5389;
wire n5390;
wire n5391;
wire n5392;
wire n5393;
wire n5394;
wire n5395;
wire n5396;
wire n5397;
wire n5398;
wire n5399;
wire n5400;
wire n5401;
wire n5402;
wire n5403;
wire n5404;
wire n5405;
wire n5406;
wire n5407;
wire n5408;
wire n5409;
wire n5410;
wire n5411;
wire n5412;
wire n5413;
wire n5414;
wire n5415;
wire n5416;
wire n5417;
wire n5418;
wire n5419;
wire n5420;
wire n5421;
wire n5422;
wire n5423;
wire n5424;
wire n5425;
wire n5426;
wire n5427;
wire n5428;
wire n5429;
wire n5430;
wire n5431;
wire n5432;
wire n5433;
wire n5434;
wire n5435;
wire n5436;
wire n5437;
wire n5438;
wire n5439;
wire n5440;
wire n5441;
wire n5442;
wire n5443;
wire n5444;
wire n5445;
wire n5446;
wire n5447;
wire n5448;
wire n5449;
wire n5450;
wire n5451;
wire n5452;
wire n5453;
wire n5454;
wire n5455;
wire n5456;
wire n5457;
wire n5458;
wire n5459;
wire n5460;
wire n5461;
wire n5462;
wire n5463;
wire n5464;
wire n5465;
wire n5466;
wire n5467;
wire n5468;
wire n5469;
wire n5470;
wire n5471;
wire n5472;
wire n5473;
wire n5474;
wire n5475;
wire n5476;
wire n5477;
wire n5478;
wire n5479;
wire n5480;
wire n5481;
wire n5482;
wire n5483;
wire n5484;
wire n5485;
wire n5486;
wire n5487;
wire n5488;
wire n5489;
wire n5490;
wire n5491;
wire n5492;
wire n5493;
wire n5494;
wire n5495;
wire n5496;
wire n5497;
wire n5498;
wire n5499;
wire n5500;
wire n5501;
wire n5502;
wire n5503;
wire n5504;
wire n5505;
wire n5506;
wire n5507;
wire n5508;
wire n5509;
wire n5510;
wire n5511;
wire n5512;
wire n5513;
wire n5514;
wire n5515;
wire n5516;
wire n5517;
wire n5518;
wire n5519;
wire n5520;
wire n5521;
wire n5522;
wire n5523;
wire n5524;
wire n5525;
wire n5526;
wire n5527;
wire n5528;
wire n5529;
wire n5530;
wire n5531;
wire n5532;
wire n5533;
wire n5534;
wire n5535;
wire n5536;
wire n5537;
wire n5538;
wire n5539;
wire n5540;
wire n5541;
wire n5542;
wire n5543;
wire n5544;
wire n5545;
wire n5546;
wire n5547;
wire n5548;
wire n5549;
wire n5550;
wire n5551;
wire n5552;
wire n5553;
wire n5554;
wire n5555;
wire n5556;
wire n5557;
wire n5558;
wire n5559;
wire n5560;
wire n5561;
wire n5562;
wire n5563;
wire n5564;
wire n5565;
wire n5566;
wire n5567;
wire n5568;
wire n5569;
wire n5570;
wire n5571;
wire n5572;
wire n5573;
wire n5574;
wire n5575;
wire n5576;
wire n5577;
wire n5578;
wire n5579;
wire n5580;
wire n5581;
wire n5582;
wire n5583;
wire n5584;
wire n5585;
wire n5586;
wire n5587;
wire n5588;
wire n5589;
wire n5590;
wire n5591;
wire n5592;
wire n5593;
wire n5594;
wire n5595;
wire n5596;
wire n5597;
wire n5598;
wire n5599;
wire n5600;
wire n5601;
wire n5602;
wire n5603;
wire n5604;
wire n5605;
wire n5606;
wire n5607;
wire n5608;
wire n5609;
wire n5610;
wire n5611;
wire n5612;
wire n5613;
wire n5614;
wire n5615;
wire n5616;
wire n5617;
wire n5618;
wire n5619;
wire n5620;
wire n5621;
wire n5622;
wire n5623;
wire n5624;
wire n5625;
wire n5626;
wire n5627;
wire n5628;
wire n5629;
wire n5630;
wire n5631;
wire n5632;
wire n5633;
wire n5634;
wire n5635;
wire n5636;
wire n5637;
wire n5638;
wire n5639;
wire n5640;
wire n5641;
wire n5642;
wire n5643;
wire n5644;
wire n5645;
wire n5646;
wire n5647;
wire n5648;
wire n5649;
wire n5650;
wire n5651;
wire n5652;
wire n5653;
wire n5654;
wire n5655;
wire n5656;
wire n5657;
wire n5658;
wire n5659;
wire n5660;
wire n5661;
wire n5662;
wire n5663;
wire n5664;
wire n5665;
wire n5666;
wire n5667;
wire n5668;
wire n5669;
wire n5670;
wire n5671;
wire n5672;
wire n5673;
wire n5674;
wire n5675;
wire n5676;
wire n5677;
wire n5678;
wire n5679;
wire n5680;
wire n5681;
wire n5682;
wire n5683;
wire n5684;
wire n5685;
wire n5686;
wire n5687;
wire n5688;
wire n5689;
wire n5690;
wire n5691;
wire n5692;
wire n5693;
wire n5694;
wire n5695;
wire n5696;
wire n5697;
wire n5698;
wire n5699;
wire n5700;
wire n5701;
wire n5702;
wire n5703;
wire n5704;
wire n5705;
wire n5706;
wire n5707;
wire n5708;
wire n5709;
wire n5710;
wire n5711;
wire n5712;
wire n5713;
wire n5714;
wire n5715;
wire n5716;
wire n5717;
wire n5718;
wire n5719;
wire n5720;
wire n5721;
wire n5722;
wire n5723;
wire n5724;
wire n5725;
wire n5726;
wire n5727;
wire n5728;
wire n5729;
wire n5730;
wire n5731;
wire n5732;
wire n5733;
wire n5734;
wire n5735;
wire n5736;
wire n5737;
wire n5738;
wire n5739;
wire n5740;
wire n5741;
wire n5742;
wire n5743;
wire n5744;
wire n5745;
wire n5746;
wire n5747;
wire n5748;
wire n5749;
wire n5750;
wire n5751;
wire n5752;
wire n5753;
wire n5754;
wire n5755;
wire n5756;
wire n5757;
wire n5758;
wire n5759;
wire n5760;
wire n5761;
wire n5762;
wire n5763;
wire n5764;
wire n5765;
wire n5766;
wire n5767;
wire n5768;
wire n5769;
wire n5770;
wire n5771;
wire n5772;
wire n5773;
wire n5774;
wire n5775;
wire n5776;
wire n5777;
wire n5778;
wire n5779;
wire n5780;
wire n5781;
wire n5782;
wire n5783;
wire n5784;
wire n5785;
wire n5786;
wire n5787;
wire n5788;
wire n5789;
wire n5790;
wire n5791;
wire n5792;
wire n5793;
wire n5794;
wire n5795;
wire n5796;
wire n5797;
wire n5798;
wire n5799;
wire n5800;
wire n5801;
wire n5802;
wire n5803;
wire n5804;
wire n5805;
wire n5806;
wire n5807;
wire n5808;
wire n5809;
wire n5810;
wire n5811;
wire n5812;
wire n5813;
wire n5814;
wire n5815;
wire n5816;
wire n5817;
wire n5818;
wire n5819;
wire n5820;
wire n5821;
wire n5822;
wire n5823;
wire n5824;
wire n5825;
wire n5826;
wire n5827;
wire n5828;
wire n5829;
wire n5830;
wire n5831;
wire n5832;
wire n5833;
wire n5834;
wire n5835;
wire n5836;
wire n5837;
wire n5838;
wire n5839;
wire n5840;
wire n5841;
wire n5842;
wire n5843;
wire n5844;
wire n5845;
wire n5846;
wire n5847;
wire n5848;
wire n5849;
wire n5850;
wire n5851;
wire n5852;
wire n5853;
wire n5854;
wire n5855;
wire n5856;
wire n5857;
wire n5858;
wire n5859;
wire n5860;
wire n5861;
wire n5862;
wire n5863;
wire n5864;
wire n5865;
wire n5866;
wire n5867;
wire n5868;
wire n5869;
wire n5870;
wire n5871;
wire n5872;
wire n5873;
wire n5874;
wire n5875;
wire n5876;
wire n5877;
wire n5878;
wire n5879;
wire n5880;
wire n5881;
wire n5882;
wire n5883;
wire n5884;
wire n5885;
wire n5886;
wire n5887;
wire n5888;
wire n5889;
wire n5890;
wire n5891;
wire n5892;
wire n5893;
wire n5894;
wire n5895;
wire n5896;
wire n5897;
wire n5898;
wire n5899;
wire n5900;
wire n5901;
wire n5902;
wire n5903;
wire n5904;
wire n5905;
wire n5906;
wire n5907;
wire n5908;
wire n5909;
wire n5910;
wire n5911;
wire n5912;
wire n5913;
wire n5914;
wire n5915;
wire n5916;
wire n5917;
wire n5918;
wire n5919;
wire n5920;
wire n5921;
wire n5922;
wire n5923;
wire n5924;
wire n5925;
wire n5926;
wire n5927;
wire n5928;
wire n5929;
wire n5930;
wire n5931;
wire n5932;
wire n5933;
wire n5934;
wire n5935;
wire n5936;
wire n5937;
wire n5938;
wire n5939;
wire n5940;
wire n5941;
wire n5942;
wire n5943;
wire n5944;
wire n5945;
wire n5946;
wire n5947;
wire n5948;
wire n5949;
wire n5950;
wire n5951;
wire n5952;
wire n5953;
wire n5954;
wire n5955;
wire n5956;
wire n5957;
wire n5958;
wire n5959;
wire n5960;
wire n5961;
wire n5962;
wire n5963;
wire n5964;
wire n5965;
wire n5966;
wire n5967;
wire n5968;
wire n5969;
wire n5970;
wire n5971;
wire n5972;
wire n5973;
wire n5974;
wire n5975;
wire n5976;
wire n5977;
wire n5978;
wire n5979;
wire n5980;
wire n5981;
wire n5982;
wire n5983;
wire n5984;
wire n5985;
wire n5986;
wire n5987;
wire n5988;
wire n5989;
wire n5990;
wire n5991;
wire n5992;
wire n5993;
wire n5994;
wire n5995;
wire n5996;
wire n5997;
wire n5998;
wire n5999;
wire n6000;
wire n6001;
wire n6002;
wire n6003;
wire n6004;
wire n6005;
wire n6006;
wire n6007;
wire n6008;
wire n6009;
wire n6010;
wire n6011;
wire n6012;
wire n6013;
wire n6014;
wire n6015;
wire n6016;
wire n6017;
wire n6018;
wire n6019;
wire n6020;
wire n6021;
wire n6022;
wire n6023;
wire n6024;
wire n6025;
wire n6026;
wire n6027;
wire n6028;
wire n6029;
wire n6030;
wire n6031;
wire n6032;
wire n6033;
wire n6034;
wire n6035;
wire n6036;
wire n6037;
wire n6038;
wire n6039;
wire n6040;
wire n6041;
wire n6042;
wire n6043;
wire n6044;
wire n6045;
wire n6046;
wire n6047;
wire n6048;
wire n6049;
wire n6050;
wire n6051;
wire n6052;
wire n6053;
wire n6054;
wire n6055;
wire n6056;
wire n6057;
wire n6058;
wire n6059;
wire n6060;
wire n6061;
wire n6062;
wire n6063;
wire n6064;
wire n6065;
wire n6066;
wire n6067;
wire n6068;
wire n6069;
wire n6070;
wire n6071;
wire n6072;
wire n6073;
wire n6074;
wire n6075;
wire n6076;
wire n6077;
wire n6078;
wire n6079;
wire n6080;
wire n6081;
wire n6082;
wire n6083;
wire n6084;
wire n6085;
wire n6086;
wire n6087;
wire n6088;
wire n6089;
wire n6090;
wire n6091;
wire n6092;
wire n6093;
wire n6094;
wire n6095;
wire n6096;
wire n6097;
wire n6098;
wire n6099;
wire n6100;
wire n6101;
wire n6102;
wire n6103;
wire n6104;
wire n6105;
wire n6106;
wire n6107;
wire n6108;
wire n6109;
wire n6110;
wire n6111;
wire n6112;
wire n6113;
wire n6114;
wire n6115;
wire n6116;
wire n6117;
wire n6118;
wire n6119;
wire n6120;
wire n6121;
wire n6122;
wire n6123;
wire n6124;
wire n6125;
wire n6126;
wire n6127;
wire n6128;
wire n6129;
wire n6130;
wire n6131;
wire n6132;
wire n6133;
wire n6134;
wire n6135;
wire n6136;
wire n6137;
wire n6138;
wire n6139;
wire n6140;
wire n6141;
wire n6142;
wire n6143;
wire n6144;
wire n6145;
wire n6146;
wire n6147;
wire n6148;
wire n6149;
wire n6150;
wire n6151;
wire n6152;
wire n6153;
wire n6154;
wire n6155;
wire n6156;
wire n6157;
wire n6158;
wire n6159;
wire n6160;
wire n6161;
wire n6162;
wire n6163;
wire n6164;
wire n6165;
wire n6166;
wire n6167;
wire n6168;
wire n6169;
wire n6170;
wire n6171;
wire n6172;
wire n6173;
wire n6174;
wire n6175;
wire n6176;
wire n6177;
wire n6178;
wire n6179;
wire n6180;
wire n6181;
wire n6182;
wire n6183;
wire n6184;
wire n6185;
wire n6186;
wire n6187;
wire n6188;
wire n6189;
wire n6190;
wire n6191;
wire n6192;
wire n6193;
wire n6194;
wire n6195;
wire n6196;
wire n6197;
wire n6198;
wire n6199;
wire n6200;
wire n6201;
wire n6202;
wire n6203;
wire n6204;
wire n6205;
wire n6206;
wire n6207;
wire n6208;
wire n6209;
wire n6210;
wire n6211;
wire n6212;
wire n6213;
wire n6214;
wire n6215;
wire n6216;
wire n6217;
wire n6218;
wire n6219;
wire n6220;
wire n6221;
wire n6222;
wire n6223;
wire n6224;
wire n6225;
wire n6226;
wire n6227;
wire n6228;
wire n6229;
wire n6230;
wire n6231;
wire n6232;
wire n6233;
wire n6234;
wire n6235;
wire n6236;
wire n6237;
wire n6238;
wire n6239;
wire n6240;
wire n6241;
wire n6242;
wire n6243;
wire n6244;
wire n6245;
wire n6246;
wire n6247;
wire n6248;
wire n6249;
wire n6250;
wire n6251;
wire n6252;
wire n6253;
wire n6254;
wire n6255;
wire n6256;
wire n6257;
wire n6258;
wire n6259;
wire n6260;
wire n6261;
wire n6262;
wire n6263;
wire n6264;
wire n6265;
wire n6266;
wire n6267;
wire n6268;
wire n6269;
wire n6270;
wire n6271;
wire n6272;
wire n6273;
wire n6274;
wire n6275;
wire n6276;
wire n6277;
wire n6278;
wire n6279;
wire n6280;
wire n6281;
wire n6282;
wire n6283;
wire n6284;
wire n6285;
wire n6286;
wire n6287;
wire n6288;
wire n6289;
wire n6290;
wire n6291;
wire n6292;
wire n6293;
wire n6294;
wire n6295;
wire n6296;
wire n6297;
wire n6298;
wire n6299;
wire n6300;
wire n6301;
wire n6302;
wire n6303;
wire n6304;
wire n6305;
wire n6306;
wire n6307;
wire n6308;
wire n6309;
wire n6310;
wire n6311;
wire n6312;
wire n6313;
wire n6314;
wire n6315;
wire n6316;
wire n6317;
wire n6318;
wire n6319;
wire n6320;
wire n6321;
wire n6322;
wire n6323;
wire n6324;
wire n6325;
wire n6326;
wire n6327;
wire n6328;
wire n6329;
wire n6330;
wire n6331;
wire n6332;
wire n6333;
wire n6334;
wire n6335;
wire n6336;
wire n6337;
wire n6338;
wire n6339;
wire n6340;
wire n6341;
wire n6342;
wire n6343;
wire n6344;
wire n6345;
wire n6346;
wire n6347;
wire n6348;
wire n6349;
wire n6350;
wire n6351;
wire n6352;
wire n6353;
wire n6354;
wire n6355;
wire n6356;
wire n6357;
wire n6358;
wire n6359;
wire n6360;
wire n6361;
wire n6362;
wire n6363;
wire n6364;
wire n6365;
wire n6366;
wire n6367;
wire n6368;
wire n6369;
wire n6370;
wire n6371;
wire n6372;
wire n6373;
wire n6374;
wire n6375;
wire n6376;
wire n6377;
wire n6378;
wire n6379;
wire n6380;
wire n6381;
wire n6382;
wire n6383;
wire n6384;
wire n6385;
wire n6386;
wire n6387;
wire n6388;
wire n6389;
wire n6390;
wire n6391;
wire n6392;
wire n6393;
wire n6394;
wire n6395;
wire n6396;
wire n6397;
wire n6398;
wire n6399;
wire n6400;
wire n6401;
wire n6402;
wire n6403;
wire n6404;
wire n6405;
wire n6406;
wire n6407;
wire n6408;
wire n6409;
wire n6410;
wire n6411;
wire n6412;
wire n6413;
wire n6414;
wire n6415;
wire n6416;
wire n6417;
wire n6418;
wire n6419;
wire n6420;
wire n6421;
wire n6422;
wire n6423;
wire n6424;
wire n6425;
wire n6426;
wire n6427;
wire n6428;
wire n6429;
wire n6430;
wire n6431;
wire n6432;
wire n6433;
wire n6434;
wire n6435;
wire n6436;
wire n6437;
wire n6438;
wire n6439;
wire n6440;
wire n6441;
wire n6442;
wire n6443;
wire n6444;
wire n6445;
wire n6446;
wire n6447;
wire n6448;
wire n6449;
wire n6450;
wire n6451;
wire n6452;
wire n6453;
wire n6454;
wire n6455;
wire n6456;
wire n6457;
wire n6458;
wire n6459;
wire n6460;
wire n6461;
wire n6462;
wire n6463;
wire n6464;
wire n6465;
wire n6466;
wire n6467;
wire n6468;
wire n6469;
wire n6470;
wire n6471;
wire n6472;
wire n6473;
wire n6474;
wire n6475;
wire n6476;
wire n6477;
wire n6478;
wire n6479;
wire n6480;
wire n6481;
wire n6482;
wire n6483;
wire n6484;
wire n6485;
wire n6486;
wire n6487;
wire n6488;
wire n6489;
wire n6490;
wire n6491;
wire n6492;
wire n6493;
wire n6494;
wire n6495;
wire n6496;
wire n6497;
wire n6498;
wire n6499;
wire n6500;
wire n6501;
wire n6502;
wire n6503;
wire n6504;
wire n6505;
wire n6506;
wire n6507;
wire n6508;
wire n6509;
wire n6510;
wire n6511;
wire n6512;
wire n6513;
wire n6514;
wire n6515;
wire n6516;
wire n6517;
wire n6518;
wire n6519;
wire n6520;
wire n6521;
wire n6522;
wire n6523;
wire n6524;
wire n6525;
wire n6526;
wire n6527;
wire n6528;
wire n6529;
wire n6530;
wire n6531;
wire n6532;
wire n6533;
wire n6534;
wire n6535;
wire n6536;
wire n6537;
wire n6538;
wire n6539;
wire n6540;
wire n6541;
wire n6542;
wire n6543;
wire n6544;
wire n6545;
wire n6546;
wire n6547;
wire n6548;
wire n6549;
wire n6550;
wire n6551;
wire n6552;
wire n6553;
wire n6554;
wire n6555;
wire n6556;
wire n6557;
wire n6558;
wire n6559;
wire n6560;
wire n6561;
wire n6562;
wire n6563;
wire n6564;
wire n6565;
wire n6566;
wire n6567;
wire n6568;
wire n6569;
wire n6570;
wire n6571;
wire n6572;
wire n6573;
wire n6574;
wire n6575;
wire n6576;
wire n6577;
wire n6578;
wire n6579;
wire n6580;
wire n6581;
wire n6582;
wire n6583;
wire n6584;
wire n6585;
wire n6586;
wire n6587;
wire n6588;
wire n6589;
wire n6590;
wire n6591;
wire n6592;
wire n6593;
wire n6594;
wire n6595;
wire n6596;
wire n6597;
wire n6598;
wire n6599;
wire n6600;
wire n6601;
wire n6602;
wire n6603;
wire n6604;
wire n6605;
wire n6606;
wire n6607;
wire n6608;
wire n6609;
wire n6610;
wire n6611;
wire n6612;
wire n6613;
wire n6614;
wire n6615;
wire n6616;
wire n6617;
wire n6618;
wire n6619;
wire n6620;
wire n6621;
wire n6622;
wire n6623;
wire n6624;
wire n6625;
wire n6626;
wire n6627;
wire n6628;
wire n6629;
wire n6630;
wire n6631;
wire n6632;
wire n6633;
wire n6634;
wire n6635;
wire n6636;
wire n6637;
wire n6638;
wire n6639;
wire n6640;
wire n6641;
wire n6642;
wire n6643;
wire n6644;
wire n6645;
wire n6646;
wire n6647;
wire n6648;
wire n6649;
wire n6650;
wire n6651;
wire n6652;
wire n6653;
wire n6654;
wire n6655;
wire n6656;
wire n6657;
wire n6658;
wire n6659;
wire n6660;
wire n6661;
wire n6662;
wire n6663;
wire n6664;
wire n6665;
wire n6666;
wire n6667;
wire n6668;
wire n6669;
wire n6670;
wire n6671;
wire n6672;
wire n6673;
wire n6674;
wire n6675;
wire n6676;
wire n6677;
wire n6678;
wire n6679;
wire n6680;
wire n6681;
wire n6682;
wire n6683;
wire n6684;
wire n6685;
wire n6686;
wire n6687;
wire n6688;
wire n6689;
wire n6690;
wire n6691;
wire n6692;
wire n6693;
wire n6694;
wire n6695;
wire n6696;
wire n6697;
wire n6698;
wire n6699;
wire n6700;
wire n6701;
wire n6702;
wire n6703;
wire n6704;
wire n6705;
wire n6706;
wire n6707;
wire n6708;
wire n6709;
wire n6710;
wire n6711;
wire n6712;
wire n6713;
wire n6714;
wire n6715;
wire n6716;
wire n6717;
wire n6718;
wire n6719;
wire n6720;
wire n6721;
wire n6722;
wire n6723;
wire n6724;
wire n6725;
wire n6726;
wire n6727;
wire n6728;
wire n6729;
wire n6730;
wire n6731;
wire n6732;
wire n6733;
wire n6734;
wire n6735;
wire n6736;
wire n6737;
wire n6738;
wire n6739;
wire n6740;
wire n6741;
wire n6742;
wire n6743;
wire n6744;
wire n6745;
wire n6746;
wire n6747;
wire n6748;
wire n6749;
wire n6750;
wire n6751;
wire n6752;
wire n6753;
wire n6754;
wire n6755;
wire n6756;
wire n6757;
wire n6758;
wire n6759;
wire n6760;
wire n6761;
wire n6762;
wire n6763;
wire n6764;
wire n6765;
wire n6766;
wire n6767;
wire n6768;
wire n6769;
wire n6770;
wire n6771;
wire n6772;
wire n6773;
wire n6774;
wire n6775;
wire n6776;
wire n6777;
wire n6778;
wire n6779;
wire n6780;
wire n6781;
wire n6782;
wire n6783;
wire n6784;
wire n6785;
wire n6786;
wire n6787;
wire n6788;
wire n6789;
wire n6790;
wire n6791;
wire n6792;
wire n6793;
wire n6794;
wire n6795;
wire n6796;
wire n6797;
wire n6798;
wire n6799;
wire n6800;
wire n6801;
wire n6802;
wire n6803;
wire n6804;
wire n6805;
wire n6806;
wire n6807;
wire n6808;
wire n6809;
wire n6810;
wire n6811;
wire n6812;
wire n6813;
wire n6814;
wire n6815;
wire n6816;
wire n6817;
wire n6818;
wire n6819;
wire n6820;
wire n6821;
wire n6822;
wire n6823;
wire n6824;
wire n6825;
wire n6826;
wire n6827;
wire n6828;
wire n6829;
wire n6830;
wire n6831;
wire n6832;
wire n6833;
wire n6834;
wire n6835;
wire n6836;
wire n6837;
wire n6838;
wire n6839;
wire n6840;
wire n6841;
wire n6842;
wire n6843;
wire n6844;
wire n6845;
wire n6846;
wire n6847;
wire n6848;
wire n6849;
wire n6850;
wire n6851;
wire n6852;
wire n6853;
wire n6854;
wire n6855;
wire n6856;
wire n6857;
wire n6858;
wire n6859;
wire n6860;
wire n6861;
wire n6862;
wire n6863;
wire n6864;
wire n6865;
wire n6866;
wire n6867;
wire n6868;
wire n6869;
wire n6870;
wire n6871;
wire n6872;
wire n6873;
wire n6874;
wire n6875;
wire n6876;
wire n6877;
wire n6878;
wire n6879;
wire n6880;
wire n6881;
wire n6882;
wire n6883;
wire n6884;
wire n6885;
wire n6886;
wire n6887;
wire n6888;
wire n6889;
wire n6890;
wire n6891;
wire n6892;
wire n6893;
wire n6894;
wire n6895;
wire n6896;
wire n6897;
wire n6898;
wire n6899;
wire n6900;
wire n6901;
wire n6902;
wire n6903;
wire n6904;
wire n6905;
wire n6906;
wire n6907;
wire n6908;
wire n6909;
wire n6910;
wire n6911;
wire n6912;
wire n6913;
wire n6914;
wire n6915;
wire n6916;
wire n6917;
wire n6918;
wire n6919;
wire n6920;
wire n6921;
wire n6922;
wire n6923;
wire n6924;
wire n6925;
wire n6926;
wire n6927;
wire n6928;
wire n6929;
wire n6930;
wire n6931;
wire n6932;
wire n6933;
wire n6934;
wire n6935;
wire n6936;
wire n6937;
wire n6938;
wire n6939;
wire n6940;
wire n6941;
wire n6942;
wire n6943;
wire n6944;
wire n6945;
wire n6946;
wire n6947;
wire n6948;
wire n6949;
wire n6950;
wire n6951;
wire n6952;
wire n6953;
wire n6954;
wire n6955;
wire n6956;
wire n6957;
wire n6958;
wire n6959;
wire n6960;
wire n6961;
wire n6962;
wire n6963;
wire n6964;
wire n6965;
wire n6966;
wire n6967;
wire n6968;
wire n6969;
wire n6970;
wire n6971;
wire n6972;
wire n6973;
wire n6974;
wire n6975;
wire n6976;
wire n6977;
wire n6978;
wire n6979;
wire n6980;
wire n6981;
wire n6982;
wire n6983;
wire n6984;
wire n6985;
wire n6986;
wire n6987;
wire n6988;
wire n6989;
wire n6990;
wire n6991;
wire n6992;
wire n6993;
wire n6994;
wire n6995;
wire n6996;
wire n6997;
wire n6998;
wire n6999;
wire n7000;
wire n7001;
wire n7002;
wire n7003;
wire n7004;
wire n7005;
wire n7006;
wire n7007;
wire n7008;
wire n7009;
wire n7010;
wire n7011;
wire n7012;
wire n7013;
wire n7014;
wire n7015;
wire n7016;
wire n7017;
wire n7018;
wire n7019;
wire n7020;
wire n7021;
wire n7022;
wire n7023;
wire n7024;
wire n7025;
wire n7026;
wire n7027;
wire n7028;
wire n7029;
wire n7030;
wire n7031;
wire n7032;
wire n7033;
wire n7034;
wire n7035;
wire n7036;
wire n7037;
wire n7038;
wire n7039;
wire n7040;
wire n7041;
wire n7042;
wire n7043;
wire n7044;
wire n7045;
wire n7046;
wire n7047;
wire n7048;
wire n7049;
wire n7050;
wire n7051;
wire n7052;
wire n7053;
wire n7054;
wire n7055;
wire n7056;
wire n7057;
wire n7058;
wire n7059;
wire n7060;
wire n7061;
wire n7062;
wire n7063;
wire n7064;
wire n7065;
wire n7066;
wire n7067;
wire n7068;
wire n7069;
wire n7070;
wire n7071;
wire n7072;
wire n7073;
wire n7074;
wire n7075;
wire n7076;
wire n7077;
wire n7078;
wire n7079;
wire n7080;
wire n7081;
wire n7082;
wire n7083;
wire n7084;
wire n7085;
wire n7086;
wire n7087;
wire n7088;
wire n7089;
wire n7090;
wire n7091;
wire n7092;
wire n7093;
wire n7094;
wire n7095;
wire n7096;
wire n7097;
wire n7098;
wire n7099;
wire n7100;
wire n7101;
wire n7102;
wire n7103;
wire n7104;
wire n7105;
wire n7106;
wire n7107;
wire n7108;
wire n7109;
wire n7110;
wire n7111;
wire n7112;
wire n7113;
wire n7114;
wire n7115;
wire n7116;
wire n7117;
wire n7118;
wire n7119;
wire n7120;
wire n7121;
wire n7122;
wire n7123;
wire n7124;
wire n7125;
wire n7126;
wire n7127;
wire n7128;
wire n7129;
wire n7130;
wire n7131;
wire n7132;
wire n7133;
wire n7134;
wire n7135;
wire n7136;
wire n7137;
wire n7138;
wire n7139;
wire n7140;
wire n7141;
wire n7142;
wire n7143;
wire n7144;
wire n7145;
wire n7146;
wire n7147;
wire n7148;
wire n7149;
wire n7150;
wire n7151;
wire n7152;
wire n7153;
wire n7154;
wire n7155;
wire n7156;
wire n7157;
wire n7158;
wire n7159;
wire n7160;
wire n7161;
wire n7162;
wire n7163;
wire n7164;
wire n7165;
wire n7166;
wire n7167;
wire n7168;
wire n7169;
wire n7170;
wire n7171;
wire n7172;
wire n7173;
wire n7174;
wire n7175;
wire n7176;
wire n7177;
wire n7178;
wire n7179;
wire n7180;
wire n7181;
wire n7182;
wire n7183;
wire n7184;
wire n7185;
wire n7186;
wire n7187;
wire n7188;
wire n7189;
wire n7190;
wire n7191;
wire n7192;
wire n7193;
wire n7194;
wire n7195;
wire n7196;
wire n7197;
wire n7198;
wire n7199;
wire n7200;
wire n7201;
wire n7202;
wire n7203;
wire n7204;
wire n7205;
wire n7206;
wire n7207;
wire n7208;
wire n7209;
wire n7210;
wire n7211;
wire n7212;
wire n7213;
wire n7214;
wire n7215;
wire n7216;
wire n7217;
wire n7218;
wire n7219;
wire n7220;
wire n7221;
wire n7222;
wire n7223;
wire n7224;
wire n7225;
wire n7226;
wire n7227;
wire n7228;
wire n7229;
wire n7230;
wire n7231;
wire n7232;
wire n7233;
wire n7234;
wire n7235;
wire n7236;
wire n7237;
wire n7238;
wire n7239;
wire n7240;
wire n7241;
wire n7242;
wire n7243;
wire n7244;
wire n7245;
wire n7246;
wire n7247;
wire n7248;
wire n7249;
wire n7250;
wire n7251;
wire n7252;
wire n7253;
wire n7254;
wire n7255;
wire n7256;
wire n7257;
wire n7258;
wire n7259;
wire n7260;
wire n7261;
wire n7262;
wire n7263;
wire n7264;
wire n7265;
wire n7266;
wire n7267;
wire n7268;
wire n7269;
wire n7270;
wire n7271;
wire n7272;
wire n7273;
wire n7274;
wire n7275;
wire n7276;
wire n7277;
wire n7278;
wire n7279;
wire n7280;
wire n7281;
wire n7282;
wire n7283;
wire n7284;
wire n7285;
wire n7286;
wire n7287;
wire n7288;
wire n7289;
wire n7290;
wire n7291;
wire n7292;
wire n7293;
wire n7294;
wire n7295;
wire n7296;
wire n7297;
wire n7298;
wire n7299;
wire n7300;
wire n7301;
wire n7302;
wire n7303;
wire n7304;
wire n7305;
wire n7306;
wire n7307;
wire n7308;
wire n7309;
wire n7310;
wire n7311;
wire n7312;
wire n7313;
wire n7314;
wire n7315;
wire n7316;
wire n7317;
wire n7318;
wire n7319;
wire n7320;
wire n7321;
wire n7322;
wire n7323;
wire n7324;
wire n7325;
wire n7326;
wire n7327;
wire n7328;
wire n7329;
wire n7330;
wire n7331;
wire n7332;
wire n7333;
wire n7334;
wire n7335;
wire n7336;
wire n7337;
wire n7338;
wire n7339;
wire n7340;
wire n7341;
wire n7342;
wire n7343;
wire n7344;
wire n7345;
wire n7346;
wire n7347;
wire n7348;
wire n7349;
wire n7350;
wire n7351;
wire n7352;
wire n7353;
wire n7354;
wire n7355;
wire n7356;
wire n7357;
wire n7358;
wire n7359;
wire n7360;
wire n7361;
wire n7362;
wire n7363;
wire n7364;
wire n7365;
wire n7366;
wire n7367;
wire n7368;
wire n7369;
wire n7370;
wire n7371;
wire n7372;
wire n7373;
wire n7374;
wire n7375;
wire n7376;
wire n7377;
wire n7378;
wire n7379;
wire n7380;
wire n7381;
wire n7382;
wire n7383;
wire n7384;
wire n7385;
wire n7386;
wire n7387;
wire n7388;
wire n7389;
wire n7390;
wire n7391;
wire n7392;
wire n7393;
wire n7394;
wire n7395;
wire n7396;
wire n7397;
wire n7398;
wire n7399;
wire n7400;
wire n7401;
wire n7402;
wire n7403;
wire n7404;
wire n7405;
wire n7406;
wire n7407;
wire n7408;
wire n7409;
wire n7410;
wire n7411;
wire n7412;
wire n7413;
wire n7414;
wire n7415;
wire n7416;
wire n7417;
wire n7418;
wire n7419;
wire n7420;
wire n7421;
wire n7422;
wire n7423;
wire n7424;
wire n7425;
wire n7426;
wire n7427;
wire n7428;
wire n7429;
wire n7430;
wire n7431;
wire n7432;
wire n7433;
wire n7434;
wire n7435;
wire n7436;
wire n7437;
wire n7438;
wire n7439;
wire n7440;
wire n7441;
wire n7442;
wire n7443;
wire n7444;
wire n7445;
wire n7446;
wire n7447;
wire n7448;
wire n7449;
wire n7450;
wire n7451;
wire n7452;
wire n7453;
wire n7454;
wire n7455;
wire n7456;
wire n7457;
wire n7458;
wire n7459;
wire n7460;
wire n7461;
wire n7462;
wire n7463;
wire n7464;
wire n7465;
wire n7466;
wire n7467;
wire n7468;
wire n7469;
wire n7470;
wire n7471;
wire n7472;
wire n7473;
wire n7474;
wire n7475;
wire n7476;
wire n7477;
wire n7478;
wire n7479;
wire n7480;
wire n7481;
wire n7482;
wire n7483;
wire n7484;
wire n7485;
wire n7486;
wire n7487;
wire n7488;
wire n7489;
wire n7490;
wire n7491;
wire n7492;
wire n7493;
wire n7494;
wire n7495;
wire n7496;
wire n7497;
wire n7498;
wire n7499;
wire n7500;
wire n7501;
wire n7502;
wire n7503;
wire n7504;
wire n7505;
wire n7506;
wire n7507;
wire n7508;
wire n7509;
wire n7510;
wire n7511;
wire n7512;
wire n7513;
wire n7514;
wire n7515;
wire n7516;
wire n7517;
wire n7518;
wire n7519;
wire n7520;
wire n7521;
wire n7522;
wire n7523;
wire n7524;
wire n7525;
wire n7526;
wire n7527;
wire n7528;
wire n7529;
wire n7530;
wire n7531;
wire n7532;
wire n7533;
wire n7534;
wire n7535;
wire n7536;
wire n7537;
wire n7538;
wire n7539;
wire n7540;
wire n7541;
wire n7542;
wire n7543;
wire n7544;
wire n7545;
wire n7546;
wire n7547;
wire n7548;
wire n7549;
wire n7550;
wire n7551;
wire n7552;
wire n7553;
wire n7554;
wire n7555;
wire n7556;
wire n7557;
wire n7558;
wire n7559;
wire n7560;
wire n7561;
wire n7562;
wire n7563;
wire n7564;
wire n7565;
wire n7566;
wire n7567;
wire n7568;
wire n7569;
wire n7570;
wire n7571;
wire n7572;
wire n7573;
wire n7574;
wire n7575;
wire n7576;
wire n7577;
wire n7578;
wire n7579;
wire n7580;
wire n7581;
wire n7582;
wire n7583;
wire n7584;
wire n7585;
wire n7586;
wire n7587;
wire n7588;
wire n7589;
wire n7590;
wire n7591;
wire n7592;
wire n7593;
wire n7594;
wire n7595;
wire n7596;
wire n7597;
wire n7598;
wire n7599;
wire n7600;
wire n7601;
wire n7602;
wire n7603;
wire n7604;
wire n7605;
wire n7606;
wire n7607;
wire n7608;
wire n7609;
wire n7610;
wire n7611;
wire n7612;
wire n7613;
wire n7614;
wire n7615;
wire n7616;
wire n7617;
wire n7618;
wire n7619;
wire n7620;
wire n7621;
wire n7622;
wire n7623;
wire n7624;
wire n7625;
wire n7626;
wire n7627;
wire n7628;
wire n7629;
wire n7630;
wire n7631;
wire n7632;
wire n7633;
wire n7634;
wire n7635;
wire n7636;
wire n7637;
wire n7638;
wire n7639;
wire n7640;
wire n7641;
wire n7642;
wire n7643;
wire n7644;
wire n7645;
wire n7646;
wire n7647;
wire n7648;
wire n7649;
wire n7650;
wire n7651;
wire n7652;
wire n7653;
wire n7654;
wire n7655;
wire n7656;
wire n7657;
wire n7658;
wire n7659;
wire n7660;
wire n7661;
wire n7662;
wire n7663;
wire n7664;
wire n7665;
wire n7666;
wire n7667;
wire n7668;
wire n7669;
wire n7670;
wire n7671;
wire n7672;
wire n7673;
wire n7674;
wire n7675;
wire n7676;
wire n7677;
wire n7678;
wire n7679;
wire n7680;
wire n7681;
wire n7682;
wire n7683;
wire n7684;
wire n7685;
wire n7686;
wire n7687;
wire n7688;
wire n7689;
wire n7690;
wire n7691;
wire n7692;
wire n7693;
wire n7694;
wire n7695;
wire n7696;
wire n7697;
wire n7698;
wire n7699;
wire n7700;
wire n7701;
wire n7702;
wire n7703;
wire n7704;
wire n7705;
wire n7706;
wire n7707;
wire n7708;
wire n7709;
wire n7710;
wire n7711;
wire n7712;
wire n7713;
wire n7714;
wire n7715;
wire n7716;
wire n7717;
wire n7718;
wire n7719;
wire n7720;
wire n7721;
wire n7722;
wire n7723;
wire n7724;
wire n7725;
wire n7726;
wire n7727;
wire n7728;
wire n7729;
wire n7730;
wire n7731;
wire n7732;
wire n7733;
wire n7734;
wire n7735;
wire n7736;
wire n7737;
wire n7738;
wire n7739;
wire n7740;
wire n7741;
wire n7742;
wire n7743;
wire n7744;
wire n7745;
wire n7746;
wire n7747;
wire n7748;
wire n7749;
wire n7750;
wire n7751;
wire n7752;
wire n7753;
wire n7754;
wire n7755;
wire n7756;
wire n7757;
wire n7758;
wire n7759;
wire n7760;
wire n7761;
wire n7762;
wire n7763;
wire n7764;
wire n7765;
wire n7766;
wire n7767;
wire n7768;
wire n7769;
wire n7770;
wire n7771;
wire n7772;
wire n7773;
wire n7774;
wire n7775;
wire n7776;
wire n7777;
wire n7778;
wire n7779;
wire n7780;
wire n7781;
wire n7782;
wire n7783;
wire n7784;
wire n7785;
wire n7786;
wire n7787;
wire n7788;
wire n7789;
wire n7790;
wire n7791;
wire n7792;
wire n7793;
wire n7794;
wire n7795;
wire n7796;
wire n7797;
wire n7798;
wire n7799;
wire n7800;
wire n7801;
wire n7802;
wire n7803;
wire n7804;
wire n7805;
wire n7806;
wire n7807;
wire n7808;
wire n7809;
wire n7810;
wire n7811;
wire n7812;
wire n7813;
wire n7814;
wire n7815;
wire n7816;
wire n7817;
wire n7818;
wire n7819;
wire n7820;
wire n7821;
wire n7822;
wire n7823;
wire n7824;
wire n7825;
wire n7826;
wire n7827;
wire n7828;
wire n7829;
wire n7830;
wire n7831;
wire n7832;
wire n7833;
wire n7834;
wire n7835;
wire n7836;
wire n7837;
wire n7838;
wire n7839;
wire n7840;
wire n7841;
wire n7842;
wire n7843;
wire n7844;
wire n7845;
wire n7846;
wire n7847;
wire n7848;
wire n7849;
wire n7850;
wire n7851;
wire n7852;
wire n7853;
wire n7854;
wire n7855;
wire n7856;
wire n7857;
wire n7858;
wire n7859;
wire n7860;
wire n7861;
wire n7862;
wire n7863;
wire n7864;
wire n7865;
wire n7866;
wire n7867;
wire n7868;
wire n7869;
wire n7870;
wire n7871;
wire n7872;
wire n7873;
wire n7874;
wire n7875;
wire n7876;
wire n7877;
wire n7878;
wire n7879;
wire n7880;
wire n7881;
wire n7882;
wire n7883;
wire n7884;
wire n7885;
wire n7886;
wire n7887;
wire n7888;
wire n7889;
wire n7890;
wire n7891;
wire n7892;
wire n7893;
wire n7894;
wire n7895;
wire n7896;
wire n7897;
wire n7898;
wire n7899;
wire n7900;
wire n7901;
wire n7902;
wire n7903;
wire n7904;
wire n7905;
wire n7906;
wire n7907;
wire n7908;
wire n7909;
wire n7910;
wire n7911;
wire n7912;
wire n7913;
wire n7914;
wire n7915;
wire n7916;
wire n7917;
wire n7918;
wire n7919;
wire n7920;
wire n7921;
wire n7922;
wire n7923;
wire n7924;
wire n7925;
wire n7926;
wire n7927;
wire n7928;
wire n7929;
wire n7930;
wire n7931;
wire n7932;
wire n7933;
wire n7934;
wire n7935;
wire n7936;
wire n7937;
wire n7938;
wire n7939;
wire n7940;
wire n7941;
wire n7942;
wire n7943;
wire n7944;
wire n7945;
wire n7946;
wire n7947;
wire n7948;
wire n7949;
wire n7950;
wire n7951;
wire n7952;
wire n7953;
wire n7954;
wire n7955;
wire n7956;
wire n7957;
wire n7958;
wire n7959;
wire n7960;
wire n7961;
wire n7962;
wire n7963;
wire n7964;
wire n7965;
wire n7966;
wire n7967;
wire n7968;
wire n7969;
wire n7970;
wire n7971;
wire n7972;
wire n7973;
wire n7974;
wire n7975;
wire n7976;
wire n7977;
wire n7978;
wire n7979;
wire n7980;
wire n7981;
wire n7982;
wire n7983;
wire n7984;
wire n7985;
wire n7986;
wire n7987;
wire n7988;
wire n7989;
wire n7990;
wire n7991;
wire n7992;
wire n7993;
wire n7994;
wire n7995;
wire n7996;
wire n7997;
wire n7998;
wire n7999;
wire n8000;
wire n8001;
wire n8002;
wire n8003;
wire n8004;
wire n8005;
wire n8006;
wire n8007;
wire n8008;
wire n8009;
wire n8010;
wire n8011;
wire n8012;
wire n8013;
wire n8014;
wire n8015;
wire n8016;
wire n8017;
wire n8018;
wire n8019;
wire n8020;
wire n8021;
wire n8022;
wire n8023;
wire n8024;
wire n8025;
wire n8026;
wire n8027;
wire n8028;
wire n8029;
wire n8030;
wire n8031;
wire n8032;
wire n8033;
wire n8034;
wire n8035;
wire n8036;
wire n8037;
wire n8038;
wire n8039;
wire n8040;
wire n8041;
wire n8042;
wire n8043;
wire n8044;
wire n8045;
wire n8046;
wire n8047;
wire n8048;
wire n8049;
wire n8050;
wire n8051;
wire n8052;
wire n8053;
wire n8054;
wire n8055;
wire n8056;
wire n8057;
wire n8058;
wire n8059;
wire n8060;
wire n8061;
wire n8062;
wire n8063;
wire n8064;
wire n8065;
wire n8066;
wire n8067;
wire n8068;
wire n8069;
wire n8070;
wire n8071;
wire n8072;
wire n8073;
wire n8074;
wire n8075;
wire n8076;
wire n8077;
wire n8078;
wire n8079;
wire n8080;
wire n8081;
wire n8082;
wire n8083;
wire n8084;
wire n8085;
wire n8086;
wire n8087;
wire n8088;
wire n8089;
wire n8090;
wire n8091;
wire n8092;
wire n8093;
wire n8094;
wire n8095;
wire n8096;
wire n8097;
wire n8098;
wire n8099;
wire n8100;
wire n8101;
wire n8102;
wire n8103;
wire n8104;
wire n8105;
wire n8106;
wire n8107;
wire n8108;
wire n8109;
wire n8110;
wire n8111;
wire n8112;
wire n8113;
wire n8114;
wire n8115;
wire n8116;
wire n8117;
wire n8118;
wire n8119;
wire n8120;
wire n8121;
wire n8122;
wire n8123;
wire n8124;
wire n8125;
wire n8126;
wire n8127;
wire n8128;
wire n8129;
wire n8130;
wire n8131;
wire n8132;
wire n8133;
wire n8134;
wire n8135;
wire n8136;
wire n8137;
wire n8138;
wire n8139;
wire n8140;
wire n8141;
wire n8142;
wire n8143;
wire n8144;
wire n8145;
wire n8146;
wire n8147;
wire n8148;
wire n8149;
wire n8150;
wire n8151;
wire n8152;
wire n8153;
wire n8154;
wire n8155;
wire n8156;
wire n8157;
wire n8158;
wire n8159;
wire n8160;
wire n8161;
wire n8162;
wire n8163;
wire n8164;
wire n8165;
wire n8166;
wire n8167;
wire n8168;
wire n8169;
wire n8170;
wire n8171;
wire n8172;
wire n8173;
wire n8174;
wire n8175;
wire n8176;
wire n8177;
wire n8178;
wire n8179;
wire n8180;
wire n8181;
wire n8182;
wire n8183;
wire n8184;
wire n8185;
wire n8186;
wire n8187;
wire n8188;
wire n8189;
wire n8190;
wire n8191;
wire n8192;
wire n8193;
wire n8194;
wire n8195;
wire n8196;
wire n8197;
wire n8198;
wire n8199;
wire n8200;
wire n8201;
wire n8202;
wire n8203;
wire n8204;
wire n8205;
wire n8206;
wire n8207;
wire n8208;
wire n8209;
wire n8210;
wire n8211;
wire n8212;
wire n8213;
wire n8214;
wire n8215;
wire n8216;
wire n8217;
wire n8218;
wire n8219;
wire n8220;
wire n8221;
wire n8222;
wire n8223;
wire n8224;
wire n8225;
wire n8226;
wire n8227;
wire n8228;
wire n8229;
wire n8230;
wire n8231;
wire n8232;
wire n8233;
wire n8234;
wire n8235;
wire n8236;
wire n8237;
wire n8238;
wire n8239;
wire n8240;
wire n8241;
wire n8242;
wire n8243;
wire n8244;
wire n8245;
wire n8246;
wire n8247;
wire n8248;
wire n8249;
wire n8250;
wire n8251;
wire n8252;
wire n8253;
wire n8254;
wire n8255;
wire n8256;
wire n8257;
wire n8258;
wire n8259;
wire n8260;
wire n8261;
wire n8262;
wire n8263;
wire n8264;
wire n8265;
wire n8266;
wire n8267;
wire n8268;
wire n8269;
wire n8270;
wire n8271;
wire n8272;
wire n8273;
wire n8274;
wire n8275;
wire n8276;
wire n8277;
wire n8278;
wire n8279;
wire n8280;
wire n8281;
wire n8282;
wire n8283;
wire n8284;
wire n8285;
wire n8286;
wire n8287;
wire n8288;
wire n8289;
wire n8290;
wire n8291;
wire n8292;
wire n8293;
wire n8294;
wire n8295;
wire n8296;
wire n8297;
wire n8298;
wire n8299;
wire n8300;
wire n8301;
wire n8302;
wire n8303;
wire n8304;
wire n8305;
wire n8306;
wire n8307;
wire n8308;
wire n8309;
wire n8310;
wire n8311;
wire n8312;
wire n8313;
wire n8314;
wire n8315;
wire n8316;
wire n8317;
wire n8318;
wire n8319;
wire n8320;
wire n8321;
wire n8322;
wire n8323;
wire n8324;
wire n8325;
wire n8326;
wire n8327;
wire n8328;
wire n8329;
wire n8330;
wire n8331;
wire n8332;
wire n8333;
wire n8334;
wire n8335;
wire n8336;
wire n8337;
wire n8338;
wire n8339;
wire n8340;
wire n8341;
wire n8342;
wire n8343;
wire n8344;
wire n8345;
wire n8346;
wire n8347;
wire n8348;
wire n8349;
wire n8350;
wire n8351;
wire n8352;
wire n8353;
wire n8354;
wire n8355;
wire n8356;
wire n8357;
wire n8358;
wire n8359;
wire n8360;
wire n8361;
wire n8362;
wire n8363;
wire n8364;
wire n8365;
wire n8366;
wire n8367;
wire n8368;
wire n8369;
wire n8370;
wire n8371;
wire n8372;
wire n8373;
wire n8374;
wire n8375;
wire n8376;
wire n8377;
wire n8378;
wire n8379;
wire n8380;
wire n8381;
wire n8382;
wire n8383;
wire n8384;
wire n8385;
wire n8386;
wire n8387;
wire n8388;
wire n8389;
wire n8390;
wire n8391;
wire n8392;
wire n8393;
wire n8394;
wire n8395;
wire n8396;
wire n8397;
wire n8398;
wire n8399;
wire n8400;
wire n8401;
wire n8402;
wire n8403;
wire n8404;
wire n8405;
wire n8406;
wire n8407;
wire n8408;
wire n8409;
wire n8410;
wire n8411;
wire n8412;
wire n8413;
wire n8414;
wire n8415;
wire n8416;
wire n8417;
wire n8418;
wire n8419;
xor (out,n0,n4392);
nand (n0,n1,n11);
or (n1,n2,n4);
not (n2,n3);
not (n4,n5);
nand (n5,n6,n8,n10);
not (n6,n7);
not (n8,n9);
nand (n11,n12,n4);
nand (n12,n13,n4391);
or (n13,n14,n1146);
not (n14,n15);
nand (n15,n16,n1145);
or (n16,n17,n1028);
xor (n17,n18,n859);
xor (n18,n19,n587);
xor (n19,n20,n510);
xor (n20,n21,n252);
xor (n21,n22,n175);
xor (n22,n23,n98);
xor (n23,n24,n70);
xor (n24,n25,n45);
nand (n25,n26,n40);
or (n26,n27,n28);
nor (n27,n28,n34);
nand (n28,n29,n33);
or (n29,n30,n31);
not (n31,n32);
nand (n33,n30,n31);
nor (n34,n35,n38);
and (n35,n30,n36);
not (n36,n37);
and (n38,n37,n39);
not (n39,n30);
nand (n40,n41,n44);
or (n41,n37,n42);
not (n42,n43);
or (n44,n36,n43);
nand (n45,n46,n64);
or (n46,n47,n58);
nand (n47,n48,n54);
not (n48,n49);
nand (n49,n50,n53);
or (n50,n37,n51);
not (n51,n52);
nand (n53,n37,n51);
nand (n54,n55,n57);
or (n55,n56,n51);
nand (n57,n56,n51);
nor (n58,n59,n62);
and (n59,n60,n61);
not (n60,n56);
and (n62,n56,n63);
not (n63,n61);
or (n64,n48,n65);
nor (n65,n66,n68);
and (n66,n60,n67);
and (n68,n56,n69);
not (n69,n67);
nand (n70,n71,n91);
or (n71,n72,n86);
not (n72,n73);
nor (n73,n74,n80);
nand (n74,n75,n79);
or (n75,n76,n77);
not (n77,n78);
nand (n79,n76,n77);
nor (n80,n81,n84);
and (n81,n82,n76);
not (n82,n83);
and (n84,n83,n85);
not (n85,n76);
nor (n86,n87,n89);
and (n87,n82,n88);
and (n89,n83,n90);
not (n90,n88);
or (n91,n92,n93);
not (n92,n74);
nor (n93,n94,n96);
and (n94,n82,n95);
and (n96,n83,n97);
not (n97,n95);
xor (n98,n99,n153);
xor (n99,n100,n128);
nand (n100,n101,n121);
or (n101,n102,n116);
not (n102,n103);
nor (n103,n104,n111);
nor (n104,n105,n109);
and (n105,n106,n107);
not (n107,n108);
and (n109,n110,n108);
not (n110,n106);
nand (n111,n112,n115);
or (n112,n113,n108);
not (n113,n114);
nand (n115,n108,n113);
nor (n116,n117,n119);
and (n117,n110,n118);
and (n119,n106,n120);
not (n120,n118);
or (n121,n122,n127);
nor (n122,n123,n125);
and (n123,n110,n124);
and (n125,n106,n126);
not (n126,n124);
not (n127,n111);
nand (n128,n129,n147);
or (n129,n130,n142);
not (n130,n131);
and (n131,n132,n137);
nor (n132,n133,n135);
and (n133,n110,n134);
and (n135,n106,n136);
not (n136,n134);
nor (n137,n138,n141);
and (n138,n139,n136);
not (n139,n140);
and (n141,n140,n134);
nor (n142,n143,n145);
and (n143,n139,n144);
and (n145,n140,n146);
not (n146,n144);
or (n147,n132,n148);
nor (n148,n149,n151);
and (n149,n139,n150);
and (n151,n140,n152);
not (n152,n150);
nand (n153,n154,n169);
or (n154,n155,n164);
nand (n155,n156,n161);
nor (n156,n157,n160);
and (n157,n56,n158);
not (n158,n159);
and (n160,n60,n159);
nand (n161,n162,n163);
or (n162,n159,n77);
nand (n163,n77,n159);
nor (n164,n165,n167);
and (n165,n77,n166);
and (n167,n78,n168);
not (n168,n166);
or (n169,n156,n170);
nor (n170,n171,n173);
and (n171,n77,n172);
and (n173,n78,n174);
not (n174,n172);
xor (n175,n176,n226);
xor (n176,n177,n204);
nand (n177,n178,n198);
or (n178,n179,n193);
nand (n179,n180,n188);
not (n180,n181);
nor (n181,n182,n186);
and (n182,n183,n185);
not (n183,n184);
and (n186,n184,n187);
not (n187,n185);
and (n188,n189,n191);
nand (n189,n183,n190);
nand (n191,n192,n184);
not (n192,n190);
nor (n193,n194,n196);
and (n194,n187,n195);
and (n196,n185,n197);
not (n197,n195);
or (n198,n188,n199);
nor (n199,n200,n202);
and (n200,n187,n201);
and (n202,n185,n203);
not (n203,n201);
nand (n204,n205,n220);
or (n205,n206,n215);
nand (n206,n207,n212);
nor (n207,n208,n210);
and (n208,n187,n209);
and (n210,n185,n211);
not (n211,n209);
nand (n212,n213,n214);
or (n213,n209,n113);
nand (n214,n113,n209);
nor (n215,n216,n218);
and (n216,n113,n217);
and (n218,n114,n219);
not (n219,n217);
or (n220,n207,n221);
nor (n221,n222,n224);
and (n222,n113,n223);
and (n224,n114,n225);
not (n225,n223);
nand (n226,n227,n246);
or (n227,n228,n241);
nand (n228,n229,n234);
not (n229,n230);
nand (n230,n231,n233);
or (n231,n82,n232);
nand (n233,n82,n232);
not (n234,n235);
nor (n235,n236,n239);
and (n236,n237,n238);
not (n237,n232);
and (n239,n232,n240);
not (n240,n238);
nor (n241,n242,n244);
and (n242,n240,n243);
and (n244,n238,n245);
not (n245,n243);
or (n246,n229,n247);
nor (n247,n248,n250);
and (n248,n240,n249);
and (n250,n238,n251);
not (n251,n249);
or (n252,n253,n509);
and (n253,n254,n454);
xor (n254,n255,n323);
or (n255,n256,n322);
and (n256,n257,n311);
xor (n257,n258,n284);
nand (n258,n259,n277);
or (n259,n260,n272);
not (n260,n261);
nor (n261,n262,n269);
nor (n262,n263,n267);
and (n263,n264,n266);
not (n264,n265);
and (n267,n265,n268);
not (n268,n266);
nor (n269,n270,n271);
and (n270,n266,n238);
and (n271,n268,n240);
nor (n272,n273,n275);
and (n273,n264,n274);
and (n275,n265,n276);
not (n276,n274);
or (n277,n278,n279);
not (n278,n269);
nor (n279,n280,n282);
and (n280,n264,n281);
and (n282,n265,n283);
not (n283,n281);
nand (n284,n285,n305);
or (n285,n286,n300);
not (n286,n287);
and (n287,n288,n295);
nor (n288,n289,n293);
and (n289,n290,n291);
not (n291,n292);
and (n293,n294,n292);
not (n294,n290);
nor (n295,n296,n299);
and (n296,n297,n291);
not (n297,n298);
and (n299,n298,n292);
nor (n300,n301,n303);
and (n301,n297,n302);
and (n303,n304,n298);
not (n304,n302);
or (n305,n288,n306);
nor (n306,n307,n309);
and (n307,n308,n297);
and (n309,n310,n298);
not (n310,n308);
nand (n311,n312,n317);
or (n312,n313,n314);
not (n313,n27);
nor (n314,n315,n316);
and (n315,n36,n172);
and (n316,n37,n174);
or (n317,n318,n319);
not (n318,n28);
nor (n319,n320,n321);
and (n320,n36,n61);
and (n321,n37,n63);
and (n322,n258,n284);
or (n323,n324,n453);
and (n324,n325,n405);
xor (n325,n326,n369);
or (n326,n327,n368);
and (n327,n328,n359);
xor (n328,n329,n338);
nand (n329,n330,n334);
or (n330,n155,n331);
nor (n331,n332,n333);
and (n332,n77,n249);
and (n333,n78,n251);
or (n334,n156,n335);
nor (n335,n336,n337);
and (n336,n77,n88);
and (n337,n78,n90);
nand (n338,n339,n354);
or (n339,n340,n344);
not (n340,n341);
nand (n341,n342,n343);
or (n342,n190,n225);
or (n343,n192,n223);
not (n344,n345);
nor (n345,n346,n350);
nand (n346,n347,n349);
or (n347,n348,n264);
nand (n349,n348,n264);
nor (n350,n351,n352);
and (n351,n192,n348);
and (n352,n190,n353);
not (n353,n348);
nand (n354,n355,n346);
not (n355,n356);
nor (n356,n357,n358);
and (n357,n192,n195);
and (n358,n190,n197);
nand (n359,n360,n364);
or (n360,n179,n361);
nor (n361,n362,n363);
and (n362,n187,n124);
and (n363,n185,n126);
or (n364,n188,n365);
nor (n365,n366,n367);
and (n366,n187,n217);
and (n367,n185,n219);
and (n368,n329,n338);
or (n369,n370,n404);
and (n370,n371,n392);
xor (n371,n372,n383);
nand (n372,n373,n379);
or (n373,n72,n374);
nor (n374,n375,n378);
and (n375,n376,n83);
not (n376,n377);
and (n378,n377,n82);
or (n379,n92,n380);
nor (n380,n381,n382);
and (n381,n82,n243);
and (n382,n83,n245);
nand (n383,n384,n388);
or (n384,n206,n385);
nor (n385,n386,n387);
and (n386,n113,n150);
and (n387,n114,n152);
or (n388,n207,n389);
nor (n389,n390,n391);
and (n390,n113,n118);
and (n391,n114,n120);
nand (n392,n393,n400);
or (n393,n102,n394);
not (n394,n395);
nor (n395,n396,n399);
and (n396,n397,n110);
not (n397,n398);
and (n399,n398,n106);
or (n400,n401,n127);
nor (n401,n402,n403);
and (n402,n110,n144);
and (n403,n106,n146);
and (n404,n372,n383);
or (n405,n406,n452);
and (n406,n407,n439);
xor (n407,n408,n428);
nand (n408,n409,n424);
or (n409,n410,n421);
nand (n410,n411,n418);
nor (n411,n412,n416);
and (n412,n413,n415);
not (n413,n414);
and (n416,n417,n414);
not (n417,n415);
nand (n418,n419,n420);
or (n419,n414,n31);
nand (n420,n414,n31);
nor (n421,n422,n423);
and (n422,n69,n32);
and (n423,n67,n31);
or (n424,n411,n425);
nor (n425,n426,n427);
and (n426,n31,n43);
and (n427,n32,n42);
nand (n428,n429,n433);
or (n429,n228,n430);
nor (n430,n431,n432);
and (n431,n240,n281);
and (n432,n238,n283);
or (n433,n229,n434);
nor (n434,n435,n437);
and (n435,n240,n436);
and (n437,n238,n438);
not (n438,n436);
nand (n439,n440,n446);
or (n440,n130,n441);
nor (n441,n442,n444);
and (n442,n139,n443);
and (n444,n140,n445);
not (n445,n443);
or (n446,n132,n447);
nor (n447,n448,n450);
and (n448,n139,n449);
and (n450,n140,n451);
not (n451,n449);
and (n452,n408,n428);
and (n453,n326,n369);
xor (n454,n455,n487);
xor (n455,n456,n464);
not (n456,n457);
nand (n457,n458,n463);
or (n458,n459,n47);
not (n459,n460);
nand (n460,n461,n462);
or (n461,n56,n174);
or (n462,n60,n172);
or (n463,n48,n58);
or (n464,n465,n486);
and (n465,n466,n480);
xor (n466,n467,n474);
nand (n467,n468,n469);
or (n468,n344,n356);
or (n469,n470,n471);
not (n470,n346);
nor (n471,n472,n473);
and (n472,n192,n201);
and (n473,n190,n203);
nand (n474,n475,n476);
or (n475,n179,n365);
or (n476,n188,n477);
nor (n477,n478,n479);
and (n478,n187,n223);
and (n479,n185,n225);
nand (n480,n481,n482);
or (n481,n72,n380);
or (n482,n92,n483);
nor (n483,n484,n485);
and (n484,n82,n249);
and (n485,n83,n251);
and (n486,n467,n474);
or (n487,n488,n508);
and (n488,n489,n502);
xor (n489,n490,n496);
nand (n490,n491,n492);
or (n491,n206,n389);
or (n492,n207,n493);
nor (n493,n494,n495);
and (n494,n113,n124);
and (n495,n114,n126);
nand (n496,n497,n498);
or (n497,n102,n401);
or (n498,n127,n499);
nor (n499,n500,n501);
and (n500,n110,n150);
and (n501,n106,n152);
nand (n502,n503,n504);
or (n503,n459,n48);
or (n504,n47,n505);
nor (n505,n506,n507);
and (n506,n60,n166);
and (n507,n56,n168);
and (n508,n490,n496);
and (n509,n255,n323);
xor (n510,n511,n584);
xor (n511,n512,n554);
xor (n512,n513,n543);
xor (n513,n514,n523);
nand (n514,n515,n519);
or (n515,n260,n516);
nor (n516,n517,n518);
and (n517,n264,n436);
and (n518,n265,n438);
or (n519,n278,n520);
nor (n520,n521,n522);
and (n521,n264,n377);
and (n522,n265,n376);
nand (n523,n524,n539);
or (n524,n525,n529);
not (n525,n526);
nand (n526,n527,n528);
or (n527,n451,n290);
or (n528,n294,n449);
nand (n529,n530,n535);
not (n530,n531);
nand (n531,n532,n534);
or (n532,n533,n139);
nand (n534,n533,n139);
nor (n535,n536,n538);
and (n536,n537,n294);
not (n537,n533);
and (n538,n533,n290);
or (n539,n530,n540);
nor (n540,n541,n542);
and (n541,n398,n294);
and (n542,n397,n290);
nand (n543,n544,n548);
or (n544,n545,n288);
nor (n545,n546,n547);
and (n546,n443,n297);
and (n547,n445,n298);
or (n548,n286,n549);
nor (n549,n550,n552);
and (n550,n551,n297);
and (n552,n553,n298);
not (n553,n551);
xor (n554,n555,n565);
xor (n555,n556,n457);
nand (n556,n557,n561);
or (n557,n344,n558);
nor (n558,n559,n560);
and (n559,n192,n274);
and (n560,n190,n276);
or (n561,n470,n562);
nor (n562,n563,n564);
and (n563,n192,n281);
and (n564,n190,n283);
or (n565,n566,n583);
and (n566,n567,n577);
xor (n567,n568,n574);
nand (n568,n569,n573);
or (n569,n228,n570);
nor (n570,n571,n572);
and (n571,n376,n238);
and (n572,n377,n240);
or (n573,n229,n241);
nand (n574,n575,n576);
or (n575,n102,n499);
or (n576,n116,n127);
nand (n577,n578,n582);
or (n578,n130,n579);
nor (n579,n580,n581);
and (n580,n139,n398);
and (n581,n140,n397);
or (n582,n132,n142);
and (n583,n568,n574);
or (n584,n585,n586);
and (n585,n455,n487);
and (n586,n456,n464);
xor (n587,n588,n729);
xor (n588,n589,n686);
or (n589,n590,n685);
and (n590,n591,n678);
xor (n591,n592,n647);
xor (n592,n593,n636);
xor (n593,n594,n614);
or (n594,n595,n613);
and (n595,n596,n604);
xor (n596,n597,n601);
nand (n597,n598,n599);
or (n598,n434,n228);
nand (n599,n600,n230);
not (n600,n570);
nand (n601,n602,n603);
or (n602,n130,n447);
or (n603,n132,n579);
nand (n604,n605,n609);
or (n605,n529,n606);
nor (n606,n607,n608);
and (n607,n551,n294);
and (n608,n290,n553);
or (n609,n530,n610);
nor (n610,n611,n612);
and (n611,n443,n294);
and (n612,n445,n290);
and (n613,n597,n601);
or (n614,n615,n635);
and (n615,n616,n629);
xor (n616,n617,n622);
nand (n617,n618,n621);
or (n618,n619,n620);
not (n619,n411);
not (n620,n410);
not (n621,n425);
nand (n622,n623,n624);
or (n623,n313,n319);
or (n624,n318,n625);
not (n625,n626);
nand (n626,n627,n628);
or (n627,n37,n69);
or (n628,n36,n67);
nand (n629,n630,n631);
or (n630,n155,n335);
or (n631,n156,n632);
nor (n632,n633,n634);
and (n633,n77,n95);
and (n634,n78,n97);
and (n635,n617,n622);
xor (n636,n637,n644);
xor (n637,n638,n641);
nand (n638,n639,n640);
or (n639,n286,n306);
or (n640,n288,n549);
nand (n641,n642,n643);
or (n642,n155,n632);
or (n643,n156,n164);
nand (n644,n645,n646);
or (n645,n344,n471);
or (n646,n470,n558);
or (n647,n648,n677);
and (n648,n649,n676);
xor (n649,n650,n675);
or (n650,n651,n674);
and (n651,n652,n666);
xor (n652,n653,n659);
nand (n653,n654,n658);
or (n654,n529,n655);
nor (n655,n656,n657);
and (n656,n308,n294);
and (n657,n290,n310);
or (n658,n530,n606);
nand (n659,n660,n664);
or (n660,n661,n47);
nor (n661,n662,n663);
and (n662,n60,n95);
and (n663,n56,n97);
nand (n664,n665,n49);
not (n665,n505);
nand (n666,n667,n673);
or (n667,n286,n668);
nor (n668,n669,n671);
and (n669,n297,n670);
and (n671,n672,n298);
not (n672,n670);
or (n673,n288,n300);
and (n674,n653,n659);
xor (n675,n466,n480);
xor (n676,n616,n629);
and (n677,n650,n675);
or (n678,n679,n684);
and (n679,n680,n683);
xor (n680,n681,n682);
xor (n681,n596,n604);
xor (n682,n489,n502);
xor (n683,n257,n311);
and (n684,n681,n682);
and (n685,n592,n647);
xor (n686,n687,n722);
xor (n687,n688,n719);
xor (n688,n689,n706);
xor (n689,n690,n703);
or (n690,n691,n702);
and (n691,n692,n699);
xor (n692,n693,n696);
nand (n693,n694,n695);
or (n694,n625,n313);
nand (n695,n28,n40);
nand (n696,n697,n698);
or (n697,n260,n279);
or (n698,n278,n516);
nand (n699,n700,n701);
or (n700,n529,n610);
or (n701,n530,n525);
and (n702,n693,n696);
or (n703,n704,n705);
and (n704,n637,n644);
and (n705,n638,n641);
or (n706,n707,n718);
and (n707,n708,n715);
xor (n708,n709,n712);
nand (n709,n710,n711);
or (n710,n72,n483);
or (n711,n92,n86);
nand (n712,n713,n714);
or (n713,n179,n477);
or (n714,n188,n193);
nand (n715,n716,n717);
or (n716,n206,n493);
or (n717,n207,n215);
and (n718,n709,n712);
or (n719,n720,n721);
and (n720,n593,n636);
and (n721,n594,n614);
or (n722,n723,n728);
and (n723,n724,n727);
xor (n724,n725,n726);
xor (n725,n708,n715);
xor (n726,n692,n699);
xor (n727,n567,n577);
and (n728,n725,n726);
or (n729,n730,n858);
and (n730,n731,n857);
xor (n731,n732,n733);
xor (n732,n724,n727);
or (n733,n734,n856);
and (n734,n735,n855);
xor (n735,n736,n771);
or (n736,n737,n770);
and (n737,n738,n746);
xor (n738,n739,n745);
nand (n739,n740,n744);
or (n740,n260,n741);
nor (n741,n742,n743);
and (n742,n264,n201);
and (n743,n265,n203);
or (n744,n278,n272);
not (n745,n311);
or (n746,n747,n769);
and (n747,n748,n762);
xor (n748,n749,n755);
nand (n749,n750,n754);
or (n750,n72,n751);
nor (n751,n752,n753);
and (n752,n436,n82);
and (n753,n83,n438);
or (n754,n92,n374);
nand (n755,n756,n761);
or (n756,n757,n102);
not (n757,n758);
nor (n758,n759,n760);
and (n759,n451,n110);
and (n760,n449,n106);
nand (n761,n395,n111);
nand (n762,n763,n768);
or (n763,n130,n764);
not (n764,n765);
nand (n765,n766,n767);
or (n766,n553,n140);
or (n767,n139,n551);
or (n768,n132,n441);
and (n769,n749,n755);
and (n770,n739,n745);
or (n771,n772,n854);
and (n772,n773,n832);
xor (n773,n774,n808);
or (n774,n775,n807);
and (n775,n776,n801);
xor (n776,n777,n793);
nand (n777,n778,n790);
or (n778,n779,n785);
nand (n779,n780,n784);
or (n780,n781,n782);
not (n782,n783);
nand (n784,n782,n781);
nor (n785,n779,n786);
nor (n786,n787,n788);
and (n787,n417,n781);
and (n788,n415,n789);
not (n789,n781);
nor (n790,n791,n792);
and (n791,n43,n415);
and (n792,n42,n417);
nand (n793,n794,n799);
or (n794,n795,n410);
not (n795,n796);
nor (n796,n797,n798);
and (n797,n61,n32);
and (n798,n63,n31);
nand (n799,n800,n619);
not (n800,n421);
nand (n801,n802,n806);
or (n802,n47,n803);
nor (n803,n804,n805);
and (n804,n60,n88);
and (n805,n56,n90);
or (n806,n48,n661);
and (n807,n777,n793);
or (n808,n809,n831);
and (n809,n810,n825);
xor (n810,n811,n818);
nand (n811,n812,n813);
or (n812,n278,n741);
nand (n813,n814,n261);
not (n814,n815);
nor (n815,n816,n817);
and (n816,n264,n195);
and (n817,n265,n197);
nand (n818,n819,n824);
or (n819,n820,n344);
not (n820,n821);
nand (n821,n822,n823);
or (n822,n190,n219);
or (n823,n192,n217);
nand (n824,n346,n341);
nand (n825,n826,n830);
or (n826,n155,n827);
nor (n827,n828,n829);
and (n828,n77,n243);
and (n829,n78,n245);
or (n830,n156,n331);
and (n831,n811,n818);
or (n832,n833,n853);
and (n833,n834,n847);
xor (n834,n835,n841);
nand (n835,n836,n840);
or (n836,n179,n837);
nor (n837,n838,n839);
and (n838,n187,n118);
and (n839,n185,n120);
or (n840,n188,n361);
nand (n841,n842,n846);
or (n842,n206,n843);
nor (n843,n844,n845);
and (n844,n144,n113);
and (n845,n114,n146);
or (n846,n207,n385);
nand (n847,n848,n852);
or (n848,n313,n849);
nor (n849,n850,n851);
and (n850,n36,n166);
and (n851,n37,n168);
or (n852,n318,n314);
and (n853,n835,n841);
and (n854,n774,n808);
xor (n855,n325,n405);
and (n856,n736,n771);
xor (n857,n254,n454);
and (n858,n732,n733);
or (n859,n860,n1027);
and (n860,n861,n900);
xor (n861,n862,n863);
xor (n862,n591,n678);
or (n863,n864,n899);
and (n864,n865,n898);
xor (n865,n866,n897);
or (n866,n867,n896);
and (n867,n868,n895);
xor (n868,n869,n894);
or (n869,n870,n893);
and (n870,n871,n885);
xor (n871,n872,n879);
nand (n872,n873,n877);
or (n873,n874,n228);
nor (n874,n875,n876);
and (n875,n240,n274);
and (n876,n238,n276);
nand (n877,n878,n230);
not (n878,n430);
nand (n879,n880,n884);
or (n880,n529,n881);
nor (n881,n882,n883);
and (n882,n302,n294);
and (n883,n290,n304);
or (n884,n530,n655);
nand (n885,n886,n892);
or (n886,n286,n887);
nor (n887,n888,n890);
and (n888,n889,n297);
and (n890,n891,n298);
not (n891,n889);
or (n892,n288,n668);
and (n893,n872,n879);
xor (n894,n652,n666);
xor (n895,n328,n359);
and (n896,n869,n894);
xor (n897,n649,n676);
xor (n898,n680,n683);
and (n899,n866,n897);
or (n900,n901,n1026);
and (n901,n902,n911);
xor (n902,n903,n910);
or (n903,n904,n909);
and (n904,n905,n908);
xor (n905,n906,n907);
xor (n906,n407,n439);
xor (n907,n371,n392);
xor (n908,n738,n746);
and (n909,n906,n907);
xor (n910,n735,n855);
or (n911,n912,n1025);
and (n912,n913,n973);
xor (n913,n914,n972);
or (n914,n915,n971);
and (n915,n916,n949);
xor (n916,n917,n925);
not (n917,n918);
nor (n918,n919,n924);
and (n919,n785,n920);
not (n920,n921);
nor (n921,n922,n923);
and (n922,n417,n67);
and (n923,n415,n69);
and (n924,n779,n790);
or (n925,n926,n948);
and (n926,n927,n942);
xor (n927,n928,n935);
nand (n928,n929,n934);
or (n929,n930,n410);
not (n930,n931);
nand (n931,n932,n933);
or (n932,n32,n174);
or (n933,n31,n172);
nand (n934,n619,n796);
nand (n935,n936,n941);
or (n936,n937,n47);
not (n937,n938);
nand (n938,n939,n940);
or (n939,n56,n251);
or (n940,n60,n249);
or (n941,n48,n803);
nand (n942,n943,n947);
or (n943,n260,n944);
nor (n944,n945,n946);
and (n945,n264,n223);
and (n946,n265,n225);
or (n947,n278,n815);
and (n948,n928,n935);
or (n949,n950,n970);
and (n950,n951,n964);
xor (n951,n952,n958);
nand (n952,n953,n957);
or (n953,n954,n344);
nor (n954,n955,n956);
and (n955,n192,n124);
and (n956,n190,n126);
nand (n957,n346,n821);
nand (n958,n959,n963);
or (n959,n155,n960);
nor (n960,n961,n962);
and (n961,n77,n377);
and (n962,n78,n376);
or (n963,n156,n827);
nand (n964,n965,n969);
or (n965,n179,n966);
nor (n966,n967,n968);
and (n967,n187,n150);
and (n968,n185,n152);
or (n969,n188,n837);
and (n970,n952,n958);
and (n971,n917,n925);
xor (n972,n773,n832);
or (n973,n974,n1024);
and (n974,n975,n1023);
xor (n975,n976,n999);
or (n976,n977,n998);
and (n977,n978,n992);
xor (n978,n979,n985);
nand (n979,n980,n984);
or (n980,n206,n981);
nor (n981,n982,n983);
and (n982,n398,n113);
and (n983,n114,n397);
or (n984,n843,n207);
nand (n985,n986,n990);
or (n986,n987,n313);
nor (n987,n988,n989);
and (n988,n97,n37);
and (n989,n95,n36);
nand (n990,n991,n28);
not (n991,n849);
nand (n992,n993,n997);
or (n993,n72,n994);
nor (n994,n995,n996);
and (n995,n82,n281);
and (n996,n83,n283);
or (n997,n92,n751);
and (n998,n979,n985);
or (n999,n1000,n1022);
and (n1000,n1001,n1016);
xor (n1001,n1002,n1008);
nand (n1002,n1003,n1004);
or (n1003,n127,n757);
or (n1004,n102,n1005);
nor (n1005,n1006,n1007);
and (n1006,n110,n443);
and (n1007,n106,n445);
nand (n1008,n1009,n1014);
or (n1009,n1010,n130);
not (n1010,n1011);
nand (n1011,n1012,n1013);
or (n1012,n310,n140);
or (n1013,n139,n308);
nand (n1014,n765,n1015);
not (n1015,n132);
nand (n1016,n1017,n1021);
or (n1017,n228,n1018);
nor (n1018,n1019,n1020);
and (n1019,n240,n201);
and (n1020,n238,n203);
or (n1021,n229,n874);
and (n1022,n1002,n1008);
xor (n1023,n810,n825);
and (n1024,n976,n999);
and (n1025,n914,n972);
and (n1026,n903,n910);
and (n1027,n862,n863);
or (n1028,n1029,n1144);
and (n1029,n1030,n1033);
xor (n1030,n1031,n1032);
xor (n1031,n731,n857);
xor (n1032,n861,n900);
or (n1033,n1034,n1143);
and (n1034,n1035,n1142);
xor (n1035,n1036,n1141);
or (n1036,n1037,n1140);
and (n1037,n1038,n1047);
xor (n1038,n1039,n1046);
or (n1039,n1040,n1045);
and (n1040,n1041,n1044);
xor (n1041,n1042,n1043);
xor (n1042,n871,n885);
xor (n1043,n776,n801);
xor (n1044,n748,n762);
and (n1045,n1042,n1043);
xor (n1046,n868,n895);
or (n1047,n1048,n1139);
and (n1048,n1049,n1069);
xor (n1049,n1050,n1051);
xor (n1050,n834,n847);
or (n1051,n1052,n1068);
and (n1052,n1053,n918);
xor (n1053,n1054,n1060);
nand (n1054,n1055,n1059);
or (n1055,n529,n1056);
nor (n1056,n1057,n1058);
and (n1057,n670,n294);
and (n1058,n672,n290);
or (n1059,n530,n881);
nand (n1060,n1061,n1067);
or (n1061,n286,n1062);
nor (n1062,n1063,n1065);
and (n1063,n1064,n297);
and (n1065,n298,n1066);
not (n1066,n1064);
or (n1067,n288,n887);
and (n1068,n1054,n1060);
or (n1069,n1070,n1138);
and (n1070,n1071,n1114);
xor (n1071,n1072,n1090);
or (n1072,n1073,n1081);
nand (n1073,n1074,n1079);
or (n1074,n1075,n1076);
not (n1075,n785);
nor (n1076,n1077,n1078);
and (n1077,n63,n415);
and (n1078,n61,n417);
or (n1079,n1080,n921);
not (n1080,n779);
nand (n1081,n1082,n1087);
or (n1082,n1083,n1086);
not (n1083,n1084);
nand (n1084,n783,n1085);
not (n1085,n1086);
nor (n1087,n1088,n1089);
and (n1088,n43,n783);
and (n1089,n42,n782);
or (n1090,n1091,n1113);
and (n1091,n1092,n1107);
xor (n1092,n1093,n1099);
nand (n1093,n1094,n1098);
or (n1094,n313,n1095);
nor (n1095,n1096,n1097);
and (n1096,n90,n37);
and (n1097,n88,n36);
or (n1098,n318,n987);
nand (n1099,n1100,n1106);
or (n1100,n286,n1101);
nor (n1101,n1102,n1104);
and (n1102,n1103,n297);
and (n1104,n298,n1105);
not (n1105,n1103);
or (n1106,n1062,n288);
nand (n1107,n1108,n1112);
or (n1108,n228,n1109);
nor (n1109,n1110,n1111);
and (n1110,n240,n195);
and (n1111,n238,n197);
or (n1112,n229,n1018);
and (n1113,n1093,n1099);
or (n1114,n1115,n1137);
and (n1115,n1116,n1131);
xor (n1116,n1117,n1123);
nand (n1117,n1118,n1122);
or (n1118,n260,n1119);
nor (n1119,n1120,n1121);
and (n1120,n264,n217);
and (n1121,n265,n219);
or (n1122,n278,n944);
nand (n1123,n1124,n1125);
or (n1124,n937,n48);
nand (n1125,n1126,n1130);
not (n1126,n1127);
nor (n1127,n1128,n1129);
and (n1128,n60,n243);
and (n1129,n56,n245);
not (n1130,n47);
nand (n1131,n1132,n1136);
or (n1132,n344,n1133);
nor (n1133,n1134,n1135);
and (n1134,n192,n118);
and (n1135,n190,n120);
or (n1136,n470,n954);
and (n1137,n1117,n1123);
and (n1138,n1072,n1090);
and (n1139,n1050,n1051);
and (n1140,n1039,n1046);
xor (n1141,n865,n898);
xor (n1142,n902,n911);
and (n1143,n1036,n1141);
and (n1144,n1031,n1032);
nand (n1145,n17,n1028);
not (n1146,n1147);
nand (n1147,n1148,n4386);
or (n1148,n1149,n1587);
not (n1149,n1150);
nor (n1150,n1151,n1582);
nor (n1151,n1152,n1235);
xor (n1152,n1153,n1216);
xor (n1153,n1154,n1215);
or (n1154,n1155,n1214);
and (n1155,n1156,n1213);
xor (n1156,n1157,n1158);
xor (n1157,n905,n908);
or (n1158,n1159,n1212);
and (n1159,n1160,n1163);
xor (n1160,n1161,n1162);
xor (n1161,n916,n949);
xor (n1162,n975,n1023);
or (n1163,n1164,n1211);
and (n1164,n1165,n1210);
xor (n1165,n1166,n1188);
or (n1166,n1167,n1187);
and (n1167,n1168,n1181);
xor (n1168,n1169,n1175);
nand (n1169,n1170,n1174);
or (n1170,n1171,n179);
nor (n1171,n1172,n1173);
and (n1172,n146,n185);
and (n1173,n144,n187);
or (n1174,n188,n966);
nand (n1175,n1176,n1180);
or (n1176,n1177,n410);
nor (n1177,n1178,n1179);
and (n1178,n31,n166);
and (n1179,n32,n168);
nand (n1180,n619,n931);
nand (n1181,n1182,n1186);
or (n1182,n155,n1183);
nor (n1183,n1184,n1185);
and (n1184,n77,n436);
and (n1185,n78,n438);
or (n1186,n156,n960);
and (n1187,n1169,n1175);
or (n1188,n1189,n1209);
and (n1189,n1190,n1203);
xor (n1190,n1191,n1197);
nand (n1191,n1192,n1196);
or (n1192,n206,n1193);
nor (n1193,n1194,n1195);
and (n1194,n113,n449);
and (n1195,n114,n451);
or (n1196,n207,n981);
nand (n1197,n1198,n1202);
or (n1198,n102,n1199);
nor (n1199,n1200,n1201);
and (n1200,n110,n551);
and (n1201,n106,n553);
or (n1202,n127,n1005);
nand (n1203,n1204,n1205);
or (n1204,n994,n92);
or (n1205,n72,n1206);
nor (n1206,n1207,n1208);
and (n1207,n82,n274);
and (n1208,n83,n276);
and (n1209,n1191,n1197);
xor (n1210,n927,n942);
and (n1211,n1166,n1188);
and (n1212,n1161,n1162);
xor (n1213,n913,n973);
and (n1214,n1157,n1158);
xor (n1215,n1035,n1142);
or (n1216,n1217,n1234);
and (n1217,n1218,n1233);
xor (n1218,n1219,n1220);
xor (n1219,n1038,n1047);
or (n1220,n1221,n1232);
and (n1221,n1222,n1231);
xor (n1222,n1223,n1230);
or (n1223,n1224,n1229);
and (n1224,n1225,n1228);
xor (n1225,n1226,n1227);
xor (n1226,n1001,n1016);
xor (n1227,n951,n964);
xor (n1228,n978,n992);
and (n1229,n1226,n1227);
xor (n1230,n1041,n1044);
xor (n1231,n1049,n1069);
and (n1232,n1223,n1230);
xor (n1233,n1156,n1213);
and (n1234,n1219,n1220);
or (n1235,n1236,n1581);
and (n1236,n1237,n1418);
xor (n1237,n1238,n1417);
or (n1238,n1239,n1416);
and (n1239,n1240,n1415);
xor (n1240,n1241,n1353);
or (n1241,n1242,n1352);
and (n1242,n1243,n1278);
xor (n1243,n1244,n1245);
xor (n1244,n1053,n918);
or (n1245,n1246,n1277);
and (n1246,n1247,n1260);
xor (n1247,n1248,n1254);
nand (n1248,n1249,n1253);
or (n1249,n130,n1250);
nor (n1250,n1251,n1252);
and (n1251,n139,n302);
and (n1252,n140,n304);
or (n1253,n132,n1010);
nand (n1254,n1255,n1259);
or (n1255,n529,n1256);
nor (n1256,n1257,n1258);
and (n1257,n889,n294);
and (n1258,n891,n290);
or (n1259,n530,n1056);
and (n1260,n1261,n1269);
nor (n1261,n1262,n297);
nor (n1262,n1263,n1267);
and (n1263,n1264,n294);
not (n1264,n1265);
and (n1265,n1266,n292);
and (n1267,n1268,n291);
not (n1268,n1266);
nand (n1269,n1270,n1272);
or (n1270,n1085,n1271);
not (n1271,n1087);
or (n1272,n1084,n1273);
not (n1273,n1274);
nand (n1274,n1275,n1276);
or (n1275,n67,n782);
nand (n1276,n782,n67);
and (n1277,n1248,n1254);
or (n1278,n1279,n1351);
and (n1279,n1280,n1329);
xor (n1280,n1281,n1307);
or (n1281,n1282,n1306);
and (n1282,n1283,n1300);
xor (n1283,n1284,n1292);
nand (n1284,n1285,n1290);
or (n1285,n1286,n1075);
not (n1286,n1287);
nor (n1287,n1288,n1289);
and (n1288,n172,n415);
and (n1289,n174,n417);
nand (n1290,n1291,n779);
not (n1291,n1076);
nand (n1292,n1293,n1298);
or (n1293,n1294,n313);
not (n1294,n1295);
nand (n1295,n1296,n1297);
or (n1296,n37,n251);
or (n1297,n36,n249);
nand (n1298,n1299,n28);
not (n1299,n1095);
nand (n1300,n1301,n1305);
or (n1301,n286,n1302);
nor (n1302,n1303,n1304);
and (n1303,n1268,n298);
and (n1304,n1266,n297);
or (n1305,n288,n1101);
and (n1306,n1284,n1292);
or (n1307,n1308,n1328);
and (n1308,n1309,n1322);
xor (n1309,n1310,n1316);
nand (n1310,n1311,n1315);
or (n1311,n228,n1312);
nor (n1312,n1313,n1314);
and (n1313,n223,n240);
and (n1314,n225,n238);
or (n1315,n229,n1109);
nand (n1316,n1317,n1321);
or (n1317,n260,n1318);
nor (n1318,n1319,n1320);
and (n1319,n264,n124);
and (n1320,n265,n126);
or (n1321,n278,n1119);
nand (n1322,n1323,n1327);
or (n1323,n47,n1324);
nor (n1324,n1325,n1326);
and (n1325,n376,n56);
and (n1326,n377,n60);
or (n1327,n48,n1127);
and (n1328,n1310,n1316);
or (n1329,n1330,n1350);
and (n1330,n1331,n1344);
xor (n1331,n1332,n1338);
nand (n1332,n1333,n1337);
or (n1333,n344,n1334);
nor (n1334,n1335,n1336);
and (n1335,n152,n190);
and (n1336,n150,n192);
or (n1337,n470,n1133);
nand (n1338,n1339,n1343);
or (n1339,n179,n1340);
nor (n1340,n1341,n1342);
and (n1341,n187,n398);
and (n1342,n185,n397);
or (n1343,n188,n1171);
nand (n1344,n1345,n1349);
or (n1345,n410,n1346);
nor (n1346,n1347,n1348);
and (n1347,n31,n95);
and (n1348,n32,n97);
or (n1349,n411,n1177);
and (n1350,n1332,n1338);
and (n1351,n1281,n1307);
and (n1352,n1244,n1245);
or (n1353,n1354,n1414);
and (n1354,n1355,n1413);
xor (n1355,n1356,n1412);
or (n1356,n1357,n1411);
and (n1357,n1358,n1407);
xor (n1358,n1359,n1383);
or (n1359,n1360,n1382);
and (n1360,n1361,n1376);
xor (n1361,n1362,n1370);
nand (n1362,n1363,n1367);
or (n1363,n1364,n155);
nor (n1364,n1365,n1366);
and (n1365,n283,n78);
and (n1366,n281,n77);
nand (n1367,n1368,n1369);
not (n1368,n1183);
not (n1369,n156);
nand (n1370,n1371,n1375);
or (n1371,n206,n1372);
nor (n1372,n1373,n1374);
and (n1373,n113,n443);
and (n1374,n114,n445);
or (n1375,n207,n1193);
nand (n1376,n1377,n1381);
or (n1377,n102,n1378);
nor (n1378,n1379,n1380);
and (n1379,n110,n308);
and (n1380,n106,n310);
or (n1381,n127,n1199);
and (n1382,n1362,n1370);
or (n1383,n1384,n1406);
and (n1384,n1385,n1400);
xor (n1385,n1386,n1394);
nand (n1386,n1387,n1392);
or (n1387,n1388,n72);
not (n1388,n1389);
nand (n1389,n1390,n1391);
or (n1390,n83,n203);
or (n1391,n82,n201);
nand (n1392,n1393,n74);
not (n1393,n1206);
nand (n1394,n1395,n1399);
or (n1395,n1396,n130);
nor (n1396,n1397,n1398);
and (n1397,n139,n670);
and (n1398,n140,n672);
or (n1399,n132,n1250);
nand (n1400,n1401,n1405);
or (n1401,n529,n1402);
nor (n1402,n1403,n1404);
and (n1403,n1064,n294);
and (n1404,n1066,n290);
or (n1405,n530,n1256);
and (n1406,n1386,n1394);
nand (n1407,n1408,n1072);
or (n1408,n1409,n1410);
not (n1409,n1081);
not (n1410,n1073);
and (n1411,n1359,n1383);
xor (n1412,n1071,n1114);
xor (n1413,n1165,n1210);
and (n1414,n1356,n1412);
xor (n1415,n1160,n1163);
and (n1416,n1241,n1353);
xor (n1417,n1218,n1233);
or (n1418,n1419,n1580);
and (n1419,n1420,n1435);
xor (n1420,n1421,n1422);
xor (n1421,n1222,n1231);
or (n1422,n1423,n1434);
and (n1423,n1424,n1433);
xor (n1424,n1425,n1432);
or (n1425,n1426,n1431);
and (n1426,n1427,n1430);
xor (n1427,n1428,n1429);
xor (n1428,n1116,n1131);
xor (n1429,n1168,n1181);
xor (n1430,n1190,n1203);
and (n1431,n1428,n1429);
xor (n1432,n1225,n1228);
xor (n1433,n1243,n1278);
and (n1434,n1425,n1432);
or (n1435,n1436,n1579);
and (n1436,n1437,n1578);
xor (n1437,n1438,n1519);
or (n1438,n1439,n1518);
and (n1439,n1440,n1443);
xor (n1440,n1441,n1442);
xor (n1441,n1092,n1107);
xor (n1442,n1247,n1260);
or (n1443,n1444,n1517);
and (n1444,n1445,n1493);
xor (n1445,n1446,n1470);
or (n1446,n1447,n1469);
and (n1447,n1448,n1463);
xor (n1448,n1449,n1457);
nand (n1449,n1450,n1455);
or (n1450,n1451,n47);
not (n1451,n1452);
nor (n1452,n1453,n1454);
and (n1453,n436,n56);
and (n1454,n438,n60);
nand (n1455,n1456,n49);
not (n1456,n1324);
nand (n1457,n1458,n1462);
or (n1458,n344,n1459);
nor (n1459,n1460,n1461);
and (n1460,n192,n144);
and (n1461,n190,n146);
or (n1462,n470,n1334);
nand (n1463,n1464,n1468);
or (n1464,n179,n1465);
nor (n1465,n1466,n1467);
and (n1466,n187,n449);
and (n1467,n185,n451);
or (n1468,n188,n1340);
and (n1469,n1449,n1457);
or (n1470,n1471,n1492);
and (n1471,n1472,n1486);
xor (n1472,n1473,n1480);
nand (n1473,n1474,n1478);
or (n1474,n1475,n410);
nor (n1475,n1476,n1477);
and (n1476,n90,n32);
and (n1477,n88,n31);
nand (n1478,n1479,n619);
not (n1479,n1346);
nand (n1480,n1481,n1485);
or (n1481,n155,n1482);
nor (n1482,n1483,n1484);
and (n1483,n77,n274);
and (n1484,n78,n276);
or (n1485,n156,n1364);
nand (n1486,n1487,n1491);
or (n1487,n206,n1488);
nor (n1488,n1489,n1490);
and (n1489,n113,n551);
and (n1490,n114,n553);
or (n1491,n207,n1372);
and (n1492,n1473,n1480);
or (n1493,n1494,n1516);
and (n1494,n1495,n1510);
xor (n1495,n1496,n1503);
nand (n1496,n1497,n1502);
or (n1497,n1498,n102);
not (n1498,n1499);
nand (n1499,n1500,n1501);
or (n1500,n106,n304);
or (n1501,n110,n302);
or (n1502,n127,n1378);
nand (n1503,n1504,n1509);
or (n1504,n1505,n72);
not (n1505,n1506);
nand (n1506,n1507,n1508);
or (n1507,n83,n197);
or (n1508,n82,n195);
nand (n1509,n74,n1389);
nand (n1510,n1511,n1515);
or (n1511,n130,n1512);
nor (n1512,n1513,n1514);
and (n1513,n139,n889);
and (n1514,n140,n891);
or (n1515,n132,n1396);
and (n1516,n1496,n1503);
and (n1517,n1446,n1470);
and (n1518,n1441,n1442);
or (n1519,n1520,n1577);
and (n1520,n1521,n1576);
xor (n1521,n1522,n1569);
or (n1522,n1523,n1568);
and (n1523,n1524,n1545);
xor (n1524,n1525,n1526);
xor (n1525,n1261,n1269);
or (n1526,n1527,n1544);
and (n1527,n1528,n1537);
xor (n1528,n1529,n1530);
nor (n1529,n288,n1268);
nand (n1530,n1531,n1536);
or (n1531,n1084,n1532);
not (n1532,n1533);
nor (n1533,n1534,n1535);
and (n1534,n63,n782);
and (n1535,n61,n783);
nand (n1536,n1274,n1086);
nand (n1537,n1538,n1543);
or (n1538,n1539,n1075);
not (n1539,n1540);
nand (n1540,n1541,n1542);
or (n1541,n415,n168);
or (n1542,n417,n166);
nand (n1543,n779,n1287);
and (n1544,n1529,n1530);
or (n1545,n1546,n1567);
and (n1546,n1547,n1561);
xor (n1547,n1548,n1555);
nand (n1548,n1549,n1554);
or (n1549,n1550,n313);
not (n1550,n1551);
nand (n1551,n1552,n1553);
or (n1552,n37,n245);
or (n1553,n36,n243);
nand (n1554,n28,n1295);
nand (n1555,n1556,n1560);
or (n1556,n228,n1557);
nor (n1557,n1558,n1559);
and (n1558,n240,n217);
and (n1559,n238,n219);
or (n1560,n229,n1312);
nand (n1561,n1562,n1566);
or (n1562,n260,n1563);
nor (n1563,n1564,n1565);
and (n1564,n264,n118);
and (n1565,n265,n120);
or (n1566,n278,n1318);
and (n1567,n1548,n1555);
and (n1568,n1525,n1526);
or (n1569,n1570,n1575);
and (n1570,n1571,n1574);
xor (n1571,n1572,n1573);
xor (n1572,n1385,n1400);
xor (n1573,n1283,n1300);
xor (n1574,n1309,n1322);
and (n1575,n1572,n1573);
xor (n1576,n1358,n1407);
and (n1577,n1522,n1569);
xor (n1578,n1355,n1413);
and (n1579,n1438,n1519);
and (n1580,n1421,n1422);
and (n1581,n1238,n1417);
nor (n1582,n1583,n1584);
xor (n1583,n1030,n1033);
or (n1584,n1585,n1586);
and (n1585,n1153,n1216);
and (n1586,n1154,n1215);
not (n1587,n1588);
nand (n1588,n1589,n4371);
or (n1589,n1590,n2228);
nand (n1590,n1591,n1798);
nor (n1591,n1592,n1783);
nor (n1592,n1593,n1594);
xor (n1593,n1237,n1418);
or (n1594,n1595,n1782);
and (n1595,n1596,n1599);
xor (n1596,n1597,n1598);
xor (n1597,n1240,n1415);
xor (n1598,n1420,n1435);
or (n1599,n1600,n1781);
and (n1600,n1601,n1690);
xor (n1601,n1602,n1603);
xor (n1602,n1424,n1433);
or (n1603,n1604,n1689);
and (n1604,n1605,n1608);
xor (n1605,n1606,n1607);
xor (n1606,n1280,n1329);
xor (n1607,n1427,n1430);
or (n1608,n1609,n1688);
and (n1609,n1610,n1613);
xor (n1610,n1611,n1612);
xor (n1611,n1331,n1344);
xor (n1612,n1361,n1376);
or (n1613,n1614,n1687);
and (n1614,n1615,n1664);
xor (n1615,n1616,n1639);
or (n1616,n1617,n1638);
and (n1617,n1618,n1631);
xor (n1618,n1619,n1625);
nand (n1619,n1620,n1624);
or (n1620,n260,n1621);
nor (n1621,n1622,n1623);
and (n1622,n264,n150);
and (n1623,n265,n152);
or (n1624,n278,n1563);
nand (n1625,n1626,n1630);
or (n1626,n47,n1627);
nor (n1627,n1628,n1629);
and (n1628,n60,n281);
and (n1629,n56,n283);
or (n1630,n48,n1451);
nand (n1631,n1632,n1637);
or (n1632,n344,n1633);
not (n1633,n1634);
nor (n1634,n1635,n1636);
and (n1635,n398,n190);
and (n1636,n397,n192);
or (n1637,n470,n1459);
and (n1638,n1619,n1625);
or (n1639,n1640,n1663);
and (n1640,n1641,n1657);
xor (n1641,n1642,n1651);
nand (n1642,n1643,n1648);
or (n1643,n1644,n179);
not (n1644,n1645);
nand (n1645,n1646,n1647);
or (n1646,n185,n445);
or (n1647,n187,n443);
nand (n1648,n1649,n1650);
not (n1649,n1465);
not (n1650,n188);
nand (n1651,n1652,n1656);
or (n1652,n410,n1653);
nor (n1653,n1654,n1655);
and (n1654,n31,n249);
and (n1655,n32,n251);
or (n1656,n411,n1475);
nand (n1657,n1658,n1662);
or (n1658,n155,n1659);
nor (n1659,n1660,n1661);
and (n1660,n77,n201);
and (n1661,n78,n203);
or (n1662,n156,n1482);
and (n1663,n1642,n1651);
or (n1664,n1665,n1686);
and (n1665,n1666,n1680);
xor (n1666,n1667,n1673);
nand (n1667,n1668,n1672);
or (n1668,n206,n1669);
nor (n1669,n1670,n1671);
and (n1670,n113,n308);
and (n1671,n114,n310);
or (n1672,n207,n1488);
nand (n1673,n1674,n1675);
or (n1674,n1498,n127);
nand (n1675,n1676,n103);
not (n1676,n1677);
nor (n1677,n1678,n1679);
and (n1678,n110,n670);
and (n1679,n672,n106);
nand (n1680,n1681,n1685);
or (n1681,n1682,n72);
nor (n1682,n1683,n1684);
and (n1683,n82,n223);
and (n1684,n83,n225);
or (n1685,n92,n1505);
and (n1686,n1667,n1673);
and (n1687,n1616,n1639);
and (n1688,n1611,n1612);
and (n1689,n1606,n1607);
or (n1690,n1691,n1780);
and (n1691,n1692,n1745);
xor (n1692,n1693,n1694);
xor (n1693,n1440,n1443);
or (n1694,n1695,n1744);
and (n1695,n1696,n1743);
xor (n1696,n1697,n1742);
or (n1697,n1698,n1741);
and (n1698,n1699,n1719);
xor (n1699,n1700,n1706);
nand (n1700,n1701,n1705);
or (n1701,n529,n1702);
nor (n1702,n1703,n1704);
and (n1703,n294,n1103);
and (n1704,n1105,n290);
or (n1705,n530,n1402);
and (n1706,n1707,n1713);
nor (n1707,n1708,n294);
nor (n1708,n1709,n1712);
and (n1709,n1710,n139);
not (n1710,n1711);
and (n1711,n1266,n533);
and (n1712,n1268,n537);
nand (n1713,n1714,n1715);
or (n1714,n1085,n1532);
or (n1715,n1084,n1716);
nor (n1716,n1717,n1718);
and (n1717,n782,n172);
and (n1718,n783,n174);
or (n1719,n1720,n1740);
and (n1720,n1721,n1734);
xor (n1721,n1722,n1728);
nand (n1722,n1723,n1724);
or (n1723,n1539,n1080);
or (n1724,n1075,n1725);
nor (n1725,n1726,n1727);
and (n1726,n97,n415);
and (n1727,n95,n417);
nand (n1728,n1729,n1730);
or (n1729,n1550,n318);
or (n1730,n313,n1731);
nor (n1731,n1732,n1733);
and (n1732,n36,n377);
and (n1733,n37,n376);
nand (n1734,n1735,n1739);
or (n1735,n228,n1736);
nor (n1736,n1737,n1738);
and (n1737,n240,n124);
and (n1738,n238,n126);
or (n1739,n229,n1557);
and (n1740,n1722,n1728);
and (n1741,n1700,n1706);
xor (n1742,n1445,n1493);
xor (n1743,n1524,n1545);
and (n1744,n1697,n1742);
or (n1745,n1746,n1779);
and (n1746,n1747,n1778);
xor (n1747,n1748,n1755);
or (n1748,n1749,n1754);
and (n1749,n1750,n1753);
xor (n1750,n1751,n1752);
xor (n1751,n1528,n1537);
xor (n1752,n1495,n1510);
xor (n1753,n1472,n1486);
and (n1754,n1751,n1752);
or (n1755,n1756,n1777);
and (n1756,n1757,n1760);
xor (n1757,n1758,n1759);
xor (n1758,n1448,n1463);
xor (n1759,n1547,n1561);
or (n1760,n1761,n1776);
and (n1761,n1762,n1775);
xor (n1762,n1763,n1769);
nand (n1763,n1764,n1768);
or (n1764,n130,n1765);
nor (n1765,n1766,n1767);
and (n1766,n139,n1064);
and (n1767,n140,n1066);
or (n1768,n132,n1512);
nand (n1769,n1770,n1774);
or (n1770,n529,n1771);
nor (n1771,n1772,n1773);
and (n1772,n1268,n290);
and (n1773,n1266,n294);
or (n1774,n530,n1702);
xor (n1775,n1707,n1713);
and (n1776,n1763,n1769);
and (n1777,n1758,n1759);
xor (n1778,n1571,n1574);
and (n1779,n1748,n1755);
and (n1780,n1693,n1694);
and (n1781,n1602,n1603);
and (n1782,n1597,n1598);
nor (n1783,n1784,n1797);
or (n1784,n1785,n1796);
and (n1785,n1786,n1789);
xor (n1786,n1787,n1788);
xor (n1787,n1437,n1578);
xor (n1788,n1601,n1690);
or (n1789,n1790,n1795);
and (n1790,n1791,n1794);
xor (n1791,n1792,n1793);
xor (n1792,n1521,n1576);
xor (n1793,n1605,n1608);
xor (n1794,n1692,n1745);
and (n1795,n1792,n1793);
and (n1796,n1787,n1788);
xor (n1797,n1596,n1599);
nor (n1798,n1799,n2091);
nor (n1799,n1800,n1801);
xor (n1800,n1786,n1789);
or (n1801,n1802,n2090);
and (n1802,n1803,n2089);
xor (n1803,n1804,n1946);
or (n1804,n1805,n1945);
and (n1805,n1806,n1889);
xor (n1806,n1807,n1808);
xor (n1807,n1610,n1613);
or (n1808,n1809,n1888);
and (n1809,n1810,n1881);
xor (n1810,n1811,n1812);
xor (n1811,n1699,n1719);
or (n1812,n1813,n1880);
and (n1813,n1814,n1857);
xor (n1814,n1815,n1838);
or (n1815,n1816,n1837);
and (n1816,n1817,n1831);
xor (n1817,n1818,n1825);
nand (n1818,n1819,n1824);
or (n1819,n1820,n344);
not (n1820,n1821);
nor (n1821,n1822,n1823);
and (n1822,n449,n190);
and (n1823,n451,n192);
nand (n1824,n1634,n346);
nand (n1825,n1826,n1830);
or (n1826,n1827,n179);
nor (n1827,n1828,n1829);
and (n1828,n553,n185);
and (n1829,n551,n187);
nand (n1830,n1645,n1650);
nand (n1831,n1832,n1836);
or (n1832,n1084,n1833);
nor (n1833,n1834,n1835);
and (n1834,n782,n166);
and (n1835,n783,n168);
or (n1836,n1716,n1085);
and (n1837,n1818,n1825);
or (n1838,n1839,n1856);
and (n1839,n1840,n1850);
xor (n1840,n1841,n1842);
nor (n1841,n530,n1268);
nand (n1842,n1843,n1848);
or (n1843,n1844,n1075);
not (n1844,n1845);
nand (n1845,n1846,n1847);
or (n1846,n415,n90);
or (n1847,n417,n88);
nand (n1848,n1849,n779);
not (n1849,n1725);
nand (n1850,n1851,n1855);
or (n1851,n313,n1852);
nor (n1852,n1853,n1854);
and (n1853,n36,n436);
and (n1854,n37,n438);
or (n1855,n318,n1731);
and (n1856,n1841,n1842);
or (n1857,n1858,n1879);
and (n1858,n1859,n1873);
xor (n1859,n1860,n1867);
nand (n1860,n1861,n1865);
or (n1861,n1862,n228);
nor (n1862,n1863,n1864);
and (n1863,n118,n240);
and (n1864,n120,n238);
nand (n1865,n1866,n230);
not (n1866,n1736);
nand (n1867,n1868,n1872);
or (n1868,n260,n1869);
nor (n1869,n1870,n1871);
and (n1870,n264,n144);
and (n1871,n265,n146);
or (n1872,n278,n1621);
nand (n1873,n1874,n1878);
or (n1874,n47,n1875);
nor (n1875,n1876,n1877);
and (n1876,n60,n274);
and (n1877,n56,n276);
or (n1878,n48,n1627);
and (n1879,n1860,n1867);
and (n1880,n1815,n1838);
or (n1881,n1882,n1887);
and (n1882,n1883,n1886);
xor (n1883,n1884,n1885);
xor (n1884,n1666,n1680);
xor (n1885,n1618,n1631);
xor (n1886,n1641,n1657);
and (n1887,n1884,n1885);
and (n1888,n1811,n1812);
or (n1889,n1890,n1944);
and (n1890,n1891,n1943);
xor (n1891,n1892,n1893);
xor (n1892,n1615,n1664);
or (n1893,n1894,n1942);
and (n1894,n1895,n1941);
xor (n1895,n1896,n1919);
or (n1896,n1897,n1918);
and (n1897,n1898,n1912);
xor (n1898,n1899,n1906);
nand (n1899,n1900,n1905);
or (n1900,n1901,n155);
not (n1901,n1902);
nor (n1902,n1903,n1904);
and (n1903,n195,n78);
and (n1904,n197,n77);
or (n1905,n156,n1659);
nand (n1906,n1907,n1911);
or (n1907,n206,n1908);
nor (n1908,n1909,n1910);
and (n1909,n113,n302);
and (n1910,n114,n304);
or (n1911,n207,n1669);
nand (n1912,n1913,n1917);
or (n1913,n102,n1914);
nor (n1914,n1915,n1916);
and (n1915,n889,n110);
and (n1916,n106,n891);
or (n1917,n1677,n127);
and (n1918,n1899,n1906);
or (n1919,n1920,n1940);
and (n1920,n1921,n1934);
xor (n1921,n1922,n1928);
nand (n1922,n1923,n1927);
or (n1923,n410,n1924);
nor (n1924,n1925,n1926);
and (n1925,n245,n32);
and (n1926,n243,n31);
or (n1927,n411,n1653);
nand (n1928,n1929,n1933);
or (n1929,n130,n1930);
nor (n1930,n1931,n1932);
and (n1931,n1103,n139);
and (n1932,n140,n1105);
or (n1933,n132,n1765);
nand (n1934,n1935,n1939);
or (n1935,n72,n1936);
nor (n1936,n1937,n1938);
and (n1937,n82,n217);
and (n1938,n83,n219);
or (n1939,n92,n1682);
and (n1940,n1922,n1928);
xor (n1941,n1721,n1734);
and (n1942,n1896,n1919);
xor (n1943,n1757,n1760);
and (n1944,n1892,n1893);
and (n1945,n1807,n1808);
or (n1946,n1947,n2088);
and (n1947,n1948,n1951);
xor (n1948,n1949,n1950);
xor (n1949,n1696,n1743);
xor (n1950,n1747,n1778);
or (n1951,n1952,n2087);
and (n1952,n1953,n2010);
xor (n1953,n1954,n1955);
xor (n1954,n1750,n1753);
or (n1955,n1956,n2009);
and (n1956,n1957,n2008);
xor (n1957,n1958,n1959);
xor (n1958,n1814,n1857);
or (n1959,n1960,n2007);
and (n1960,n1961,n2006);
xor (n1961,n1962,n1984);
or (n1962,n1963,n1983);
and (n1963,n1964,n1977);
xor (n1964,n1965,n1971);
nand (n1965,n1966,n1970);
or (n1966,n102,n1967);
nor (n1967,n1968,n1969);
and (n1968,n1066,n106);
and (n1969,n1064,n110);
or (n1970,n1914,n127);
nand (n1971,n1972,n1976);
or (n1972,n410,n1973);
nor (n1973,n1974,n1975);
and (n1974,n31,n377);
and (n1975,n32,n376);
or (n1976,n411,n1924);
nand (n1977,n1978,n1982);
or (n1978,n130,n1979);
nor (n1979,n1980,n1981);
and (n1980,n1268,n140);
and (n1981,n1266,n139);
or (n1982,n1930,n132);
and (n1983,n1965,n1971);
or (n1984,n1985,n2005);
and (n1985,n1986,n1999);
xor (n1986,n1987,n1993);
nand (n1987,n1988,n1992);
or (n1988,n1084,n1989);
nor (n1989,n1990,n1991);
and (n1990,n97,n783);
and (n1991,n95,n782);
or (n1992,n1833,n1085);
nand (n1993,n1994,n1998);
or (n1994,n1995,n155);
nor (n1995,n1996,n1997);
and (n1996,n77,n223);
and (n1997,n78,n225);
nand (n1998,n1369,n1902);
nand (n1999,n2000,n2004);
or (n2000,n206,n2001);
nor (n2001,n2002,n2003);
and (n2002,n113,n670);
and (n2003,n114,n672);
or (n2004,n207,n1908);
and (n2005,n1987,n1993);
xor (n2006,n1859,n1873);
and (n2007,n1962,n1984);
xor (n2008,n1895,n1941);
and (n2009,n1958,n1959);
or (n2010,n2011,n2086);
and (n2011,n2012,n2079);
xor (n2012,n2013,n2014);
xor (n2013,n1762,n1775);
or (n2014,n2015,n2078);
and (n2015,n2016,n2054);
xor (n2016,n2017,n2031);
and (n2017,n2018,n2024);
nand (n2018,n2019,n2023);
or (n2019,n2020,n1075);
nor (n2020,n2021,n2022);
and (n2021,n417,n249);
and (n2022,n415,n251);
nand (n2023,n779,n1845);
not (n2024,n2025);
nand (n2025,n2026,n140);
nand (n2026,n2027,n2028);
or (n2027,n1266,n134);
nand (n2028,n2029,n110);
not (n2029,n2030);
and (n2030,n1266,n134);
or (n2031,n2032,n2053);
and (n2032,n2033,n2047);
xor (n2033,n2034,n2041);
nand (n2034,n2035,n2039);
or (n2035,n2036,n313);
nor (n2036,n2037,n2038);
and (n2037,n36,n281);
and (n2038,n37,n283);
nand (n2039,n2040,n28);
not (n2040,n1852);
nand (n2041,n2042,n2046);
or (n2042,n228,n2043);
nor (n2043,n2044,n2045);
and (n2044,n240,n150);
and (n2045,n238,n152);
or (n2046,n229,n1862);
nand (n2047,n2048,n2052);
or (n2048,n260,n2049);
nor (n2049,n2050,n2051);
and (n2050,n398,n264);
and (n2051,n265,n397);
or (n2052,n278,n1869);
and (n2053,n2034,n2041);
or (n2054,n2055,n2077);
and (n2055,n2056,n2071);
xor (n2056,n2057,n2064);
nand (n2057,n2058,n2062);
or (n2058,n2059,n47);
nor (n2059,n2060,n2061);
and (n2060,n60,n201);
and (n2061,n56,n203);
nand (n2062,n2063,n49);
not (n2063,n1875);
nand (n2064,n2065,n2070);
or (n2065,n2066,n344);
not (n2066,n2067);
nand (n2067,n2068,n2069);
or (n2068,n190,n445);
or (n2069,n192,n443);
nand (n2070,n346,n1821);
nand (n2071,n2072,n2076);
or (n2072,n179,n2073);
nor (n2073,n2074,n2075);
and (n2074,n187,n308);
and (n2075,n185,n310);
or (n2076,n188,n1827);
and (n2077,n2057,n2064);
and (n2078,n2017,n2031);
or (n2079,n2080,n2085);
and (n2080,n2081,n2084);
xor (n2081,n2082,n2083);
xor (n2082,n1921,n1934);
xor (n2083,n1840,n1850);
xor (n2084,n1817,n1831);
and (n2085,n2082,n2083);
and (n2086,n2013,n2014);
and (n2087,n1954,n1955);
and (n2088,n1949,n1950);
xor (n2089,n1791,n1794);
and (n2090,n1804,n1946);
nor (n2091,n2092,n2227);
or (n2092,n2093,n2226);
and (n2093,n2094,n2097);
xor (n2094,n2095,n2096);
xor (n2095,n1806,n1889);
xor (n2096,n1948,n1951);
or (n2097,n2098,n2225);
and (n2098,n2099,n2102);
xor (n2099,n2100,n2101);
xor (n2100,n1810,n1881);
xor (n2101,n1891,n1943);
or (n2102,n2103,n2224);
and (n2103,n2104,n2211);
xor (n2104,n2105,n2106);
xor (n2105,n1883,n1886);
or (n2106,n2107,n2210);
and (n2107,n2108,n2180);
xor (n2108,n2109,n2110);
xor (n2109,n1898,n1912);
or (n2110,n2111,n2179);
and (n2111,n2112,n2157);
xor (n2112,n2113,n2135);
or (n2113,n2114,n2134);
and (n2114,n2115,n2128);
xor (n2115,n2116,n2122);
nand (n2116,n2117,n2121);
or (n2117,n228,n2118);
nor (n2118,n2119,n2120);
and (n2119,n146,n238);
and (n2120,n144,n240);
or (n2121,n2043,n229);
nand (n2122,n2123,n2127);
or (n2123,n260,n2124);
nor (n2124,n2125,n2126);
and (n2125,n449,n264);
and (n2126,n265,n451);
or (n2127,n278,n2049);
nand (n2128,n2129,n2133);
or (n2129,n47,n2130);
nor (n2130,n2131,n2132);
and (n2131,n60,n195);
and (n2132,n56,n197);
or (n2133,n48,n2059);
and (n2134,n2116,n2122);
or (n2135,n2136,n2156);
and (n2136,n2137,n2150);
xor (n2137,n2138,n2144);
nand (n2138,n2139,n2140);
or (n2139,n470,n2066);
nand (n2140,n345,n2141);
nand (n2141,n2142,n2143);
or (n2142,n190,n553);
or (n2143,n192,n551);
nand (n2144,n2145,n2149);
or (n2145,n179,n2146);
nor (n2146,n2147,n2148);
and (n2147,n187,n302);
and (n2148,n185,n304);
or (n2149,n188,n2073);
nand (n2150,n2151,n2155);
or (n2151,n1084,n2152);
nor (n2152,n2153,n2154);
and (n2153,n782,n88);
and (n2154,n783,n90);
or (n2155,n1989,n1085);
and (n2156,n2138,n2144);
or (n2157,n2158,n2178);
and (n2158,n2159,n2172);
xor (n2159,n2160,n2166);
nand (n2160,n2161,n2165);
or (n2161,n155,n2162);
nor (n2162,n2163,n2164);
and (n2163,n77,n217);
and (n2164,n78,n219);
or (n2165,n156,n1995);
nand (n2166,n2167,n2171);
or (n2167,n206,n2168);
nor (n2168,n2169,n2170);
and (n2169,n113,n889);
and (n2170,n114,n891);
or (n2171,n207,n2001);
nand (n2172,n2173,n2177);
or (n2173,n102,n2174);
nor (n2174,n2175,n2176);
and (n2175,n110,n1103);
and (n2176,n106,n1105);
or (n2177,n127,n1967);
and (n2178,n2160,n2166);
and (n2179,n2113,n2135);
or (n2180,n2181,n2209);
and (n2181,n2182,n2192);
xor (n2182,n2183,n2189);
nand (n2183,n2184,n2188);
or (n2184,n72,n2185);
nor (n2185,n2186,n2187);
and (n2186,n82,n124);
and (n2187,n83,n126);
or (n2188,n92,n1936);
nor (n2189,n2017,n2190);
and (n2190,n2191,n2025);
not (n2191,n2018);
or (n2192,n2193,n2208);
and (n2193,n2194,n2202);
xor (n2194,n2195,n2196);
nor (n2195,n132,n1268);
nand (n2196,n2197,n2201);
or (n2197,n1075,n2198);
nor (n2198,n2199,n2200);
and (n2199,n417,n243);
and (n2200,n415,n245);
or (n2201,n1080,n2020);
nand (n2202,n2203,n2207);
or (n2203,n313,n2204);
nor (n2204,n2205,n2206);
and (n2205,n36,n274);
and (n2206,n37,n276);
or (n2207,n318,n2036);
and (n2208,n2195,n2196);
and (n2209,n2183,n2189);
and (n2210,n2109,n2110);
or (n2211,n2212,n2223);
and (n2212,n2213,n2216);
xor (n2213,n2214,n2215);
xor (n2214,n2016,n2054);
xor (n2215,n1961,n2006);
or (n2216,n2217,n2222);
and (n2217,n2218,n2221);
xor (n2218,n2219,n2220);
xor (n2219,n1964,n1977);
xor (n2220,n2033,n2047);
xor (n2221,n1986,n1999);
and (n2222,n2219,n2220);
and (n2223,n2214,n2215);
and (n2224,n2105,n2106);
and (n2225,n2100,n2101);
and (n2226,n2095,n2096);
xor (n2227,n1803,n2089);
not (n2228,n2229);
nand (n2229,n2230,n4348,n4361);
nand (n2230,n2231,n2418,n4127,n4331);
nor (n2231,n2232,n2247);
nor (n2232,n2233,n2234);
xor (n2233,n2094,n2097);
or (n2234,n2235,n2246);
and (n2235,n2236,n2239);
xor (n2236,n2237,n2238);
xor (n2237,n1953,n2010);
xor (n2238,n2099,n2102);
or (n2239,n2240,n2245);
and (n2240,n2241,n2244);
xor (n2241,n2242,n2243);
xor (n2242,n2012,n2079);
xor (n2243,n1957,n2008);
xor (n2244,n2104,n2211);
and (n2245,n2242,n2243);
and (n2246,n2237,n2238);
nor (n2247,n2248,n2249);
xor (n2248,n2236,n2239);
or (n2249,n2250,n2417);
and (n2250,n2251,n2416);
xor (n2251,n2252,n2397);
or (n2252,n2253,n2396);
and (n2253,n2254,n2291);
xor (n2254,n2255,n2256);
xor (n2255,n2081,n2084);
or (n2256,n2257,n2290);
and (n2257,n2258,n2289);
xor (n2258,n2259,n2260);
xor (n2259,n2056,n2071);
or (n2260,n2261,n2288);
and (n2261,n2262,n2275);
xor (n2262,n2263,n2269);
nand (n2263,n2264,n2268);
or (n2264,n410,n2265);
nor (n2265,n2266,n2267);
and (n2266,n31,n436);
and (n2267,n32,n438);
or (n2268,n411,n1973);
nand (n2269,n2270,n2274);
or (n2270,n72,n2271);
nor (n2271,n2272,n2273);
and (n2272,n82,n118);
and (n2273,n83,n120);
or (n2274,n92,n2185);
and (n2275,n2276,n2282);
nor (n2276,n2277,n110);
nor (n2277,n2278,n2281);
and (n2278,n2279,n113);
not (n2279,n2280);
and (n2280,n1266,n108);
and (n2281,n1268,n107);
nand (n2282,n2283,n2287);
or (n2283,n1075,n2284);
nor (n2284,n2285,n2286);
and (n2285,n417,n377);
and (n2286,n415,n376);
or (n2287,n1080,n2198);
and (n2288,n2263,n2269);
xor (n2289,n2182,n2192);
and (n2290,n2259,n2260);
or (n2291,n2292,n2395);
and (n2292,n2293,n2394);
xor (n2293,n2294,n2366);
or (n2294,n2295,n2365);
and (n2295,n2296,n2343);
xor (n2296,n2297,n2320);
or (n2297,n2298,n2319);
and (n2298,n2299,n2313);
xor (n2299,n2300,n2307);
nand (n2300,n2301,n2305);
or (n2301,n2302,n313);
nor (n2302,n2303,n2304);
and (n2303,n36,n201);
and (n2304,n37,n203);
nand (n2305,n2306,n28);
not (n2306,n2204);
nand (n2307,n2308,n2312);
or (n2308,n228,n2309);
nor (n2309,n2310,n2311);
and (n2310,n240,n398);
and (n2311,n238,n397);
or (n2312,n229,n2118);
nand (n2313,n2314,n2318);
or (n2314,n260,n2315);
nor (n2315,n2316,n2317);
and (n2316,n264,n443);
and (n2317,n265,n445);
or (n2318,n278,n2124);
and (n2319,n2300,n2307);
or (n2320,n2321,n2342);
and (n2321,n2322,n2336);
xor (n2322,n2323,n2329);
nand (n2323,n2324,n2328);
or (n2324,n47,n2325);
nor (n2325,n2326,n2327);
and (n2326,n60,n223);
and (n2327,n56,n225);
or (n2328,n48,n2130);
nand (n2329,n2330,n2334);
or (n2330,n344,n2331);
nor (n2331,n2332,n2333);
and (n2332,n192,n308);
and (n2333,n190,n310);
or (n2334,n470,n2335);
not (n2335,n2141);
nand (n2336,n2337,n2341);
or (n2337,n179,n2338);
nor (n2338,n2339,n2340);
and (n2339,n187,n670);
and (n2340,n185,n672);
or (n2341,n188,n2146);
and (n2342,n2323,n2329);
or (n2343,n2344,n2364);
and (n2344,n2345,n2358);
xor (n2345,n2346,n2352);
nand (n2346,n2347,n2351);
or (n2347,n1084,n2348);
nor (n2348,n2349,n2350);
and (n2349,n782,n249);
and (n2350,n783,n251);
or (n2351,n2152,n1085);
nand (n2352,n2353,n2357);
or (n2353,n155,n2354);
nor (n2354,n2355,n2356);
and (n2355,n77,n124);
and (n2356,n78,n126);
or (n2357,n156,n2162);
nand (n2358,n2359,n2360);
or (n2359,n2168,n207);
or (n2360,n206,n2361);
nor (n2361,n2362,n2363);
and (n2362,n1064,n113);
and (n2363,n114,n1066);
and (n2364,n2346,n2352);
and (n2365,n2297,n2320);
or (n2366,n2367,n2393);
and (n2367,n2368,n2392);
xor (n2368,n2369,n2391);
or (n2369,n2370,n2390);
and (n2370,n2371,n2384);
xor (n2371,n2372,n2378);
nand (n2372,n2373,n2377);
or (n2373,n102,n2374);
nor (n2374,n2375,n2376);
and (n2375,n1268,n106);
and (n2376,n1266,n110);
or (n2377,n2174,n127);
nand (n2378,n2379,n2383);
or (n2379,n410,n2380);
nor (n2380,n2381,n2382);
and (n2381,n31,n281);
and (n2382,n32,n283);
or (n2383,n411,n2265);
nand (n2384,n2385,n2389);
or (n2385,n72,n2386);
nor (n2386,n2387,n2388);
and (n2387,n82,n150);
and (n2388,n83,n152);
or (n2389,n92,n2271);
and (n2390,n2372,n2378);
xor (n2391,n2194,n2202);
xor (n2392,n2137,n2150);
and (n2393,n2369,n2391);
xor (n2394,n2112,n2157);
and (n2395,n2294,n2366);
and (n2396,n2255,n2256);
or (n2397,n2398,n2415);
and (n2398,n2399,n2402);
xor (n2399,n2400,n2401);
xor (n2400,n2108,n2180);
xor (n2401,n2213,n2216);
or (n2402,n2403,n2414);
and (n2403,n2404,n2413);
xor (n2404,n2405,n2412);
or (n2405,n2406,n2411);
and (n2406,n2407,n2410);
xor (n2407,n2408,n2409);
xor (n2408,n2115,n2128);
xor (n2409,n2159,n2172);
xor (n2410,n2262,n2275);
and (n2411,n2408,n2409);
xor (n2412,n2218,n2221);
xor (n2413,n2258,n2289);
and (n2414,n2405,n2412);
and (n2415,n2400,n2401);
xor (n2416,n2241,n2244);
and (n2417,n2252,n2397);
nand (n2418,n2419,n3612);
nor (n2419,n2420,n3598);
and (n2420,n2421,n3009,n3331);
nor (n2421,n2422,n2924);
nor (n2422,n2423,n2811);
xor (n2423,n2424,n2804);
xor (n2424,n2425,n2597);
or (n2425,n2426,n2596);
and (n2426,n2427,n2521);
xor (n2427,n2428,n2464);
xor (n2428,n2429,n2448);
xor (n2429,n2430,n2439);
nand (n2430,n2431,n2435);
or (n2431,n155,n2432);
nor (n2432,n2433,n2434);
and (n2433,n77,n449);
and (n2434,n78,n451);
or (n2435,n156,n2436);
nor (n2436,n2437,n2438);
and (n2437,n77,n398);
and (n2438,n78,n397);
nand (n2439,n2440,n2444);
or (n2440,n72,n2441);
nor (n2441,n2442,n2443);
and (n2442,n551,n82);
and (n2443,n83,n553);
or (n2444,n92,n2445);
nor (n2445,n2446,n2447);
and (n2446,n82,n443);
and (n2447,n83,n445);
and (n2448,n2449,n2455);
nor (n2449,n2450,n192);
nor (n2450,n2451,n2454);
and (n2451,n2452,n264);
not (n2452,n2453);
and (n2453,n1266,n348);
and (n2454,n1268,n353);
nand (n2455,n2456,n2460);
or (n2456,n1084,n2457);
nor (n2457,n2458,n2459);
and (n2458,n782,n201);
and (n2459,n783,n203);
or (n2460,n2461,n1085);
nor (n2461,n2462,n2463);
and (n2462,n782,n274);
and (n2463,n783,n276);
or (n2464,n2465,n2520);
and (n2465,n2466,n2489);
xor (n2466,n2467,n2468);
xor (n2467,n2449,n2455);
or (n2468,n2469,n2488);
and (n2469,n2470,n2478);
xor (n2470,n2471,n2472);
and (n2471,n346,n1266);
nand (n2472,n2473,n2477);
or (n2473,n1084,n2474);
nor (n2474,n2475,n2476);
and (n2475,n782,n195);
and (n2476,n783,n197);
or (n2477,n2457,n1085);
nand (n2478,n2479,n2483);
or (n2479,n313,n2480);
nor (n2480,n2481,n2482);
and (n2481,n36,n144);
and (n2482,n37,n146);
or (n2483,n318,n2484);
not (n2484,n2485);
nor (n2485,n2486,n2487);
and (n2486,n150,n37);
and (n2487,n152,n36);
and (n2488,n2471,n2472);
or (n2489,n2490,n2519);
and (n2490,n2491,n2510);
xor (n2491,n2492,n2501);
nand (n2492,n2493,n2497);
or (n2493,n228,n2494);
nor (n2494,n2495,n2496);
and (n2495,n240,n889);
and (n2496,n238,n891);
or (n2497,n229,n2498);
nor (n2498,n2499,n2500);
and (n2499,n670,n240);
and (n2500,n672,n238);
nand (n2501,n2502,n2506);
or (n2502,n260,n2503);
nor (n2503,n2504,n2505);
and (n2504,n264,n1103);
and (n2505,n265,n1105);
or (n2506,n278,n2507);
nor (n2507,n2508,n2509);
and (n2508,n264,n1064);
and (n2509,n265,n1066);
nand (n2510,n2511,n2515);
or (n2511,n1075,n2512);
nor (n2512,n2513,n2514);
and (n2513,n417,n217);
and (n2514,n415,n219);
or (n2515,n1080,n2516);
nor (n2516,n2517,n2518);
and (n2517,n223,n417);
and (n2518,n225,n415);
and (n2519,n2492,n2501);
and (n2520,n2467,n2468);
or (n2521,n2522,n2595);
and (n2522,n2523,n2575);
xor (n2523,n2524,n2556);
or (n2524,n2525,n2555);
and (n2525,n2526,n2546);
xor (n2526,n2527,n2537);
nand (n2527,n2528,n2533);
or (n2528,n2529,n47);
not (n2529,n2530);
nand (n2530,n2531,n2532);
or (n2531,n56,n451);
or (n2532,n60,n449);
nand (n2533,n49,n2534);
nor (n2534,n2535,n2536);
and (n2535,n397,n60);
and (n2536,n398,n56);
nand (n2537,n2538,n2542);
or (n2538,n2539,n410);
nor (n2539,n2540,n2541);
and (n2540,n31,n118);
and (n2541,n32,n120);
nand (n2542,n619,n2543);
nand (n2543,n2544,n2545);
or (n2544,n32,n126);
or (n2545,n31,n124);
nand (n2546,n2547,n2551);
or (n2547,n155,n2548);
nor (n2548,n2549,n2550);
and (n2549,n77,n551);
and (n2550,n78,n553);
or (n2551,n156,n2552);
nor (n2552,n2553,n2554);
and (n2553,n443,n77);
and (n2554,n78,n445);
and (n2555,n2527,n2537);
xor (n2556,n2557,n2569);
xor (n2557,n2558,n2566);
nand (n2558,n2559,n2561);
or (n2559,n2560,n410);
not (n2560,n2543);
nand (n2561,n2562,n619);
not (n2562,n2563);
nor (n2563,n2564,n2565);
and (n2564,n219,n32);
and (n2565,n217,n31);
nand (n2566,n2567,n2568);
or (n2567,n155,n2552);
or (n2568,n2432,n156);
nand (n2569,n2570,n2574);
or (n2570,n72,n2571);
nor (n2571,n2572,n2573);
and (n2572,n308,n82);
and (n2573,n83,n310);
or (n2574,n92,n2441);
xor (n2575,n2576,n2589);
xor (n2576,n2577,n2583);
nand (n2577,n2578,n2579);
or (n2578,n2484,n313);
nand (n2579,n2580,n28);
nor (n2580,n2581,n2582);
and (n2581,n120,n36);
and (n2582,n118,n37);
nand (n2583,n2584,n2585);
or (n2584,n2498,n228);
nand (n2585,n2586,n230);
nor (n2586,n2587,n2588);
and (n2587,n304,n240);
and (n2588,n302,n238);
nand (n2589,n2590,n2591);
or (n2590,n260,n2507);
or (n2591,n2592,n278);
nor (n2592,n2593,n2594);
and (n2593,n264,n889);
and (n2594,n265,n891);
and (n2595,n2524,n2556);
and (n2596,n2428,n2464);
xor (n2597,n2598,n2722);
xor (n2598,n2599,n2673);
or (n2599,n2600,n2672);
and (n2600,n2601,n2643);
xor (n2601,n2602,n2619);
xor (n2602,n2603,n2611);
xor (n2603,n2604,n2605);
and (n2604,n1650,n1266);
nand (n2605,n2606,n2607);
or (n2606,n1084,n2461);
or (n2607,n2608,n1085);
nor (n2608,n2609,n2610);
and (n2609,n283,n783);
and (n2610,n281,n782);
nand (n2611,n2612,n2614);
or (n2612,n313,n2613);
not (n2613,n2580);
or (n2614,n318,n2615);
not (n2615,n2616);
nor (n2616,n2617,n2618);
and (n2617,n124,n37);
and (n2618,n126,n36);
xor (n2619,n2620,n2634);
xor (n2620,n2621,n2628);
nand (n2621,n2622,n2624);
or (n2622,n2623,n228);
not (n2623,n2586);
or (n2624,n229,n2625);
nor (n2625,n2626,n2627);
and (n2626,n310,n238);
and (n2627,n308,n240);
nand (n2628,n2629,n2630);
or (n2629,n260,n2592);
or (n2630,n278,n2631);
nor (n2631,n2632,n2633);
and (n2632,n264,n670);
and (n2633,n265,n672);
nand (n2634,n2635,n2639);
or (n2635,n1075,n2636);
nor (n2636,n2637,n2638);
and (n2637,n417,n195);
and (n2638,n415,n197);
or (n2639,n1080,n2640);
nor (n2640,n2641,n2642);
and (n2641,n417,n201);
and (n2642,n415,n203);
xor (n2643,n2644,n2666);
xor (n2644,n2645,n2655);
nand (n2645,n2646,n2651);
or (n2646,n2647,n344);
not (n2647,n2648);
nand (n2648,n2649,n2650);
or (n2649,n190,n1105);
or (n2650,n192,n1103);
or (n2651,n470,n2652);
nor (n2652,n2653,n2654);
and (n2653,n1066,n190);
and (n2654,n1064,n192);
nand (n2655,n2656,n2661);
or (n2656,n2657,n48);
not (n2657,n2658);
nand (n2658,n2659,n2660);
or (n2659,n56,n152);
or (n2660,n60,n150);
nand (n2661,n2662,n1130);
not (n2662,n2663);
nor (n2663,n2664,n2665);
and (n2664,n60,n144);
and (n2665,n56,n146);
nand (n2666,n2667,n2668);
or (n2667,n410,n2563);
or (n2668,n411,n2669);
nor (n2669,n2670,n2671);
and (n2670,n31,n223);
and (n2671,n32,n225);
and (n2672,n2602,n2619);
xor (n2673,n2674,n2719);
xor (n2674,n2675,n2695);
xor (n2675,n2676,n2689);
xor (n2676,n2677,n2683);
nand (n2677,n2678,n2679);
or (n2678,n2615,n313);
nand (n2679,n28,n2680);
nor (n2680,n2681,n2682);
and (n2681,n217,n37);
and (n2682,n219,n36);
nand (n2683,n2684,n2685);
or (n2684,n2625,n228);
nand (n2685,n230,n2686);
nand (n2686,n2687,n2688);
or (n2687,n238,n553);
or (n2688,n240,n551);
nand (n2689,n2690,n2691);
or (n2690,n260,n2631);
or (n2691,n278,n2692);
nor (n2692,n2693,n2694);
and (n2693,n264,n302);
and (n2694,n265,n304);
xor (n2695,n2696,n2710);
xor (n2696,n2697,n2704);
nand (n2697,n2698,n2699);
or (n2698,n2657,n47);
nand (n2699,n2700,n49);
not (n2700,n2701);
nor (n2701,n2702,n2703);
and (n2702,n120,n56);
and (n2703,n118,n60);
nand (n2704,n2705,n2706);
or (n2705,n344,n2652);
nand (n2706,n346,n2707);
nor (n2707,n2708,n2709);
and (n2708,n891,n192);
and (n2709,n889,n190);
nand (n2710,n2711,n2715);
or (n2711,n179,n2712);
nor (n2712,n2713,n2714);
and (n2713,n1268,n185);
and (n2714,n187,n1266);
or (n2715,n188,n2716);
nor (n2716,n2717,n2718);
and (n2717,n187,n1103);
and (n2718,n185,n1105);
or (n2719,n2720,n2721);
and (n2720,n2429,n2448);
and (n2721,n2430,n2439);
xor (n2722,n2723,n2776);
xor (n2723,n2724,n2752);
or (n2724,n2725,n2751);
and (n2725,n2726,n2733);
xor (n2726,n2727,n2730);
or (n2727,n2728,n2729);
and (n2728,n2576,n2589);
and (n2729,n2577,n2583);
or (n2730,n2731,n2732);
and (n2731,n2557,n2569);
and (n2732,n2558,n2566);
or (n2733,n2734,n2750);
and (n2734,n2735,n2746);
xor (n2735,n2736,n2740);
nand (n2736,n2737,n2738);
or (n2737,n2516,n1075);
nand (n2738,n2739,n779);
not (n2739,n2636);
nand (n2740,n2741,n2742);
or (n2741,n2647,n470);
or (n2742,n344,n2743);
nor (n2743,n2744,n2745);
and (n2744,n190,n1268);
and (n2745,n192,n1266);
nand (n2746,n2747,n2749);
or (n2747,n47,n2748);
not (n2748,n2534);
or (n2749,n48,n2663);
and (n2750,n2736,n2740);
and (n2751,n2727,n2730);
xor (n2752,n2753,n2773);
xor (n2753,n2754,n2760);
nand (n2754,n2755,n2756);
or (n2755,n72,n2445);
or (n2756,n92,n2757);
nor (n2757,n2758,n2759);
and (n2758,n82,n449);
and (n2759,n83,n451);
xor (n2760,n2761,n2767);
and (n2761,n2762,n185);
nand (n2762,n2763,n2764);
or (n2763,n1266,n184);
nand (n2764,n2765,n192);
not (n2765,n2766);
and (n2766,n1266,n184);
nand (n2767,n2768,n2769);
or (n2768,n2640,n1075);
nand (n2769,n779,n2770);
nor (n2770,n2771,n2772);
and (n2771,n274,n415);
and (n2772,n276,n417);
or (n2773,n2774,n2775);
and (n2774,n2620,n2634);
and (n2775,n2621,n2628);
xor (n2776,n2777,n2784);
xor (n2777,n2778,n2781);
or (n2778,n2779,n2780);
and (n2779,n2603,n2611);
and (n2780,n2604,n2605);
or (n2781,n2782,n2783);
and (n2782,n2644,n2666);
and (n2783,n2645,n2655);
xor (n2784,n2785,n2798);
xor (n2785,n2786,n2792);
nand (n2786,n2787,n2788);
or (n2787,n1084,n2608);
or (n2788,n2789,n1085);
nor (n2789,n2790,n2791);
and (n2790,n782,n436);
and (n2791,n783,n438);
nand (n2792,n2793,n2794);
or (n2793,n410,n2669);
nand (n2794,n619,n2795);
nor (n2795,n2796,n2797);
and (n2796,n195,n32);
and (n2797,n197,n31);
nand (n2798,n2799,n2800);
or (n2799,n155,n2436);
or (n2800,n156,n2801);
nor (n2801,n2802,n2803);
and (n2802,n77,n144);
and (n2803,n78,n146);
or (n2804,n2805,n2810);
and (n2805,n2806,n2809);
xor (n2806,n2807,n2808);
xor (n2807,n2726,n2733);
xor (n2808,n2601,n2643);
xor (n2809,n2427,n2521);
and (n2810,n2807,n2808);
or (n2811,n2812,n2923);
and (n2812,n2813,n2922);
xor (n2813,n2814,n2866);
or (n2814,n2815,n2865);
and (n2815,n2816,n2864);
xor (n2816,n2817,n2818);
xor (n2817,n2735,n2746);
or (n2818,n2819,n2863);
and (n2819,n2820,n2840);
xor (n2820,n2821,n2827);
nand (n2821,n2822,n2826);
or (n2822,n72,n2823);
nor (n2823,n2824,n2825);
and (n2824,n82,n302);
and (n2825,n83,n304);
or (n2826,n92,n2571);
and (n2827,n2828,n2834);
nor (n2828,n2829,n264);
nor (n2829,n2830,n2833);
and (n2830,n2831,n240);
not (n2831,n2832);
and (n2832,n1266,n266);
and (n2833,n1268,n268);
nand (n2834,n2835,n2839);
or (n2835,n1084,n2836);
nor (n2836,n2837,n2838);
and (n2837,n782,n223);
and (n2838,n783,n225);
or (n2839,n2474,n1085);
or (n2840,n2841,n2862);
and (n2841,n2842,n2856);
xor (n2842,n2843,n2850);
nand (n2843,n2844,n2848);
or (n2844,n2845,n313);
nor (n2845,n2846,n2847);
and (n2846,n36,n398);
and (n2847,n37,n397);
nand (n2848,n2849,n28);
not (n2849,n2480);
nand (n2850,n2851,n2855);
or (n2851,n228,n2852);
nor (n2852,n2853,n2854);
and (n2853,n240,n1064);
and (n2854,n238,n1066);
or (n2855,n229,n2494);
nand (n2856,n2857,n2861);
or (n2857,n260,n2858);
nor (n2858,n2859,n2860);
and (n2859,n1268,n265);
and (n2860,n264,n1266);
or (n2861,n278,n2503);
and (n2862,n2843,n2850);
and (n2863,n2821,n2827);
xor (n2864,n2466,n2489);
and (n2865,n2817,n2818);
or (n2866,n2867,n2921);
and (n2867,n2868,n2898);
xor (n2868,n2869,n2897);
or (n2869,n2870,n2896);
and (n2870,n2871,n2895);
xor (n2871,n2872,n2894);
or (n2872,n2873,n2893);
and (n2873,n2874,n2887);
xor (n2874,n2875,n2881);
nand (n2875,n2876,n2880);
or (n2876,n1075,n2877);
nor (n2877,n2878,n2879);
and (n2878,n417,n124);
and (n2879,n415,n126);
or (n2880,n1080,n2512);
nand (n2881,n2882,n2886);
or (n2882,n47,n2883);
nor (n2883,n2884,n2885);
and (n2884,n60,n443);
and (n2885,n56,n445);
or (n2886,n48,n2529);
nand (n2887,n2888,n2892);
or (n2888,n410,n2889);
nor (n2889,n2890,n2891);
and (n2890,n31,n150);
and (n2891,n32,n152);
or (n2892,n411,n2539);
and (n2893,n2875,n2881);
xor (n2894,n2526,n2546);
xor (n2895,n2470,n2478);
and (n2896,n2872,n2894);
xor (n2897,n2523,n2575);
or (n2898,n2899,n2920);
and (n2899,n2900,n2919);
xor (n2900,n2901,n2902);
xor (n2901,n2491,n2510);
or (n2902,n2903,n2918);
and (n2903,n2904,n2917);
xor (n2904,n2905,n2911);
nand (n2905,n2906,n2910);
or (n2906,n155,n2907);
nor (n2907,n2908,n2909);
and (n2908,n77,n308);
and (n2909,n78,n310);
or (n2910,n156,n2548);
nand (n2911,n2912,n2916);
or (n2912,n72,n2913);
nor (n2913,n2914,n2915);
and (n2914,n82,n670);
and (n2915,n83,n672);
or (n2916,n92,n2823);
xor (n2917,n2828,n2834);
and (n2918,n2905,n2911);
xor (n2919,n2820,n2840);
and (n2920,n2901,n2902);
and (n2921,n2869,n2897);
xor (n2922,n2806,n2809);
and (n2923,n2814,n2866);
nor (n2924,n2925,n2926);
xor (n2925,n2813,n2922);
or (n2926,n2927,n3008);
and (n2927,n2928,n3007);
xor (n2928,n2929,n2930);
xor (n2929,n2816,n2864);
or (n2930,n2931,n3006);
and (n2931,n2932,n3005);
xor (n2932,n2933,n2998);
or (n2933,n2934,n2997);
and (n2934,n2935,n2975);
xor (n2935,n2936,n2953);
or (n2936,n2937,n2952);
and (n2937,n2938,n2946);
xor (n2938,n2939,n2940);
and (n2939,n269,n1266);
nand (n2940,n2941,n2945);
or (n2941,n1084,n2942);
nor (n2942,n2943,n2944);
and (n2943,n782,n217);
and (n2944,n783,n219);
or (n2945,n2836,n1085);
nand (n2946,n2947,n2951);
or (n2947,n1075,n2948);
nor (n2948,n2949,n2950);
and (n2949,n417,n118);
and (n2950,n415,n120);
or (n2951,n1080,n2877);
and (n2952,n2939,n2940);
or (n2953,n2954,n2974);
and (n2954,n2955,n2968);
xor (n2955,n2956,n2962);
nand (n2956,n2957,n2961);
or (n2957,n410,n2958);
nor (n2958,n2959,n2960);
and (n2959,n31,n144);
and (n2960,n32,n146);
or (n2961,n411,n2889);
nand (n2962,n2963,n2967);
or (n2963,n155,n2964);
nor (n2964,n2965,n2966);
and (n2965,n77,n302);
and (n2966,n78,n304);
or (n2967,n156,n2907);
nand (n2968,n2969,n2973);
or (n2969,n72,n2970);
nor (n2970,n2971,n2972);
and (n2971,n82,n889);
and (n2972,n83,n891);
or (n2973,n92,n2913);
and (n2974,n2956,n2962);
or (n2975,n2976,n2996);
and (n2976,n2977,n2990);
xor (n2977,n2978,n2984);
nand (n2978,n2979,n2983);
or (n2979,n228,n2980);
nor (n2980,n2981,n2982);
and (n2981,n240,n1103);
and (n2982,n238,n1105);
or (n2983,n229,n2852);
nand (n2984,n2985,n2989);
or (n2985,n313,n2986);
nor (n2986,n2987,n2988);
and (n2987,n36,n449);
and (n2988,n37,n451);
or (n2989,n318,n2845);
nand (n2990,n2991,n2995);
or (n2991,n47,n2992);
nor (n2992,n2993,n2994);
and (n2993,n551,n60);
and (n2994,n56,n553);
or (n2995,n48,n2883);
and (n2996,n2978,n2984);
and (n2997,n2936,n2953);
or (n2998,n2999,n3004);
and (n2999,n3000,n3003);
xor (n3000,n3001,n3002);
xor (n3001,n2842,n2856);
xor (n3002,n2874,n2887);
xor (n3003,n2904,n2917);
and (n3004,n3001,n3002);
xor (n3005,n2871,n2895);
and (n3006,n2933,n2998);
xor (n3007,n2868,n2898);
and (n3008,n2929,n2930);
nand (n3009,n3010,n3330);
or (n3010,n3011,n3325);
nor (n3011,n3012,n3324);
and (n3012,n3013,n3312);
not (n3013,n3014);
nand (n3014,n3015,n3309);
or (n3015,n3016,n3289);
not (n3016,n3017);
nand (n3017,n3018,n3231);
xor (n3018,n3019,n3162);
xor (n3019,n3020,n3025);
xor (n3020,n3021,n3024);
xor (n3021,n3022,n3023);
xor (n3022,n2955,n2968);
xor (n3023,n2938,n2946);
xor (n3024,n2977,n2990);
or (n3025,n3026,n3161);
and (n3026,n3027,n3102);
xor (n3027,n3028,n3067);
or (n3028,n3029,n3066);
and (n3029,n3030,n3050);
xor (n3030,n3031,n3040);
nand (n3031,n3032,n3036);
or (n3032,n155,n3033);
nor (n3033,n3034,n3035);
and (n3034,n77,n889);
and (n3035,n78,n891);
or (n3036,n156,n3037);
nor (n3037,n3038,n3039);
and (n3038,n77,n670);
and (n3039,n78,n672);
nand (n3040,n3041,n3046);
or (n3041,n3042,n72);
not (n3042,n3043);
nand (n3043,n3044,n3045);
or (n3044,n1105,n83);
or (n3045,n82,n1103);
or (n3046,n92,n3047);
nor (n3047,n3048,n3049);
and (n3048,n82,n1064);
and (n3049,n83,n1066);
and (n3050,n3051,n3057);
nor (n3051,n3052,n82);
nor (n3052,n3053,n3056);
and (n3053,n3054,n77);
not (n3054,n3055);
and (n3055,n1266,n76);
and (n3056,n1268,n85);
nand (n3057,n3058,n3062);
or (n3058,n3059,n1084);
nor (n3059,n3060,n3061);
and (n3060,n782,n150);
and (n3061,n783,n152);
or (n3062,n3063,n1085);
nor (n3063,n3064,n3065);
and (n3064,n782,n118);
and (n3065,n783,n120);
and (n3066,n3031,n3040);
xor (n3067,n3068,n3085);
xor (n3068,n3069,n3072);
nand (n3069,n3070,n3071);
or (n3070,n72,n3047);
or (n3071,n92,n2970);
xor (n3072,n3073,n3079);
nor (n3073,n3074,n240);
nor (n3074,n3075,n3078);
and (n3075,n3076,n82);
not (n3076,n3077);
and (n3077,n1266,n232);
and (n3078,n1268,n237);
nand (n3079,n3080,n3084);
or (n3080,n1084,n3081);
nor (n3081,n3082,n3083);
and (n3082,n782,n124);
and (n3083,n783,n126);
or (n3084,n2942,n1085);
or (n3085,n3086,n3101);
and (n3086,n3087,n3092);
xor (n3087,n3088,n3089);
nor (n3088,n229,n1268);
nand (n3089,n3090,n3091);
or (n3090,n1084,n3063);
or (n3091,n3081,n1085);
nand (n3092,n3093,n3097);
or (n3093,n1075,n3094);
nor (n3094,n3095,n3096);
and (n3095,n417,n144);
and (n3096,n415,n146);
or (n3097,n1080,n3098);
nor (n3098,n3099,n3100);
and (n3099,n417,n150);
and (n3100,n415,n152);
and (n3101,n3088,n3089);
or (n3102,n3103,n3160);
and (n3103,n3104,n3159);
xor (n3104,n3105,n3134);
or (n3105,n3106,n3133);
and (n3106,n3107,n3124);
xor (n3107,n3108,n3114);
nand (n3108,n3109,n3113);
or (n3109,n1075,n3110);
nor (n3110,n3111,n3112);
and (n3111,n417,n398);
and (n3112,n415,n397);
or (n3113,n1080,n3094);
nand (n3114,n3115,n3119);
or (n3115,n313,n3116);
nor (n3116,n3117,n3118);
and (n3117,n36,n308);
and (n3118,n37,n310);
or (n3119,n318,n3120);
not (n3120,n3121);
nor (n3121,n3122,n3123);
and (n3122,n551,n37);
and (n3123,n553,n36);
nand (n3124,n3125,n3129);
or (n3125,n47,n3126);
nor (n3126,n3127,n3128);
and (n3127,n60,n670);
and (n3128,n56,n672);
or (n3129,n48,n3130);
nor (n3130,n3131,n3132);
and (n3131,n60,n302);
and (n3132,n56,n304);
and (n3133,n3108,n3114);
or (n3134,n3135,n3158);
and (n3135,n3136,n3152);
xor (n3136,n3137,n3146);
nand (n3137,n3138,n3142);
or (n3138,n410,n3139);
nor (n3139,n3140,n3141);
and (n3140,n31,n443);
and (n3141,n32,n445);
or (n3142,n411,n3143);
nor (n3143,n3144,n3145);
and (n3144,n31,n449);
and (n3145,n32,n451);
nand (n3146,n3147,n3151);
or (n3147,n155,n3148);
nor (n3148,n3149,n3150);
and (n3149,n77,n1064);
and (n3150,n78,n1066);
or (n3151,n156,n3033);
nand (n3152,n3153,n3154);
or (n3153,n3042,n92);
or (n3154,n72,n3155);
nor (n3155,n3156,n3157);
and (n3156,n1268,n83);
and (n3157,n1266,n82);
and (n3158,n3137,n3146);
xor (n3159,n3087,n3092);
and (n3160,n3105,n3134);
and (n3161,n3028,n3067);
xor (n3162,n3163,n3211);
xor (n3163,n3164,n3167);
or (n3164,n3165,n3166);
and (n3165,n3068,n3085);
and (n3166,n3069,n3072);
xor (n3167,n3168,n3190);
xor (n3168,n3169,n3170);
and (n3169,n3073,n3079);
or (n3170,n3171,n3189);
and (n3171,n3172,n3183);
xor (n3172,n3173,n3177);
nand (n3173,n3174,n3175);
or (n3174,n2948,n1080);
nand (n3175,n3176,n785);
not (n3176,n3098);
nand (n3177,n3178,n3182);
or (n3178,n228,n3179);
nor (n3179,n3180,n3181);
and (n3180,n238,n1268);
and (n3181,n240,n1266);
or (n3182,n229,n2980);
nand (n3183,n3184,n3188);
or (n3184,n313,n3185);
nor (n3185,n3186,n3187);
and (n3186,n36,n443);
and (n3187,n37,n445);
or (n3188,n318,n2986);
and (n3189,n3173,n3177);
or (n3190,n3191,n3210);
and (n3191,n3192,n3207);
xor (n3192,n3193,n3200);
nand (n3193,n3194,n3198);
or (n3194,n3195,n47);
nor (n3195,n3196,n3197);
and (n3196,n310,n56);
and (n3197,n308,n60);
nand (n3198,n3199,n49);
not (n3199,n2992);
nand (n3200,n3201,n3205);
or (n3201,n3202,n410);
nor (n3202,n3203,n3204);
and (n3203,n31,n398);
and (n3204,n32,n397);
nand (n3205,n3206,n619);
not (n3206,n2958);
nand (n3207,n3208,n3209);
or (n3208,n155,n3037);
or (n3209,n156,n2964);
and (n3210,n3193,n3200);
or (n3211,n3212,n3230);
and (n3212,n3213,n3229);
xor (n3213,n3214,n3228);
or (n3214,n3215,n3227);
and (n3215,n3216,n3224);
xor (n3216,n3217,n3221);
nand (n3217,n3218,n3219);
or (n3218,n3120,n313);
nand (n3219,n3220,n28);
not (n3220,n3185);
nand (n3221,n3222,n3223);
or (n3222,n47,n3130);
or (n3223,n48,n3195);
nand (n3224,n3225,n3226);
or (n3225,n410,n3143);
or (n3226,n411,n3202);
and (n3227,n3217,n3221);
xor (n3228,n3192,n3207);
xor (n3229,n3172,n3183);
and (n3230,n3214,n3228);
or (n3231,n3232,n3288);
and (n3232,n3233,n3287);
xor (n3233,n3234,n3235);
xor (n3234,n3213,n3229);
or (n3235,n3236,n3286);
and (n3236,n3237,n3240);
xor (n3237,n3238,n3239);
xor (n3238,n3216,n3224);
xor (n3239,n3030,n3050);
or (n3240,n3241,n3285);
and (n3241,n3242,n3262);
xor (n3242,n3243,n3244);
xor (n3243,n3051,n3057);
or (n3244,n3245,n3261);
and (n3245,n3246,n3255);
xor (n3246,n3247,n3248);
nor (n3247,n92,n1268);
nand (n3248,n3249,n3254);
or (n3249,n3250,n1075);
not (n3250,n3251);
nand (n3251,n3252,n3253);
or (n3252,n415,n451);
or (n3253,n417,n449);
or (n3254,n1080,n3110);
nand (n3255,n3256,n3260);
or (n3256,n313,n3257);
nor (n3257,n3258,n3259);
and (n3258,n36,n302);
and (n3259,n37,n304);
or (n3260,n318,n3116);
and (n3261,n3247,n3248);
or (n3262,n3263,n3284);
and (n3263,n3264,n3278);
xor (n3264,n3265,n3271);
nand (n3265,n3266,n3270);
or (n3266,n47,n3267);
nor (n3267,n3268,n3269);
and (n3268,n60,n889);
and (n3269,n56,n891);
or (n3270,n48,n3126);
nand (n3271,n3272,n3277);
or (n3272,n1084,n3273);
not (n3273,n3274);
nor (n3274,n3275,n3276);
and (n3275,n144,n783);
and (n3276,n146,n782);
or (n3277,n3059,n1085);
nand (n3278,n3279,n3283);
or (n3279,n155,n3280);
nor (n3280,n3281,n3282);
and (n3281,n77,n1103);
and (n3282,n78,n1105);
or (n3283,n156,n3148);
and (n3284,n3265,n3271);
and (n3285,n3243,n3244);
and (n3286,n3238,n3239);
xor (n3287,n3027,n3102);
and (n3288,n3234,n3235);
not (n3289,n3290);
nand (n3290,n3291,n3306);
xor (n3291,n3292,n3297);
xor (n3292,n3293,n3294);
xor (n3293,n3000,n3003);
or (n3294,n3295,n3296);
and (n3295,n3163,n3211);
and (n3296,n3164,n3167);
xor (n3297,n3298,n3303);
xor (n3298,n3299,n3302);
or (n3299,n3300,n3301);
and (n3300,n3168,n3190);
and (n3301,n3169,n3170);
xor (n3302,n2935,n2975);
or (n3303,n3304,n3305);
and (n3304,n3021,n3024);
and (n3305,n3022,n3023);
or (n3306,n3307,n3308);
and (n3307,n3019,n3162);
and (n3308,n3020,n3025);
nand (n3309,n3310,n3311);
not (n3310,n3291);
not (n3311,n3306);
not (n3312,n3313);
nor (n3313,n3314,n3321);
xor (n3314,n3315,n3320);
xor (n3315,n3316,n3317);
xor (n3316,n2900,n2919);
or (n3317,n3318,n3319);
and (n3318,n3298,n3303);
and (n3319,n3299,n3302);
xor (n3320,n2932,n3005);
or (n3321,n3322,n3323);
and (n3322,n3292,n3297);
and (n3323,n3293,n3294);
and (n3324,n3314,n3321);
nor (n3325,n3326,n3327);
xor (n3326,n2928,n3007);
or (n3327,n3328,n3329);
and (n3328,n3315,n3320);
and (n3329,n3316,n3317);
nand (n3330,n3326,n3327);
nor (n3331,n3332,n3458);
nor (n3332,n3333,n3455);
xor (n3333,n3334,n3452);
xor (n3334,n3335,n3352);
xor (n3335,n3336,n3349);
xor (n3336,n3337,n3340);
or (n3337,n3338,n3339);
and (n3338,n2777,n2784);
and (n3339,n2778,n2781);
xor (n3340,n3341,n3346);
xor (n3341,n3342,n3343);
and (n3342,n2761,n2767);
or (n3343,n3344,n3345);
and (n3344,n2785,n2798);
and (n3345,n2786,n2792);
or (n3346,n3347,n3348);
and (n3347,n2696,n2710);
and (n3348,n2697,n2704);
or (n3349,n3350,n3351);
and (n3350,n2674,n2719);
and (n3351,n2675,n2695);
xor (n3352,n3353,n3449);
xor (n3353,n3354,n3402);
xor (n3354,n3355,n3380);
xor (n3355,n3356,n3359);
or (n3356,n3357,n3358);
and (n3357,n2676,n2689);
and (n3358,n2677,n2683);
xor (n3359,n3360,n3374);
xor (n3360,n3361,n3368);
nand (n3361,n3362,n3364);
or (n3362,n3363,n410);
not (n3363,n2795);
nand (n3364,n619,n3365);
nor (n3365,n3366,n3367);
and (n3366,n201,n32);
and (n3367,n203,n31);
nand (n3368,n3369,n3370);
or (n3369,n155,n2801);
or (n3370,n3371,n156);
nor (n3371,n3372,n3373);
and (n3372,n77,n150);
and (n3373,n78,n152);
nand (n3374,n3375,n3376);
or (n3375,n72,n2757);
or (n3376,n92,n3377);
nor (n3377,n3378,n3379);
and (n3378,n82,n398);
and (n3379,n83,n397);
xor (n3380,n3381,n3395);
xor (n3381,n3382,n3389);
nand (n3382,n3383,n3385);
or (n3383,n3384,n228);
not (n3384,n2686);
nand (n3385,n3386,n230);
nor (n3386,n3387,n3388);
and (n3387,n443,n238);
and (n3388,n445,n240);
nand (n3389,n3390,n3391);
or (n3390,n260,n2692);
or (n3391,n278,n3392);
nor (n3392,n3393,n3394);
and (n3393,n264,n308);
and (n3394,n265,n310);
nand (n3395,n3396,n3397);
or (n3396,n47,n2701);
or (n3397,n48,n3398);
not (n3398,n3399);
nand (n3399,n3400,n3401);
or (n3400,n56,n126);
or (n3401,n60,n124);
xor (n3402,n3403,n3446);
xor (n3403,n3404,n3428);
xor (n3404,n3405,n3422);
xor (n3405,n3406,n3413);
nand (n3406,n3407,n3409);
or (n3407,n3408,n344);
not (n3408,n2707);
nand (n3409,n3410,n346);
nor (n3410,n3411,n3412);
and (n3411,n672,n192);
and (n3412,n670,n190);
nand (n3413,n3414,n3419);
or (n3414,n3415,n188);
not (n3415,n3416);
nand (n3416,n3417,n3418);
or (n3417,n185,n1066);
or (n3418,n187,n1064);
nand (n3419,n3420,n3421);
not (n3420,n2716);
not (n3421,n179);
nand (n3422,n3423,n3424);
or (n3423,n1084,n2789);
or (n3424,n3425,n1085);
nor (n3425,n3426,n3427);
and (n3426,n376,n783);
and (n3427,n377,n782);
xor (n3428,n3429,n3439);
xor (n3429,n3430,n3431);
nor (n3430,n207,n1268);
nand (n3431,n3432,n3434);
or (n3432,n3433,n1075);
not (n3433,n2770);
nand (n3434,n3435,n779);
not (n3435,n3436);
nor (n3436,n3437,n3438);
and (n3437,n283,n415);
and (n3438,n281,n417);
nand (n3439,n3440,n3442);
or (n3440,n3441,n313);
not (n3441,n2680);
nand (n3442,n28,n3443);
nand (n3443,n3444,n3445);
or (n3444,n37,n225);
or (n3445,n36,n223);
or (n3446,n3447,n3448);
and (n3447,n2753,n2773);
and (n3448,n2754,n2760);
or (n3449,n3450,n3451);
and (n3450,n2723,n2776);
and (n3451,n2724,n2752);
or (n3452,n3453,n3454);
and (n3453,n2598,n2722);
and (n3454,n2599,n2673);
or (n3455,n3456,n3457);
and (n3456,n2424,n2804);
and (n3457,n2425,n2597);
nor (n3458,n3459,n3462);
or (n3459,n3460,n3461);
and (n3460,n3334,n3452);
and (n3461,n3335,n3352);
xor (n3462,n3463,n3470);
xor (n3463,n3464,n3467);
or (n3464,n3465,n3466);
and (n3465,n3336,n3349);
and (n3466,n3337,n3340);
or (n3467,n3468,n3469);
and (n3468,n3353,n3449);
and (n3469,n3354,n3402);
xor (n3470,n3471,n3531);
xor (n3471,n3472,n3528);
xor (n3472,n3473,n3525);
xor (n3473,n3474,n3497);
xor (n3474,n3475,n3491);
xor (n3475,n3476,n3484);
nand (n3476,n3477,n3479);
or (n3477,n3478,n313);
not (n3478,n3443);
nand (n3479,n3480,n28);
not (n3480,n3481);
nor (n3481,n3482,n3483);
and (n3482,n36,n195);
and (n3483,n37,n197);
nand (n3484,n3485,n3487);
or (n3485,n228,n3486);
not (n3486,n3386);
or (n3487,n229,n3488);
nor (n3488,n3489,n3490);
and (n3489,n240,n449);
and (n3490,n238,n451);
nand (n3491,n3492,n3493);
or (n3492,n260,n3392);
or (n3493,n278,n3494);
nor (n3494,n3495,n3496);
and (n3495,n264,n551);
and (n3496,n265,n553);
xor (n3497,n3498,n3511);
xor (n3498,n3499,n3505);
nand (n3499,n3500,n3501);
or (n3500,n155,n3371);
or (n3501,n156,n3502);
nor (n3502,n3503,n3504);
and (n3503,n77,n118);
and (n3504,n78,n120);
nand (n3505,n3506,n3507);
or (n3506,n72,n3377);
or (n3507,n92,n3508);
nor (n3508,n3509,n3510);
and (n3509,n82,n144);
and (n3510,n83,n146);
xor (n3511,n3512,n3518);
nor (n3512,n3513,n113);
nor (n3513,n3514,n3517);
and (n3514,n3515,n187);
not (n3515,n3516);
and (n3516,n1266,n209);
and (n3517,n1268,n211);
nand (n3518,n3519,n3524);
or (n3519,n3520,n1080);
not (n3520,n3521);
nand (n3521,n3522,n3523);
or (n3522,n415,n438);
or (n3523,n417,n436);
or (n3524,n1075,n3436);
or (n3525,n3526,n3527);
and (n3526,n3341,n3346);
and (n3527,n3342,n3343);
or (n3528,n3529,n3530);
and (n3529,n3403,n3446);
and (n3530,n3404,n3428);
xor (n3531,n3532,n3547);
xor (n3532,n3533,n3544);
xor (n3533,n3534,n3541);
xor (n3534,n3535,n3538);
or (n3535,n3536,n3537);
and (n3536,n3405,n3422);
and (n3537,n3406,n3413);
or (n3538,n3539,n3540);
and (n3539,n3360,n3374);
and (n3540,n3361,n3368);
or (n3541,n3542,n3543);
and (n3542,n3429,n3439);
and (n3543,n3430,n3431);
or (n3544,n3545,n3546);
and (n3545,n3355,n3380);
and (n3546,n3356,n3359);
xor (n3547,n3548,n3576);
xor (n3548,n3549,n3552);
or (n3549,n3550,n3551);
and (n3550,n3381,n3395);
and (n3551,n3382,n3389);
xor (n3552,n3553,n3567);
xor (n3553,n3554,n3560);
nand (n3554,n3555,n3556);
or (n3555,n1084,n3425);
or (n3556,n3557,n1085);
nor (n3557,n3558,n3559);
and (n3558,n243,n782);
and (n3559,n245,n783);
nand (n3560,n3561,n3563);
or (n3561,n3562,n410);
not (n3562,n3365);
nand (n3563,n619,n3564);
nand (n3564,n3565,n3566);
or (n3565,n32,n276);
or (n3566,n31,n274);
nand (n3567,n3568,n3572);
or (n3568,n206,n3569);
nor (n3569,n3570,n3571);
and (n3570,n1268,n114);
and (n3571,n1266,n113);
or (n3572,n207,n3573);
nor (n3573,n3574,n3575);
and (n3574,n1103,n113);
and (n3575,n114,n1105);
xor (n3576,n3577,n3592);
xor (n3577,n3578,n3585);
nand (n3578,n3579,n3584);
or (n3579,n3580,n48);
not (n3580,n3581);
nand (n3581,n3582,n3583);
or (n3582,n56,n219);
or (n3583,n60,n217);
nand (n3584,n1130,n3399);
nand (n3585,n3586,n3588);
or (n3586,n344,n3587);
not (n3587,n3410);
or (n3588,n470,n3589);
nor (n3589,n3590,n3591);
and (n3590,n192,n302);
and (n3591,n190,n304);
nand (n3592,n3593,n3594);
or (n3593,n179,n3415);
or (n3594,n188,n3595);
nor (n3595,n3596,n3597);
and (n3596,n187,n889);
and (n3597,n185,n891);
nand (n3598,n3599,n3606);
or (n3599,n3600,n3601);
not (n3600,n3331);
not (n3601,n3602);
nand (n3602,n3603,n3605);
or (n3603,n2422,n3604);
nand (n3604,n2925,n2926);
nand (n3605,n2423,n2811);
nor (n3606,n3607,n3611);
and (n3607,n3608,n3610);
not (n3608,n3609);
nand (n3609,n3333,n3455);
not (n3610,n3458);
and (n3611,n3459,n3462);
nand (n3612,n2421,n3331,n3613,n3617);
and (n3613,n3614,n3615,n3312);
not (n3614,n3325);
and (n3615,n3309,n3616);
or (n3616,n3231,n3018);
nand (n3617,n3618,n4117,n4126);
nand (n3618,n3619,n4055,n4112);
or (n3619,n3620,n4054);
and (n3620,n3621,n3797);
xor (n3621,n3622,n3745);
or (n3622,n3623,n3744);
and (n3623,n3624,n3705);
xor (n3624,n3625,n3654);
xor (n3625,n3626,n3645);
xor (n3626,n3627,n3636);
nand (n3627,n3628,n3632);
or (n3628,n47,n3629);
nor (n3629,n3630,n3631);
and (n3630,n60,n1103);
and (n3631,n56,n1105);
or (n3632,n48,n3633);
nor (n3633,n3634,n3635);
and (n3634,n60,n1064);
and (n3635,n56,n1066);
nand (n3636,n3637,n3641);
or (n3637,n3638,n1084);
nor (n3638,n3639,n3640);
and (n3639,n782,n449);
and (n3640,n783,n451);
or (n3641,n3642,n1085);
nor (n3642,n3643,n3644);
and (n3643,n782,n398);
and (n3644,n783,n397);
nand (n3645,n3646,n3650);
or (n3646,n410,n3647);
nor (n3647,n3648,n3649);
and (n3648,n31,n302);
and (n3649,n32,n304);
or (n3650,n411,n3651);
nor (n3651,n3652,n3653);
and (n3652,n31,n308);
and (n3653,n32,n310);
or (n3654,n3655,n3704);
and (n3655,n3656,n3679);
xor (n3656,n3657,n3663);
nand (n3657,n3658,n3662);
or (n3658,n410,n3659);
nor (n3659,n3660,n3661);
and (n3660,n31,n670);
and (n3661,n32,n672);
or (n3662,n411,n3647);
xor (n3663,n3664,n3670);
and (n3664,n3665,n56);
nand (n3665,n3666,n3667);
or (n3666,n1266,n52);
nand (n3667,n3668,n36);
not (n3668,n3669);
and (n3669,n1266,n52);
nand (n3670,n3671,n3675);
or (n3671,n1075,n3672);
nor (n3672,n3673,n3674);
and (n3673,n417,n308);
and (n3674,n415,n310);
or (n3675,n1080,n3676);
nor (n3676,n3677,n3678);
and (n3677,n417,n551);
and (n3678,n415,n553);
or (n3679,n3680,n3703);
and (n3680,n3681,n3692);
xor (n3681,n3682,n3683);
and (n3682,n49,n1266);
nand (n3683,n3684,n3688);
or (n3684,n1084,n3685);
nor (n3685,n3686,n3687);
and (n3686,n782,n551);
and (n3687,n783,n553);
or (n3688,n3689,n1085);
nor (n3689,n3690,n3691);
and (n3690,n782,n443);
and (n3691,n783,n445);
nand (n3692,n3693,n3698);
or (n3693,n3694,n313);
not (n3694,n3695);
nor (n3695,n3696,n3697);
and (n3696,n1103,n37);
and (n3697,n1105,n36);
nand (n3698,n3699,n28);
not (n3699,n3700);
nor (n3700,n3701,n3702);
and (n3701,n36,n1064);
and (n3702,n37,n1066);
and (n3703,n3682,n3683);
and (n3704,n3657,n3663);
xor (n3705,n3706,n3729);
xor (n3706,n3707,n3708);
and (n3707,n3664,n3670);
or (n3708,n3709,n3728);
and (n3709,n3710,n3725);
xor (n3710,n3711,n3717);
nand (n3711,n3712,n3713);
or (n3712,n313,n3700);
or (n3713,n318,n3714);
nor (n3714,n3715,n3716);
and (n3715,n36,n889);
and (n3716,n37,n891);
nand (n3717,n3718,n3723);
or (n3718,n3719,n47);
not (n3719,n3720);
nand (n3720,n3721,n3722);
or (n3721,n60,n1266);
or (n3722,n1268,n56);
nand (n3723,n3724,n49);
not (n3724,n3629);
nand (n3725,n3726,n3727);
or (n3726,n1084,n3689);
or (n3727,n3638,n1085);
and (n3728,n3711,n3717);
xor (n3729,n3730,n3738);
xor (n3730,n3731,n3732);
nor (n3731,n156,n1268);
nand (n3732,n3733,n3734);
or (n3733,n1075,n3676);
or (n3734,n1080,n3735);
nor (n3735,n3736,n3737);
and (n3736,n417,n443);
and (n3737,n415,n445);
nand (n3738,n3739,n3740);
or (n3739,n313,n3714);
or (n3740,n318,n3741);
nor (n3741,n3742,n3743);
and (n3742,n36,n670);
and (n3743,n37,n672);
and (n3744,n3625,n3654);
xor (n3745,n3746,n3794);
xor (n3746,n3747,n3775);
xor (n3747,n3748,n3761);
xor (n3748,n3749,n3755);
nand (n3749,n3750,n3754);
or (n3750,n155,n3751);
nor (n3751,n3752,n3753);
and (n3752,n1268,n78);
and (n3753,n77,n1266);
or (n3754,n156,n3280);
nand (n3755,n3756,n3757);
or (n3756,n410,n3651);
or (n3757,n411,n3758);
nor (n3758,n3759,n3760);
and (n3759,n31,n551);
and (n3760,n32,n553);
nand (n3761,n3762,n3774);
or (n3762,n3763,n3770);
not (n3763,n3764);
nand (n3764,n3765,n78);
nand (n3765,n3766,n3767);
or (n3766,n1266,n159);
nand (n3767,n3768,n60);
not (n3768,n3769);
and (n3769,n1266,n159);
not (n3770,n3771);
nand (n3771,n3772,n3773);
or (n3772,n1075,n3735);
or (n3773,n1080,n3250);
or (n3774,n3771,n3764);
xor (n3775,n3776,n3783);
xor (n3776,n3777,n3780);
or (n3777,n3778,n3779);
and (n3778,n3730,n3738);
and (n3779,n3731,n3732);
or (n3780,n3781,n3782);
and (n3781,n3626,n3645);
and (n3782,n3627,n3636);
xor (n3783,n3784,n3791);
xor (n3784,n3785,n3788);
nand (n3785,n3786,n3787);
or (n3786,n313,n3741);
or (n3787,n318,n3257);
nand (n3788,n3789,n3790);
or (n3789,n47,n3633);
or (n3790,n48,n3267);
nand (n3791,n3792,n3793);
or (n3792,n1085,n3273);
or (n3793,n3642,n1084);
or (n3794,n3795,n3796);
and (n3795,n3706,n3729);
and (n3796,n3707,n3708);
or (n3797,n3798,n4053);
and (n3798,n3799,n3839);
xor (n3799,n3800,n3838);
or (n3800,n3801,n3837);
and (n3801,n3802,n3836);
xor (n3802,n3803,n3804);
xor (n3803,n3710,n3725);
or (n3804,n3805,n3835);
and (n3805,n3806,n3821);
xor (n3806,n3807,n3813);
nand (n3807,n3808,n3812);
or (n3808,n1075,n3809);
nor (n3809,n3810,n3811);
and (n3810,n304,n415);
and (n3811,n302,n417);
or (n3812,n1080,n3672);
nand (n3813,n3814,n3819);
or (n3814,n3815,n410);
not (n3815,n3816);
nand (n3816,n3817,n3818);
or (n3817,n32,n891);
or (n3818,n31,n889);
nand (n3819,n3820,n619);
not (n3820,n3659);
and (n3821,n3822,n3828);
nor (n3822,n3823,n36);
nor (n3823,n3824,n3827);
and (n3824,n3825,n31);
not (n3825,n3826);
and (n3826,n1266,n30);
and (n3827,n1268,n39);
nand (n3828,n3829,n3834);
or (n3829,n1084,n3830);
not (n3830,n3831);
nor (n3831,n3832,n3833);
and (n3832,n310,n782);
and (n3833,n308,n783);
or (n3834,n3685,n1085);
and (n3835,n3807,n3813);
xor (n3836,n3656,n3679);
and (n3837,n3803,n3804);
xor (n3838,n3624,n3705);
or (n3839,n3840,n4052);
and (n3840,n3841,n3875);
xor (n3841,n3842,n3874);
or (n3842,n3843,n3873);
and (n3843,n3844,n3872);
xor (n3844,n3845,n3871);
or (n3845,n3846,n3870);
and (n3846,n3847,n3863);
xor (n3847,n3848,n3855);
nand (n3848,n3849,n3854);
or (n3849,n3850,n313);
not (n3850,n3851);
nand (n3851,n3852,n3853);
or (n3852,n36,n1266);
or (n3853,n1268,n37);
nand (n3854,n28,n3695);
nand (n3855,n3856,n3861);
or (n3856,n3857,n1075);
not (n3857,n3858);
nor (n3858,n3859,n3860);
and (n3859,n672,n417);
and (n3860,n670,n415);
nand (n3861,n3862,n779);
not (n3862,n3809);
nand (n3863,n3864,n3869);
or (n3864,n3865,n410);
not (n3865,n3866);
nor (n3866,n3867,n3868);
and (n3867,n1064,n32);
and (n3868,n1066,n31);
nand (n3869,n619,n3816);
and (n3870,n3848,n3855);
xor (n3871,n3681,n3692);
xor (n3872,n3806,n3821);
and (n3873,n3845,n3871);
xor (n3874,n3802,n3836);
nand (n3875,n3876,n4051);
or (n3876,n3877,n3907);
not (n3877,n3878);
nand (n3878,n3879,n3881);
not (n3879,n3880);
xor (n3880,n3844,n3872);
not (n3881,n3882);
or (n3882,n3883,n3906);
and (n3883,n3884,n3905);
xor (n3884,n3885,n3886);
xor (n3885,n3822,n3828);
or (n3886,n3887,n3904);
and (n3887,n3888,n3897);
xor (n3888,n3889,n3890);
and (n3889,n28,n1266);
nand (n3890,n3891,n3896);
or (n3891,n1084,n3892);
not (n3892,n3893);
nor (n3893,n3894,n3895);
and (n3894,n302,n783);
and (n3895,n304,n782);
nand (n3896,n3831,n1086);
nand (n3897,n3898,n3903);
or (n3898,n3899,n1075);
not (n3899,n3900);
nor (n3900,n3901,n3902);
and (n3901,n891,n417);
and (n3902,n889,n415);
nand (n3903,n779,n3858);
and (n3904,n3889,n3890);
xor (n3905,n3847,n3863);
and (n3906,n3885,n3886);
not (n3907,n3908);
nand (n3908,n3909,n4050);
or (n3909,n3910,n3940);
not (n3910,n3911);
nand (n3911,n3912,n3914);
not (n3912,n3913);
xor (n3913,n3884,n3905);
not (n3914,n3915);
or (n3915,n3916,n3939);
and (n3916,n3917,n3938);
xor (n3917,n3918,n3925);
nand (n3918,n3919,n3924);
or (n3919,n3920,n410);
not (n3920,n3921);
nor (n3921,n3922,n3923);
and (n3922,n1103,n32);
and (n3923,n1105,n31);
nand (n3924,n619,n3866);
and (n3925,n3926,n3931);
and (n3926,n3927,n32);
nand (n3927,n3928,n3930);
or (n3928,n3929,n415);
and (n3929,n1266,n414);
or (n3930,n1266,n414);
nand (n3931,n3932,n3933);
or (n3932,n1085,n3892);
nand (n3933,n3934,n1083);
not (n3934,n3935);
nor (n3935,n3936,n3937);
and (n3936,n670,n782);
and (n3937,n672,n783);
xor (n3938,n3888,n3897);
and (n3939,n3918,n3925);
not (n3940,n3941);
nand (n3941,n3942,n4049);
or (n3942,n3943,n3967);
not (n3943,n3944);
nand (n3944,n3945,n3947);
not (n3945,n3946);
xor (n3946,n3917,n3938);
not (n3947,n3948);
or (n3948,n3949,n3966);
and (n3949,n3950,n3965);
xor (n3950,n3951,n3958);
nand (n3951,n3952,n3957);
or (n3952,n3953,n1075);
not (n3953,n3954);
nor (n3954,n3955,n3956);
and (n3955,n1066,n417);
and (n3956,n1064,n415);
nand (n3957,n779,n3900);
nand (n3958,n3959,n3964);
or (n3959,n3960,n410);
not (n3960,n3961);
nand (n3961,n3962,n3963);
or (n3962,n31,n1266);
or (n3963,n32,n1268);
nand (n3964,n619,n3921);
xor (n3965,n3926,n3931);
and (n3966,n3951,n3958);
not (n3967,n3968);
nand (n3968,n3969,n4048);
or (n3969,n3970,n3994);
not (n3970,n3971);
nand (n3971,n3972,n3974);
not (n3972,n3973);
xor (n3973,n3950,n3965);
not (n3974,n3975);
or (n3975,n3976,n3993);
and (n3976,n3977,n3986);
xor (n3977,n3978,n3979);
and (n3978,n619,n1266);
nand (n3979,n3980,n3985);
or (n3980,n3981,n1075);
not (n3981,n3982);
nor (n3982,n3983,n3984);
and (n3983,n1103,n415);
and (n3984,n1105,n417);
nand (n3985,n779,n3954);
nand (n3986,n3987,n3992);
or (n3987,n1084,n3988);
not (n3988,n3989);
nor (n3989,n3990,n3991);
and (n3990,n891,n782);
and (n3991,n889,n783);
or (n3992,n3935,n1085);
and (n3993,n3978,n3979);
not (n3994,n3995);
nand (n3995,n3996,n4047);
or (n3996,n3997,n4013);
nor (n3997,n3998,n3999);
xor (n3998,n3977,n3986);
and (n3999,n4000,n4006);
nor (n4000,n4001,n417);
nor (n4001,n4002,n4003);
and (n4002,n789,n1268);
and (n4003,n4004,n782);
not (n4004,n4005);
and (n4005,n1266,n781);
nand (n4006,n4007,n4008);
or (n4007,n1085,n3988);
nand (n4008,n4009,n1083);
not (n4009,n4010);
nor (n4010,n4011,n4012);
and (n4011,n782,n1064);
and (n4012,n783,n1066);
not (n4013,n4014);
or (n4014,n4015,n4046);
and (n4015,n4016,n4025);
xor (n4016,n4017,n4024);
nand (n4017,n4018,n4023);
or (n4018,n4019,n1075);
not (n4019,n4020);
nand (n4020,n4021,n4022);
or (n4021,n417,n1266);
or (n4022,n415,n1268);
nand (n4023,n779,n3982);
xor (n4024,n4000,n4006);
or (n4025,n4026,n4045);
and (n4026,n4027,n4035);
xor (n4027,n4028,n4029);
nor (n4028,n1080,n1268);
nand (n4029,n4030,n4034);
or (n4030,n4031,n1084);
nor (n4031,n4032,n4033);
and (n4032,n782,n1103);
and (n4033,n783,n1105);
or (n4034,n4010,n1085);
nor (n4035,n4036,n4043);
nor (n4036,n4037,n4039);
and (n4037,n4038,n1086);
not (n4038,n4031);
nor (n4039,n4040,n1084);
nor (n4040,n4041,n4042);
and (n4041,n1266,n782);
and (n4042,n1268,n783);
or (n4043,n4044,n782);
and (n4044,n1266,n1086);
and (n4045,n4028,n4029);
and (n4046,n4017,n4024);
nand (n4047,n3998,n3999);
nand (n4048,n3973,n3975);
nand (n4049,n3946,n3948);
nand (n4050,n3913,n3915);
nand (n4051,n3880,n3882);
and (n4052,n3842,n3874);
and (n4053,n3800,n3838);
and (n4054,n3622,n3745);
nor (n4055,n4056,n4094);
not (n4056,n4057);
or (n4057,n4058,n4079);
xor (n4058,n4059,n4062);
xor (n4059,n4060,n4061);
xor (n4060,n3104,n3159);
xor (n4061,n3237,n3240);
or (n4062,n4063,n4078);
and (n4063,n4064,n4067);
xor (n4064,n4065,n4066);
xor (n4065,n3136,n3152);
xor (n4066,n3107,n3124);
or (n4067,n4068,n4077);
and (n4068,n4069,n4074);
xor (n4069,n4070,n4073);
nand (n4070,n4071,n4072);
or (n4071,n410,n3758);
or (n4072,n411,n3139);
nor (n4073,n3770,n3764);
or (n4074,n4075,n4076);
and (n4075,n3784,n3791);
and (n4076,n3785,n3788);
and (n4077,n4070,n4073);
and (n4078,n4065,n4066);
or (n4079,n4080,n4093);
and (n4080,n4081,n4092);
xor (n4081,n4082,n4083);
xor (n4082,n3242,n3262);
or (n4083,n4084,n4091);
and (n4084,n4085,n4088);
xor (n4085,n4086,n4087);
xor (n4086,n3264,n3278);
xor (n4087,n3246,n3255);
or (n4088,n4089,n4090);
and (n4089,n3748,n3761);
and (n4090,n3749,n3755);
and (n4091,n4086,n4087);
xor (n4092,n4064,n4067);
and (n4093,n4082,n4083);
nand (n4094,n4095,n4107);
not (n4095,n4096);
nor (n4096,n4097,n4098);
xor (n4097,n4081,n4092);
or (n4098,n4099,n4106);
and (n4099,n4100,n4105);
xor (n4100,n4101,n4102);
xor (n4101,n4069,n4074);
or (n4102,n4103,n4104);
and (n4103,n3776,n3783);
and (n4104,n3777,n3780);
xor (n4105,n4085,n4088);
and (n4106,n4101,n4102);
or (n4107,n4108,n4111);
or (n4108,n4109,n4110);
and (n4109,n3746,n3794);
and (n4110,n3747,n3775);
xor (n4111,n4100,n4105);
or (n4112,n4113,n4114);
xor (n4113,n3233,n3287);
or (n4114,n4115,n4116);
and (n4115,n4059,n4062);
and (n4116,n4060,n4061);
nand (n4117,n4118,n4112);
nand (n4118,n4119,n4125);
or (n4119,n4056,n4120);
not (n4120,n4121);
nand (n4121,n4122,n4124);
or (n4122,n4096,n4123);
nand (n4123,n4108,n4111);
nand (n4124,n4097,n4098);
nand (n4125,n4058,n4079);
nand (n4126,n4113,n4114);
and (n4127,n4128,n4294,n4325);
nand (n4128,n4129,n4262);
not (n4129,n4130);
xor (n4130,n4131,n4249);
xor (n4131,n4132,n4133);
xor (n4132,n2404,n2413);
or (n4133,n4134,n4248);
and (n4134,n4135,n4231);
xor (n4135,n4136,n4208);
or (n4136,n4137,n4207);
and (n4137,n4138,n4179);
xor (n4138,n4139,n4150);
or (n4139,n4140,n4149);
and (n4140,n4141,n4146);
xor (n4141,n4142,n4145);
nand (n4142,n4143,n4144);
or (n4143,n72,n3508);
or (n4144,n92,n2386);
and (n4145,n3512,n3518);
or (n4146,n4147,n4148);
and (n4147,n3577,n3592);
and (n4148,n3578,n3585);
and (n4149,n4142,n4145);
xor (n4150,n4151,n4178);
xor (n4151,n4152,n4167);
or (n4152,n4153,n4166);
and (n4153,n4154,n4163);
xor (n4154,n4155,n4160);
nand (n4155,n4156,n4158);
or (n4156,n4157,n410);
not (n4157,n3564);
nand (n4158,n4159,n619);
not (n4159,n2380);
nand (n4160,n4161,n4162);
or (n4161,n206,n3573);
or (n4162,n207,n2361);
nand (n4163,n4164,n4165);
or (n4164,n155,n3502);
or (n4165,n156,n2354);
and (n4166,n4155,n4160);
or (n4167,n4168,n4177);
and (n4168,n4169,n4174);
xor (n4169,n4170,n4171);
nor (n4170,n127,n1268);
nand (n4171,n4172,n4173);
or (n4172,n3520,n1075);
or (n4173,n1080,n2284);
nand (n4174,n4175,n4176);
or (n4175,n313,n3481);
or (n4176,n318,n2302);
and (n4177,n4170,n4171);
xor (n4178,n2371,n2384);
or (n4179,n4180,n4206);
and (n4180,n4181,n4195);
xor (n4181,n4182,n4194);
xor (n4182,n4183,n4191);
xor (n4183,n4184,n4188);
nand (n4184,n4185,n4186);
or (n4185,n3589,n344);
nand (n4186,n4187,n346);
not (n4187,n2331);
nand (n4188,n4189,n4190);
or (n4189,n179,n3595);
or (n4190,n188,n2338);
nand (n4191,n4192,n4193);
or (n4192,n1084,n3557);
or (n4193,n2348,n1085);
xor (n4194,n4169,n4174);
xor (n4195,n4196,n4203);
xor (n4196,n4197,n4200);
nand (n4197,n4198,n4199);
or (n4198,n228,n3488);
or (n4199,n229,n2309);
nand (n4200,n4201,n4202);
or (n4201,n260,n3494);
or (n4202,n278,n2315);
nand (n4203,n4204,n4205);
or (n4204,n47,n3580);
or (n4205,n48,n2325);
and (n4206,n4182,n4194);
and (n4207,n4139,n4150);
xor (n4208,n4209,n4224);
xor (n4209,n4210,n4221);
or (n4210,n4211,n4220);
and (n4211,n4212,n4217);
xor (n4212,n4213,n4214);
xor (n4213,n2276,n2282);
or (n4214,n4215,n4216);
and (n4215,n4196,n4203);
and (n4216,n4197,n4200);
or (n4217,n4218,n4219);
and (n4218,n4183,n4191);
and (n4219,n4184,n4188);
and (n4220,n4213,n4214);
or (n4221,n4222,n4223);
and (n4222,n4151,n4178);
and (n4223,n4152,n4167);
or (n4224,n4225,n4230);
and (n4225,n4226,n4229);
xor (n4226,n4227,n4228);
xor (n4227,n2299,n2313);
xor (n4228,n2322,n2336);
xor (n4229,n2345,n2358);
and (n4230,n4227,n4228);
or (n4231,n4232,n4247);
and (n4232,n4233,n4246);
xor (n4233,n4234,n4245);
or (n4234,n4235,n4244);
and (n4235,n4236,n4243);
xor (n4236,n4237,n4240);
or (n4237,n4238,n4239);
and (n4238,n3553,n3567);
and (n4239,n3554,n3560);
or (n4240,n4241,n4242);
and (n4241,n3475,n3491);
and (n4242,n3476,n3484);
xor (n4243,n4154,n4163);
and (n4244,n4237,n4240);
xor (n4245,n4212,n4217);
xor (n4246,n4226,n4229);
and (n4247,n4234,n4245);
and (n4248,n4136,n4208);
xor (n4249,n4250,n4261);
xor (n4250,n4251,n4254);
or (n4251,n4252,n4253);
and (n4252,n4209,n4224);
and (n4253,n4210,n4221);
or (n4254,n4255,n4260);
and (n4255,n4256,n4259);
xor (n4256,n4257,n4258);
xor (n4257,n2296,n2343);
xor (n4258,n2407,n2410);
xor (n4259,n2368,n2392);
and (n4260,n4257,n4258);
xor (n4261,n2293,n2394);
not (n4262,n4263);
or (n4263,n4264,n4293);
and (n4264,n4265,n4292);
xor (n4265,n4266,n4267);
xor (n4266,n4256,n4259);
or (n4267,n4268,n4291);
and (n4268,n4269,n4290);
xor (n4269,n4270,n4281);
or (n4270,n4271,n4280);
and (n4271,n4272,n4279);
xor (n4272,n4273,n4276);
or (n4273,n4274,n4275);
and (n4274,n3498,n3511);
and (n4275,n3499,n3505);
or (n4276,n4277,n4278);
and (n4277,n3534,n3541);
and (n4278,n3535,n3538);
xor (n4279,n4141,n4146);
and (n4280,n4273,n4276);
or (n4281,n4282,n4289);
and (n4282,n4283,n4288);
xor (n4283,n4284,n4285);
xor (n4284,n4236,n4243);
or (n4285,n4286,n4287);
and (n4286,n3548,n3576);
and (n4287,n3549,n3552);
xor (n4288,n4181,n4195);
and (n4289,n4284,n4285);
xor (n4290,n4138,n4179);
and (n4291,n4270,n4281);
xor (n4292,n4135,n4231);
and (n4293,n4266,n4267);
nor (n4294,n4295,n4314);
nor (n4295,n4296,n4311);
xor (n4296,n4297,n4308);
xor (n4297,n4298,n4299);
xor (n4298,n4283,n4288);
xor (n4299,n4300,n4305);
xor (n4300,n4301,n4304);
or (n4301,n4302,n4303);
and (n4302,n3473,n3525);
and (n4303,n3474,n3497);
xor (n4304,n4272,n4279);
or (n4305,n4306,n4307);
and (n4306,n3532,n3547);
and (n4307,n3533,n3544);
or (n4308,n4309,n4310);
and (n4309,n3471,n3531);
and (n4310,n3472,n3528);
or (n4311,n4312,n4313);
and (n4312,n3463,n3470);
and (n4313,n3464,n3467);
nor (n4314,n4315,n4318);
or (n4315,n4316,n4317);
and (n4316,n4297,n4308);
and (n4317,n4298,n4299);
xor (n4318,n4319,n4324);
xor (n4319,n4320,n4321);
xor (n4320,n4233,n4246);
or (n4321,n4322,n4323);
and (n4322,n4300,n4305);
and (n4323,n4301,n4304);
xor (n4324,n4269,n4290);
not (n4325,n4326);
nor (n4326,n4327,n4328);
xor (n4327,n4265,n4292);
or (n4328,n4329,n4330);
and (n4329,n4319,n4324);
and (n4330,n4320,n4321);
nor (n4331,n4332,n4343);
nor (n4332,n4333,n4334);
xor (n4333,n2251,n2416);
or (n4334,n4335,n4342);
and (n4335,n4336,n4341);
xor (n4336,n4337,n4338);
xor (n4337,n2254,n2291);
or (n4338,n4339,n4340);
and (n4339,n4250,n4261);
and (n4340,n4251,n4254);
xor (n4341,n2399,n2402);
and (n4342,n4337,n4338);
nor (n4343,n4344,n4345);
xor (n4344,n4336,n4341);
or (n4345,n4346,n4347);
and (n4346,n4131,n4249);
and (n4347,n4132,n4133);
nand (n4348,n4349,n2231,n4331);
nand (n4349,n4350,n4360);
or (n4350,n4351,n4352);
not (n4351,n4128);
not (n4352,n4353);
nand (n4353,n4354,n4359);
or (n4354,n4355,n4326);
nor (n4355,n4356,n4358);
nor (n4356,n4314,n4357);
nand (n4357,n4296,n4311);
and (n4358,n4315,n4318);
nand (n4359,n4327,n4328);
nand (n4360,n4130,n4263);
nor (n4361,n4362,n4367);
and (n4362,n2231,n4363);
nand (n4363,n4364,n4366);
or (n4364,n4332,n4365);
nand (n4365,n4344,n4345);
nand (n4366,n4333,n4334);
nand (n4367,n4368,n4370);
or (n4368,n2232,n4369);
nand (n4369,n2248,n2249);
nand (n4370,n2233,n2234);
not (n4371,n4372);
nand (n4372,n4373,n4380);
or (n4373,n4374,n4379);
not (n4374,n4375);
nand (n4375,n4376,n4378);
or (n4376,n1799,n4377);
nand (n4377,n2092,n2227);
nand (n4378,n1800,n1801);
not (n4379,n1591);
nor (n4380,n4381,n4385);
and (n4381,n4382,n4383);
not (n4382,n1592);
not (n4383,n4384);
nand (n4384,n1784,n1797);
and (n4385,n1593,n1594);
not (n4386,n4387);
nand (n4387,n4388,n4390);
or (n4388,n1582,n4389);
nand (n4389,n1152,n1235);
nand (n4390,n1583,n1584);
or (n4391,n1147,n15);
or (n4392,n4393,n8418);
and (n4393,n4394,n8417);
wire s0n4394,s1n4394,notn4394;
or (n4394,s0n4394,s1n4394);
not(notn4394,n10);
and (s0n4394,notn4394,n3);
and (s1n4394,n10,n4395);
xor (n4395,n4396,n8329);
xor (n4396,n4397,n8415);
xor (n4397,n4398,n8324);
xor (n4398,n4399,n8408);
xor (n4399,n4400,n8318);
xor (n4400,n4401,n8396);
xor (n4401,n4402,n8312);
xor (n4402,n4403,n8379);
xor (n4403,n4404,n8306);
xor (n4404,n4405,n8357);
xor (n4405,n4406,n8300);
xor (n4406,n4407,n8330);
xor (n4407,n4408,n8294);
xor (n4408,n4409,n8291);
xor (n4409,n4410,n8290);
xor (n4410,n4411,n8246);
xor (n4411,n4412,n8245);
xor (n4412,n4413,n8194);
xor (n4413,n4414,n8193);
xor (n4414,n4415,n8137);
xor (n4415,n4416,n8136);
xor (n4416,n4417,n8073);
xor (n4417,n4418,n8072);
xor (n4418,n4419,n8004);
xor (n4419,n4420,n8003);
xor (n4420,n4421,n7930);
xor (n4421,n4422,n7929);
xor (n4422,n4423,n7849);
xor (n4423,n4424,n7848);
xor (n4424,n4425,n7761);
xor (n4425,n4426,n7760);
xor (n4426,n4427,n7668);
xor (n4427,n4428,n7667);
xor (n4428,n4429,n7568);
xor (n4429,n4430,n7567);
xor (n4430,n4431,n7463);
xor (n4431,n4432,n7462);
xor (n4432,n4433,n7355);
xor (n4433,n4434,n7354);
xor (n4434,n4435,n7238);
xor (n4435,n4436,n7237);
xor (n4436,n4437,n7114);
xor (n4437,n4438,n7113);
xor (n4438,n4439,n6985);
xor (n4439,n4440,n6984);
xor (n4440,n4441,n6851);
xor (n4441,n4442,n6850);
xor (n4442,n4443,n6710);
xor (n4443,n4444,n6709);
xor (n4444,n4445,n6562);
xor (n4445,n4446,n6561);
xor (n4446,n4447,n6409);
xor (n4447,n4448,n6408);
xor (n4448,n4449,n6250);
xor (n4449,n4450,n6249);
xor (n4450,n4451,n6085);
xor (n4451,n4452,n6084);
xor (n4452,n4453,n5915);
xor (n4453,n4454,n5914);
xor (n4454,n4455,n5738);
xor (n4455,n4456,n5737);
xor (n4456,n4457,n4482);
xor (n4457,n4458,n4481);
xor (n4458,n4459,n4480);
xor (n4459,n4460,n4479);
xor (n4460,n4461,n4478);
xor (n4461,n4462,n4477);
xor (n4462,n4463,n4476);
xor (n4463,n4464,n4475);
xor (n4464,n4465,n4474);
xor (n4465,n4466,n791);
xor (n4466,n4467,n4473);
xor (n4467,n4468,n4472);
xor (n4468,n4469,n4471);
xor (n4469,n4470,n1088);
and (n4470,n43,n1086);
and (n4471,n4470,n1088);
and (n4472,n43,n781);
and (n4473,n4468,n4472);
and (n4474,n4466,n791);
and (n4475,n43,n414);
and (n4476,n4464,n4475);
and (n4477,n43,n32);
and (n4478,n4462,n4477);
and (n4479,n43,n30);
and (n4480,n4460,n4479);
and (n4481,n43,n37);
or (n4482,n4483,n5564);
and (n4483,n4484,n5563);
xor (n4484,n4459,n4485);
or (n4485,n4486,n5385);
and (n4486,n4487,n5384);
xor (n4487,n4461,n4488);
or (n4488,n4489,n5210);
and (n4489,n4490,n5209);
xor (n4490,n4463,n4491);
or (n4491,n4492,n5031);
and (n4492,n4493,n5030);
xor (n4493,n4465,n4494);
or (n4494,n4495,n4857);
and (n4495,n4496,n4856);
xor (n4496,n4467,n4497);
or (n4497,n4498,n4678);
and (n4498,n4499,n4677);
xor (n4499,n4469,n4500);
or (n4500,n4501,n4503);
and (n4501,n4470,n4502);
and (n4502,n67,n783);
and (n4503,n4504,n4505);
xor (n4504,n4470,n4502);
or (n4505,n4506,n4508);
and (n4506,n4507,n1535);
and (n4507,n67,n1086);
and (n4508,n4509,n4510);
xor (n4509,n4507,n1535);
or (n4510,n4511,n4514);
and (n4511,n4512,n4513);
and (n4512,n61,n1086);
and (n4513,n172,n783);
and (n4514,n4515,n4516);
xor (n4515,n4512,n4513);
or (n4516,n4517,n4520);
and (n4517,n4518,n4519);
and (n4518,n172,n1086);
and (n4519,n166,n783);
and (n4520,n4521,n4522);
xor (n4521,n4518,n4519);
or (n4522,n4523,n4526);
and (n4523,n4524,n4525);
and (n4524,n166,n1086);
and (n4525,n95,n783);
and (n4526,n4527,n4528);
xor (n4527,n4524,n4525);
or (n4528,n4529,n4532);
and (n4529,n4530,n4531);
and (n4530,n95,n1086);
and (n4531,n88,n783);
and (n4532,n4533,n4534);
xor (n4533,n4530,n4531);
or (n4534,n4535,n4538);
and (n4535,n4536,n4537);
and (n4536,n88,n1086);
and (n4537,n249,n783);
and (n4538,n4539,n4540);
xor (n4539,n4536,n4537);
or (n4540,n4541,n4544);
and (n4541,n4542,n4543);
and (n4542,n249,n1086);
and (n4543,n243,n783);
and (n4544,n4545,n4546);
xor (n4545,n4542,n4543);
or (n4546,n4547,n4550);
and (n4547,n4548,n4549);
and (n4548,n243,n1086);
and (n4549,n377,n783);
and (n4550,n4551,n4552);
xor (n4551,n4548,n4549);
or (n4552,n4553,n4556);
and (n4553,n4554,n4555);
and (n4554,n377,n1086);
and (n4555,n436,n783);
and (n4556,n4557,n4558);
xor (n4557,n4554,n4555);
or (n4558,n4559,n4562);
and (n4559,n4560,n4561);
and (n4560,n436,n1086);
and (n4561,n281,n783);
and (n4562,n4563,n4564);
xor (n4563,n4560,n4561);
or (n4564,n4565,n4568);
and (n4565,n4566,n4567);
and (n4566,n281,n1086);
and (n4567,n274,n783);
and (n4568,n4569,n4570);
xor (n4569,n4566,n4567);
or (n4570,n4571,n4574);
and (n4571,n4572,n4573);
and (n4572,n274,n1086);
and (n4573,n201,n783);
and (n4574,n4575,n4576);
xor (n4575,n4572,n4573);
or (n4576,n4577,n4580);
and (n4577,n4578,n4579);
and (n4578,n201,n1086);
and (n4579,n195,n783);
and (n4580,n4581,n4582);
xor (n4581,n4578,n4579);
or (n4582,n4583,n4586);
and (n4583,n4584,n4585);
and (n4584,n195,n1086);
and (n4585,n223,n783);
and (n4586,n4587,n4588);
xor (n4587,n4584,n4585);
or (n4588,n4589,n4592);
and (n4589,n4590,n4591);
and (n4590,n223,n1086);
and (n4591,n217,n783);
and (n4592,n4593,n4594);
xor (n4593,n4590,n4591);
or (n4594,n4595,n4598);
and (n4595,n4596,n4597);
and (n4596,n217,n1086);
and (n4597,n124,n783);
and (n4598,n4599,n4600);
xor (n4599,n4596,n4597);
or (n4600,n4601,n4604);
and (n4601,n4602,n4603);
and (n4602,n124,n1086);
and (n4603,n118,n783);
and (n4604,n4605,n4606);
xor (n4605,n4602,n4603);
or (n4606,n4607,n4610);
and (n4607,n4608,n4609);
and (n4608,n118,n1086);
and (n4609,n150,n783);
and (n4610,n4611,n4612);
xor (n4611,n4608,n4609);
or (n4612,n4613,n4615);
and (n4613,n4614,n3275);
and (n4614,n150,n1086);
and (n4615,n4616,n4617);
xor (n4616,n4614,n3275);
or (n4617,n4618,n4621);
and (n4618,n4619,n4620);
and (n4619,n144,n1086);
and (n4620,n398,n783);
and (n4621,n4622,n4623);
xor (n4622,n4619,n4620);
or (n4623,n4624,n4627);
and (n4624,n4625,n4626);
and (n4625,n398,n1086);
and (n4626,n449,n783);
and (n4627,n4628,n4629);
xor (n4628,n4625,n4626);
or (n4629,n4630,n4633);
and (n4630,n4631,n4632);
and (n4631,n449,n1086);
and (n4632,n443,n783);
and (n4633,n4634,n4635);
xor (n4634,n4631,n4632);
or (n4635,n4636,n4639);
and (n4636,n4637,n4638);
and (n4637,n443,n1086);
and (n4638,n551,n783);
and (n4639,n4640,n4641);
xor (n4640,n4637,n4638);
or (n4641,n4642,n4644);
and (n4642,n4643,n3833);
and (n4643,n551,n1086);
and (n4644,n4645,n4646);
xor (n4645,n4643,n3833);
or (n4646,n4647,n4649);
and (n4647,n4648,n3894);
and (n4648,n308,n1086);
and (n4649,n4650,n4651);
xor (n4650,n4648,n3894);
or (n4651,n4652,n4655);
and (n4652,n4653,n4654);
and (n4653,n302,n1086);
and (n4654,n670,n783);
and (n4655,n4656,n4657);
xor (n4656,n4653,n4654);
or (n4657,n4658,n4660);
and (n4658,n4659,n3991);
and (n4659,n670,n1086);
and (n4660,n4661,n4662);
xor (n4661,n4659,n3991);
or (n4662,n4663,n4666);
and (n4663,n4664,n4665);
and (n4664,n889,n1086);
and (n4665,n1064,n783);
and (n4666,n4667,n4668);
xor (n4667,n4664,n4665);
or (n4668,n4669,n4672);
and (n4669,n4670,n4671);
and (n4670,n1064,n1086);
and (n4671,n1103,n783);
and (n4672,n4673,n4674);
xor (n4673,n4670,n4671);
and (n4674,n4675,n4676);
and (n4675,n1103,n1086);
and (n4676,n1266,n783);
and (n4677,n67,n781);
and (n4678,n4679,n4680);
xor (n4679,n4499,n4677);
or (n4680,n4681,n4684);
and (n4681,n4682,n4683);
xor (n4682,n4504,n4505);
and (n4683,n61,n781);
and (n4684,n4685,n4686);
xor (n4685,n4682,n4683);
or (n4686,n4687,n4690);
and (n4687,n4688,n4689);
xor (n4688,n4509,n4510);
and (n4689,n172,n781);
and (n4690,n4691,n4692);
xor (n4691,n4688,n4689);
or (n4692,n4693,n4696);
and (n4693,n4694,n4695);
xor (n4694,n4515,n4516);
and (n4695,n166,n781);
and (n4696,n4697,n4698);
xor (n4697,n4694,n4695);
or (n4698,n4699,n4702);
and (n4699,n4700,n4701);
xor (n4700,n4521,n4522);
and (n4701,n95,n781);
and (n4702,n4703,n4704);
xor (n4703,n4700,n4701);
or (n4704,n4705,n4708);
and (n4705,n4706,n4707);
xor (n4706,n4527,n4528);
and (n4707,n88,n781);
and (n4708,n4709,n4710);
xor (n4709,n4706,n4707);
or (n4710,n4711,n4714);
and (n4711,n4712,n4713);
xor (n4712,n4533,n4534);
and (n4713,n249,n781);
and (n4714,n4715,n4716);
xor (n4715,n4712,n4713);
or (n4716,n4717,n4720);
and (n4717,n4718,n4719);
xor (n4718,n4539,n4540);
and (n4719,n243,n781);
and (n4720,n4721,n4722);
xor (n4721,n4718,n4719);
or (n4722,n4723,n4726);
and (n4723,n4724,n4725);
xor (n4724,n4545,n4546);
and (n4725,n377,n781);
and (n4726,n4727,n4728);
xor (n4727,n4724,n4725);
or (n4728,n4729,n4732);
and (n4729,n4730,n4731);
xor (n4730,n4551,n4552);
and (n4731,n436,n781);
and (n4732,n4733,n4734);
xor (n4733,n4730,n4731);
or (n4734,n4735,n4738);
and (n4735,n4736,n4737);
xor (n4736,n4557,n4558);
and (n4737,n281,n781);
and (n4738,n4739,n4740);
xor (n4739,n4736,n4737);
or (n4740,n4741,n4744);
and (n4741,n4742,n4743);
xor (n4742,n4563,n4564);
and (n4743,n274,n781);
and (n4744,n4745,n4746);
xor (n4745,n4742,n4743);
or (n4746,n4747,n4750);
and (n4747,n4748,n4749);
xor (n4748,n4569,n4570);
and (n4749,n201,n781);
and (n4750,n4751,n4752);
xor (n4751,n4748,n4749);
or (n4752,n4753,n4756);
and (n4753,n4754,n4755);
xor (n4754,n4575,n4576);
and (n4755,n195,n781);
and (n4756,n4757,n4758);
xor (n4757,n4754,n4755);
or (n4758,n4759,n4762);
and (n4759,n4760,n4761);
xor (n4760,n4581,n4582);
and (n4761,n223,n781);
and (n4762,n4763,n4764);
xor (n4763,n4760,n4761);
or (n4764,n4765,n4768);
and (n4765,n4766,n4767);
xor (n4766,n4587,n4588);
and (n4767,n217,n781);
and (n4768,n4769,n4770);
xor (n4769,n4766,n4767);
or (n4770,n4771,n4774);
and (n4771,n4772,n4773);
xor (n4772,n4593,n4594);
and (n4773,n124,n781);
and (n4774,n4775,n4776);
xor (n4775,n4772,n4773);
or (n4776,n4777,n4780);
and (n4777,n4778,n4779);
xor (n4778,n4599,n4600);
and (n4779,n118,n781);
and (n4780,n4781,n4782);
xor (n4781,n4778,n4779);
or (n4782,n4783,n4786);
and (n4783,n4784,n4785);
xor (n4784,n4605,n4606);
and (n4785,n150,n781);
and (n4786,n4787,n4788);
xor (n4787,n4784,n4785);
or (n4788,n4789,n4792);
and (n4789,n4790,n4791);
xor (n4790,n4611,n4612);
and (n4791,n144,n781);
and (n4792,n4793,n4794);
xor (n4793,n4790,n4791);
or (n4794,n4795,n4798);
and (n4795,n4796,n4797);
xor (n4796,n4616,n4617);
and (n4797,n398,n781);
and (n4798,n4799,n4800);
xor (n4799,n4796,n4797);
or (n4800,n4801,n4804);
and (n4801,n4802,n4803);
xor (n4802,n4622,n4623);
and (n4803,n449,n781);
and (n4804,n4805,n4806);
xor (n4805,n4802,n4803);
or (n4806,n4807,n4810);
and (n4807,n4808,n4809);
xor (n4808,n4628,n4629);
and (n4809,n443,n781);
and (n4810,n4811,n4812);
xor (n4811,n4808,n4809);
or (n4812,n4813,n4816);
and (n4813,n4814,n4815);
xor (n4814,n4634,n4635);
and (n4815,n551,n781);
and (n4816,n4817,n4818);
xor (n4817,n4814,n4815);
or (n4818,n4819,n4822);
and (n4819,n4820,n4821);
xor (n4820,n4640,n4641);
and (n4821,n308,n781);
and (n4822,n4823,n4824);
xor (n4823,n4820,n4821);
or (n4824,n4825,n4828);
and (n4825,n4826,n4827);
xor (n4826,n4645,n4646);
and (n4827,n302,n781);
and (n4828,n4829,n4830);
xor (n4829,n4826,n4827);
or (n4830,n4831,n4834);
and (n4831,n4832,n4833);
xor (n4832,n4650,n4651);
and (n4833,n670,n781);
and (n4834,n4835,n4836);
xor (n4835,n4832,n4833);
or (n4836,n4837,n4840);
and (n4837,n4838,n4839);
xor (n4838,n4656,n4657);
and (n4839,n889,n781);
and (n4840,n4841,n4842);
xor (n4841,n4838,n4839);
or (n4842,n4843,n4846);
and (n4843,n4844,n4845);
xor (n4844,n4661,n4662);
and (n4845,n1064,n781);
and (n4846,n4847,n4848);
xor (n4847,n4844,n4845);
or (n4848,n4849,n4852);
and (n4849,n4850,n4851);
xor (n4850,n4667,n4668);
and (n4851,n1103,n781);
and (n4852,n4853,n4854);
xor (n4853,n4850,n4851);
and (n4854,n4855,n4005);
xor (n4855,n4673,n4674);
and (n4856,n67,n415);
and (n4857,n4858,n4859);
xor (n4858,n4496,n4856);
or (n4859,n4860,n4863);
and (n4860,n4861,n4862);
xor (n4861,n4679,n4680);
and (n4862,n61,n415);
and (n4863,n4864,n4865);
xor (n4864,n4861,n4862);
or (n4865,n4866,n4868);
and (n4866,n4867,n1288);
xor (n4867,n4685,n4686);
and (n4868,n4869,n4870);
xor (n4869,n4867,n1288);
or (n4870,n4871,n4874);
and (n4871,n4872,n4873);
xor (n4872,n4691,n4692);
and (n4873,n166,n415);
and (n4874,n4875,n4876);
xor (n4875,n4872,n4873);
or (n4876,n4877,n4880);
and (n4877,n4878,n4879);
xor (n4878,n4697,n4698);
and (n4879,n95,n415);
and (n4880,n4881,n4882);
xor (n4881,n4878,n4879);
or (n4882,n4883,n4886);
and (n4883,n4884,n4885);
xor (n4884,n4703,n4704);
and (n4885,n88,n415);
and (n4886,n4887,n4888);
xor (n4887,n4884,n4885);
or (n4888,n4889,n4892);
and (n4889,n4890,n4891);
xor (n4890,n4709,n4710);
and (n4891,n249,n415);
and (n4892,n4893,n4894);
xor (n4893,n4890,n4891);
or (n4894,n4895,n4898);
and (n4895,n4896,n4897);
xor (n4896,n4715,n4716);
and (n4897,n243,n415);
and (n4898,n4899,n4900);
xor (n4899,n4896,n4897);
or (n4900,n4901,n4904);
and (n4901,n4902,n4903);
xor (n4902,n4721,n4722);
and (n4903,n377,n415);
and (n4904,n4905,n4906);
xor (n4905,n4902,n4903);
or (n4906,n4907,n4910);
and (n4907,n4908,n4909);
xor (n4908,n4727,n4728);
and (n4909,n436,n415);
and (n4910,n4911,n4912);
xor (n4911,n4908,n4909);
or (n4912,n4913,n4916);
and (n4913,n4914,n4915);
xor (n4914,n4733,n4734);
and (n4915,n281,n415);
and (n4916,n4917,n4918);
xor (n4917,n4914,n4915);
or (n4918,n4919,n4921);
and (n4919,n4920,n2771);
xor (n4920,n4739,n4740);
and (n4921,n4922,n4923);
xor (n4922,n4920,n2771);
or (n4923,n4924,n4927);
and (n4924,n4925,n4926);
xor (n4925,n4745,n4746);
and (n4926,n201,n415);
and (n4927,n4928,n4929);
xor (n4928,n4925,n4926);
or (n4929,n4930,n4933);
and (n4930,n4931,n4932);
xor (n4931,n4751,n4752);
and (n4932,n195,n415);
and (n4933,n4934,n4935);
xor (n4934,n4931,n4932);
or (n4935,n4936,n4939);
and (n4936,n4937,n4938);
xor (n4937,n4757,n4758);
and (n4938,n223,n415);
and (n4939,n4940,n4941);
xor (n4940,n4937,n4938);
or (n4941,n4942,n4945);
and (n4942,n4943,n4944);
xor (n4943,n4763,n4764);
and (n4944,n217,n415);
and (n4945,n4946,n4947);
xor (n4946,n4943,n4944);
or (n4947,n4948,n4951);
and (n4948,n4949,n4950);
xor (n4949,n4769,n4770);
and (n4950,n124,n415);
and (n4951,n4952,n4953);
xor (n4952,n4949,n4950);
or (n4953,n4954,n4957);
and (n4954,n4955,n4956);
xor (n4955,n4775,n4776);
and (n4956,n118,n415);
and (n4957,n4958,n4959);
xor (n4958,n4955,n4956);
or (n4959,n4960,n4963);
and (n4960,n4961,n4962);
xor (n4961,n4781,n4782);
and (n4962,n150,n415);
and (n4963,n4964,n4965);
xor (n4964,n4961,n4962);
or (n4965,n4966,n4969);
and (n4966,n4967,n4968);
xor (n4967,n4787,n4788);
and (n4968,n144,n415);
and (n4969,n4970,n4971);
xor (n4970,n4967,n4968);
or (n4971,n4972,n4975);
and (n4972,n4973,n4974);
xor (n4973,n4793,n4794);
and (n4974,n398,n415);
and (n4975,n4976,n4977);
xor (n4976,n4973,n4974);
or (n4977,n4978,n4981);
and (n4978,n4979,n4980);
xor (n4979,n4799,n4800);
and (n4980,n449,n415);
and (n4981,n4982,n4983);
xor (n4982,n4979,n4980);
or (n4983,n4984,n4987);
and (n4984,n4985,n4986);
xor (n4985,n4805,n4806);
and (n4986,n443,n415);
and (n4987,n4988,n4989);
xor (n4988,n4985,n4986);
or (n4989,n4990,n4993);
and (n4990,n4991,n4992);
xor (n4991,n4811,n4812);
and (n4992,n551,n415);
and (n4993,n4994,n4995);
xor (n4994,n4991,n4992);
or (n4995,n4996,n4999);
and (n4996,n4997,n4998);
xor (n4997,n4817,n4818);
and (n4998,n308,n415);
and (n4999,n5000,n5001);
xor (n5000,n4997,n4998);
or (n5001,n5002,n5005);
and (n5002,n5003,n5004);
xor (n5003,n4823,n4824);
and (n5004,n302,n415);
and (n5005,n5006,n5007);
xor (n5006,n5003,n5004);
or (n5007,n5008,n5010);
and (n5008,n5009,n3860);
xor (n5009,n4829,n4830);
and (n5010,n5011,n5012);
xor (n5011,n5009,n3860);
or (n5012,n5013,n5015);
and (n5013,n5014,n3902);
xor (n5014,n4835,n4836);
and (n5015,n5016,n5017);
xor (n5016,n5014,n3902);
or (n5017,n5018,n5020);
and (n5018,n5019,n3956);
xor (n5019,n4841,n4842);
and (n5020,n5021,n5022);
xor (n5021,n5019,n3956);
or (n5022,n5023,n5025);
and (n5023,n5024,n3983);
xor (n5024,n4847,n4848);
and (n5025,n5026,n5027);
xor (n5026,n5024,n3983);
and (n5027,n5028,n5029);
xor (n5028,n4853,n4854);
and (n5029,n1266,n415);
and (n5030,n67,n414);
and (n5031,n5032,n5033);
xor (n5032,n4493,n5030);
or (n5033,n5034,n5037);
and (n5034,n5035,n5036);
xor (n5035,n4858,n4859);
and (n5036,n61,n414);
and (n5037,n5038,n5039);
xor (n5038,n5035,n5036);
or (n5039,n5040,n5043);
and (n5040,n5041,n5042);
xor (n5041,n4864,n4865);
and (n5042,n172,n414);
and (n5043,n5044,n5045);
xor (n5044,n5041,n5042);
or (n5045,n5046,n5049);
and (n5046,n5047,n5048);
xor (n5047,n4869,n4870);
and (n5048,n166,n414);
and (n5049,n5050,n5051);
xor (n5050,n5047,n5048);
or (n5051,n5052,n5055);
and (n5052,n5053,n5054);
xor (n5053,n4875,n4876);
and (n5054,n95,n414);
and (n5055,n5056,n5057);
xor (n5056,n5053,n5054);
or (n5057,n5058,n5061);
and (n5058,n5059,n5060);
xor (n5059,n4881,n4882);
and (n5060,n88,n414);
and (n5061,n5062,n5063);
xor (n5062,n5059,n5060);
or (n5063,n5064,n5067);
and (n5064,n5065,n5066);
xor (n5065,n4887,n4888);
and (n5066,n249,n414);
and (n5067,n5068,n5069);
xor (n5068,n5065,n5066);
or (n5069,n5070,n5073);
and (n5070,n5071,n5072);
xor (n5071,n4893,n4894);
and (n5072,n243,n414);
and (n5073,n5074,n5075);
xor (n5074,n5071,n5072);
or (n5075,n5076,n5079);
and (n5076,n5077,n5078);
xor (n5077,n4899,n4900);
and (n5078,n377,n414);
and (n5079,n5080,n5081);
xor (n5080,n5077,n5078);
or (n5081,n5082,n5085);
and (n5082,n5083,n5084);
xor (n5083,n4905,n4906);
and (n5084,n436,n414);
and (n5085,n5086,n5087);
xor (n5086,n5083,n5084);
or (n5087,n5088,n5091);
and (n5088,n5089,n5090);
xor (n5089,n4911,n4912);
and (n5090,n281,n414);
and (n5091,n5092,n5093);
xor (n5092,n5089,n5090);
or (n5093,n5094,n5097);
and (n5094,n5095,n5096);
xor (n5095,n4917,n4918);
and (n5096,n274,n414);
and (n5097,n5098,n5099);
xor (n5098,n5095,n5096);
or (n5099,n5100,n5103);
and (n5100,n5101,n5102);
xor (n5101,n4922,n4923);
and (n5102,n201,n414);
and (n5103,n5104,n5105);
xor (n5104,n5101,n5102);
or (n5105,n5106,n5109);
and (n5106,n5107,n5108);
xor (n5107,n4928,n4929);
and (n5108,n195,n414);
and (n5109,n5110,n5111);
xor (n5110,n5107,n5108);
or (n5111,n5112,n5115);
and (n5112,n5113,n5114);
xor (n5113,n4934,n4935);
and (n5114,n223,n414);
and (n5115,n5116,n5117);
xor (n5116,n5113,n5114);
or (n5117,n5118,n5121);
and (n5118,n5119,n5120);
xor (n5119,n4940,n4941);
and (n5120,n217,n414);
and (n5121,n5122,n5123);
xor (n5122,n5119,n5120);
or (n5123,n5124,n5127);
and (n5124,n5125,n5126);
xor (n5125,n4946,n4947);
and (n5126,n124,n414);
and (n5127,n5128,n5129);
xor (n5128,n5125,n5126);
or (n5129,n5130,n5133);
and (n5130,n5131,n5132);
xor (n5131,n4952,n4953);
and (n5132,n118,n414);
and (n5133,n5134,n5135);
xor (n5134,n5131,n5132);
or (n5135,n5136,n5139);
and (n5136,n5137,n5138);
xor (n5137,n4958,n4959);
and (n5138,n150,n414);
and (n5139,n5140,n5141);
xor (n5140,n5137,n5138);
or (n5141,n5142,n5145);
and (n5142,n5143,n5144);
xor (n5143,n4964,n4965);
and (n5144,n144,n414);
and (n5145,n5146,n5147);
xor (n5146,n5143,n5144);
or (n5147,n5148,n5151);
and (n5148,n5149,n5150);
xor (n5149,n4970,n4971);
and (n5150,n398,n414);
and (n5151,n5152,n5153);
xor (n5152,n5149,n5150);
or (n5153,n5154,n5157);
and (n5154,n5155,n5156);
xor (n5155,n4976,n4977);
and (n5156,n449,n414);
and (n5157,n5158,n5159);
xor (n5158,n5155,n5156);
or (n5159,n5160,n5163);
and (n5160,n5161,n5162);
xor (n5161,n4982,n4983);
and (n5162,n443,n414);
and (n5163,n5164,n5165);
xor (n5164,n5161,n5162);
or (n5165,n5166,n5169);
and (n5166,n5167,n5168);
xor (n5167,n4988,n4989);
and (n5168,n551,n414);
and (n5169,n5170,n5171);
xor (n5170,n5167,n5168);
or (n5171,n5172,n5175);
and (n5172,n5173,n5174);
xor (n5173,n4994,n4995);
and (n5174,n308,n414);
and (n5175,n5176,n5177);
xor (n5176,n5173,n5174);
or (n5177,n5178,n5181);
and (n5178,n5179,n5180);
xor (n5179,n5000,n5001);
and (n5180,n302,n414);
and (n5181,n5182,n5183);
xor (n5182,n5179,n5180);
or (n5183,n5184,n5187);
and (n5184,n5185,n5186);
xor (n5185,n5006,n5007);
and (n5186,n670,n414);
and (n5187,n5188,n5189);
xor (n5188,n5185,n5186);
or (n5189,n5190,n5193);
and (n5190,n5191,n5192);
xor (n5191,n5011,n5012);
and (n5192,n889,n414);
and (n5193,n5194,n5195);
xor (n5194,n5191,n5192);
or (n5195,n5196,n5199);
and (n5196,n5197,n5198);
xor (n5197,n5016,n5017);
and (n5198,n1064,n414);
and (n5199,n5200,n5201);
xor (n5200,n5197,n5198);
or (n5201,n5202,n5205);
and (n5202,n5203,n5204);
xor (n5203,n5021,n5022);
and (n5204,n1103,n414);
and (n5205,n5206,n5207);
xor (n5206,n5203,n5204);
and (n5207,n5208,n3929);
xor (n5208,n5026,n5027);
and (n5209,n67,n32);
and (n5210,n5211,n5212);
xor (n5211,n4490,n5209);
or (n5212,n5213,n5215);
and (n5213,n5214,n797);
xor (n5214,n5032,n5033);
and (n5215,n5216,n5217);
xor (n5216,n5214,n797);
or (n5217,n5218,n5221);
and (n5218,n5219,n5220);
xor (n5219,n5038,n5039);
and (n5220,n172,n32);
and (n5221,n5222,n5223);
xor (n5222,n5219,n5220);
or (n5223,n5224,n5227);
and (n5224,n5225,n5226);
xor (n5225,n5044,n5045);
and (n5226,n166,n32);
and (n5227,n5228,n5229);
xor (n5228,n5225,n5226);
or (n5229,n5230,n5233);
and (n5230,n5231,n5232);
xor (n5231,n5050,n5051);
and (n5232,n95,n32);
and (n5233,n5234,n5235);
xor (n5234,n5231,n5232);
or (n5235,n5236,n5239);
and (n5236,n5237,n5238);
xor (n5237,n5056,n5057);
and (n5238,n88,n32);
and (n5239,n5240,n5241);
xor (n5240,n5237,n5238);
or (n5241,n5242,n5245);
and (n5242,n5243,n5244);
xor (n5243,n5062,n5063);
and (n5244,n249,n32);
and (n5245,n5246,n5247);
xor (n5246,n5243,n5244);
or (n5247,n5248,n5251);
and (n5248,n5249,n5250);
xor (n5249,n5068,n5069);
and (n5250,n243,n32);
and (n5251,n5252,n5253);
xor (n5252,n5249,n5250);
or (n5253,n5254,n5257);
and (n5254,n5255,n5256);
xor (n5255,n5074,n5075);
and (n5256,n377,n32);
and (n5257,n5258,n5259);
xor (n5258,n5255,n5256);
or (n5259,n5260,n5263);
and (n5260,n5261,n5262);
xor (n5261,n5080,n5081);
and (n5262,n436,n32);
and (n5263,n5264,n5265);
xor (n5264,n5261,n5262);
or (n5265,n5266,n5269);
and (n5266,n5267,n5268);
xor (n5267,n5086,n5087);
and (n5268,n281,n32);
and (n5269,n5270,n5271);
xor (n5270,n5267,n5268);
or (n5271,n5272,n5275);
and (n5272,n5273,n5274);
xor (n5273,n5092,n5093);
and (n5274,n274,n32);
and (n5275,n5276,n5277);
xor (n5276,n5273,n5274);
or (n5277,n5278,n5280);
and (n5278,n5279,n3366);
xor (n5279,n5098,n5099);
and (n5280,n5281,n5282);
xor (n5281,n5279,n3366);
or (n5282,n5283,n5285);
and (n5283,n5284,n2796);
xor (n5284,n5104,n5105);
and (n5285,n5286,n5287);
xor (n5286,n5284,n2796);
or (n5287,n5288,n5291);
and (n5288,n5289,n5290);
xor (n5289,n5110,n5111);
and (n5290,n223,n32);
and (n5291,n5292,n5293);
xor (n5292,n5289,n5290);
or (n5293,n5294,n5297);
and (n5294,n5295,n5296);
xor (n5295,n5116,n5117);
and (n5296,n217,n32);
and (n5297,n5298,n5299);
xor (n5298,n5295,n5296);
or (n5299,n5300,n5303);
and (n5300,n5301,n5302);
xor (n5301,n5122,n5123);
and (n5302,n124,n32);
and (n5303,n5304,n5305);
xor (n5304,n5301,n5302);
or (n5305,n5306,n5309);
and (n5306,n5307,n5308);
xor (n5307,n5128,n5129);
and (n5308,n118,n32);
and (n5309,n5310,n5311);
xor (n5310,n5307,n5308);
or (n5311,n5312,n5315);
and (n5312,n5313,n5314);
xor (n5313,n5134,n5135);
and (n5314,n150,n32);
and (n5315,n5316,n5317);
xor (n5316,n5313,n5314);
or (n5317,n5318,n5321);
and (n5318,n5319,n5320);
xor (n5319,n5140,n5141);
and (n5320,n144,n32);
and (n5321,n5322,n5323);
xor (n5322,n5319,n5320);
or (n5323,n5324,n5327);
and (n5324,n5325,n5326);
xor (n5325,n5146,n5147);
and (n5326,n398,n32);
and (n5327,n5328,n5329);
xor (n5328,n5325,n5326);
or (n5329,n5330,n5333);
and (n5330,n5331,n5332);
xor (n5331,n5152,n5153);
and (n5332,n449,n32);
and (n5333,n5334,n5335);
xor (n5334,n5331,n5332);
or (n5335,n5336,n5339);
and (n5336,n5337,n5338);
xor (n5337,n5158,n5159);
and (n5338,n443,n32);
and (n5339,n5340,n5341);
xor (n5340,n5337,n5338);
or (n5341,n5342,n5345);
and (n5342,n5343,n5344);
xor (n5343,n5164,n5165);
and (n5344,n551,n32);
and (n5345,n5346,n5347);
xor (n5346,n5343,n5344);
or (n5347,n5348,n5351);
and (n5348,n5349,n5350);
xor (n5349,n5170,n5171);
and (n5350,n308,n32);
and (n5351,n5352,n5353);
xor (n5352,n5349,n5350);
or (n5353,n5354,n5357);
and (n5354,n5355,n5356);
xor (n5355,n5176,n5177);
and (n5356,n302,n32);
and (n5357,n5358,n5359);
xor (n5358,n5355,n5356);
or (n5359,n5360,n5363);
and (n5360,n5361,n5362);
xor (n5361,n5182,n5183);
and (n5362,n670,n32);
and (n5363,n5364,n5365);
xor (n5364,n5361,n5362);
or (n5365,n5366,n5369);
and (n5366,n5367,n5368);
xor (n5367,n5188,n5189);
and (n5368,n889,n32);
and (n5369,n5370,n5371);
xor (n5370,n5367,n5368);
or (n5371,n5372,n5374);
and (n5372,n5373,n3867);
xor (n5373,n5194,n5195);
and (n5374,n5375,n5376);
xor (n5375,n5373,n3867);
or (n5376,n5377,n5379);
and (n5377,n5378,n3922);
xor (n5378,n5200,n5201);
and (n5379,n5380,n5381);
xor (n5380,n5378,n3922);
and (n5381,n5382,n5383);
xor (n5382,n5206,n5207);
and (n5383,n1266,n32);
and (n5384,n67,n30);
and (n5385,n5386,n5387);
xor (n5386,n4487,n5384);
or (n5387,n5388,n5391);
and (n5388,n5389,n5390);
xor (n5389,n5211,n5212);
and (n5390,n61,n30);
and (n5391,n5392,n5393);
xor (n5392,n5389,n5390);
or (n5393,n5394,n5397);
and (n5394,n5395,n5396);
xor (n5395,n5216,n5217);
and (n5396,n172,n30);
and (n5397,n5398,n5399);
xor (n5398,n5395,n5396);
or (n5399,n5400,n5403);
and (n5400,n5401,n5402);
xor (n5401,n5222,n5223);
and (n5402,n166,n30);
and (n5403,n5404,n5405);
xor (n5404,n5401,n5402);
or (n5405,n5406,n5409);
and (n5406,n5407,n5408);
xor (n5407,n5228,n5229);
and (n5408,n95,n30);
and (n5409,n5410,n5411);
xor (n5410,n5407,n5408);
or (n5411,n5412,n5415);
and (n5412,n5413,n5414);
xor (n5413,n5234,n5235);
and (n5414,n88,n30);
and (n5415,n5416,n5417);
xor (n5416,n5413,n5414);
or (n5417,n5418,n5421);
and (n5418,n5419,n5420);
xor (n5419,n5240,n5241);
and (n5420,n249,n30);
and (n5421,n5422,n5423);
xor (n5422,n5419,n5420);
or (n5423,n5424,n5427);
and (n5424,n5425,n5426);
xor (n5425,n5246,n5247);
and (n5426,n243,n30);
and (n5427,n5428,n5429);
xor (n5428,n5425,n5426);
or (n5429,n5430,n5433);
and (n5430,n5431,n5432);
xor (n5431,n5252,n5253);
and (n5432,n377,n30);
and (n5433,n5434,n5435);
xor (n5434,n5431,n5432);
or (n5435,n5436,n5439);
and (n5436,n5437,n5438);
xor (n5437,n5258,n5259);
and (n5438,n436,n30);
and (n5439,n5440,n5441);
xor (n5440,n5437,n5438);
or (n5441,n5442,n5445);
and (n5442,n5443,n5444);
xor (n5443,n5264,n5265);
and (n5444,n281,n30);
and (n5445,n5446,n5447);
xor (n5446,n5443,n5444);
or (n5447,n5448,n5451);
and (n5448,n5449,n5450);
xor (n5449,n5270,n5271);
and (n5450,n274,n30);
and (n5451,n5452,n5453);
xor (n5452,n5449,n5450);
or (n5453,n5454,n5457);
and (n5454,n5455,n5456);
xor (n5455,n5276,n5277);
and (n5456,n201,n30);
and (n5457,n5458,n5459);
xor (n5458,n5455,n5456);
or (n5459,n5460,n5463);
and (n5460,n5461,n5462);
xor (n5461,n5281,n5282);
and (n5462,n195,n30);
and (n5463,n5464,n5465);
xor (n5464,n5461,n5462);
or (n5465,n5466,n5469);
and (n5466,n5467,n5468);
xor (n5467,n5286,n5287);
and (n5468,n223,n30);
and (n5469,n5470,n5471);
xor (n5470,n5467,n5468);
or (n5471,n5472,n5475);
and (n5472,n5473,n5474);
xor (n5473,n5292,n5293);
and (n5474,n217,n30);
and (n5475,n5476,n5477);
xor (n5476,n5473,n5474);
or (n5477,n5478,n5481);
and (n5478,n5479,n5480);
xor (n5479,n5298,n5299);
and (n5480,n124,n30);
and (n5481,n5482,n5483);
xor (n5482,n5479,n5480);
or (n5483,n5484,n5487);
and (n5484,n5485,n5486);
xor (n5485,n5304,n5305);
and (n5486,n118,n30);
and (n5487,n5488,n5489);
xor (n5488,n5485,n5486);
or (n5489,n5490,n5493);
and (n5490,n5491,n5492);
xor (n5491,n5310,n5311);
and (n5492,n150,n30);
and (n5493,n5494,n5495);
xor (n5494,n5491,n5492);
or (n5495,n5496,n5499);
and (n5496,n5497,n5498);
xor (n5497,n5316,n5317);
and (n5498,n144,n30);
and (n5499,n5500,n5501);
xor (n5500,n5497,n5498);
or (n5501,n5502,n5505);
and (n5502,n5503,n5504);
xor (n5503,n5322,n5323);
and (n5504,n398,n30);
and (n5505,n5506,n5507);
xor (n5506,n5503,n5504);
or (n5507,n5508,n5511);
and (n5508,n5509,n5510);
xor (n5509,n5328,n5329);
and (n5510,n449,n30);
and (n5511,n5512,n5513);
xor (n5512,n5509,n5510);
or (n5513,n5514,n5517);
and (n5514,n5515,n5516);
xor (n5515,n5334,n5335);
and (n5516,n443,n30);
and (n5517,n5518,n5519);
xor (n5518,n5515,n5516);
or (n5519,n5520,n5523);
and (n5520,n5521,n5522);
xor (n5521,n5340,n5341);
and (n5522,n551,n30);
and (n5523,n5524,n5525);
xor (n5524,n5521,n5522);
or (n5525,n5526,n5529);
and (n5526,n5527,n5528);
xor (n5527,n5346,n5347);
and (n5528,n308,n30);
and (n5529,n5530,n5531);
xor (n5530,n5527,n5528);
or (n5531,n5532,n5535);
and (n5532,n5533,n5534);
xor (n5533,n5352,n5353);
and (n5534,n302,n30);
and (n5535,n5536,n5537);
xor (n5536,n5533,n5534);
or (n5537,n5538,n5541);
and (n5538,n5539,n5540);
xor (n5539,n5358,n5359);
and (n5540,n670,n30);
and (n5541,n5542,n5543);
xor (n5542,n5539,n5540);
or (n5543,n5544,n5547);
and (n5544,n5545,n5546);
xor (n5545,n5364,n5365);
and (n5546,n889,n30);
and (n5547,n5548,n5549);
xor (n5548,n5545,n5546);
or (n5549,n5550,n5553);
and (n5550,n5551,n5552);
xor (n5551,n5370,n5371);
and (n5552,n1064,n30);
and (n5553,n5554,n5555);
xor (n5554,n5551,n5552);
or (n5555,n5556,n5559);
and (n5556,n5557,n5558);
xor (n5557,n5375,n5376);
and (n5558,n1103,n30);
and (n5559,n5560,n5561);
xor (n5560,n5557,n5558);
and (n5561,n5562,n3826);
xor (n5562,n5380,n5381);
and (n5563,n67,n37);
and (n5564,n5565,n5566);
xor (n5565,n4484,n5563);
or (n5566,n5567,n5570);
and (n5567,n5568,n5569);
xor (n5568,n5386,n5387);
and (n5569,n61,n37);
and (n5570,n5571,n5572);
xor (n5571,n5568,n5569);
or (n5572,n5573,n5576);
and (n5573,n5574,n5575);
xor (n5574,n5392,n5393);
and (n5575,n172,n37);
and (n5576,n5577,n5578);
xor (n5577,n5574,n5575);
or (n5578,n5579,n5582);
and (n5579,n5580,n5581);
xor (n5580,n5398,n5399);
and (n5581,n166,n37);
and (n5582,n5583,n5584);
xor (n5583,n5580,n5581);
or (n5584,n5585,n5588);
and (n5585,n5586,n5587);
xor (n5586,n5404,n5405);
and (n5587,n95,n37);
and (n5588,n5589,n5590);
xor (n5589,n5586,n5587);
or (n5590,n5591,n5594);
and (n5591,n5592,n5593);
xor (n5592,n5410,n5411);
and (n5593,n88,n37);
and (n5594,n5595,n5596);
xor (n5595,n5592,n5593);
or (n5596,n5597,n5600);
and (n5597,n5598,n5599);
xor (n5598,n5416,n5417);
and (n5599,n249,n37);
and (n5600,n5601,n5602);
xor (n5601,n5598,n5599);
or (n5602,n5603,n5606);
and (n5603,n5604,n5605);
xor (n5604,n5422,n5423);
and (n5605,n243,n37);
and (n5606,n5607,n5608);
xor (n5607,n5604,n5605);
or (n5608,n5609,n5612);
and (n5609,n5610,n5611);
xor (n5610,n5428,n5429);
and (n5611,n377,n37);
and (n5612,n5613,n5614);
xor (n5613,n5610,n5611);
or (n5614,n5615,n5618);
and (n5615,n5616,n5617);
xor (n5616,n5434,n5435);
and (n5617,n436,n37);
and (n5618,n5619,n5620);
xor (n5619,n5616,n5617);
or (n5620,n5621,n5624);
and (n5621,n5622,n5623);
xor (n5622,n5440,n5441);
and (n5623,n281,n37);
and (n5624,n5625,n5626);
xor (n5625,n5622,n5623);
or (n5626,n5627,n5630);
and (n5627,n5628,n5629);
xor (n5628,n5446,n5447);
and (n5629,n274,n37);
and (n5630,n5631,n5632);
xor (n5631,n5628,n5629);
or (n5632,n5633,n5636);
and (n5633,n5634,n5635);
xor (n5634,n5452,n5453);
and (n5635,n201,n37);
and (n5636,n5637,n5638);
xor (n5637,n5634,n5635);
or (n5638,n5639,n5642);
and (n5639,n5640,n5641);
xor (n5640,n5458,n5459);
and (n5641,n195,n37);
and (n5642,n5643,n5644);
xor (n5643,n5640,n5641);
or (n5644,n5645,n5648);
and (n5645,n5646,n5647);
xor (n5646,n5464,n5465);
and (n5647,n223,n37);
and (n5648,n5649,n5650);
xor (n5649,n5646,n5647);
or (n5650,n5651,n5653);
and (n5651,n5652,n2681);
xor (n5652,n5470,n5471);
and (n5653,n5654,n5655);
xor (n5654,n5652,n2681);
or (n5655,n5656,n5658);
and (n5656,n5657,n2617);
xor (n5657,n5476,n5477);
and (n5658,n5659,n5660);
xor (n5659,n5657,n2617);
or (n5660,n5661,n5663);
and (n5661,n5662,n2582);
xor (n5662,n5482,n5483);
and (n5663,n5664,n5665);
xor (n5664,n5662,n2582);
or (n5665,n5666,n5668);
and (n5666,n5667,n2486);
xor (n5667,n5488,n5489);
and (n5668,n5669,n5670);
xor (n5669,n5667,n2486);
or (n5670,n5671,n5674);
and (n5671,n5672,n5673);
xor (n5672,n5494,n5495);
and (n5673,n144,n37);
and (n5674,n5675,n5676);
xor (n5675,n5672,n5673);
or (n5676,n5677,n5680);
and (n5677,n5678,n5679);
xor (n5678,n5500,n5501);
and (n5679,n398,n37);
and (n5680,n5681,n5682);
xor (n5681,n5678,n5679);
or (n5682,n5683,n5686);
and (n5683,n5684,n5685);
xor (n5684,n5506,n5507);
and (n5685,n449,n37);
and (n5686,n5687,n5688);
xor (n5687,n5684,n5685);
or (n5688,n5689,n5692);
and (n5689,n5690,n5691);
xor (n5690,n5512,n5513);
and (n5691,n443,n37);
and (n5692,n5693,n5694);
xor (n5693,n5690,n5691);
or (n5694,n5695,n5697);
and (n5695,n5696,n3122);
xor (n5696,n5518,n5519);
and (n5697,n5698,n5699);
xor (n5698,n5696,n3122);
or (n5699,n5700,n5703);
and (n5700,n5701,n5702);
xor (n5701,n5524,n5525);
and (n5702,n308,n37);
and (n5703,n5704,n5705);
xor (n5704,n5701,n5702);
or (n5705,n5706,n5709);
and (n5706,n5707,n5708);
xor (n5707,n5530,n5531);
and (n5708,n302,n37);
and (n5709,n5710,n5711);
xor (n5710,n5707,n5708);
or (n5711,n5712,n5715);
and (n5712,n5713,n5714);
xor (n5713,n5536,n5537);
and (n5714,n670,n37);
and (n5715,n5716,n5717);
xor (n5716,n5713,n5714);
or (n5717,n5718,n5721);
and (n5718,n5719,n5720);
xor (n5719,n5542,n5543);
and (n5720,n889,n37);
and (n5721,n5722,n5723);
xor (n5722,n5719,n5720);
or (n5723,n5724,n5727);
and (n5724,n5725,n5726);
xor (n5725,n5548,n5549);
and (n5726,n1064,n37);
and (n5727,n5728,n5729);
xor (n5728,n5725,n5726);
or (n5729,n5730,n5732);
and (n5730,n5731,n3696);
xor (n5731,n5554,n5555);
and (n5732,n5733,n5734);
xor (n5733,n5731,n3696);
and (n5734,n5735,n5736);
xor (n5735,n5560,n5561);
and (n5736,n1266,n37);
and (n5737,n67,n52);
or (n5738,n5739,n5742);
and (n5739,n5740,n5741);
xor (n5740,n5565,n5566);
and (n5741,n61,n52);
and (n5742,n5743,n5744);
xor (n5743,n5740,n5741);
or (n5744,n5745,n5748);
and (n5745,n5746,n5747);
xor (n5746,n5571,n5572);
and (n5747,n172,n52);
and (n5748,n5749,n5750);
xor (n5749,n5746,n5747);
or (n5750,n5751,n5754);
and (n5751,n5752,n5753);
xor (n5752,n5577,n5578);
and (n5753,n166,n52);
and (n5754,n5755,n5756);
xor (n5755,n5752,n5753);
or (n5756,n5757,n5760);
and (n5757,n5758,n5759);
xor (n5758,n5583,n5584);
and (n5759,n95,n52);
and (n5760,n5761,n5762);
xor (n5761,n5758,n5759);
or (n5762,n5763,n5766);
and (n5763,n5764,n5765);
xor (n5764,n5589,n5590);
and (n5765,n88,n52);
and (n5766,n5767,n5768);
xor (n5767,n5764,n5765);
or (n5768,n5769,n5772);
and (n5769,n5770,n5771);
xor (n5770,n5595,n5596);
and (n5771,n249,n52);
and (n5772,n5773,n5774);
xor (n5773,n5770,n5771);
or (n5774,n5775,n5778);
and (n5775,n5776,n5777);
xor (n5776,n5601,n5602);
and (n5777,n243,n52);
and (n5778,n5779,n5780);
xor (n5779,n5776,n5777);
or (n5780,n5781,n5784);
and (n5781,n5782,n5783);
xor (n5782,n5607,n5608);
and (n5783,n377,n52);
and (n5784,n5785,n5786);
xor (n5785,n5782,n5783);
or (n5786,n5787,n5790);
and (n5787,n5788,n5789);
xor (n5788,n5613,n5614);
and (n5789,n436,n52);
and (n5790,n5791,n5792);
xor (n5791,n5788,n5789);
or (n5792,n5793,n5796);
and (n5793,n5794,n5795);
xor (n5794,n5619,n5620);
and (n5795,n281,n52);
and (n5796,n5797,n5798);
xor (n5797,n5794,n5795);
or (n5798,n5799,n5802);
and (n5799,n5800,n5801);
xor (n5800,n5625,n5626);
and (n5801,n274,n52);
and (n5802,n5803,n5804);
xor (n5803,n5800,n5801);
or (n5804,n5805,n5808);
and (n5805,n5806,n5807);
xor (n5806,n5631,n5632);
and (n5807,n201,n52);
and (n5808,n5809,n5810);
xor (n5809,n5806,n5807);
or (n5810,n5811,n5814);
and (n5811,n5812,n5813);
xor (n5812,n5637,n5638);
and (n5813,n195,n52);
and (n5814,n5815,n5816);
xor (n5815,n5812,n5813);
or (n5816,n5817,n5820);
and (n5817,n5818,n5819);
xor (n5818,n5643,n5644);
and (n5819,n223,n52);
and (n5820,n5821,n5822);
xor (n5821,n5818,n5819);
or (n5822,n5823,n5826);
and (n5823,n5824,n5825);
xor (n5824,n5649,n5650);
and (n5825,n217,n52);
and (n5826,n5827,n5828);
xor (n5827,n5824,n5825);
or (n5828,n5829,n5832);
and (n5829,n5830,n5831);
xor (n5830,n5654,n5655);
and (n5831,n124,n52);
and (n5832,n5833,n5834);
xor (n5833,n5830,n5831);
or (n5834,n5835,n5838);
and (n5835,n5836,n5837);
xor (n5836,n5659,n5660);
and (n5837,n118,n52);
and (n5838,n5839,n5840);
xor (n5839,n5836,n5837);
or (n5840,n5841,n5844);
and (n5841,n5842,n5843);
xor (n5842,n5664,n5665);
and (n5843,n150,n52);
and (n5844,n5845,n5846);
xor (n5845,n5842,n5843);
or (n5846,n5847,n5850);
and (n5847,n5848,n5849);
xor (n5848,n5669,n5670);
and (n5849,n144,n52);
and (n5850,n5851,n5852);
xor (n5851,n5848,n5849);
or (n5852,n5853,n5856);
and (n5853,n5854,n5855);
xor (n5854,n5675,n5676);
and (n5855,n398,n52);
and (n5856,n5857,n5858);
xor (n5857,n5854,n5855);
or (n5858,n5859,n5862);
and (n5859,n5860,n5861);
xor (n5860,n5681,n5682);
and (n5861,n449,n52);
and (n5862,n5863,n5864);
xor (n5863,n5860,n5861);
or (n5864,n5865,n5868);
and (n5865,n5866,n5867);
xor (n5866,n5687,n5688);
and (n5867,n443,n52);
and (n5868,n5869,n5870);
xor (n5869,n5866,n5867);
or (n5870,n5871,n5874);
and (n5871,n5872,n5873);
xor (n5872,n5693,n5694);
and (n5873,n551,n52);
and (n5874,n5875,n5876);
xor (n5875,n5872,n5873);
or (n5876,n5877,n5880);
and (n5877,n5878,n5879);
xor (n5878,n5698,n5699);
and (n5879,n308,n52);
and (n5880,n5881,n5882);
xor (n5881,n5878,n5879);
or (n5882,n5883,n5886);
and (n5883,n5884,n5885);
xor (n5884,n5704,n5705);
and (n5885,n302,n52);
and (n5886,n5887,n5888);
xor (n5887,n5884,n5885);
or (n5888,n5889,n5892);
and (n5889,n5890,n5891);
xor (n5890,n5710,n5711);
and (n5891,n670,n52);
and (n5892,n5893,n5894);
xor (n5893,n5890,n5891);
or (n5894,n5895,n5898);
and (n5895,n5896,n5897);
xor (n5896,n5716,n5717);
and (n5897,n889,n52);
and (n5898,n5899,n5900);
xor (n5899,n5896,n5897);
or (n5900,n5901,n5904);
and (n5901,n5902,n5903);
xor (n5902,n5722,n5723);
and (n5903,n1064,n52);
and (n5904,n5905,n5906);
xor (n5905,n5902,n5903);
or (n5906,n5907,n5910);
and (n5907,n5908,n5909);
xor (n5908,n5728,n5729);
and (n5909,n1103,n52);
and (n5910,n5911,n5912);
xor (n5911,n5908,n5909);
and (n5912,n5913,n3669);
xor (n5913,n5733,n5734);
and (n5914,n61,n56);
or (n5915,n5916,n5919);
and (n5916,n5917,n5918);
xor (n5917,n5743,n5744);
and (n5918,n172,n56);
and (n5919,n5920,n5921);
xor (n5920,n5917,n5918);
or (n5921,n5922,n5925);
and (n5922,n5923,n5924);
xor (n5923,n5749,n5750);
and (n5924,n166,n56);
and (n5925,n5926,n5927);
xor (n5926,n5923,n5924);
or (n5927,n5928,n5931);
and (n5928,n5929,n5930);
xor (n5929,n5755,n5756);
and (n5930,n95,n56);
and (n5931,n5932,n5933);
xor (n5932,n5929,n5930);
or (n5933,n5934,n5937);
and (n5934,n5935,n5936);
xor (n5935,n5761,n5762);
and (n5936,n88,n56);
and (n5937,n5938,n5939);
xor (n5938,n5935,n5936);
or (n5939,n5940,n5943);
and (n5940,n5941,n5942);
xor (n5941,n5767,n5768);
and (n5942,n249,n56);
and (n5943,n5944,n5945);
xor (n5944,n5941,n5942);
or (n5945,n5946,n5949);
and (n5946,n5947,n5948);
xor (n5947,n5773,n5774);
and (n5948,n243,n56);
and (n5949,n5950,n5951);
xor (n5950,n5947,n5948);
or (n5951,n5952,n5955);
and (n5952,n5953,n5954);
xor (n5953,n5779,n5780);
and (n5954,n377,n56);
and (n5955,n5956,n5957);
xor (n5956,n5953,n5954);
or (n5957,n5958,n5960);
and (n5958,n5959,n1453);
xor (n5959,n5785,n5786);
and (n5960,n5961,n5962);
xor (n5961,n5959,n1453);
or (n5962,n5963,n5966);
and (n5963,n5964,n5965);
xor (n5964,n5791,n5792);
and (n5965,n281,n56);
and (n5966,n5967,n5968);
xor (n5967,n5964,n5965);
or (n5968,n5969,n5972);
and (n5969,n5970,n5971);
xor (n5970,n5797,n5798);
and (n5971,n274,n56);
and (n5972,n5973,n5974);
xor (n5973,n5970,n5971);
or (n5974,n5975,n5978);
and (n5975,n5976,n5977);
xor (n5976,n5803,n5804);
and (n5977,n201,n56);
and (n5978,n5979,n5980);
xor (n5979,n5976,n5977);
or (n5980,n5981,n5984);
and (n5981,n5982,n5983);
xor (n5982,n5809,n5810);
and (n5983,n195,n56);
and (n5984,n5985,n5986);
xor (n5985,n5982,n5983);
or (n5986,n5987,n5990);
and (n5987,n5988,n5989);
xor (n5988,n5815,n5816);
and (n5989,n223,n56);
and (n5990,n5991,n5992);
xor (n5991,n5988,n5989);
or (n5992,n5993,n5996);
and (n5993,n5994,n5995);
xor (n5994,n5821,n5822);
and (n5995,n217,n56);
and (n5996,n5997,n5998);
xor (n5997,n5994,n5995);
or (n5998,n5999,n6002);
and (n5999,n6000,n6001);
xor (n6000,n5827,n5828);
and (n6001,n124,n56);
and (n6002,n6003,n6004);
xor (n6003,n6000,n6001);
or (n6004,n6005,n6008);
and (n6005,n6006,n6007);
xor (n6006,n5833,n5834);
and (n6007,n118,n56);
and (n6008,n6009,n6010);
xor (n6009,n6006,n6007);
or (n6010,n6011,n6014);
and (n6011,n6012,n6013);
xor (n6012,n5839,n5840);
and (n6013,n150,n56);
and (n6014,n6015,n6016);
xor (n6015,n6012,n6013);
or (n6016,n6017,n6020);
and (n6017,n6018,n6019);
xor (n6018,n5845,n5846);
and (n6019,n144,n56);
and (n6020,n6021,n6022);
xor (n6021,n6018,n6019);
or (n6022,n6023,n6025);
and (n6023,n6024,n2536);
xor (n6024,n5851,n5852);
and (n6025,n6026,n6027);
xor (n6026,n6024,n2536);
or (n6027,n6028,n6031);
and (n6028,n6029,n6030);
xor (n6029,n5857,n5858);
and (n6030,n449,n56);
and (n6031,n6032,n6033);
xor (n6032,n6029,n6030);
or (n6033,n6034,n6037);
and (n6034,n6035,n6036);
xor (n6035,n5863,n5864);
and (n6036,n443,n56);
and (n6037,n6038,n6039);
xor (n6038,n6035,n6036);
or (n6039,n6040,n6043);
and (n6040,n6041,n6042);
xor (n6041,n5869,n5870);
and (n6042,n551,n56);
and (n6043,n6044,n6045);
xor (n6044,n6041,n6042);
or (n6045,n6046,n6049);
and (n6046,n6047,n6048);
xor (n6047,n5875,n5876);
and (n6048,n308,n56);
and (n6049,n6050,n6051);
xor (n6050,n6047,n6048);
or (n6051,n6052,n6055);
and (n6052,n6053,n6054);
xor (n6053,n5881,n5882);
and (n6054,n302,n56);
and (n6055,n6056,n6057);
xor (n6056,n6053,n6054);
or (n6057,n6058,n6061);
and (n6058,n6059,n6060);
xor (n6059,n5887,n5888);
and (n6060,n670,n56);
and (n6061,n6062,n6063);
xor (n6062,n6059,n6060);
or (n6063,n6064,n6067);
and (n6064,n6065,n6066);
xor (n6065,n5893,n5894);
and (n6066,n889,n56);
and (n6067,n6068,n6069);
xor (n6068,n6065,n6066);
or (n6069,n6070,n6073);
and (n6070,n6071,n6072);
xor (n6071,n5899,n5900);
and (n6072,n1064,n56);
and (n6073,n6074,n6075);
xor (n6074,n6071,n6072);
or (n6075,n6076,n6079);
and (n6076,n6077,n6078);
xor (n6077,n5905,n5906);
and (n6078,n1103,n56);
and (n6079,n6080,n6081);
xor (n6080,n6077,n6078);
and (n6081,n6082,n6083);
xor (n6082,n5911,n5912);
and (n6083,n1266,n56);
and (n6084,n172,n159);
or (n6085,n6086,n6089);
and (n6086,n6087,n6088);
xor (n6087,n5920,n5921);
and (n6088,n166,n159);
and (n6089,n6090,n6091);
xor (n6090,n6087,n6088);
or (n6091,n6092,n6095);
and (n6092,n6093,n6094);
xor (n6093,n5926,n5927);
and (n6094,n95,n159);
and (n6095,n6096,n6097);
xor (n6096,n6093,n6094);
or (n6097,n6098,n6101);
and (n6098,n6099,n6100);
xor (n6099,n5932,n5933);
and (n6100,n88,n159);
and (n6101,n6102,n6103);
xor (n6102,n6099,n6100);
or (n6103,n6104,n6107);
and (n6104,n6105,n6106);
xor (n6105,n5938,n5939);
and (n6106,n249,n159);
and (n6107,n6108,n6109);
xor (n6108,n6105,n6106);
or (n6109,n6110,n6113);
and (n6110,n6111,n6112);
xor (n6111,n5944,n5945);
and (n6112,n243,n159);
and (n6113,n6114,n6115);
xor (n6114,n6111,n6112);
or (n6115,n6116,n6119);
and (n6116,n6117,n6118);
xor (n6117,n5950,n5951);
and (n6118,n377,n159);
and (n6119,n6120,n6121);
xor (n6120,n6117,n6118);
or (n6121,n6122,n6125);
and (n6122,n6123,n6124);
xor (n6123,n5956,n5957);
and (n6124,n436,n159);
and (n6125,n6126,n6127);
xor (n6126,n6123,n6124);
or (n6127,n6128,n6131);
and (n6128,n6129,n6130);
xor (n6129,n5961,n5962);
and (n6130,n281,n159);
and (n6131,n6132,n6133);
xor (n6132,n6129,n6130);
or (n6133,n6134,n6137);
and (n6134,n6135,n6136);
xor (n6135,n5967,n5968);
and (n6136,n274,n159);
and (n6137,n6138,n6139);
xor (n6138,n6135,n6136);
or (n6139,n6140,n6143);
and (n6140,n6141,n6142);
xor (n6141,n5973,n5974);
and (n6142,n201,n159);
and (n6143,n6144,n6145);
xor (n6144,n6141,n6142);
or (n6145,n6146,n6149);
and (n6146,n6147,n6148);
xor (n6147,n5979,n5980);
and (n6148,n195,n159);
and (n6149,n6150,n6151);
xor (n6150,n6147,n6148);
or (n6151,n6152,n6155);
and (n6152,n6153,n6154);
xor (n6153,n5985,n5986);
and (n6154,n223,n159);
and (n6155,n6156,n6157);
xor (n6156,n6153,n6154);
or (n6157,n6158,n6161);
and (n6158,n6159,n6160);
xor (n6159,n5991,n5992);
and (n6160,n217,n159);
and (n6161,n6162,n6163);
xor (n6162,n6159,n6160);
or (n6163,n6164,n6167);
and (n6164,n6165,n6166);
xor (n6165,n5997,n5998);
and (n6166,n124,n159);
and (n6167,n6168,n6169);
xor (n6168,n6165,n6166);
or (n6169,n6170,n6173);
and (n6170,n6171,n6172);
xor (n6171,n6003,n6004);
and (n6172,n118,n159);
and (n6173,n6174,n6175);
xor (n6174,n6171,n6172);
or (n6175,n6176,n6179);
and (n6176,n6177,n6178);
xor (n6177,n6009,n6010);
and (n6178,n150,n159);
and (n6179,n6180,n6181);
xor (n6180,n6177,n6178);
or (n6181,n6182,n6185);
and (n6182,n6183,n6184);
xor (n6183,n6015,n6016);
and (n6184,n144,n159);
and (n6185,n6186,n6187);
xor (n6186,n6183,n6184);
or (n6187,n6188,n6191);
and (n6188,n6189,n6190);
xor (n6189,n6021,n6022);
and (n6190,n398,n159);
and (n6191,n6192,n6193);
xor (n6192,n6189,n6190);
or (n6193,n6194,n6197);
and (n6194,n6195,n6196);
xor (n6195,n6026,n6027);
and (n6196,n449,n159);
and (n6197,n6198,n6199);
xor (n6198,n6195,n6196);
or (n6199,n6200,n6203);
and (n6200,n6201,n6202);
xor (n6201,n6032,n6033);
and (n6202,n443,n159);
and (n6203,n6204,n6205);
xor (n6204,n6201,n6202);
or (n6205,n6206,n6209);
and (n6206,n6207,n6208);
xor (n6207,n6038,n6039);
and (n6208,n551,n159);
and (n6209,n6210,n6211);
xor (n6210,n6207,n6208);
or (n6211,n6212,n6215);
and (n6212,n6213,n6214);
xor (n6213,n6044,n6045);
and (n6214,n308,n159);
and (n6215,n6216,n6217);
xor (n6216,n6213,n6214);
or (n6217,n6218,n6221);
and (n6218,n6219,n6220);
xor (n6219,n6050,n6051);
and (n6220,n302,n159);
and (n6221,n6222,n6223);
xor (n6222,n6219,n6220);
or (n6223,n6224,n6227);
and (n6224,n6225,n6226);
xor (n6225,n6056,n6057);
and (n6226,n670,n159);
and (n6227,n6228,n6229);
xor (n6228,n6225,n6226);
or (n6229,n6230,n6233);
and (n6230,n6231,n6232);
xor (n6231,n6062,n6063);
and (n6232,n889,n159);
and (n6233,n6234,n6235);
xor (n6234,n6231,n6232);
or (n6235,n6236,n6239);
and (n6236,n6237,n6238);
xor (n6237,n6068,n6069);
and (n6238,n1064,n159);
and (n6239,n6240,n6241);
xor (n6240,n6237,n6238);
or (n6241,n6242,n6245);
and (n6242,n6243,n6244);
xor (n6243,n6074,n6075);
and (n6244,n1103,n159);
and (n6245,n6246,n6247);
xor (n6246,n6243,n6244);
and (n6247,n6248,n3769);
xor (n6248,n6080,n6081);
and (n6249,n166,n78);
or (n6250,n6251,n6254);
and (n6251,n6252,n6253);
xor (n6252,n6090,n6091);
and (n6253,n95,n78);
and (n6254,n6255,n6256);
xor (n6255,n6252,n6253);
or (n6256,n6257,n6260);
and (n6257,n6258,n6259);
xor (n6258,n6096,n6097);
and (n6259,n88,n78);
and (n6260,n6261,n6262);
xor (n6261,n6258,n6259);
or (n6262,n6263,n6266);
and (n6263,n6264,n6265);
xor (n6264,n6102,n6103);
and (n6265,n249,n78);
and (n6266,n6267,n6268);
xor (n6267,n6264,n6265);
or (n6268,n6269,n6272);
and (n6269,n6270,n6271);
xor (n6270,n6108,n6109);
and (n6271,n243,n78);
and (n6272,n6273,n6274);
xor (n6273,n6270,n6271);
or (n6274,n6275,n6278);
and (n6275,n6276,n6277);
xor (n6276,n6114,n6115);
and (n6277,n377,n78);
and (n6278,n6279,n6280);
xor (n6279,n6276,n6277);
or (n6280,n6281,n6284);
and (n6281,n6282,n6283);
xor (n6282,n6120,n6121);
and (n6283,n436,n78);
and (n6284,n6285,n6286);
xor (n6285,n6282,n6283);
or (n6286,n6287,n6290);
and (n6287,n6288,n6289);
xor (n6288,n6126,n6127);
and (n6289,n281,n78);
and (n6290,n6291,n6292);
xor (n6291,n6288,n6289);
or (n6292,n6293,n6296);
and (n6293,n6294,n6295);
xor (n6294,n6132,n6133);
and (n6295,n274,n78);
and (n6296,n6297,n6298);
xor (n6297,n6294,n6295);
or (n6298,n6299,n6302);
and (n6299,n6300,n6301);
xor (n6300,n6138,n6139);
and (n6301,n201,n78);
and (n6302,n6303,n6304);
xor (n6303,n6300,n6301);
or (n6304,n6305,n6307);
and (n6305,n6306,n1903);
xor (n6306,n6144,n6145);
and (n6307,n6308,n6309);
xor (n6308,n6306,n1903);
or (n6309,n6310,n6313);
and (n6310,n6311,n6312);
xor (n6311,n6150,n6151);
and (n6312,n223,n78);
and (n6313,n6314,n6315);
xor (n6314,n6311,n6312);
or (n6315,n6316,n6319);
and (n6316,n6317,n6318);
xor (n6317,n6156,n6157);
and (n6318,n217,n78);
and (n6319,n6320,n6321);
xor (n6320,n6317,n6318);
or (n6321,n6322,n6325);
and (n6322,n6323,n6324);
xor (n6323,n6162,n6163);
and (n6324,n124,n78);
and (n6325,n6326,n6327);
xor (n6326,n6323,n6324);
or (n6327,n6328,n6331);
and (n6328,n6329,n6330);
xor (n6329,n6168,n6169);
and (n6330,n118,n78);
and (n6331,n6332,n6333);
xor (n6332,n6329,n6330);
or (n6333,n6334,n6337);
and (n6334,n6335,n6336);
xor (n6335,n6174,n6175);
and (n6336,n150,n78);
and (n6337,n6338,n6339);
xor (n6338,n6335,n6336);
or (n6339,n6340,n6343);
and (n6340,n6341,n6342);
xor (n6341,n6180,n6181);
and (n6342,n144,n78);
and (n6343,n6344,n6345);
xor (n6344,n6341,n6342);
or (n6345,n6346,n6349);
and (n6346,n6347,n6348);
xor (n6347,n6186,n6187);
and (n6348,n398,n78);
and (n6349,n6350,n6351);
xor (n6350,n6347,n6348);
or (n6351,n6352,n6355);
and (n6352,n6353,n6354);
xor (n6353,n6192,n6193);
and (n6354,n449,n78);
and (n6355,n6356,n6357);
xor (n6356,n6353,n6354);
or (n6357,n6358,n6361);
and (n6358,n6359,n6360);
xor (n6359,n6198,n6199);
and (n6360,n443,n78);
and (n6361,n6362,n6363);
xor (n6362,n6359,n6360);
or (n6363,n6364,n6367);
and (n6364,n6365,n6366);
xor (n6365,n6204,n6205);
and (n6366,n551,n78);
and (n6367,n6368,n6369);
xor (n6368,n6365,n6366);
or (n6369,n6370,n6373);
and (n6370,n6371,n6372);
xor (n6371,n6210,n6211);
and (n6372,n308,n78);
and (n6373,n6374,n6375);
xor (n6374,n6371,n6372);
or (n6375,n6376,n6379);
and (n6376,n6377,n6378);
xor (n6377,n6216,n6217);
and (n6378,n302,n78);
and (n6379,n6380,n6381);
xor (n6380,n6377,n6378);
or (n6381,n6382,n6385);
and (n6382,n6383,n6384);
xor (n6383,n6222,n6223);
and (n6384,n670,n78);
and (n6385,n6386,n6387);
xor (n6386,n6383,n6384);
or (n6387,n6388,n6391);
and (n6388,n6389,n6390);
xor (n6389,n6228,n6229);
and (n6390,n889,n78);
and (n6391,n6392,n6393);
xor (n6392,n6389,n6390);
or (n6393,n6394,n6397);
and (n6394,n6395,n6396);
xor (n6395,n6234,n6235);
and (n6396,n1064,n78);
and (n6397,n6398,n6399);
xor (n6398,n6395,n6396);
or (n6399,n6400,n6403);
and (n6400,n6401,n6402);
xor (n6401,n6240,n6241);
and (n6402,n1103,n78);
and (n6403,n6404,n6405);
xor (n6404,n6401,n6402);
and (n6405,n6406,n6407);
xor (n6406,n6246,n6247);
and (n6407,n1266,n78);
and (n6408,n95,n76);
or (n6409,n6410,n6413);
and (n6410,n6411,n6412);
xor (n6411,n6255,n6256);
and (n6412,n88,n76);
and (n6413,n6414,n6415);
xor (n6414,n6411,n6412);
or (n6415,n6416,n6419);
and (n6416,n6417,n6418);
xor (n6417,n6261,n6262);
and (n6418,n249,n76);
and (n6419,n6420,n6421);
xor (n6420,n6417,n6418);
or (n6421,n6422,n6425);
and (n6422,n6423,n6424);
xor (n6423,n6267,n6268);
and (n6424,n243,n76);
and (n6425,n6426,n6427);
xor (n6426,n6423,n6424);
or (n6427,n6428,n6431);
and (n6428,n6429,n6430);
xor (n6429,n6273,n6274);
and (n6430,n377,n76);
and (n6431,n6432,n6433);
xor (n6432,n6429,n6430);
or (n6433,n6434,n6437);
and (n6434,n6435,n6436);
xor (n6435,n6279,n6280);
and (n6436,n436,n76);
and (n6437,n6438,n6439);
xor (n6438,n6435,n6436);
or (n6439,n6440,n6443);
and (n6440,n6441,n6442);
xor (n6441,n6285,n6286);
and (n6442,n281,n76);
and (n6443,n6444,n6445);
xor (n6444,n6441,n6442);
or (n6445,n6446,n6449);
and (n6446,n6447,n6448);
xor (n6447,n6291,n6292);
and (n6448,n274,n76);
and (n6449,n6450,n6451);
xor (n6450,n6447,n6448);
or (n6451,n6452,n6455);
and (n6452,n6453,n6454);
xor (n6453,n6297,n6298);
and (n6454,n201,n76);
and (n6455,n6456,n6457);
xor (n6456,n6453,n6454);
or (n6457,n6458,n6461);
and (n6458,n6459,n6460);
xor (n6459,n6303,n6304);
and (n6460,n195,n76);
and (n6461,n6462,n6463);
xor (n6462,n6459,n6460);
or (n6463,n6464,n6467);
and (n6464,n6465,n6466);
xor (n6465,n6308,n6309);
and (n6466,n223,n76);
and (n6467,n6468,n6469);
xor (n6468,n6465,n6466);
or (n6469,n6470,n6473);
and (n6470,n6471,n6472);
xor (n6471,n6314,n6315);
and (n6472,n217,n76);
and (n6473,n6474,n6475);
xor (n6474,n6471,n6472);
or (n6475,n6476,n6479);
and (n6476,n6477,n6478);
xor (n6477,n6320,n6321);
and (n6478,n124,n76);
and (n6479,n6480,n6481);
xor (n6480,n6477,n6478);
or (n6481,n6482,n6485);
and (n6482,n6483,n6484);
xor (n6483,n6326,n6327);
and (n6484,n118,n76);
and (n6485,n6486,n6487);
xor (n6486,n6483,n6484);
or (n6487,n6488,n6491);
and (n6488,n6489,n6490);
xor (n6489,n6332,n6333);
and (n6490,n150,n76);
and (n6491,n6492,n6493);
xor (n6492,n6489,n6490);
or (n6493,n6494,n6497);
and (n6494,n6495,n6496);
xor (n6495,n6338,n6339);
and (n6496,n144,n76);
and (n6497,n6498,n6499);
xor (n6498,n6495,n6496);
or (n6499,n6500,n6503);
and (n6500,n6501,n6502);
xor (n6501,n6344,n6345);
and (n6502,n398,n76);
and (n6503,n6504,n6505);
xor (n6504,n6501,n6502);
or (n6505,n6506,n6509);
and (n6506,n6507,n6508);
xor (n6507,n6350,n6351);
and (n6508,n449,n76);
and (n6509,n6510,n6511);
xor (n6510,n6507,n6508);
or (n6511,n6512,n6515);
and (n6512,n6513,n6514);
xor (n6513,n6356,n6357);
and (n6514,n443,n76);
and (n6515,n6516,n6517);
xor (n6516,n6513,n6514);
or (n6517,n6518,n6521);
and (n6518,n6519,n6520);
xor (n6519,n6362,n6363);
and (n6520,n551,n76);
and (n6521,n6522,n6523);
xor (n6522,n6519,n6520);
or (n6523,n6524,n6527);
and (n6524,n6525,n6526);
xor (n6525,n6368,n6369);
and (n6526,n308,n76);
and (n6527,n6528,n6529);
xor (n6528,n6525,n6526);
or (n6529,n6530,n6533);
and (n6530,n6531,n6532);
xor (n6531,n6374,n6375);
and (n6532,n302,n76);
and (n6533,n6534,n6535);
xor (n6534,n6531,n6532);
or (n6535,n6536,n6539);
and (n6536,n6537,n6538);
xor (n6537,n6380,n6381);
and (n6538,n670,n76);
and (n6539,n6540,n6541);
xor (n6540,n6537,n6538);
or (n6541,n6542,n6545);
and (n6542,n6543,n6544);
xor (n6543,n6386,n6387);
and (n6544,n889,n76);
and (n6545,n6546,n6547);
xor (n6546,n6543,n6544);
or (n6547,n6548,n6551);
and (n6548,n6549,n6550);
xor (n6549,n6392,n6393);
and (n6550,n1064,n76);
and (n6551,n6552,n6553);
xor (n6552,n6549,n6550);
or (n6553,n6554,n6557);
and (n6554,n6555,n6556);
xor (n6555,n6398,n6399);
and (n6556,n1103,n76);
and (n6557,n6558,n6559);
xor (n6558,n6555,n6556);
and (n6559,n6560,n3055);
xor (n6560,n6404,n6405);
and (n6561,n88,n83);
or (n6562,n6563,n6566);
and (n6563,n6564,n6565);
xor (n6564,n6414,n6415);
and (n6565,n249,n83);
and (n6566,n6567,n6568);
xor (n6567,n6564,n6565);
or (n6568,n6569,n6572);
and (n6569,n6570,n6571);
xor (n6570,n6420,n6421);
and (n6571,n243,n83);
and (n6572,n6573,n6574);
xor (n6573,n6570,n6571);
or (n6574,n6575,n6578);
and (n6575,n6576,n6577);
xor (n6576,n6426,n6427);
and (n6577,n377,n83);
and (n6578,n6579,n6580);
xor (n6579,n6576,n6577);
or (n6580,n6581,n6584);
and (n6581,n6582,n6583);
xor (n6582,n6432,n6433);
and (n6583,n436,n83);
and (n6584,n6585,n6586);
xor (n6585,n6582,n6583);
or (n6586,n6587,n6590);
and (n6587,n6588,n6589);
xor (n6588,n6438,n6439);
and (n6589,n281,n83);
and (n6590,n6591,n6592);
xor (n6591,n6588,n6589);
or (n6592,n6593,n6596);
and (n6593,n6594,n6595);
xor (n6594,n6444,n6445);
and (n6595,n274,n83);
and (n6596,n6597,n6598);
xor (n6597,n6594,n6595);
or (n6598,n6599,n6602);
and (n6599,n6600,n6601);
xor (n6600,n6450,n6451);
and (n6601,n201,n83);
and (n6602,n6603,n6604);
xor (n6603,n6600,n6601);
or (n6604,n6605,n6608);
and (n6605,n6606,n6607);
xor (n6606,n6456,n6457);
and (n6607,n195,n83);
and (n6608,n6609,n6610);
xor (n6609,n6606,n6607);
or (n6610,n6611,n6614);
and (n6611,n6612,n6613);
xor (n6612,n6462,n6463);
and (n6613,n223,n83);
and (n6614,n6615,n6616);
xor (n6615,n6612,n6613);
or (n6616,n6617,n6620);
and (n6617,n6618,n6619);
xor (n6618,n6468,n6469);
and (n6619,n217,n83);
and (n6620,n6621,n6622);
xor (n6621,n6618,n6619);
or (n6622,n6623,n6626);
and (n6623,n6624,n6625);
xor (n6624,n6474,n6475);
and (n6625,n124,n83);
and (n6626,n6627,n6628);
xor (n6627,n6624,n6625);
or (n6628,n6629,n6632);
and (n6629,n6630,n6631);
xor (n6630,n6480,n6481);
and (n6631,n118,n83);
and (n6632,n6633,n6634);
xor (n6633,n6630,n6631);
or (n6634,n6635,n6638);
and (n6635,n6636,n6637);
xor (n6636,n6486,n6487);
and (n6637,n150,n83);
and (n6638,n6639,n6640);
xor (n6639,n6636,n6637);
or (n6640,n6641,n6644);
and (n6641,n6642,n6643);
xor (n6642,n6492,n6493);
and (n6643,n144,n83);
and (n6644,n6645,n6646);
xor (n6645,n6642,n6643);
or (n6646,n6647,n6650);
and (n6647,n6648,n6649);
xor (n6648,n6498,n6499);
and (n6649,n398,n83);
and (n6650,n6651,n6652);
xor (n6651,n6648,n6649);
or (n6652,n6653,n6656);
and (n6653,n6654,n6655);
xor (n6654,n6504,n6505);
and (n6655,n449,n83);
and (n6656,n6657,n6658);
xor (n6657,n6654,n6655);
or (n6658,n6659,n6662);
and (n6659,n6660,n6661);
xor (n6660,n6510,n6511);
and (n6661,n443,n83);
and (n6662,n6663,n6664);
xor (n6663,n6660,n6661);
or (n6664,n6665,n6668);
and (n6665,n6666,n6667);
xor (n6666,n6516,n6517);
and (n6667,n551,n83);
and (n6668,n6669,n6670);
xor (n6669,n6666,n6667);
or (n6670,n6671,n6674);
and (n6671,n6672,n6673);
xor (n6672,n6522,n6523);
and (n6673,n308,n83);
and (n6674,n6675,n6676);
xor (n6675,n6672,n6673);
or (n6676,n6677,n6680);
and (n6677,n6678,n6679);
xor (n6678,n6528,n6529);
and (n6679,n302,n83);
and (n6680,n6681,n6682);
xor (n6681,n6678,n6679);
or (n6682,n6683,n6686);
and (n6683,n6684,n6685);
xor (n6684,n6534,n6535);
and (n6685,n670,n83);
and (n6686,n6687,n6688);
xor (n6687,n6684,n6685);
or (n6688,n6689,n6692);
and (n6689,n6690,n6691);
xor (n6690,n6540,n6541);
and (n6691,n889,n83);
and (n6692,n6693,n6694);
xor (n6693,n6690,n6691);
or (n6694,n6695,n6698);
and (n6695,n6696,n6697);
xor (n6696,n6546,n6547);
and (n6697,n1064,n83);
and (n6698,n6699,n6700);
xor (n6699,n6696,n6697);
or (n6700,n6701,n6704);
and (n6701,n6702,n6703);
xor (n6702,n6552,n6553);
and (n6703,n1103,n83);
and (n6704,n6705,n6706);
xor (n6705,n6702,n6703);
and (n6706,n6707,n6708);
xor (n6707,n6558,n6559);
and (n6708,n1266,n83);
and (n6709,n249,n232);
or (n6710,n6711,n6714);
and (n6711,n6712,n6713);
xor (n6712,n6567,n6568);
and (n6713,n243,n232);
and (n6714,n6715,n6716);
xor (n6715,n6712,n6713);
or (n6716,n6717,n6720);
and (n6717,n6718,n6719);
xor (n6718,n6573,n6574);
and (n6719,n377,n232);
and (n6720,n6721,n6722);
xor (n6721,n6718,n6719);
or (n6722,n6723,n6726);
and (n6723,n6724,n6725);
xor (n6724,n6579,n6580);
and (n6725,n436,n232);
and (n6726,n6727,n6728);
xor (n6727,n6724,n6725);
or (n6728,n6729,n6732);
and (n6729,n6730,n6731);
xor (n6730,n6585,n6586);
and (n6731,n281,n232);
and (n6732,n6733,n6734);
xor (n6733,n6730,n6731);
or (n6734,n6735,n6738);
and (n6735,n6736,n6737);
xor (n6736,n6591,n6592);
and (n6737,n274,n232);
and (n6738,n6739,n6740);
xor (n6739,n6736,n6737);
or (n6740,n6741,n6744);
and (n6741,n6742,n6743);
xor (n6742,n6597,n6598);
and (n6743,n201,n232);
and (n6744,n6745,n6746);
xor (n6745,n6742,n6743);
or (n6746,n6747,n6750);
and (n6747,n6748,n6749);
xor (n6748,n6603,n6604);
and (n6749,n195,n232);
and (n6750,n6751,n6752);
xor (n6751,n6748,n6749);
or (n6752,n6753,n6756);
and (n6753,n6754,n6755);
xor (n6754,n6609,n6610);
and (n6755,n223,n232);
and (n6756,n6757,n6758);
xor (n6757,n6754,n6755);
or (n6758,n6759,n6762);
and (n6759,n6760,n6761);
xor (n6760,n6615,n6616);
and (n6761,n217,n232);
and (n6762,n6763,n6764);
xor (n6763,n6760,n6761);
or (n6764,n6765,n6768);
and (n6765,n6766,n6767);
xor (n6766,n6621,n6622);
and (n6767,n124,n232);
and (n6768,n6769,n6770);
xor (n6769,n6766,n6767);
or (n6770,n6771,n6774);
and (n6771,n6772,n6773);
xor (n6772,n6627,n6628);
and (n6773,n118,n232);
and (n6774,n6775,n6776);
xor (n6775,n6772,n6773);
or (n6776,n6777,n6780);
and (n6777,n6778,n6779);
xor (n6778,n6633,n6634);
and (n6779,n150,n232);
and (n6780,n6781,n6782);
xor (n6781,n6778,n6779);
or (n6782,n6783,n6786);
and (n6783,n6784,n6785);
xor (n6784,n6639,n6640);
and (n6785,n144,n232);
and (n6786,n6787,n6788);
xor (n6787,n6784,n6785);
or (n6788,n6789,n6792);
and (n6789,n6790,n6791);
xor (n6790,n6645,n6646);
and (n6791,n398,n232);
and (n6792,n6793,n6794);
xor (n6793,n6790,n6791);
or (n6794,n6795,n6798);
and (n6795,n6796,n6797);
xor (n6796,n6651,n6652);
and (n6797,n449,n232);
and (n6798,n6799,n6800);
xor (n6799,n6796,n6797);
or (n6800,n6801,n6804);
and (n6801,n6802,n6803);
xor (n6802,n6657,n6658);
and (n6803,n443,n232);
and (n6804,n6805,n6806);
xor (n6805,n6802,n6803);
or (n6806,n6807,n6810);
and (n6807,n6808,n6809);
xor (n6808,n6663,n6664);
and (n6809,n551,n232);
and (n6810,n6811,n6812);
xor (n6811,n6808,n6809);
or (n6812,n6813,n6816);
and (n6813,n6814,n6815);
xor (n6814,n6669,n6670);
and (n6815,n308,n232);
and (n6816,n6817,n6818);
xor (n6817,n6814,n6815);
or (n6818,n6819,n6822);
and (n6819,n6820,n6821);
xor (n6820,n6675,n6676);
and (n6821,n302,n232);
and (n6822,n6823,n6824);
xor (n6823,n6820,n6821);
or (n6824,n6825,n6828);
and (n6825,n6826,n6827);
xor (n6826,n6681,n6682);
and (n6827,n670,n232);
and (n6828,n6829,n6830);
xor (n6829,n6826,n6827);
or (n6830,n6831,n6834);
and (n6831,n6832,n6833);
xor (n6832,n6687,n6688);
and (n6833,n889,n232);
and (n6834,n6835,n6836);
xor (n6835,n6832,n6833);
or (n6836,n6837,n6840);
and (n6837,n6838,n6839);
xor (n6838,n6693,n6694);
and (n6839,n1064,n232);
and (n6840,n6841,n6842);
xor (n6841,n6838,n6839);
or (n6842,n6843,n6846);
and (n6843,n6844,n6845);
xor (n6844,n6699,n6700);
and (n6845,n1103,n232);
and (n6846,n6847,n6848);
xor (n6847,n6844,n6845);
and (n6848,n6849,n3077);
xor (n6849,n6705,n6706);
and (n6850,n243,n238);
or (n6851,n6852,n6855);
and (n6852,n6853,n6854);
xor (n6853,n6715,n6716);
and (n6854,n377,n238);
and (n6855,n6856,n6857);
xor (n6856,n6853,n6854);
or (n6857,n6858,n6861);
and (n6858,n6859,n6860);
xor (n6859,n6721,n6722);
and (n6860,n436,n238);
and (n6861,n6862,n6863);
xor (n6862,n6859,n6860);
or (n6863,n6864,n6867);
and (n6864,n6865,n6866);
xor (n6865,n6727,n6728);
and (n6866,n281,n238);
and (n6867,n6868,n6869);
xor (n6868,n6865,n6866);
or (n6869,n6870,n6873);
and (n6870,n6871,n6872);
xor (n6871,n6733,n6734);
and (n6872,n274,n238);
and (n6873,n6874,n6875);
xor (n6874,n6871,n6872);
or (n6875,n6876,n6879);
and (n6876,n6877,n6878);
xor (n6877,n6739,n6740);
and (n6878,n201,n238);
and (n6879,n6880,n6881);
xor (n6880,n6877,n6878);
or (n6881,n6882,n6885);
and (n6882,n6883,n6884);
xor (n6883,n6745,n6746);
and (n6884,n195,n238);
and (n6885,n6886,n6887);
xor (n6886,n6883,n6884);
or (n6887,n6888,n6891);
and (n6888,n6889,n6890);
xor (n6889,n6751,n6752);
and (n6890,n223,n238);
and (n6891,n6892,n6893);
xor (n6892,n6889,n6890);
or (n6893,n6894,n6897);
and (n6894,n6895,n6896);
xor (n6895,n6757,n6758);
and (n6896,n217,n238);
and (n6897,n6898,n6899);
xor (n6898,n6895,n6896);
or (n6899,n6900,n6903);
and (n6900,n6901,n6902);
xor (n6901,n6763,n6764);
and (n6902,n124,n238);
and (n6903,n6904,n6905);
xor (n6904,n6901,n6902);
or (n6905,n6906,n6909);
and (n6906,n6907,n6908);
xor (n6907,n6769,n6770);
and (n6908,n118,n238);
and (n6909,n6910,n6911);
xor (n6910,n6907,n6908);
or (n6911,n6912,n6915);
and (n6912,n6913,n6914);
xor (n6913,n6775,n6776);
and (n6914,n150,n238);
and (n6915,n6916,n6917);
xor (n6916,n6913,n6914);
or (n6917,n6918,n6921);
and (n6918,n6919,n6920);
xor (n6919,n6781,n6782);
and (n6920,n144,n238);
and (n6921,n6922,n6923);
xor (n6922,n6919,n6920);
or (n6923,n6924,n6927);
and (n6924,n6925,n6926);
xor (n6925,n6787,n6788);
and (n6926,n398,n238);
and (n6927,n6928,n6929);
xor (n6928,n6925,n6926);
or (n6929,n6930,n6933);
and (n6930,n6931,n6932);
xor (n6931,n6793,n6794);
and (n6932,n449,n238);
and (n6933,n6934,n6935);
xor (n6934,n6931,n6932);
or (n6935,n6936,n6938);
and (n6936,n6937,n3387);
xor (n6937,n6799,n6800);
and (n6938,n6939,n6940);
xor (n6939,n6937,n3387);
or (n6940,n6941,n6944);
and (n6941,n6942,n6943);
xor (n6942,n6805,n6806);
and (n6943,n551,n238);
and (n6944,n6945,n6946);
xor (n6945,n6942,n6943);
or (n6946,n6947,n6950);
and (n6947,n6948,n6949);
xor (n6948,n6811,n6812);
and (n6949,n308,n238);
and (n6950,n6951,n6952);
xor (n6951,n6948,n6949);
or (n6952,n6953,n6955);
and (n6953,n6954,n2588);
xor (n6954,n6817,n6818);
and (n6955,n6956,n6957);
xor (n6956,n6954,n2588);
or (n6957,n6958,n6961);
and (n6958,n6959,n6960);
xor (n6959,n6823,n6824);
and (n6960,n670,n238);
and (n6961,n6962,n6963);
xor (n6962,n6959,n6960);
or (n6963,n6964,n6967);
and (n6964,n6965,n6966);
xor (n6965,n6829,n6830);
and (n6966,n889,n238);
and (n6967,n6968,n6969);
xor (n6968,n6965,n6966);
or (n6969,n6970,n6973);
and (n6970,n6971,n6972);
xor (n6971,n6835,n6836);
and (n6972,n1064,n238);
and (n6973,n6974,n6975);
xor (n6974,n6971,n6972);
or (n6975,n6976,n6979);
and (n6976,n6977,n6978);
xor (n6977,n6841,n6842);
and (n6978,n1103,n238);
and (n6979,n6980,n6981);
xor (n6980,n6977,n6978);
and (n6981,n6982,n6983);
xor (n6982,n6847,n6848);
and (n6983,n1266,n238);
and (n6984,n377,n266);
or (n6985,n6986,n6989);
and (n6986,n6987,n6988);
xor (n6987,n6856,n6857);
and (n6988,n436,n266);
and (n6989,n6990,n6991);
xor (n6990,n6987,n6988);
or (n6991,n6992,n6995);
and (n6992,n6993,n6994);
xor (n6993,n6862,n6863);
and (n6994,n281,n266);
and (n6995,n6996,n6997);
xor (n6996,n6993,n6994);
or (n6997,n6998,n7001);
and (n6998,n6999,n7000);
xor (n6999,n6868,n6869);
and (n7000,n274,n266);
and (n7001,n7002,n7003);
xor (n7002,n6999,n7000);
or (n7003,n7004,n7007);
and (n7004,n7005,n7006);
xor (n7005,n6874,n6875);
and (n7006,n201,n266);
and (n7007,n7008,n7009);
xor (n7008,n7005,n7006);
or (n7009,n7010,n7013);
and (n7010,n7011,n7012);
xor (n7011,n6880,n6881);
and (n7012,n195,n266);
and (n7013,n7014,n7015);
xor (n7014,n7011,n7012);
or (n7015,n7016,n7019);
and (n7016,n7017,n7018);
xor (n7017,n6886,n6887);
and (n7018,n223,n266);
and (n7019,n7020,n7021);
xor (n7020,n7017,n7018);
or (n7021,n7022,n7025);
and (n7022,n7023,n7024);
xor (n7023,n6892,n6893);
and (n7024,n217,n266);
and (n7025,n7026,n7027);
xor (n7026,n7023,n7024);
or (n7027,n7028,n7031);
and (n7028,n7029,n7030);
xor (n7029,n6898,n6899);
and (n7030,n124,n266);
and (n7031,n7032,n7033);
xor (n7032,n7029,n7030);
or (n7033,n7034,n7037);
and (n7034,n7035,n7036);
xor (n7035,n6904,n6905);
and (n7036,n118,n266);
and (n7037,n7038,n7039);
xor (n7038,n7035,n7036);
or (n7039,n7040,n7043);
and (n7040,n7041,n7042);
xor (n7041,n6910,n6911);
and (n7042,n150,n266);
and (n7043,n7044,n7045);
xor (n7044,n7041,n7042);
or (n7045,n7046,n7049);
and (n7046,n7047,n7048);
xor (n7047,n6916,n6917);
and (n7048,n144,n266);
and (n7049,n7050,n7051);
xor (n7050,n7047,n7048);
or (n7051,n7052,n7055);
and (n7052,n7053,n7054);
xor (n7053,n6922,n6923);
and (n7054,n398,n266);
and (n7055,n7056,n7057);
xor (n7056,n7053,n7054);
or (n7057,n7058,n7061);
and (n7058,n7059,n7060);
xor (n7059,n6928,n6929);
and (n7060,n449,n266);
and (n7061,n7062,n7063);
xor (n7062,n7059,n7060);
or (n7063,n7064,n7067);
and (n7064,n7065,n7066);
xor (n7065,n6934,n6935);
and (n7066,n443,n266);
and (n7067,n7068,n7069);
xor (n7068,n7065,n7066);
or (n7069,n7070,n7073);
and (n7070,n7071,n7072);
xor (n7071,n6939,n6940);
and (n7072,n551,n266);
and (n7073,n7074,n7075);
xor (n7074,n7071,n7072);
or (n7075,n7076,n7079);
and (n7076,n7077,n7078);
xor (n7077,n6945,n6946);
and (n7078,n308,n266);
and (n7079,n7080,n7081);
xor (n7080,n7077,n7078);
or (n7081,n7082,n7085);
and (n7082,n7083,n7084);
xor (n7083,n6951,n6952);
and (n7084,n302,n266);
and (n7085,n7086,n7087);
xor (n7086,n7083,n7084);
or (n7087,n7088,n7091);
and (n7088,n7089,n7090);
xor (n7089,n6956,n6957);
and (n7090,n670,n266);
and (n7091,n7092,n7093);
xor (n7092,n7089,n7090);
or (n7093,n7094,n7097);
and (n7094,n7095,n7096);
xor (n7095,n6962,n6963);
and (n7096,n889,n266);
and (n7097,n7098,n7099);
xor (n7098,n7095,n7096);
or (n7099,n7100,n7103);
and (n7100,n7101,n7102);
xor (n7101,n6968,n6969);
and (n7102,n1064,n266);
and (n7103,n7104,n7105);
xor (n7104,n7101,n7102);
or (n7105,n7106,n7109);
and (n7106,n7107,n7108);
xor (n7107,n6974,n6975);
and (n7108,n1103,n266);
and (n7109,n7110,n7111);
xor (n7110,n7107,n7108);
and (n7111,n7112,n2832);
xor (n7112,n6980,n6981);
and (n7113,n436,n265);
or (n7114,n7115,n7118);
and (n7115,n7116,n7117);
xor (n7116,n6990,n6991);
and (n7117,n281,n265);
and (n7118,n7119,n7120);
xor (n7119,n7116,n7117);
or (n7120,n7121,n7124);
and (n7121,n7122,n7123);
xor (n7122,n6996,n6997);
and (n7123,n274,n265);
and (n7124,n7125,n7126);
xor (n7125,n7122,n7123);
or (n7126,n7127,n7130);
and (n7127,n7128,n7129);
xor (n7128,n7002,n7003);
and (n7129,n201,n265);
and (n7130,n7131,n7132);
xor (n7131,n7128,n7129);
or (n7132,n7133,n7136);
and (n7133,n7134,n7135);
xor (n7134,n7008,n7009);
and (n7135,n195,n265);
and (n7136,n7137,n7138);
xor (n7137,n7134,n7135);
or (n7138,n7139,n7142);
and (n7139,n7140,n7141);
xor (n7140,n7014,n7015);
and (n7141,n223,n265);
and (n7142,n7143,n7144);
xor (n7143,n7140,n7141);
or (n7144,n7145,n7148);
and (n7145,n7146,n7147);
xor (n7146,n7020,n7021);
and (n7147,n217,n265);
and (n7148,n7149,n7150);
xor (n7149,n7146,n7147);
or (n7150,n7151,n7154);
and (n7151,n7152,n7153);
xor (n7152,n7026,n7027);
and (n7153,n124,n265);
and (n7154,n7155,n7156);
xor (n7155,n7152,n7153);
or (n7156,n7157,n7160);
and (n7157,n7158,n7159);
xor (n7158,n7032,n7033);
and (n7159,n118,n265);
and (n7160,n7161,n7162);
xor (n7161,n7158,n7159);
or (n7162,n7163,n7166);
and (n7163,n7164,n7165);
xor (n7164,n7038,n7039);
and (n7165,n150,n265);
and (n7166,n7167,n7168);
xor (n7167,n7164,n7165);
or (n7168,n7169,n7172);
and (n7169,n7170,n7171);
xor (n7170,n7044,n7045);
and (n7171,n144,n265);
and (n7172,n7173,n7174);
xor (n7173,n7170,n7171);
or (n7174,n7175,n7178);
and (n7175,n7176,n7177);
xor (n7176,n7050,n7051);
and (n7177,n398,n265);
and (n7178,n7179,n7180);
xor (n7179,n7176,n7177);
or (n7180,n7181,n7184);
and (n7181,n7182,n7183);
xor (n7182,n7056,n7057);
and (n7183,n449,n265);
and (n7184,n7185,n7186);
xor (n7185,n7182,n7183);
or (n7186,n7187,n7190);
and (n7187,n7188,n7189);
xor (n7188,n7062,n7063);
and (n7189,n443,n265);
and (n7190,n7191,n7192);
xor (n7191,n7188,n7189);
or (n7192,n7193,n7196);
and (n7193,n7194,n7195);
xor (n7194,n7068,n7069);
and (n7195,n551,n265);
and (n7196,n7197,n7198);
xor (n7197,n7194,n7195);
or (n7198,n7199,n7202);
and (n7199,n7200,n7201);
xor (n7200,n7074,n7075);
and (n7201,n308,n265);
and (n7202,n7203,n7204);
xor (n7203,n7200,n7201);
or (n7204,n7205,n7208);
and (n7205,n7206,n7207);
xor (n7206,n7080,n7081);
and (n7207,n302,n265);
and (n7208,n7209,n7210);
xor (n7209,n7206,n7207);
or (n7210,n7211,n7214);
and (n7211,n7212,n7213);
xor (n7212,n7086,n7087);
and (n7213,n670,n265);
and (n7214,n7215,n7216);
xor (n7215,n7212,n7213);
or (n7216,n7217,n7220);
and (n7217,n7218,n7219);
xor (n7218,n7092,n7093);
and (n7219,n889,n265);
and (n7220,n7221,n7222);
xor (n7221,n7218,n7219);
or (n7222,n7223,n7226);
and (n7223,n7224,n7225);
xor (n7224,n7098,n7099);
and (n7225,n1064,n265);
and (n7226,n7227,n7228);
xor (n7227,n7224,n7225);
or (n7228,n7229,n7232);
and (n7229,n7230,n7231);
xor (n7230,n7104,n7105);
and (n7231,n1103,n265);
and (n7232,n7233,n7234);
xor (n7233,n7230,n7231);
and (n7234,n7235,n7236);
xor (n7235,n7110,n7111);
and (n7236,n1266,n265);
and (n7237,n281,n348);
or (n7238,n7239,n7242);
and (n7239,n7240,n7241);
xor (n7240,n7119,n7120);
and (n7241,n274,n348);
and (n7242,n7243,n7244);
xor (n7243,n7240,n7241);
or (n7244,n7245,n7248);
and (n7245,n7246,n7247);
xor (n7246,n7125,n7126);
and (n7247,n201,n348);
and (n7248,n7249,n7250);
xor (n7249,n7246,n7247);
or (n7250,n7251,n7254);
and (n7251,n7252,n7253);
xor (n7252,n7131,n7132);
and (n7253,n195,n348);
and (n7254,n7255,n7256);
xor (n7255,n7252,n7253);
or (n7256,n7257,n7260);
and (n7257,n7258,n7259);
xor (n7258,n7137,n7138);
and (n7259,n223,n348);
and (n7260,n7261,n7262);
xor (n7261,n7258,n7259);
or (n7262,n7263,n7266);
and (n7263,n7264,n7265);
xor (n7264,n7143,n7144);
and (n7265,n217,n348);
and (n7266,n7267,n7268);
xor (n7267,n7264,n7265);
or (n7268,n7269,n7272);
and (n7269,n7270,n7271);
xor (n7270,n7149,n7150);
and (n7271,n124,n348);
and (n7272,n7273,n7274);
xor (n7273,n7270,n7271);
or (n7274,n7275,n7278);
and (n7275,n7276,n7277);
xor (n7276,n7155,n7156);
and (n7277,n118,n348);
and (n7278,n7279,n7280);
xor (n7279,n7276,n7277);
or (n7280,n7281,n7284);
and (n7281,n7282,n7283);
xor (n7282,n7161,n7162);
and (n7283,n150,n348);
and (n7284,n7285,n7286);
xor (n7285,n7282,n7283);
or (n7286,n7287,n7290);
and (n7287,n7288,n7289);
xor (n7288,n7167,n7168);
and (n7289,n144,n348);
and (n7290,n7291,n7292);
xor (n7291,n7288,n7289);
or (n7292,n7293,n7296);
and (n7293,n7294,n7295);
xor (n7294,n7173,n7174);
and (n7295,n398,n348);
and (n7296,n7297,n7298);
xor (n7297,n7294,n7295);
or (n7298,n7299,n7302);
and (n7299,n7300,n7301);
xor (n7300,n7179,n7180);
and (n7301,n449,n348);
and (n7302,n7303,n7304);
xor (n7303,n7300,n7301);
or (n7304,n7305,n7308);
and (n7305,n7306,n7307);
xor (n7306,n7185,n7186);
and (n7307,n443,n348);
and (n7308,n7309,n7310);
xor (n7309,n7306,n7307);
or (n7310,n7311,n7314);
and (n7311,n7312,n7313);
xor (n7312,n7191,n7192);
and (n7313,n551,n348);
and (n7314,n7315,n7316);
xor (n7315,n7312,n7313);
or (n7316,n7317,n7320);
and (n7317,n7318,n7319);
xor (n7318,n7197,n7198);
and (n7319,n308,n348);
and (n7320,n7321,n7322);
xor (n7321,n7318,n7319);
or (n7322,n7323,n7326);
and (n7323,n7324,n7325);
xor (n7324,n7203,n7204);
and (n7325,n302,n348);
and (n7326,n7327,n7328);
xor (n7327,n7324,n7325);
or (n7328,n7329,n7332);
and (n7329,n7330,n7331);
xor (n7330,n7209,n7210);
and (n7331,n670,n348);
and (n7332,n7333,n7334);
xor (n7333,n7330,n7331);
or (n7334,n7335,n7338);
and (n7335,n7336,n7337);
xor (n7336,n7215,n7216);
and (n7337,n889,n348);
and (n7338,n7339,n7340);
xor (n7339,n7336,n7337);
or (n7340,n7341,n7344);
and (n7341,n7342,n7343);
xor (n7342,n7221,n7222);
and (n7343,n1064,n348);
and (n7344,n7345,n7346);
xor (n7345,n7342,n7343);
or (n7346,n7347,n7350);
and (n7347,n7348,n7349);
xor (n7348,n7227,n7228);
and (n7349,n1103,n348);
and (n7350,n7351,n7352);
xor (n7351,n7348,n7349);
and (n7352,n7353,n2453);
xor (n7353,n7233,n7234);
and (n7354,n274,n190);
or (n7355,n7356,n7359);
and (n7356,n7357,n7358);
xor (n7357,n7243,n7244);
and (n7358,n201,n190);
and (n7359,n7360,n7361);
xor (n7360,n7357,n7358);
or (n7361,n7362,n7365);
and (n7362,n7363,n7364);
xor (n7363,n7249,n7250);
and (n7364,n195,n190);
and (n7365,n7366,n7367);
xor (n7366,n7363,n7364);
or (n7367,n7368,n7371);
and (n7368,n7369,n7370);
xor (n7369,n7255,n7256);
and (n7370,n223,n190);
and (n7371,n7372,n7373);
xor (n7372,n7369,n7370);
or (n7373,n7374,n7377);
and (n7374,n7375,n7376);
xor (n7375,n7261,n7262);
and (n7376,n217,n190);
and (n7377,n7378,n7379);
xor (n7378,n7375,n7376);
or (n7379,n7380,n7383);
and (n7380,n7381,n7382);
xor (n7381,n7267,n7268);
and (n7382,n124,n190);
and (n7383,n7384,n7385);
xor (n7384,n7381,n7382);
or (n7385,n7386,n7389);
and (n7386,n7387,n7388);
xor (n7387,n7273,n7274);
and (n7388,n118,n190);
and (n7389,n7390,n7391);
xor (n7390,n7387,n7388);
or (n7391,n7392,n7395);
and (n7392,n7393,n7394);
xor (n7393,n7279,n7280);
and (n7394,n150,n190);
and (n7395,n7396,n7397);
xor (n7396,n7393,n7394);
or (n7397,n7398,n7401);
and (n7398,n7399,n7400);
xor (n7399,n7285,n7286);
and (n7400,n144,n190);
and (n7401,n7402,n7403);
xor (n7402,n7399,n7400);
or (n7403,n7404,n7406);
and (n7404,n7405,n1635);
xor (n7405,n7291,n7292);
and (n7406,n7407,n7408);
xor (n7407,n7405,n1635);
or (n7408,n7409,n7411);
and (n7409,n7410,n1822);
xor (n7410,n7297,n7298);
and (n7411,n7412,n7413);
xor (n7412,n7410,n1822);
or (n7413,n7414,n7417);
and (n7414,n7415,n7416);
xor (n7415,n7303,n7304);
and (n7416,n443,n190);
and (n7417,n7418,n7419);
xor (n7418,n7415,n7416);
or (n7419,n7420,n7423);
and (n7420,n7421,n7422);
xor (n7421,n7309,n7310);
and (n7422,n551,n190);
and (n7423,n7424,n7425);
xor (n7424,n7421,n7422);
or (n7425,n7426,n7429);
and (n7426,n7427,n7428);
xor (n7427,n7315,n7316);
and (n7428,n308,n190);
and (n7429,n7430,n7431);
xor (n7430,n7427,n7428);
or (n7431,n7432,n7435);
and (n7432,n7433,n7434);
xor (n7433,n7321,n7322);
and (n7434,n302,n190);
and (n7435,n7436,n7437);
xor (n7436,n7433,n7434);
or (n7437,n7438,n7440);
and (n7438,n7439,n3412);
xor (n7439,n7327,n7328);
and (n7440,n7441,n7442);
xor (n7441,n7439,n3412);
or (n7442,n7443,n7445);
and (n7443,n7444,n2709);
xor (n7444,n7333,n7334);
and (n7445,n7446,n7447);
xor (n7446,n7444,n2709);
or (n7447,n7448,n7451);
and (n7448,n7449,n7450);
xor (n7449,n7339,n7340);
and (n7450,n1064,n190);
and (n7451,n7452,n7453);
xor (n7452,n7449,n7450);
or (n7453,n7454,n7457);
and (n7454,n7455,n7456);
xor (n7455,n7345,n7346);
and (n7456,n1103,n190);
and (n7457,n7458,n7459);
xor (n7458,n7455,n7456);
and (n7459,n7460,n7461);
xor (n7460,n7351,n7352);
and (n7461,n1266,n190);
and (n7462,n201,n184);
or (n7463,n7464,n7467);
and (n7464,n7465,n7466);
xor (n7465,n7360,n7361);
and (n7466,n195,n184);
and (n7467,n7468,n7469);
xor (n7468,n7465,n7466);
or (n7469,n7470,n7473);
and (n7470,n7471,n7472);
xor (n7471,n7366,n7367);
and (n7472,n223,n184);
and (n7473,n7474,n7475);
xor (n7474,n7471,n7472);
or (n7475,n7476,n7479);
and (n7476,n7477,n7478);
xor (n7477,n7372,n7373);
and (n7478,n217,n184);
and (n7479,n7480,n7481);
xor (n7480,n7477,n7478);
or (n7481,n7482,n7485);
and (n7482,n7483,n7484);
xor (n7483,n7378,n7379);
and (n7484,n124,n184);
and (n7485,n7486,n7487);
xor (n7486,n7483,n7484);
or (n7487,n7488,n7491);
and (n7488,n7489,n7490);
xor (n7489,n7384,n7385);
and (n7490,n118,n184);
and (n7491,n7492,n7493);
xor (n7492,n7489,n7490);
or (n7493,n7494,n7497);
and (n7494,n7495,n7496);
xor (n7495,n7390,n7391);
and (n7496,n150,n184);
and (n7497,n7498,n7499);
xor (n7498,n7495,n7496);
or (n7499,n7500,n7503);
and (n7500,n7501,n7502);
xor (n7501,n7396,n7397);
and (n7502,n144,n184);
and (n7503,n7504,n7505);
xor (n7504,n7501,n7502);
or (n7505,n7506,n7509);
and (n7506,n7507,n7508);
xor (n7507,n7402,n7403);
and (n7508,n398,n184);
and (n7509,n7510,n7511);
xor (n7510,n7507,n7508);
or (n7511,n7512,n7515);
and (n7512,n7513,n7514);
xor (n7513,n7407,n7408);
and (n7514,n449,n184);
and (n7515,n7516,n7517);
xor (n7516,n7513,n7514);
or (n7517,n7518,n7521);
and (n7518,n7519,n7520);
xor (n7519,n7412,n7413);
and (n7520,n443,n184);
and (n7521,n7522,n7523);
xor (n7522,n7519,n7520);
or (n7523,n7524,n7527);
and (n7524,n7525,n7526);
xor (n7525,n7418,n7419);
and (n7526,n551,n184);
and (n7527,n7528,n7529);
xor (n7528,n7525,n7526);
or (n7529,n7530,n7533);
and (n7530,n7531,n7532);
xor (n7531,n7424,n7425);
and (n7532,n308,n184);
and (n7533,n7534,n7535);
xor (n7534,n7531,n7532);
or (n7535,n7536,n7539);
and (n7536,n7537,n7538);
xor (n7537,n7430,n7431);
and (n7538,n302,n184);
and (n7539,n7540,n7541);
xor (n7540,n7537,n7538);
or (n7541,n7542,n7545);
and (n7542,n7543,n7544);
xor (n7543,n7436,n7437);
and (n7544,n670,n184);
and (n7545,n7546,n7547);
xor (n7546,n7543,n7544);
or (n7547,n7548,n7551);
and (n7548,n7549,n7550);
xor (n7549,n7441,n7442);
and (n7550,n889,n184);
and (n7551,n7552,n7553);
xor (n7552,n7549,n7550);
or (n7553,n7554,n7557);
and (n7554,n7555,n7556);
xor (n7555,n7446,n7447);
and (n7556,n1064,n184);
and (n7557,n7558,n7559);
xor (n7558,n7555,n7556);
or (n7559,n7560,n7563);
and (n7560,n7561,n7562);
xor (n7561,n7452,n7453);
and (n7562,n1103,n184);
and (n7563,n7564,n7565);
xor (n7564,n7561,n7562);
and (n7565,n7566,n2766);
xor (n7566,n7458,n7459);
and (n7567,n195,n185);
or (n7568,n7569,n7572);
and (n7569,n7570,n7571);
xor (n7570,n7468,n7469);
and (n7571,n223,n185);
and (n7572,n7573,n7574);
xor (n7573,n7570,n7571);
or (n7574,n7575,n7578);
and (n7575,n7576,n7577);
xor (n7576,n7474,n7475);
and (n7577,n217,n185);
and (n7578,n7579,n7580);
xor (n7579,n7576,n7577);
or (n7580,n7581,n7584);
and (n7581,n7582,n7583);
xor (n7582,n7480,n7481);
and (n7583,n124,n185);
and (n7584,n7585,n7586);
xor (n7585,n7582,n7583);
or (n7586,n7587,n7590);
and (n7587,n7588,n7589);
xor (n7588,n7486,n7487);
and (n7589,n118,n185);
and (n7590,n7591,n7592);
xor (n7591,n7588,n7589);
or (n7592,n7593,n7596);
and (n7593,n7594,n7595);
xor (n7594,n7492,n7493);
and (n7595,n150,n185);
and (n7596,n7597,n7598);
xor (n7597,n7594,n7595);
or (n7598,n7599,n7602);
and (n7599,n7600,n7601);
xor (n7600,n7498,n7499);
and (n7601,n144,n185);
and (n7602,n7603,n7604);
xor (n7603,n7600,n7601);
or (n7604,n7605,n7608);
and (n7605,n7606,n7607);
xor (n7606,n7504,n7505);
and (n7607,n398,n185);
and (n7608,n7609,n7610);
xor (n7609,n7606,n7607);
or (n7610,n7611,n7614);
and (n7611,n7612,n7613);
xor (n7612,n7510,n7511);
and (n7613,n449,n185);
and (n7614,n7615,n7616);
xor (n7615,n7612,n7613);
or (n7616,n7617,n7620);
and (n7617,n7618,n7619);
xor (n7618,n7516,n7517);
and (n7619,n443,n185);
and (n7620,n7621,n7622);
xor (n7621,n7618,n7619);
or (n7622,n7623,n7626);
and (n7623,n7624,n7625);
xor (n7624,n7522,n7523);
and (n7625,n551,n185);
and (n7626,n7627,n7628);
xor (n7627,n7624,n7625);
or (n7628,n7629,n7632);
and (n7629,n7630,n7631);
xor (n7630,n7528,n7529);
and (n7631,n308,n185);
and (n7632,n7633,n7634);
xor (n7633,n7630,n7631);
or (n7634,n7635,n7638);
and (n7635,n7636,n7637);
xor (n7636,n7534,n7535);
and (n7637,n302,n185);
and (n7638,n7639,n7640);
xor (n7639,n7636,n7637);
or (n7640,n7641,n7644);
and (n7641,n7642,n7643);
xor (n7642,n7540,n7541);
and (n7643,n670,n185);
and (n7644,n7645,n7646);
xor (n7645,n7642,n7643);
or (n7646,n7647,n7650);
and (n7647,n7648,n7649);
xor (n7648,n7546,n7547);
and (n7649,n889,n185);
and (n7650,n7651,n7652);
xor (n7651,n7648,n7649);
or (n7652,n7653,n7656);
and (n7653,n7654,n7655);
xor (n7654,n7552,n7553);
and (n7655,n1064,n185);
and (n7656,n7657,n7658);
xor (n7657,n7654,n7655);
or (n7658,n7659,n7662);
and (n7659,n7660,n7661);
xor (n7660,n7558,n7559);
and (n7661,n1103,n185);
and (n7662,n7663,n7664);
xor (n7663,n7660,n7661);
and (n7664,n7665,n7666);
xor (n7665,n7564,n7565);
and (n7666,n1266,n185);
and (n7667,n223,n209);
or (n7668,n7669,n7672);
and (n7669,n7670,n7671);
xor (n7670,n7573,n7574);
and (n7671,n217,n209);
and (n7672,n7673,n7674);
xor (n7673,n7670,n7671);
or (n7674,n7675,n7678);
and (n7675,n7676,n7677);
xor (n7676,n7579,n7580);
and (n7677,n124,n209);
and (n7678,n7679,n7680);
xor (n7679,n7676,n7677);
or (n7680,n7681,n7684);
and (n7681,n7682,n7683);
xor (n7682,n7585,n7586);
and (n7683,n118,n209);
and (n7684,n7685,n7686);
xor (n7685,n7682,n7683);
or (n7686,n7687,n7690);
and (n7687,n7688,n7689);
xor (n7688,n7591,n7592);
and (n7689,n150,n209);
and (n7690,n7691,n7692);
xor (n7691,n7688,n7689);
or (n7692,n7693,n7696);
and (n7693,n7694,n7695);
xor (n7694,n7597,n7598);
and (n7695,n144,n209);
and (n7696,n7697,n7698);
xor (n7697,n7694,n7695);
or (n7698,n7699,n7702);
and (n7699,n7700,n7701);
xor (n7700,n7603,n7604);
and (n7701,n398,n209);
and (n7702,n7703,n7704);
xor (n7703,n7700,n7701);
or (n7704,n7705,n7708);
and (n7705,n7706,n7707);
xor (n7706,n7609,n7610);
and (n7707,n449,n209);
and (n7708,n7709,n7710);
xor (n7709,n7706,n7707);
or (n7710,n7711,n7714);
and (n7711,n7712,n7713);
xor (n7712,n7615,n7616);
and (n7713,n443,n209);
and (n7714,n7715,n7716);
xor (n7715,n7712,n7713);
or (n7716,n7717,n7720);
and (n7717,n7718,n7719);
xor (n7718,n7621,n7622);
and (n7719,n551,n209);
and (n7720,n7721,n7722);
xor (n7721,n7718,n7719);
or (n7722,n7723,n7726);
and (n7723,n7724,n7725);
xor (n7724,n7627,n7628);
and (n7725,n308,n209);
and (n7726,n7727,n7728);
xor (n7727,n7724,n7725);
or (n7728,n7729,n7732);
and (n7729,n7730,n7731);
xor (n7730,n7633,n7634);
and (n7731,n302,n209);
and (n7732,n7733,n7734);
xor (n7733,n7730,n7731);
or (n7734,n7735,n7738);
and (n7735,n7736,n7737);
xor (n7736,n7639,n7640);
and (n7737,n670,n209);
and (n7738,n7739,n7740);
xor (n7739,n7736,n7737);
or (n7740,n7741,n7744);
and (n7741,n7742,n7743);
xor (n7742,n7645,n7646);
and (n7743,n889,n209);
and (n7744,n7745,n7746);
xor (n7745,n7742,n7743);
or (n7746,n7747,n7750);
and (n7747,n7748,n7749);
xor (n7748,n7651,n7652);
and (n7749,n1064,n209);
and (n7750,n7751,n7752);
xor (n7751,n7748,n7749);
or (n7752,n7753,n7756);
and (n7753,n7754,n7755);
xor (n7754,n7657,n7658);
and (n7755,n1103,n209);
and (n7756,n7757,n7758);
xor (n7757,n7754,n7755);
and (n7758,n7759,n3516);
xor (n7759,n7663,n7664);
and (n7760,n217,n114);
or (n7761,n7762,n7765);
and (n7762,n7763,n7764);
xor (n7763,n7673,n7674);
and (n7764,n124,n114);
and (n7765,n7766,n7767);
xor (n7766,n7763,n7764);
or (n7767,n7768,n7771);
and (n7768,n7769,n7770);
xor (n7769,n7679,n7680);
and (n7770,n118,n114);
and (n7771,n7772,n7773);
xor (n7772,n7769,n7770);
or (n7773,n7774,n7777);
and (n7774,n7775,n7776);
xor (n7775,n7685,n7686);
and (n7776,n150,n114);
and (n7777,n7778,n7779);
xor (n7778,n7775,n7776);
or (n7779,n7780,n7783);
and (n7780,n7781,n7782);
xor (n7781,n7691,n7692);
and (n7782,n144,n114);
and (n7783,n7784,n7785);
xor (n7784,n7781,n7782);
or (n7785,n7786,n7789);
and (n7786,n7787,n7788);
xor (n7787,n7697,n7698);
and (n7788,n398,n114);
and (n7789,n7790,n7791);
xor (n7790,n7787,n7788);
or (n7791,n7792,n7795);
and (n7792,n7793,n7794);
xor (n7793,n7703,n7704);
and (n7794,n449,n114);
and (n7795,n7796,n7797);
xor (n7796,n7793,n7794);
or (n7797,n7798,n7801);
and (n7798,n7799,n7800);
xor (n7799,n7709,n7710);
and (n7800,n443,n114);
and (n7801,n7802,n7803);
xor (n7802,n7799,n7800);
or (n7803,n7804,n7807);
and (n7804,n7805,n7806);
xor (n7805,n7715,n7716);
and (n7806,n551,n114);
and (n7807,n7808,n7809);
xor (n7808,n7805,n7806);
or (n7809,n7810,n7813);
and (n7810,n7811,n7812);
xor (n7811,n7721,n7722);
and (n7812,n308,n114);
and (n7813,n7814,n7815);
xor (n7814,n7811,n7812);
or (n7815,n7816,n7819);
and (n7816,n7817,n7818);
xor (n7817,n7727,n7728);
and (n7818,n302,n114);
and (n7819,n7820,n7821);
xor (n7820,n7817,n7818);
or (n7821,n7822,n7825);
and (n7822,n7823,n7824);
xor (n7823,n7733,n7734);
and (n7824,n670,n114);
and (n7825,n7826,n7827);
xor (n7826,n7823,n7824);
or (n7827,n7828,n7831);
and (n7828,n7829,n7830);
xor (n7829,n7739,n7740);
and (n7830,n889,n114);
and (n7831,n7832,n7833);
xor (n7832,n7829,n7830);
or (n7833,n7834,n7837);
and (n7834,n7835,n7836);
xor (n7835,n7745,n7746);
and (n7836,n1064,n114);
and (n7837,n7838,n7839);
xor (n7838,n7835,n7836);
or (n7839,n7840,n7843);
and (n7840,n7841,n7842);
xor (n7841,n7751,n7752);
and (n7842,n1103,n114);
and (n7843,n7844,n7845);
xor (n7844,n7841,n7842);
and (n7845,n7846,n7847);
xor (n7846,n7757,n7758);
and (n7847,n1266,n114);
and (n7848,n124,n108);
or (n7849,n7850,n7853);
and (n7850,n7851,n7852);
xor (n7851,n7766,n7767);
and (n7852,n118,n108);
and (n7853,n7854,n7855);
xor (n7854,n7851,n7852);
or (n7855,n7856,n7859);
and (n7856,n7857,n7858);
xor (n7857,n7772,n7773);
and (n7858,n150,n108);
and (n7859,n7860,n7861);
xor (n7860,n7857,n7858);
or (n7861,n7862,n7865);
and (n7862,n7863,n7864);
xor (n7863,n7778,n7779);
and (n7864,n144,n108);
and (n7865,n7866,n7867);
xor (n7866,n7863,n7864);
or (n7867,n7868,n7871);
and (n7868,n7869,n7870);
xor (n7869,n7784,n7785);
and (n7870,n398,n108);
and (n7871,n7872,n7873);
xor (n7872,n7869,n7870);
or (n7873,n7874,n7877);
and (n7874,n7875,n7876);
xor (n7875,n7790,n7791);
and (n7876,n449,n108);
and (n7877,n7878,n7879);
xor (n7878,n7875,n7876);
or (n7879,n7880,n7883);
and (n7880,n7881,n7882);
xor (n7881,n7796,n7797);
and (n7882,n443,n108);
and (n7883,n7884,n7885);
xor (n7884,n7881,n7882);
or (n7885,n7886,n7889);
and (n7886,n7887,n7888);
xor (n7887,n7802,n7803);
and (n7888,n551,n108);
and (n7889,n7890,n7891);
xor (n7890,n7887,n7888);
or (n7891,n7892,n7895);
and (n7892,n7893,n7894);
xor (n7893,n7808,n7809);
and (n7894,n308,n108);
and (n7895,n7896,n7897);
xor (n7896,n7893,n7894);
or (n7897,n7898,n7901);
and (n7898,n7899,n7900);
xor (n7899,n7814,n7815);
and (n7900,n302,n108);
and (n7901,n7902,n7903);
xor (n7902,n7899,n7900);
or (n7903,n7904,n7907);
and (n7904,n7905,n7906);
xor (n7905,n7820,n7821);
and (n7906,n670,n108);
and (n7907,n7908,n7909);
xor (n7908,n7905,n7906);
or (n7909,n7910,n7913);
and (n7910,n7911,n7912);
xor (n7911,n7826,n7827);
and (n7912,n889,n108);
and (n7913,n7914,n7915);
xor (n7914,n7911,n7912);
or (n7915,n7916,n7919);
and (n7916,n7917,n7918);
xor (n7917,n7832,n7833);
and (n7918,n1064,n108);
and (n7919,n7920,n7921);
xor (n7920,n7917,n7918);
or (n7921,n7922,n7925);
and (n7922,n7923,n7924);
xor (n7923,n7838,n7839);
and (n7924,n1103,n108);
and (n7925,n7926,n7927);
xor (n7926,n7923,n7924);
and (n7927,n7928,n2280);
xor (n7928,n7844,n7845);
and (n7929,n118,n106);
or (n7930,n7931,n7934);
and (n7931,n7932,n7933);
xor (n7932,n7854,n7855);
and (n7933,n150,n106);
and (n7934,n7935,n7936);
xor (n7935,n7932,n7933);
or (n7936,n7937,n7940);
and (n7937,n7938,n7939);
xor (n7938,n7860,n7861);
and (n7939,n144,n106);
and (n7940,n7941,n7942);
xor (n7941,n7938,n7939);
or (n7942,n7943,n7945);
and (n7943,n7944,n399);
xor (n7944,n7866,n7867);
and (n7945,n7946,n7947);
xor (n7946,n7944,n399);
or (n7947,n7948,n7950);
and (n7948,n7949,n760);
xor (n7949,n7872,n7873);
and (n7950,n7951,n7952);
xor (n7951,n7949,n760);
or (n7952,n7953,n7956);
and (n7953,n7954,n7955);
xor (n7954,n7878,n7879);
and (n7955,n443,n106);
and (n7956,n7957,n7958);
xor (n7957,n7954,n7955);
or (n7958,n7959,n7962);
and (n7959,n7960,n7961);
xor (n7960,n7884,n7885);
and (n7961,n551,n106);
and (n7962,n7963,n7964);
xor (n7963,n7960,n7961);
or (n7964,n7965,n7968);
and (n7965,n7966,n7967);
xor (n7966,n7890,n7891);
and (n7967,n308,n106);
and (n7968,n7969,n7970);
xor (n7969,n7966,n7967);
or (n7970,n7971,n7974);
and (n7971,n7972,n7973);
xor (n7972,n7896,n7897);
and (n7973,n302,n106);
and (n7974,n7975,n7976);
xor (n7975,n7972,n7973);
or (n7976,n7977,n7980);
and (n7977,n7978,n7979);
xor (n7978,n7902,n7903);
and (n7979,n670,n106);
and (n7980,n7981,n7982);
xor (n7981,n7978,n7979);
or (n7982,n7983,n7986);
and (n7983,n7984,n7985);
xor (n7984,n7908,n7909);
and (n7985,n889,n106);
and (n7986,n7987,n7988);
xor (n7987,n7984,n7985);
or (n7988,n7989,n7992);
and (n7989,n7990,n7991);
xor (n7990,n7914,n7915);
and (n7991,n1064,n106);
and (n7992,n7993,n7994);
xor (n7993,n7990,n7991);
or (n7994,n7995,n7998);
and (n7995,n7996,n7997);
xor (n7996,n7920,n7921);
and (n7997,n1103,n106);
and (n7998,n7999,n8000);
xor (n7999,n7996,n7997);
and (n8000,n8001,n8002);
xor (n8001,n7926,n7927);
and (n8002,n1266,n106);
and (n8003,n150,n134);
or (n8004,n8005,n8008);
and (n8005,n8006,n8007);
xor (n8006,n7935,n7936);
and (n8007,n144,n134);
and (n8008,n8009,n8010);
xor (n8009,n8006,n8007);
or (n8010,n8011,n8014);
and (n8011,n8012,n8013);
xor (n8012,n7941,n7942);
and (n8013,n398,n134);
and (n8014,n8015,n8016);
xor (n8015,n8012,n8013);
or (n8016,n8017,n8020);
and (n8017,n8018,n8019);
xor (n8018,n7946,n7947);
and (n8019,n449,n134);
and (n8020,n8021,n8022);
xor (n8021,n8018,n8019);
or (n8022,n8023,n8026);
and (n8023,n8024,n8025);
xor (n8024,n7951,n7952);
and (n8025,n443,n134);
and (n8026,n8027,n8028);
xor (n8027,n8024,n8025);
or (n8028,n8029,n8032);
and (n8029,n8030,n8031);
xor (n8030,n7957,n7958);
and (n8031,n551,n134);
and (n8032,n8033,n8034);
xor (n8033,n8030,n8031);
or (n8034,n8035,n8038);
and (n8035,n8036,n8037);
xor (n8036,n7963,n7964);
and (n8037,n308,n134);
and (n8038,n8039,n8040);
xor (n8039,n8036,n8037);
or (n8040,n8041,n8044);
and (n8041,n8042,n8043);
xor (n8042,n7969,n7970);
and (n8043,n302,n134);
and (n8044,n8045,n8046);
xor (n8045,n8042,n8043);
or (n8046,n8047,n8050);
and (n8047,n8048,n8049);
xor (n8048,n7975,n7976);
and (n8049,n670,n134);
and (n8050,n8051,n8052);
xor (n8051,n8048,n8049);
or (n8052,n8053,n8056);
and (n8053,n8054,n8055);
xor (n8054,n7981,n7982);
and (n8055,n889,n134);
and (n8056,n8057,n8058);
xor (n8057,n8054,n8055);
or (n8058,n8059,n8062);
and (n8059,n8060,n8061);
xor (n8060,n7987,n7988);
and (n8061,n1064,n134);
and (n8062,n8063,n8064);
xor (n8063,n8060,n8061);
or (n8064,n8065,n8068);
and (n8065,n8066,n8067);
xor (n8066,n7993,n7994);
and (n8067,n1103,n134);
and (n8068,n8069,n8070);
xor (n8069,n8066,n8067);
and (n8070,n8071,n2030);
xor (n8071,n7999,n8000);
and (n8072,n144,n140);
or (n8073,n8074,n8077);
and (n8074,n8075,n8076);
xor (n8075,n8009,n8010);
and (n8076,n398,n140);
and (n8077,n8078,n8079);
xor (n8078,n8075,n8076);
or (n8079,n8080,n8083);
and (n8080,n8081,n8082);
xor (n8081,n8015,n8016);
and (n8082,n449,n140);
and (n8083,n8084,n8085);
xor (n8084,n8081,n8082);
or (n8085,n8086,n8089);
and (n8086,n8087,n8088);
xor (n8087,n8021,n8022);
and (n8088,n443,n140);
and (n8089,n8090,n8091);
xor (n8090,n8087,n8088);
or (n8091,n8092,n8095);
and (n8092,n8093,n8094);
xor (n8093,n8027,n8028);
and (n8094,n551,n140);
and (n8095,n8096,n8097);
xor (n8096,n8093,n8094);
or (n8097,n8098,n8101);
and (n8098,n8099,n8100);
xor (n8099,n8033,n8034);
and (n8100,n308,n140);
and (n8101,n8102,n8103);
xor (n8102,n8099,n8100);
or (n8103,n8104,n8107);
and (n8104,n8105,n8106);
xor (n8105,n8039,n8040);
and (n8106,n302,n140);
and (n8107,n8108,n8109);
xor (n8108,n8105,n8106);
or (n8109,n8110,n8113);
and (n8110,n8111,n8112);
xor (n8111,n8045,n8046);
and (n8112,n670,n140);
and (n8113,n8114,n8115);
xor (n8114,n8111,n8112);
or (n8115,n8116,n8119);
and (n8116,n8117,n8118);
xor (n8117,n8051,n8052);
and (n8118,n889,n140);
and (n8119,n8120,n8121);
xor (n8120,n8117,n8118);
or (n8121,n8122,n8125);
and (n8122,n8123,n8124);
xor (n8123,n8057,n8058);
and (n8124,n1064,n140);
and (n8125,n8126,n8127);
xor (n8126,n8123,n8124);
or (n8127,n8128,n8131);
and (n8128,n8129,n8130);
xor (n8129,n8063,n8064);
and (n8130,n1103,n140);
and (n8131,n8132,n8133);
xor (n8132,n8129,n8130);
and (n8133,n8134,n8135);
xor (n8134,n8069,n8070);
and (n8135,n1266,n140);
and (n8136,n398,n533);
or (n8137,n8138,n8141);
and (n8138,n8139,n8140);
xor (n8139,n8078,n8079);
and (n8140,n449,n533);
and (n8141,n8142,n8143);
xor (n8142,n8139,n8140);
or (n8143,n8144,n8147);
and (n8144,n8145,n8146);
xor (n8145,n8084,n8085);
and (n8146,n443,n533);
and (n8147,n8148,n8149);
xor (n8148,n8145,n8146);
or (n8149,n8150,n8153);
and (n8150,n8151,n8152);
xor (n8151,n8090,n8091);
and (n8152,n551,n533);
and (n8153,n8154,n8155);
xor (n8154,n8151,n8152);
or (n8155,n8156,n8159);
and (n8156,n8157,n8158);
xor (n8157,n8096,n8097);
and (n8158,n308,n533);
and (n8159,n8160,n8161);
xor (n8160,n8157,n8158);
or (n8161,n8162,n8165);
and (n8162,n8163,n8164);
xor (n8163,n8102,n8103);
and (n8164,n302,n533);
and (n8165,n8166,n8167);
xor (n8166,n8163,n8164);
or (n8167,n8168,n8171);
and (n8168,n8169,n8170);
xor (n8169,n8108,n8109);
and (n8170,n670,n533);
and (n8171,n8172,n8173);
xor (n8172,n8169,n8170);
or (n8173,n8174,n8177);
and (n8174,n8175,n8176);
xor (n8175,n8114,n8115);
and (n8176,n889,n533);
and (n8177,n8178,n8179);
xor (n8178,n8175,n8176);
or (n8179,n8180,n8183);
and (n8180,n8181,n8182);
xor (n8181,n8120,n8121);
and (n8182,n1064,n533);
and (n8183,n8184,n8185);
xor (n8184,n8181,n8182);
or (n8185,n8186,n8189);
and (n8186,n8187,n8188);
xor (n8187,n8126,n8127);
and (n8188,n1103,n533);
and (n8189,n8190,n8191);
xor (n8190,n8187,n8188);
and (n8191,n8192,n1711);
xor (n8192,n8132,n8133);
and (n8193,n449,n290);
or (n8194,n8195,n8198);
and (n8195,n8196,n8197);
xor (n8196,n8142,n8143);
and (n8197,n443,n290);
and (n8198,n8199,n8200);
xor (n8199,n8196,n8197);
or (n8200,n8201,n8204);
and (n8201,n8202,n8203);
xor (n8202,n8148,n8149);
and (n8203,n551,n290);
and (n8204,n8205,n8206);
xor (n8205,n8202,n8203);
or (n8206,n8207,n8210);
and (n8207,n8208,n8209);
xor (n8208,n8154,n8155);
and (n8209,n308,n290);
and (n8210,n8211,n8212);
xor (n8211,n8208,n8209);
or (n8212,n8213,n8216);
and (n8213,n8214,n8215);
xor (n8214,n8160,n8161);
and (n8215,n302,n290);
and (n8216,n8217,n8218);
xor (n8217,n8214,n8215);
or (n8218,n8219,n8222);
and (n8219,n8220,n8221);
xor (n8220,n8166,n8167);
and (n8221,n670,n290);
and (n8222,n8223,n8224);
xor (n8223,n8220,n8221);
or (n8224,n8225,n8228);
and (n8225,n8226,n8227);
xor (n8226,n8172,n8173);
and (n8227,n889,n290);
and (n8228,n8229,n8230);
xor (n8229,n8226,n8227);
or (n8230,n8231,n8234);
and (n8231,n8232,n8233);
xor (n8232,n8178,n8179);
and (n8233,n1064,n290);
and (n8234,n8235,n8236);
xor (n8235,n8232,n8233);
or (n8236,n8237,n8240);
and (n8237,n8238,n8239);
xor (n8238,n8184,n8185);
and (n8239,n1103,n290);
and (n8240,n8241,n8242);
xor (n8241,n8238,n8239);
and (n8242,n8243,n8244);
xor (n8243,n8190,n8191);
and (n8244,n1266,n290);
and (n8245,n443,n292);
or (n8246,n8247,n8250);
and (n8247,n8248,n8249);
xor (n8248,n8199,n8200);
and (n8249,n551,n292);
and (n8250,n8251,n8252);
xor (n8251,n8248,n8249);
or (n8252,n8253,n8256);
and (n8253,n8254,n8255);
xor (n8254,n8205,n8206);
and (n8255,n308,n292);
and (n8256,n8257,n8258);
xor (n8257,n8254,n8255);
or (n8258,n8259,n8262);
and (n8259,n8260,n8261);
xor (n8260,n8211,n8212);
and (n8261,n302,n292);
and (n8262,n8263,n8264);
xor (n8263,n8260,n8261);
or (n8264,n8265,n8268);
and (n8265,n8266,n8267);
xor (n8266,n8217,n8218);
and (n8267,n670,n292);
and (n8268,n8269,n8270);
xor (n8269,n8266,n8267);
or (n8270,n8271,n8274);
and (n8271,n8272,n8273);
xor (n8272,n8223,n8224);
and (n8273,n889,n292);
and (n8274,n8275,n8276);
xor (n8275,n8272,n8273);
or (n8276,n8277,n8280);
and (n8277,n8278,n8279);
xor (n8278,n8229,n8230);
and (n8279,n1064,n292);
and (n8280,n8281,n8282);
xor (n8281,n8278,n8279);
or (n8282,n8283,n8286);
and (n8283,n8284,n8285);
xor (n8284,n8235,n8236);
and (n8285,n1103,n292);
and (n8286,n8287,n8288);
xor (n8287,n8284,n8285);
and (n8288,n8289,n1265);
xor (n8289,n8241,n8242);
and (n8290,n551,n298);
or (n8291,n8292,n8295);
and (n8292,n8293,n8294);
xor (n8293,n8251,n8252);
and (n8294,n308,n298);
and (n8295,n8296,n8297);
xor (n8296,n8293,n8294);
or (n8297,n8298,n8301);
and (n8298,n8299,n8300);
xor (n8299,n8257,n8258);
and (n8300,n302,n298);
and (n8301,n8302,n8303);
xor (n8302,n8299,n8300);
or (n8303,n8304,n8307);
and (n8304,n8305,n8306);
xor (n8305,n8263,n8264);
and (n8306,n670,n298);
and (n8307,n8308,n8309);
xor (n8308,n8305,n8306);
or (n8309,n8310,n8313);
and (n8310,n8311,n8312);
xor (n8311,n8269,n8270);
and (n8312,n889,n298);
and (n8313,n8314,n8315);
xor (n8314,n8311,n8312);
or (n8315,n8316,n8319);
and (n8316,n8317,n8318);
xor (n8317,n8275,n8276);
and (n8318,n1064,n298);
and (n8319,n8320,n8321);
xor (n8320,n8317,n8318);
or (n8321,n8322,n8325);
and (n8322,n8323,n8324);
xor (n8323,n8281,n8282);
and (n8324,n1103,n298);
and (n8325,n8326,n8327);
xor (n8326,n8323,n8324);
and (n8327,n8328,n8329);
xor (n8328,n8287,n8288);
and (n8329,n1266,n298);
or (n8330,n8331,n8333);
and (n8331,n8332,n8300);
xor (n8332,n8296,n8297);
and (n8333,n8334,n8335);
xor (n8334,n8332,n8300);
or (n8335,n8336,n8338);
and (n8336,n8337,n8306);
xor (n8337,n8302,n8303);
and (n8338,n8339,n8340);
xor (n8339,n8337,n8306);
or (n8340,n8341,n8343);
and (n8341,n8342,n8312);
xor (n8342,n8308,n8309);
and (n8343,n8344,n8345);
xor (n8344,n8342,n8312);
or (n8345,n8346,n8348);
and (n8346,n8347,n8318);
xor (n8347,n8314,n8315);
and (n8348,n8349,n8350);
xor (n8349,n8347,n8318);
or (n8350,n8351,n8353);
and (n8351,n8352,n8324);
xor (n8352,n8320,n8321);
and (n8353,n8354,n8355);
xor (n8354,n8352,n8324);
and (n8355,n8356,n8329);
xor (n8356,n8326,n8327);
or (n8357,n8358,n8360);
and (n8358,n8359,n8306);
xor (n8359,n8334,n8335);
and (n8360,n8361,n8362);
xor (n8361,n8359,n8306);
or (n8362,n8363,n8365);
and (n8363,n8364,n8312);
xor (n8364,n8339,n8340);
and (n8365,n8366,n8367);
xor (n8366,n8364,n8312);
or (n8367,n8368,n8370);
and (n8368,n8369,n8318);
xor (n8369,n8344,n8345);
and (n8370,n8371,n8372);
xor (n8371,n8369,n8318);
or (n8372,n8373,n8375);
and (n8373,n8374,n8324);
xor (n8374,n8349,n8350);
and (n8375,n8376,n8377);
xor (n8376,n8374,n8324);
and (n8377,n8378,n8329);
xor (n8378,n8354,n8355);
or (n8379,n8380,n8382);
and (n8380,n8381,n8312);
xor (n8381,n8361,n8362);
and (n8382,n8383,n8384);
xor (n8383,n8381,n8312);
or (n8384,n8385,n8387);
and (n8385,n8386,n8318);
xor (n8386,n8366,n8367);
and (n8387,n8388,n8389);
xor (n8388,n8386,n8318);
or (n8389,n8390,n8392);
and (n8390,n8391,n8324);
xor (n8391,n8371,n8372);
and (n8392,n8393,n8394);
xor (n8393,n8391,n8324);
and (n8394,n8395,n8329);
xor (n8395,n8376,n8377);
or (n8396,n8397,n8399);
and (n8397,n8398,n8318);
xor (n8398,n8383,n8384);
and (n8399,n8400,n8401);
xor (n8400,n8398,n8318);
or (n8401,n8402,n8404);
and (n8402,n8403,n8324);
xor (n8403,n8388,n8389);
and (n8404,n8405,n8406);
xor (n8405,n8403,n8324);
and (n8406,n8407,n8329);
xor (n8407,n8393,n8394);
or (n8408,n8409,n8411);
and (n8409,n8410,n8324);
xor (n8410,n8400,n8401);
and (n8411,n8412,n8413);
xor (n8412,n8410,n8324);
and (n8413,n8414,n8329);
xor (n8414,n8405,n8406);
and (n8415,n8416,n8329);
xor (n8416,n8412,n8413);
nor (n8417,n9,n7);
and (n8418,n3,n8419);
not (n8419,n8417);
endmodule
