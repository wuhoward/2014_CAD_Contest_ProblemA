module top (out,n1,n20,n21,n23,n24,n29,n36,n43,n50
        ,n57,n63,n65,n94,n117,n134,n145,n150,n166,n167
        ,n169,n170,n175,n182,n189,n196,n203,n209,n211,n240
        ,n263,n280,n291,n296,n344,n350,n357,n364,n371,n378
        ,n385,n391,n393,n409,n410,n412,n413,n415,n416,n418
        ,n419,n421,n422);
output out;
input n1;
input n20;
input n21;
input n23;
input n24;
input n29;
input n36;
input n43;
input n50;
input n57;
input n63;
input n65;
input n94;
input n117;
input n134;
input n145;
input n150;
input n166;
input n167;
input n169;
input n170;
input n175;
input n182;
input n189;
input n196;
input n203;
input n209;
input n211;
input n240;
input n263;
input n280;
input n291;
input n296;
input n344;
input n350;
input n357;
input n364;
input n371;
input n378;
input n385;
input n391;
input n393;
input n409;
input n410;
input n412;
input n413;
input n415;
input n416;
input n418;
input n419;
input n421;
input n422;
wire n0;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n22;
wire n25;
wire n26;
wire n27;
wire n28;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n64;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n146;
wire n147;
wire n148;
wire n149;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n168;
wire n171;
wire n172;
wire n173;
wire n174;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n210;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n292;
wire n293;
wire n294;
wire n295;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n392;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n411;
wire n414;
wire n417;
wire n420;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
xor (out,n0,n423);
wire s0n0,s1n0,notn0;
or (n0,s0n0,s1n0);
not(notn0,n402);
and (s0n0,notn0,n1);
and (s1n0,n402,n2);
xor (n2,n3,n345);
xor (n3,n4,n343);
xor (n4,n5,n297);
xor (n5,n6,n151);
xor (n6,n7,n149);
xor (n7,n8,n146);
xor (n8,n9,n144);
xor (n9,n10,n135);
xor (n10,n11,n133);
xor (n11,n12,n118);
xor (n12,n13,n116);
xor (n13,n14,n95);
xor (n14,n15,n93);
xor (n15,n16,n66);
xor (n16,n17,n64);
xor (n17,n18,n25);
xor (n18,n19,n22);
and (n19,n20,n21);
and (n22,n23,n24);
or (n25,n26,n30);
and (n26,n27,n28);
and (n27,n23,n21);
and (n28,n29,n24);
and (n30,n31,n32);
xor (n31,n27,n28);
or (n32,n33,n37);
and (n33,n34,n35);
and (n34,n29,n21);
and (n35,n36,n24);
and (n37,n38,n39);
xor (n38,n34,n35);
or (n39,n40,n44);
and (n40,n41,n42);
and (n41,n36,n21);
and (n42,n43,n24);
and (n44,n45,n46);
xor (n45,n41,n42);
or (n46,n47,n51);
and (n47,n48,n49);
and (n48,n43,n21);
and (n49,n50,n24);
and (n51,n52,n53);
xor (n52,n48,n49);
or (n53,n54,n58);
and (n54,n55,n56);
and (n55,n50,n21);
and (n56,n57,n24);
and (n58,n59,n60);
xor (n59,n55,n56);
and (n60,n61,n62);
and (n61,n57,n21);
and (n62,n63,n24);
and (n64,n29,n65);
or (n66,n67,n70);
and (n67,n68,n69);
xor (n68,n31,n32);
and (n69,n36,n65);
and (n70,n71,n72);
xor (n71,n68,n69);
or (n72,n73,n76);
and (n73,n74,n75);
xor (n74,n38,n39);
and (n75,n43,n65);
and (n76,n77,n78);
xor (n77,n74,n75);
or (n78,n79,n82);
and (n79,n80,n81);
xor (n80,n45,n46);
and (n81,n50,n65);
and (n82,n83,n84);
xor (n83,n80,n81);
or (n84,n85,n88);
and (n85,n86,n87);
xor (n86,n52,n53);
and (n87,n57,n65);
and (n88,n89,n90);
xor (n89,n86,n87);
and (n90,n91,n92);
xor (n91,n59,n60);
and (n92,n63,n65);
and (n93,n36,n94);
or (n95,n96,n99);
and (n96,n97,n98);
xor (n97,n71,n72);
and (n98,n43,n94);
and (n99,n100,n101);
xor (n100,n97,n98);
or (n101,n102,n105);
and (n102,n103,n104);
xor (n103,n77,n78);
and (n104,n50,n94);
and (n105,n106,n107);
xor (n106,n103,n104);
or (n107,n108,n111);
and (n108,n109,n110);
xor (n109,n83,n84);
and (n110,n57,n94);
and (n111,n112,n113);
xor (n112,n109,n110);
and (n113,n114,n115);
xor (n114,n89,n90);
and (n115,n63,n94);
and (n116,n43,n117);
or (n118,n119,n122);
and (n119,n120,n121);
xor (n120,n100,n101);
and (n121,n50,n117);
and (n122,n123,n124);
xor (n123,n120,n121);
or (n124,n125,n128);
and (n125,n126,n127);
xor (n126,n106,n107);
and (n127,n57,n117);
and (n128,n129,n130);
xor (n129,n126,n127);
and (n130,n131,n132);
xor (n131,n112,n113);
and (n132,n63,n117);
and (n133,n50,n134);
or (n135,n136,n139);
and (n136,n137,n138);
xor (n137,n123,n124);
and (n138,n57,n134);
and (n139,n140,n141);
xor (n140,n137,n138);
and (n141,n142,n143);
xor (n142,n129,n130);
and (n143,n63,n134);
and (n144,n57,n145);
and (n146,n147,n148);
xor (n147,n140,n141);
and (n148,n63,n145);
and (n149,n63,n150);
not (n151,n152);
xor (n152,n153,n295);
xor (n153,n154,n292);
xor (n154,n155,n290);
xor (n155,n156,n281);
xor (n156,n157,n279);
xor (n157,n158,n264);
xor (n158,n159,n262);
xor (n159,n160,n241);
xor (n160,n161,n239);
xor (n161,n162,n212);
xor (n162,n163,n210);
xor (n163,n164,n171);
xor (n164,n165,n168);
and (n165,n166,n167);
and (n168,n169,n170);
or (n171,n172,n176);
and (n172,n173,n174);
and (n173,n170,n167);
and (n174,n175,n169);
and (n176,n177,n178);
xor (n177,n173,n174);
or (n178,n179,n183);
and (n179,n180,n181);
and (n180,n175,n167);
and (n181,n182,n169);
and (n183,n184,n185);
xor (n184,n180,n181);
or (n185,n186,n190);
and (n186,n187,n188);
and (n187,n182,n167);
and (n188,n189,n169);
and (n190,n191,n192);
xor (n191,n187,n188);
or (n192,n193,n197);
and (n193,n194,n195);
and (n194,n189,n167);
and (n195,n196,n169);
and (n197,n198,n199);
xor (n198,n194,n195);
or (n199,n200,n204);
and (n200,n201,n202);
and (n201,n196,n167);
and (n202,n203,n169);
and (n204,n205,n206);
xor (n205,n201,n202);
and (n206,n207,n208);
and (n207,n203,n167);
and (n208,n209,n169);
and (n210,n175,n211);
or (n212,n213,n216);
and (n213,n214,n215);
xor (n214,n177,n178);
and (n215,n182,n211);
and (n216,n217,n218);
xor (n217,n214,n215);
or (n218,n219,n222);
and (n219,n220,n221);
xor (n220,n184,n185);
and (n221,n189,n211);
and (n222,n223,n224);
xor (n223,n220,n221);
or (n224,n225,n228);
and (n225,n226,n227);
xor (n226,n191,n192);
and (n227,n196,n211);
and (n228,n229,n230);
xor (n229,n226,n227);
or (n230,n231,n234);
and (n231,n232,n233);
xor (n232,n198,n199);
and (n233,n203,n211);
and (n234,n235,n236);
xor (n235,n232,n233);
and (n236,n237,n238);
xor (n237,n205,n206);
and (n238,n209,n211);
and (n239,n182,n240);
or (n241,n242,n245);
and (n242,n243,n244);
xor (n243,n217,n218);
and (n244,n189,n240);
and (n245,n246,n247);
xor (n246,n243,n244);
or (n247,n248,n251);
and (n248,n249,n250);
xor (n249,n223,n224);
and (n250,n196,n240);
and (n251,n252,n253);
xor (n252,n249,n250);
or (n253,n254,n257);
and (n254,n255,n256);
xor (n255,n229,n230);
and (n256,n203,n240);
and (n257,n258,n259);
xor (n258,n255,n256);
and (n259,n260,n261);
xor (n260,n235,n236);
and (n261,n209,n240);
and (n262,n189,n263);
or (n264,n265,n268);
and (n265,n266,n267);
xor (n266,n246,n247);
and (n267,n196,n263);
and (n268,n269,n270);
xor (n269,n266,n267);
or (n270,n271,n274);
and (n271,n272,n273);
xor (n272,n252,n253);
and (n273,n203,n263);
and (n274,n275,n276);
xor (n275,n272,n273);
and (n276,n277,n278);
xor (n277,n258,n259);
and (n278,n209,n263);
and (n279,n196,n280);
or (n281,n282,n285);
and (n282,n283,n284);
xor (n283,n269,n270);
and (n284,n203,n280);
and (n285,n286,n287);
xor (n286,n283,n284);
and (n287,n288,n289);
xor (n288,n275,n276);
and (n289,n209,n280);
and (n290,n203,n291);
and (n292,n293,n294);
xor (n293,n286,n287);
and (n294,n209,n291);
and (n295,n209,n296);
or (n297,n298,n302,n342);
and (n298,n299,n300);
xor (n299,n147,n148);
not (n300,n301);
xor (n301,n293,n294);
and (n302,n300,n303);
or (n303,n304,n308,n341);
and (n304,n305,n306);
xor (n305,n142,n143);
not (n306,n307);
xor (n307,n288,n289);
and (n308,n306,n309);
or (n309,n310,n314,n340);
and (n310,n311,n312);
xor (n311,n131,n132);
not (n312,n313);
xor (n313,n277,n278);
and (n314,n312,n315);
or (n315,n316,n320,n339);
and (n316,n317,n318);
xor (n317,n114,n115);
not (n318,n319);
xor (n319,n260,n261);
and (n320,n318,n321);
or (n321,n322,n326,n338);
and (n322,n323,n324);
xor (n323,n91,n92);
not (n324,n325);
xor (n325,n237,n238);
and (n326,n324,n327);
or (n327,n328,n332,n337);
and (n328,n329,n330);
xor (n329,n61,n62);
not (n330,n331);
xor (n331,n207,n208);
and (n332,n330,n333);
or (n333,n334,n335);
and (n334,n63,n21);
not (n335,n336);
and (n336,n209,n167);
and (n337,n329,n333);
and (n338,n323,n327);
and (n339,n317,n321);
and (n340,n311,n315);
and (n341,n305,n309);
and (n342,n299,n303);
not (n343,n344);
or (n345,n346,n351,n401);
and (n346,n347,n349);
xor (n347,n348,n303);
xor (n348,n299,n300);
not (n349,n350);
and (n351,n349,n352);
or (n352,n353,n358,n400);
and (n353,n354,n356);
xor (n354,n355,n309);
xor (n355,n305,n306);
not (n356,n357);
and (n358,n356,n359);
or (n359,n360,n365,n399);
and (n360,n361,n363);
xor (n361,n362,n315);
xor (n362,n311,n312);
not (n363,n364);
and (n365,n363,n366);
or (n366,n367,n372,n398);
and (n367,n368,n370);
xor (n368,n369,n321);
xor (n369,n317,n318);
not (n370,n371);
and (n372,n370,n373);
or (n373,n374,n379,n397);
and (n374,n375,n377);
xor (n375,n376,n327);
xor (n376,n323,n324);
not (n377,n378);
and (n379,n377,n380);
or (n380,n381,n386,n396);
and (n381,n382,n384);
xor (n382,n383,n333);
xor (n383,n329,n330);
not (n384,n385);
and (n386,n387,n384);
or (n387,n388,n395);
and (n388,n389,n394);
xor (n389,n390,n392);
not (n390,n391);
not (n392,n393);
xor (n394,n334,n336);
and (n395,n392,n390);
and (n396,n382,n387);
and (n397,n375,n380);
and (n398,n368,n373);
and (n399,n361,n366);
and (n400,n354,n359);
and (n401,n347,n352);
not (n402,n403);
and (n403,n404,n420);
not (n404,n405);
or (n405,n406,n417);
or (n406,n407,n414);
or (n407,n408,n411);
xor (n408,n409,n410);
xor (n411,n412,n413);
xor (n414,n415,n416);
xor (n417,n418,n419);
xor (n420,n421,n422);
not (n423,n424);
nor (n424,n425,n963);
and (n425,n426,n402);
nand (n426,n427,n962);
or (n427,n428,n830);
not (n428,n429);
or (n429,n430,n829);
and (n430,n431,n352);
xor (n431,n349,n432);
nand (n432,n433,n828);
or (n433,n434,n743);
not (n434,n435);
nand (n435,n436,n742);
or (n436,n437,n649);
not (n437,n438);
nand (n438,n439,n648);
or (n439,n440,n608);
not (n440,n441);
nand (n441,n442,n569);
not (n442,n443);
xor (n443,n444,n536);
xor (n444,n445,n504);
or (n445,n446,n503);
and (n446,n447,n483);
xor (n447,n448,n468);
nand (n448,n449,n461);
or (n449,n450,n455);
not (n450,n451);
nand (n451,n452,n454);
or (n452,n63,n453);
not (n453,n94);
nand (n454,n453,n63);
not (n455,n456);
nand (n456,n457,n458);
nand (n457,n65,n24,n453);
nand (n458,n459,n460,n94);
not (n459,n65);
not (n460,n24);
nand (n461,n462,n465);
nand (n462,n463,n464);
or (n463,n57,n453);
nand (n464,n453,n57);
nand (n465,n466,n467);
or (n466,n459,n24);
nand (n467,n459,n24);
nand (n468,n469,n478);
or (n469,n470,n476);
not (n470,n471);
nand (n471,n472,n473);
not (n472,n195);
nand (n473,n474,n475);
not (n474,n169);
not (n475,n196);
nand (n476,n477,n169);
not (n477,n167);
nand (n478,n479,n167);
nand (n479,n480,n481);
not (n480,n188);
nand (n481,n474,n482);
not (n482,n189);
nand (n483,n484,n499);
or (n484,n485,n496);
nand (n485,n486,n493);
or (n486,n487,n490);
not (n487,n488);
nand (n488,n489,n211);
not (n489,n240);
not (n490,n491);
nand (n491,n240,n492);
not (n492,n211);
nor (n493,n494,n495);
and (n494,n474,n211);
and (n495,n169,n492);
nor (n496,n497,n261);
and (n497,n489,n498);
not (n498,n209);
or (n499,n493,n500);
nor (n500,n501,n256);
and (n501,n502,n489);
not (n502,n203);
and (n503,n448,n468);
xor (n504,n505,n522);
xor (n505,n506,n513);
nand (n506,n507,n509);
or (n507,n508,n455);
not (n508,n462);
nand (n509,n510,n465);
nand (n510,n511,n512);
or (n511,n50,n453);
nand (n512,n453,n50);
nand (n513,n514,n520);
or (n514,n477,n515);
not (n515,n516);
nand (n516,n517,n518);
not (n517,n181);
nand (n518,n474,n519);
not (n519,n182);
nand (n520,n479,n521);
not (n521,n476);
nand (n522,n523,n535);
or (n523,n524,n530);
not (n524,n525);
nand (n525,n63,n526);
nand (n526,n527,n529);
or (n527,n528,n94);
not (n528,n117);
nand (n529,n528,n94);
not (n530,n531);
and (n531,n532,n209);
nand (n532,n533,n534);
or (n533,n263,n489);
nand (n534,n489,n263);
or (n535,n531,n525);
xor (n536,n537,n557);
xor (n537,n538,n545);
nand (n538,n539,n540);
or (n539,n500,n485);
nand (n540,n541,n544);
nor (n541,n542,n543);
and (n542,n196,n489);
and (n543,n475,n240);
not (n544,n493);
nand (n545,n546,n553);
or (n546,n547,n549);
nand (n547,n548,n24);
not (n548,n21);
not (n549,n550);
nor (n550,n42,n551);
and (n551,n552,n460);
not (n552,n43);
nand (n553,n554,n21);
nor (n554,n35,n555);
and (n555,n556,n460);
not (n556,n36);
and (n557,n558,n564);
nor (n558,n559,n453);
and (n559,n560,n562);
nand (n560,n561,n460);
not (n561,n92);
nand (n562,n459,n563);
not (n563,n63);
nor (n564,n565,n240);
and (n565,n566,n568);
nand (n566,n567,n169);
or (n567,n498,n211);
nand (n568,n498,n211);
not (n569,n570);
or (n570,n571,n607);
and (n571,n572,n585);
xor (n572,n573,n580);
nand (n573,n574,n575);
or (n574,n548,n549);
or (n575,n547,n576);
not (n576,n577);
nor (n577,n49,n578);
and (n578,n579,n460);
not (n579,n50);
xor (n580,n581,n582);
xor (n581,n558,n564);
nor (n582,n583,n584);
nand (n583,n544,n209);
nand (n584,n465,n63);
or (n585,n586,n606);
and (n586,n587,n599);
xor (n587,n588,n595);
nand (n588,n589,n594);
or (n589,n547,n590);
not (n590,n591);
nor (n591,n592,n56);
and (n592,n593,n460);
not (n593,n57);
nand (n594,n577,n21);
nand (n595,n596,n598);
or (n596,n584,n597);
not (n597,n583);
nand (n598,n597,n584);
nand (n599,n600,n605);
or (n600,n476,n601);
not (n601,n602);
nor (n602,n603,n604);
and (n603,n502,n169);
and (n604,n203,n474);
nand (n605,n471,n167);
and (n606,n588,n595);
and (n607,n573,n580);
not (n608,n609);
nand (n609,n610,n647);
or (n610,n611,n614);
nor (n611,n612,n613);
xor (n612,n572,n585);
xor (n613,n447,n483);
nor (n614,n615,n645);
and (n615,n616,n632);
nand (n616,n617,n619);
not (n617,n618);
xor (n618,n587,n599);
not (n619,n620);
or (n620,n621,n631);
and (n621,n622,n625);
xor (n622,n623,n624);
nor (n623,n334,n460);
and (n624,n474,n498,n167);
nand (n625,n626,n627);
or (n626,n477,n601);
nand (n627,n628,n521);
nor (n628,n629,n630);
and (n629,n498,n169);
and (n630,n209,n474);
and (n631,n623,n624);
or (n632,n633,n644);
and (n633,n634,n643);
xor (n634,n635,n636);
and (n635,n334,n336);
nand (n636,n637,n638);
or (n637,n548,n590);
nand (n638,n639,n642);
nand (n639,n640,n641);
or (n640,n460,n63);
or (n641,n563,n24);
not (n642,n547);
xor (n643,n622,n625);
and (n644,n635,n636);
not (n645,n646);
nand (n646,n618,n620);
nand (n647,n612,n613);
nand (n648,n443,n570);
not (n649,n650);
nand (n650,n651,n738);
not (n651,n652);
xor (n652,n653,n697);
xor (n653,n654,n694);
xor (n654,n655,n677);
xor (n655,n656,n670);
nand (n656,n657,n667);
or (n657,n658,n662);
not (n658,n659);
nor (n659,n660,n143);
and (n660,n661,n563);
not (n661,n134);
nand (n662,n663,n664);
not (n663,n526);
nand (n664,n665,n666);
or (n665,n117,n661);
nand (n666,n661,n117);
nand (n667,n668,n526);
nor (n668,n669,n138);
and (n669,n593,n661);
nand (n670,n671,n673);
or (n671,n672,n485);
not (n672,n541);
nand (n673,n544,n674);
nand (n674,n675,n676);
or (n675,n189,n240);
not (n676,n244);
nand (n677,n678,n689);
or (n678,n679,n683);
not (n679,n680);
nand (n680,n681,n682);
or (n681,n209,n280);
not (n682,n289);
nand (n683,n684,n685);
not (n684,n532);
nand (n685,n686,n688);
or (n686,n687,n280);
not (n687,n263);
nand (n688,n280,n687);
nand (n689,n532,n690);
nor (n690,n691,n692);
and (n691,n502,n280);
and (n692,n203,n693);
not (n693,n280);
or (n694,n695,n696);
and (n695,n537,n557);
and (n696,n538,n545);
xor (n697,n698,n721);
xor (n698,n699,n702);
or (n699,n700,n701);
and (n700,n505,n522);
and (n701,n506,n513);
xor (n702,n703,n714);
xor (n703,n704,n709);
nor (n704,n705,n661);
and (n705,n706,n708);
nand (n706,n707,n453);
not (n707,n132);
nand (n708,n563,n528);
nor (n709,n710,n280);
nor (n710,n711,n713);
and (n711,n712,n240);
nand (n712,n209,n687);
and (n713,n498,n263);
nand (n714,n715,n720);
or (n715,n548,n716);
not (n716,n717);
nor (n717,n28,n718);
and (n718,n719,n460);
not (n719,n29);
nand (n720,n554,n642);
xor (n721,n722,n730);
xor (n722,n723,n729);
nand (n723,n724,n726);
or (n724,n725,n455);
not (n725,n510);
nand (n726,n727,n465);
nor (n727,n728,n98);
and (n728,n552,n453);
nor (n729,n530,n525);
nand (n730,n731,n732);
or (n731,n476,n515);
nand (n732,n733,n167);
not (n733,n734);
or (n734,n735,n736);
and (n735,n175,n474);
and (n736,n737,n169);
not (n737,n175);
not (n738,n739);
or (n739,n740,n741);
and (n740,n444,n536);
and (n741,n445,n504);
nand (n742,n652,n739);
not (n743,n744);
nand (n744,n745,n827);
nand (n745,n746,n823);
not (n746,n747);
xor (n747,n748,n767);
xor (n748,n749,n764);
xor (n749,n750,n761);
xor (n750,n751,n758);
nand (n751,n752,n754);
or (n752,n753,n683);
not (n753,n690);
nand (n754,n532,n755);
nor (n755,n756,n757);
and (n756,n475,n280);
and (n757,n196,n693);
or (n758,n759,n760);
and (n759,n722,n730);
and (n760,n723,n729);
or (n761,n762,n763);
and (n762,n703,n714);
and (n763,n704,n709);
or (n764,n765,n766);
and (n765,n698,n721);
and (n766,n699,n702);
xor (n767,n768,n794);
xor (n768,n769,n772);
or (n769,n770,n771);
and (n770,n655,n677);
and (n771,n656,n670);
xor (n772,n773,n787);
xor (n773,n774,n780);
nand (n774,n775,n776);
or (n775,n734,n476);
or (n776,n777,n477);
nor (n777,n778,n168);
and (n778,n474,n779);
not (n779,n170);
nand (n780,n781,n783);
or (n781,n782,n662);
not (n782,n668);
nand (n783,n784,n526);
nand (n784,n785,n786);
or (n785,n50,n661);
nand (n786,n50,n661);
nand (n787,n788,n790);
or (n788,n789,n485);
not (n789,n674);
nand (n790,n544,n791);
nor (n791,n792,n793);
and (n792,n519,n240);
and (n793,n182,n489);
xor (n794,n795,n814);
xor (n795,n796,n802);
nand (n796,n797,n798);
or (n797,n716,n547);
nand (n798,n799,n21);
nand (n799,n800,n801);
or (n800,n23,n460);
nand (n801,n460,n23);
nand (n802,n803,n813);
or (n803,n804,n809);
not (n804,n805);
nand (n805,n806,n63);
nand (n806,n807,n808);
or (n807,n661,n145);
nand (n808,n661,n145);
nand (n809,n810,n209);
nand (n810,n811,n812);
or (n811,n693,n291);
nand (n812,n693,n291);
nand (n813,n804,n809);
nand (n814,n815,n817);
or (n815,n816,n455);
not (n816,n727);
or (n817,n818,n819);
not (n818,n465);
not (n819,n820);
nand (n820,n821,n822);
or (n821,n556,n94);
nand (n822,n94,n556);
not (n823,n824);
or (n824,n825,n826);
and (n825,n653,n697);
and (n826,n654,n694);
nand (n827,n747,n824);
or (n828,n435,n744);
and (n829,n349,n432);
not (n830,n831);
nand (n831,n832,n961);
nand (n832,n833,n344);
not (n833,n834);
xnor (n834,n835,n838);
nand (n835,n836,n827);
or (n836,n837,n434);
not (n837,n745);
nand (n838,n839,n960);
nand (n839,n840,n956);
not (n840,n841);
xor (n841,n842,n914);
xor (n842,n843,n846);
or (n843,n844,n845);
and (n844,n768,n794);
and (n845,n769,n772);
xor (n846,n847,n880);
xor (n847,n848,n877);
xor (n848,n849,n863);
xor (n849,n850,n857);
nor (n850,n851,n856);
and (n851,n852,n854);
nand (n852,n853,n661);
not (n853,n148);
nand (n854,n563,n855);
not (n855,n145);
not (n856,n150);
nor (n857,n858,n296);
nor (n858,n859,n862);
and (n859,n860,n280);
nand (n860,n209,n861);
not (n861,n291);
nor (n862,n209,n861);
nand (n863,n864,n873);
or (n864,n865,n868);
not (n865,n866);
nor (n866,n867,n149);
and (n867,n856,n563);
nand (n868,n869,n872);
nand (n869,n870,n871);
or (n870,n145,n856);
nand (n871,n856,n145);
not (n872,n806);
nand (n873,n874,n806);
nand (n874,n875,n876);
or (n875,n57,n856);
nand (n876,n856,n57);
or (n877,n878,n879);
and (n878,n773,n787);
and (n879,n774,n780);
xor (n880,n881,n906);
xor (n881,n882,n889);
nand (n882,n883,n885);
or (n883,n884,n683);
not (n884,n755);
nand (n885,n532,n886);
nor (n886,n887,n888);
and (n887,n482,n280);
and (n888,n189,n693);
nand (n889,n890,n897);
or (n890,n891,n892);
not (n891,n810);
not (n892,n893);
nor (n893,n894,n895);
and (n894,n502,n296);
and (n895,n203,n896);
not (n896,n296);
nand (n897,n898,n901);
not (n898,n899);
nor (n899,n900,n295);
and (n900,n498,n896);
not (n901,n902);
nand (n902,n891,n903);
nand (n903,n904,n905);
or (n904,n291,n896);
nand (n905,n896,n291);
nand (n906,n907,n909);
or (n907,n547,n908);
not (n908,n799);
or (n909,n910,n548);
nor (n910,n911,n912);
and (n911,n20,n460);
and (n912,n913,n24);
not (n913,n20);
xor (n914,n915,n935);
xor (n915,n916,n932);
xor (n916,n917,n925);
xor (n917,n918,n924);
nand (n918,n919,n920);
or (n919,n819,n455);
nand (n920,n921,n465);
nor (n921,n922,n923);
and (n922,n719,n453);
and (n923,n29,n94);
nor (n924,n805,n809);
nand (n925,n926,n928);
or (n926,n927,n662);
not (n927,n784);
nand (n928,n526,n929);
nand (n929,n930,n931);
or (n930,n43,n661);
nand (n931,n661,n43);
or (n932,n933,n934);
and (n933,n750,n761);
and (n934,n751,n758);
xor (n935,n936,n953);
xor (n936,n937,n946);
nand (n937,n938,n939);
or (n938,n777,n476);
or (n939,n940,n477);
not (n940,n941);
nand (n941,n942,n944);
not (n942,n943);
and (n943,n166,n169);
nand (n944,n945,n474);
not (n945,n166);
nand (n946,n947,n949);
or (n947,n948,n485);
not (n948,n791);
nand (n949,n544,n950);
nor (n950,n951,n952);
and (n951,n737,n240);
and (n952,n175,n489);
or (n953,n954,n955);
and (n954,n795,n814);
and (n955,n796,n802);
not (n956,n957);
or (n957,n958,n959);
and (n958,n748,n767);
and (n959,n749,n764);
nand (n960,n841,n957);
nand (n961,n343,n834);
or (n962,n831,n429);
and (n963,n1,n403);
endmodule
