module top (out,n17,n18,n19,n21,n22,n27,n28,n34,n42
        ,n55,n56,n61,n62,n67,n83,n98,n137,n138,n144
        ,n145,n161,n186,n227,n232,n233,n282,n294,n352,n391
        ,n497,n503,n512,n522,n528);
output out;
input n17;
input n18;
input n19;
input n21;
input n22;
input n27;
input n28;
input n34;
input n42;
input n55;
input n56;
input n61;
input n62;
input n67;
input n83;
input n98;
input n137;
input n138;
input n144;
input n145;
input n161;
input n186;
input n227;
input n232;
input n233;
input n282;
input n294;
input n352;
input n391;
input n497;
input n503;
input n512;
input n522;
input n528;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n20;
wire n23;
wire n24;
wire n25;
wire n26;
wire n29;
wire n30;
wire n31;
wire n32;
wire n33;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n57;
wire n58;
wire n59;
wire n60;
wire n63;
wire n64;
wire n65;
wire n66;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n79;
wire n80;
wire n81;
wire n82;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n228;
wire n229;
wire n230;
wire n231;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
xor (out,n0,n996);
nand (n0,n1,n995);
or (n1,n2,n120);
nand (n2,n3,n119);
or (n3,n4,n102);
or (n4,n5,n101);
and (n5,n6,n85);
xor (n6,n7,n44);
not (n7,n8);
nor (n8,n9,n37);
and (n9,n10,n30);
not (n10,n11);
nand (n11,n12,n24);
not (n12,n13);
nand (n13,n14,n23);
or (n14,n15,n20);
not (n15,n16);
wire s0n16,s1n16,notn16;
or (n16,s0n16,s1n16);
not(notn16,n19);
and (s0n16,notn16,n17);
and (s1n16,n19,n18);
wire s0n20,s1n20,notn20;
or (n20,s0n20,s1n20);
not(notn20,n19);
and (s0n20,notn20,n21);
and (s1n20,n19,n22);
nand (n23,n20,n15);
nand (n24,n25,n29);
or (n25,n15,n26);
wire s0n26,s1n26,notn26;
or (n26,s0n26,s1n26);
not(notn26,n19);
and (s0n26,notn26,n27);
and (s1n26,n19,n28);
nand (n29,n26,n15);
not (n30,n31);
nor (n31,n32,n35);
and (n32,n33,n34);
not (n33,n26);
and (n35,n26,n36);
not (n36,n34);
and (n37,n13,n38);
nand (n38,n39,n43);
or (n39,n26,n40);
not (n40,n41);
and (n41,n42,n34);
or (n43,n33,n41);
xor (n44,n45,n74);
xor (n45,n46,n48);
nand (n46,n47,n38);
or (n47,n10,n13);
nand (n48,n49,n70);
or (n49,n50,n64);
nand (n50,n51,n58);
nor (n51,n52,n57);
and (n52,n53,n26);
not (n53,n54);
wire s0n54,s1n54,notn54;
or (n54,s0n54,s1n54);
not(notn54,n19);
and (s0n54,notn54,n55);
and (s1n54,n19,n56);
and (n57,n54,n33);
nand (n58,n59,n63);
or (n59,n53,n60);
wire s0n60,s1n60,notn60;
or (n60,s0n60,s1n60);
not(notn60,n19);
and (s0n60,notn60,n61);
and (s1n60,n19,n62);
nand (n63,n60,n53);
nor (n64,n65,n68);
and (n65,n66,n67);
not (n66,n60);
and (n68,n60,n69);
not (n69,n67);
or (n70,n51,n71);
nor (n71,n72,n73);
and (n72,n66,n34);
and (n73,n60,n36);
nor (n74,n75,n80);
nand (n75,n60,n76);
not (n76,n77);
wire s0n77,s1n77,notn77;
or (n77,s0n77,s1n77);
not(notn77,n19);
and (s0n77,notn77,1'b0);
and (s1n77,n19,n79);
and (n79,n42,n62);
nor (n80,n81,n84);
and (n81,n77,n82);
not (n82,n83);
and (n84,n76,n83);
or (n85,n86,n100);
and (n86,n87,n8);
xor (n87,n88,n94);
nand (n88,n89,n93);
or (n89,n50,n90);
nor (n90,n91,n92);
and (n91,n66,n83);
and (n92,n60,n82);
or (n93,n51,n64);
nor (n94,n75,n95);
nor (n95,n96,n99);
and (n96,n77,n97);
not (n97,n98);
and (n99,n76,n98);
and (n100,n88,n94);
and (n101,n7,n44);
xor (n102,n103,n116);
xor (n103,n104,n111);
nand (n104,n105,n110);
or (n105,n106,n51);
not (n106,n107);
nand (n107,n108,n109);
or (n108,n60,n40);
or (n109,n66,n41);
or (n110,n50,n71);
nand (n111,n112,n113,n115);
or (n112,n77,n67);
not (n113,n114);
and (n114,n67,n77);
not (n115,n75);
or (n116,n117,n118);
and (n117,n45,n74);
and (n118,n46,n48);
nand (n119,n4,n102);
nand (n120,n121,n989);
or (n121,n122,n265);
not (n122,n123);
nor (n123,n124,n258);
nor (n124,n125,n249);
or (n125,n126,n248);
and (n126,n127,n201);
xor (n127,n128,n163);
xor (n128,n129,n157);
xor (n129,n130,n151);
nand (n130,n131,n147);
or (n131,n132,n141);
and (n132,n133,n140);
nand (n133,n134,n139);
or (n134,n135,n20);
not (n135,n136);
wire s0n136,s1n136,notn136;
or (n136,s0n136,s1n136);
not(notn136,n19);
and (s0n136,notn136,n137);
and (s1n136,n19,n138);
nand (n139,n20,n135);
not (n140,n141);
nand (n141,n142,n146);
or (n142,n135,n143);
wire s0n143,s1n143,notn143;
or (n143,s0n143,s1n143);
not(notn143,n19);
and (s0n143,notn143,n144);
and (s1n143,n19,n145);
nand (n146,n143,n135);
nand (n147,n148,n149);
or (n148,n20,n40);
or (n149,n150,n41);
not (n150,n20);
nand (n151,n152,n156);
or (n152,n11,n153);
nor (n153,n154,n155);
and (n154,n33,n67);
and (n155,n26,n69);
or (n156,n12,n31);
nor (n157,n75,n158);
nor (n158,n159,n162);
and (n159,n77,n160);
not (n160,n161);
and (n162,n76,n161);
xor (n163,n164,n179);
xor (n164,n165,n171);
nand (n165,n166,n170);
or (n166,n50,n167);
nor (n167,n168,n169);
and (n168,n66,n98);
and (n169,n60,n97);
or (n170,n51,n90);
nand (n171,n172,n174);
or (n172,n173,n140);
not (n173,n147);
nand (n174,n175,n132);
not (n175,n176);
nor (n176,n177,n178);
and (n177,n150,n34);
and (n178,n20,n36);
or (n179,n180,n200);
and (n180,n181,n194);
xor (n181,n182,n188);
nor (n182,n75,n183);
nor (n183,n184,n187);
and (n184,n77,n185);
not (n185,n186);
and (n187,n76,n186);
nand (n188,n189,n193);
or (n189,n11,n190);
nor (n190,n191,n192);
and (n191,n83,n33);
and (n192,n82,n26);
or (n193,n12,n153);
nand (n194,n195,n199);
or (n195,n50,n196);
nor (n196,n197,n198);
and (n197,n66,n161);
and (n198,n60,n160);
or (n199,n51,n167);
and (n200,n182,n188);
or (n201,n202,n247);
and (n202,n203,n220);
xor (n203,n204,n205);
not (n204,n171);
or (n205,n206,n212);
nand (n206,n207,n211);
or (n207,n50,n208);
nor (n208,n209,n210);
and (n209,n66,n186);
and (n210,n60,n185);
or (n211,n51,n196);
nand (n212,n213,n219);
or (n213,n214,n215);
not (n214,n132);
not (n215,n216);
nand (n216,n217,n218);
or (n217,n20,n69);
or (n218,n150,n67);
or (n219,n140,n176);
or (n220,n221,n246);
and (n221,n222,n240);
xor (n222,n223,n229);
nor (n223,n75,n224);
nor (n224,n225,n228);
and (n225,n77,n226);
not (n226,n227);
and (n228,n76,n227);
nand (n229,n230,n236);
or (n230,n231,n234);
wire s0n231,s1n231,notn231;
or (n231,s0n231,s1n231);
not(notn231,n19);
and (s0n231,notn231,n232);
and (s1n231,n19,n233);
nor (n234,n235,n231);
not (n235,n143);
not (n236,n237);
nor (n237,n238,n239);
and (n238,n235,n41);
and (n239,n143,n40);
nand (n240,n241,n242);
or (n241,n190,n12);
or (n242,n11,n243);
nor (n243,n244,n245);
and (n244,n33,n98);
and (n245,n26,n97);
and (n246,n223,n229);
and (n247,n204,n205);
and (n248,n128,n163);
xor (n249,n250,n255);
xor (n250,n251,n254);
or (n251,n252,n253);
and (n252,n129,n157);
and (n253,n130,n151);
xor (n254,n87,n8);
or (n255,n256,n257);
and (n256,n164,n179);
and (n257,n165,n171);
and (n258,n259,n263);
not (n259,n260);
or (n260,n261,n262);
and (n261,n250,n255);
and (n262,n251,n254);
not (n263,n264);
xor (n264,n6,n85);
not (n265,n266);
nand (n266,n267,n976);
or (n267,n268,n475);
not (n268,n269);
and (n269,n270,n456,n469);
nor (n270,n271,n433);
nor (n271,n272,n402);
or (n272,n273,n401);
and (n273,n274,n361);
xor (n274,n275,n305);
xor (n275,n276,n296);
xor (n276,n277,n290);
nand (n277,n278,n285);
or (n278,n279,n50);
not (n279,n280);
nor (n280,n281,n283);
and (n281,n282,n60);
and (n283,n284,n66);
not (n284,n282);
nand (n285,n286,n287);
not (n286,n51);
nor (n287,n288,n289);
and (n288,n227,n60);
and (n289,n226,n66);
nor (n290,n75,n291);
nor (n291,n292,n295);
and (n292,n77,n293);
not (n293,n294);
and (n295,n76,n294);
nand (n296,n297,n301);
or (n297,n11,n298);
nor (n298,n299,n300);
and (n299,n33,n186);
and (n300,n26,n185);
or (n301,n12,n302);
nor (n302,n303,n304);
and (n303,n33,n161);
and (n304,n26,n160);
xor (n305,n306,n339);
xor (n306,n307,n326);
xor (n307,n308,n319);
nand (n308,n309,n314);
or (n309,n310,n311);
not (n310,n234);
nor (n311,n312,n313);
and (n312,n235,n67);
and (n313,n143,n69);
or (n314,n315,n318);
nor (n315,n316,n317);
and (n316,n235,n34);
and (n317,n143,n36);
not (n318,n231);
nand (n319,n320,n324);
or (n320,n214,n321);
nor (n321,n322,n323);
and (n322,n150,n98);
and (n323,n20,n97);
or (n324,n325,n140);
xor (n325,n83,n150);
and (n326,n327,n333);
nand (n327,n328,n332);
or (n328,n310,n329);
nor (n329,n330,n331);
and (n330,n235,n83);
and (n331,n143,n82);
or (n332,n311,n318);
nand (n333,n334,n338);
or (n334,n214,n335);
nor (n335,n336,n337);
and (n336,n150,n161);
and (n337,n20,n160);
or (n338,n140,n321);
or (n339,n340,n360);
and (n340,n341,n354);
xor (n341,n342,n348);
nand (n342,n343,n347);
or (n343,n344,n50);
nor (n344,n345,n346);
and (n345,n294,n66);
and (n346,n293,n60);
nand (n347,n286,n280);
nor (n348,n75,n349);
nor (n349,n350,n353);
and (n350,n77,n351);
not (n351,n352);
and (n353,n76,n352);
nand (n354,n355,n359);
or (n355,n11,n356);
nor (n356,n357,n358);
and (n357,n33,n227);
and (n358,n26,n226);
or (n359,n12,n298);
and (n360,n342,n348);
or (n361,n362,n400);
and (n362,n363,n378);
xor (n363,n364,n365);
xor (n364,n327,n333);
and (n365,n366,n372);
nand (n366,n367,n371);
or (n367,n310,n368);
nor (n368,n369,n370);
and (n369,n235,n98);
and (n370,n143,n97);
or (n371,n329,n318);
nand (n372,n373,n377);
or (n373,n214,n374);
nor (n374,n375,n376);
and (n375,n150,n186);
and (n376,n20,n185);
or (n377,n335,n140);
or (n378,n379,n399);
and (n379,n380,n393);
xor (n380,n381,n387);
nand (n381,n382,n386);
or (n382,n50,n383);
nor (n383,n384,n385);
and (n384,n66,n352);
and (n385,n60,n351);
or (n386,n51,n344);
nor (n387,n75,n388);
nor (n388,n389,n392);
and (n389,n77,n390);
not (n390,n391);
and (n392,n76,n391);
nand (n393,n394,n395);
or (n394,n356,n12);
or (n395,n11,n396);
nor (n396,n397,n398);
and (n397,n33,n282);
and (n398,n26,n284);
and (n399,n381,n387);
and (n400,n364,n365);
and (n401,n275,n305);
xor (n402,n403,n430);
xor (n403,n404,n417);
xor (n404,n405,n414);
xor (n405,n406,n410);
nand (n406,n407,n409);
or (n407,n408,n50);
not (n408,n287);
or (n409,n51,n208);
nor (n410,n75,n411);
nor (n411,n412,n413);
and (n412,n77,n284);
and (n413,n76,n282);
nand (n414,n415,n416);
or (n415,n11,n302);
or (n416,n12,n243);
xor (n417,n418,n427);
xor (n418,n419,n426);
xor (n419,n420,n423);
nand (n420,n421,n422);
or (n421,n310,n315);
or (n422,n237,n318);
nand (n423,n424,n425);
or (n424,n325,n214);
nand (n425,n141,n216);
and (n426,n308,n319);
or (n427,n428,n429);
and (n428,n276,n296);
and (n429,n277,n290);
or (n430,n431,n432);
and (n431,n306,n339);
and (n432,n307,n326);
not (n433,n434);
nand (n434,n435,n452);
not (n435,n436);
xor (n436,n437,n442);
xor (n437,n438,n439);
xor (n438,n222,n240);
or (n439,n440,n441);
and (n440,n418,n427);
and (n441,n419,n426);
xor (n442,n443,n448);
xor (n443,n444,n445);
and (n444,n420,n423);
or (n445,n446,n447);
and (n446,n405,n414);
and (n447,n406,n410);
nand (n448,n449,n205);
or (n449,n450,n451);
not (n450,n212);
not (n451,n206);
not (n452,n453);
or (n453,n454,n455);
and (n454,n403,n430);
and (n455,n404,n417);
nand (n456,n457,n459);
not (n457,n458);
xor (n458,n127,n201);
not (n459,n460);
or (n460,n461,n468);
and (n461,n462,n465);
xor (n462,n463,n464);
xor (n463,n181,n194);
xor (n464,n203,n220);
or (n465,n466,n467);
and (n466,n443,n448);
and (n467,n444,n445);
and (n468,n463,n464);
not (n469,n470);
nor (n470,n471,n472);
xor (n471,n462,n465);
or (n472,n473,n474);
and (n473,n437,n442);
and (n474,n438,n439);
not (n475,n476);
nand (n476,n477,n965,n975);
nand (n477,n478,n886);
nand (n478,n479,n742,n885);
nand (n479,n480,n695);
nand (n480,n481,n694);
or (n481,n482,n649);
nor (n482,n483,n648);
and (n483,n484,n620);
not (n484,n485);
nor (n485,n486,n580);
or (n486,n487,n579);
and (n487,n488,n550);
xor (n488,n489,n532);
or (n489,n490,n531);
and (n490,n491,n518);
xor (n491,n492,n506);
nand (n492,n493,n500);
or (n493,n494,n50);
not (n494,n495);
nand (n495,n496,n498);
or (n496,n66,n497);
or (n498,n60,n499);
not (n499,n497);
or (n500,n51,n501);
nor (n501,n502,n504);
and (n502,n503,n66);
and (n504,n505,n60);
not (n505,n503);
nand (n506,n507,n514);
or (n507,n508,n214);
not (n508,n509);
nand (n509,n510,n513);
or (n510,n20,n511);
not (n511,n512);
or (n513,n150,n512);
nand (n514,n141,n515);
nor (n515,n516,n517);
and (n516,n391,n20);
and (n517,n390,n150);
nand (n518,n519,n525);
or (n519,n11,n520);
nor (n520,n521,n523);
and (n521,n33,n522);
and (n523,n26,n524);
not (n524,n522);
or (n525,n12,n526);
nor (n526,n527,n529);
and (n527,n33,n528);
and (n529,n26,n530);
not (n530,n528);
and (n531,n492,n506);
xor (n532,n533,n544);
xor (n533,n534,n535);
and (n534,n115,n497);
nand (n535,n536,n540);
or (n536,n310,n537);
nor (n537,n538,n539);
and (n538,n293,n143);
and (n539,n294,n235);
or (n540,n541,n318);
nor (n541,n542,n543);
and (n542,n235,n282);
and (n543,n143,n284);
nand (n544,n545,n546);
or (n545,n50,n501);
or (n546,n51,n547);
nor (n547,n548,n549);
and (n548,n522,n66);
and (n549,n524,n60);
xor (n550,n551,n565);
xor (n551,n552,n559);
nand (n552,n553,n555);
or (n553,n214,n554);
not (n554,n515);
or (n555,n140,n556);
nor (n556,n557,n558);
and (n557,n150,n352);
and (n558,n20,n351);
nand (n559,n560,n561);
or (n560,n11,n526);
or (n561,n12,n562);
nor (n562,n563,n564);
and (n563,n33,n512);
and (n564,n26,n511);
and (n565,n566,n571);
nor (n566,n567,n66);
nor (n567,n568,n570);
and (n568,n33,n569);
nand (n569,n54,n497);
and (n570,n53,n499);
nand (n571,n572,n577);
or (n572,n573,n310);
not (n573,n574);
nor (n574,n575,n576);
and (n575,n352,n143);
and (n576,n351,n235);
nand (n577,n578,n231);
not (n578,n537);
and (n579,n489,n532);
xor (n580,n581,n603);
xor (n581,n582,n600);
xor (n582,n583,n594);
xor (n583,n584,n590);
nand (n584,n585,n586);
or (n585,n547,n50);
nand (n586,n587,n286);
nor (n587,n588,n589);
and (n588,n528,n60);
and (n589,n530,n66);
nor (n590,n75,n591);
nor (n591,n592,n593);
and (n592,n77,n505);
and (n593,n76,n503);
nand (n594,n595,n596);
or (n595,n310,n541);
or (n596,n597,n318);
nor (n597,n598,n599);
and (n598,n235,n227);
and (n599,n143,n226);
or (n600,n601,n602);
and (n601,n551,n565);
and (n602,n552,n559);
xor (n603,n604,n617);
xor (n604,n605,n611);
nand (n605,n606,n607);
or (n606,n11,n562);
or (n607,n12,n608);
nor (n608,n609,n610);
and (n609,n33,n391);
and (n610,n26,n390);
nand (n611,n612,n613);
or (n612,n214,n556);
or (n613,n614,n140);
nor (n614,n615,n616);
and (n615,n150,n294);
and (n616,n20,n293);
or (n617,n618,n619);
and (n618,n533,n544);
and (n619,n534,n535);
not (n620,n621);
nand (n621,n622,n623);
xor (n622,n488,n550);
or (n623,n624,n647);
and (n624,n625,n646);
xor (n625,n626,n627);
xor (n626,n566,n571);
or (n627,n628,n645);
and (n628,n629,n638);
xor (n629,n630,n631);
and (n630,n286,n497);
nand (n631,n632,n633);
or (n632,n318,n573);
nand (n633,n634,n234);
not (n634,n635);
nor (n635,n636,n637);
and (n636,n391,n235);
and (n637,n390,n143);
nand (n638,n639,n644);
or (n639,n640,n214);
not (n640,n641);
nor (n641,n642,n643);
and (n642,n528,n20);
and (n643,n150,n530);
nand (n644,n141,n509);
and (n645,n630,n631);
xor (n646,n491,n518);
and (n647,n626,n627);
and (n648,n486,n580);
nor (n649,n650,n691);
xor (n650,n651,n688);
xor (n651,n652,n671);
xor (n652,n653,n665);
xor (n653,n654,n661);
nand (n654,n655,n657);
or (n655,n656,n50);
not (n656,n587);
nand (n657,n286,n658);
nor (n658,n659,n660);
and (n659,n512,n60);
and (n660,n511,n66);
nor (n661,n75,n662);
nor (n662,n663,n664);
and (n663,n77,n524);
and (n664,n76,n522);
nand (n665,n666,n667);
or (n666,n11,n608);
or (n667,n12,n668);
nor (n668,n669,n670);
and (n669,n33,n352);
and (n670,n26,n351);
xor (n671,n672,n685);
xor (n672,n673,n679);
nand (n673,n674,n675);
or (n674,n310,n597);
or (n675,n676,n318);
nor (n676,n677,n678);
and (n677,n235,n186);
and (n678,n143,n185);
nand (n679,n680,n681);
or (n680,n214,n614);
or (n681,n682,n140);
nor (n682,n683,n684);
and (n683,n150,n282);
and (n684,n20,n284);
or (n685,n686,n687);
and (n686,n583,n594);
and (n687,n584,n590);
or (n688,n689,n690);
and (n689,n604,n617);
and (n690,n605,n611);
or (n691,n692,n693);
and (n692,n581,n603);
and (n693,n582,n600);
nand (n694,n650,n691);
nand (n695,n696,n738);
not (n696,n697);
xor (n697,n698,n737);
xor (n698,n699,n718);
xor (n699,n700,n712);
xor (n700,n701,n708);
nand (n701,n702,n704);
or (n702,n703,n50);
not (n703,n658);
nand (n704,n286,n705);
nor (n705,n706,n707);
and (n706,n391,n60);
and (n707,n390,n66);
nor (n708,n75,n709);
nor (n709,n710,n711);
and (n710,n77,n530);
and (n711,n76,n528);
nand (n712,n713,n714);
or (n713,n11,n668);
or (n714,n12,n715);
nor (n715,n716,n717);
and (n716,n33,n294);
and (n717,n26,n293);
xor (n718,n719,n734);
xor (n719,n720,n733);
xor (n720,n721,n727);
nand (n721,n722,n723);
or (n722,n310,n676);
or (n723,n724,n318);
nor (n724,n725,n726);
and (n725,n235,n161);
and (n726,n143,n160);
nand (n727,n728,n729);
or (n728,n214,n682);
or (n729,n140,n730);
nor (n730,n731,n732);
and (n731,n150,n227);
and (n732,n20,n226);
and (n733,n673,n679);
or (n734,n735,n736);
and (n735,n653,n665);
and (n736,n654,n661);
and (n737,n672,n685);
not (n738,n739);
or (n739,n740,n741);
and (n740,n651,n688);
and (n741,n652,n671);
nand (n742,n695,n743,n884);
nor (n743,n744,n881);
nor (n744,n745,n879);
and (n745,n746,n874);
or (n746,n747,n873);
and (n747,n748,n789);
xor (n748,n749,n782);
or (n749,n750,n781);
and (n750,n751,n769);
xor (n751,n752,n759);
nand (n752,n753,n758);
or (n753,n754,n214);
not (n754,n755);
nor (n755,n756,n757);
and (n756,n524,n150);
and (n757,n522,n20);
nand (n758,n141,n641);
nand (n759,n760,n765);
or (n760,n761,n12);
not (n761,n762);
nor (n762,n763,n764);
and (n763,n503,n26);
and (n764,n505,n33);
nand (n765,n10,n766);
nand (n766,n767,n768);
or (n767,n33,n497);
or (n768,n26,n499);
xor (n769,n770,n775);
and (n770,n771,n26);
nand (n771,n772,n774);
or (n772,n20,n773);
and (n773,n497,n16);
or (n774,n16,n497);
nand (n775,n776,n780);
or (n776,n310,n777);
nor (n777,n778,n779);
and (n778,n235,n512);
and (n779,n143,n511);
or (n780,n635,n318);
and (n781,n752,n759);
xor (n782,n783,n788);
xor (n783,n784,n787);
nand (n784,n785,n786);
or (n785,n761,n11);
or (n786,n12,n520);
and (n787,n770,n775);
xor (n788,n629,n638);
or (n789,n790,n872);
and (n790,n791,n812);
xor (n791,n792,n811);
or (n792,n793,n810);
and (n793,n794,n803);
xor (n794,n795,n796);
and (n795,n13,n497);
nand (n796,n797,n802);
or (n797,n798,n214);
not (n798,n799);
nor (n799,n800,n801);
and (n800,n503,n20);
and (n801,n505,n150);
nand (n802,n755,n141);
nand (n803,n804,n809);
or (n804,n310,n805);
not (n805,n806);
nor (n806,n807,n808);
and (n807,n530,n235);
and (n808,n528,n143);
or (n809,n777,n318);
and (n810,n795,n796);
xor (n811,n751,n769);
or (n812,n813,n871);
and (n813,n814,n870);
xor (n814,n815,n829);
nor (n815,n816,n824);
not (n816,n817);
nand (n817,n818,n823);
or (n818,n819,n310);
not (n819,n820);
nand (n820,n821,n822);
or (n821,n524,n143);
nand (n822,n143,n524);
nand (n823,n806,n231);
nand (n824,n825,n20);
nand (n825,n826,n828);
or (n826,n143,n827);
and (n827,n497,n136);
or (n828,n136,n497);
nand (n829,n830,n868);
or (n830,n831,n854);
not (n831,n832);
nand (n832,n833,n853);
or (n833,n834,n843);
nor (n834,n835,n842);
nand (n835,n836,n841);
or (n836,n837,n310);
not (n837,n838);
nand (n838,n839,n840);
or (n839,n505,n143);
nand (n840,n143,n505);
nand (n841,n820,n231);
nor (n842,n140,n499);
nand (n843,n844,n851);
nand (n844,n845,n850);
or (n845,n846,n310);
not (n846,n847);
nand (n847,n848,n849);
or (n848,n235,n497);
or (n849,n143,n499);
nand (n850,n838,n231);
nor (n851,n852,n235);
and (n852,n497,n231);
nand (n853,n835,n842);
not (n854,n855);
nand (n855,n856,n864);
not (n856,n857);
nand (n857,n858,n863);
or (n858,n859,n214);
not (n859,n860);
nand (n860,n861,n862);
or (n861,n150,n497);
or (n862,n20,n499);
nand (n863,n141,n799);
nor (n864,n865,n867);
and (n865,n816,n866);
not (n866,n824);
and (n867,n817,n824);
nand (n868,n869,n857);
not (n869,n864);
xor (n870,n794,n803);
and (n871,n815,n829);
and (n872,n792,n811);
and (n873,n749,n782);
or (n874,n875,n876);
xor (n875,n625,n646);
or (n876,n877,n878);
and (n877,n783,n788);
and (n878,n784,n787);
not (n879,n880);
nand (n880,n875,n876);
nand (n881,n882,n484);
not (n882,n883);
nor (n883,n622,n623);
not (n884,n649);
nand (n885,n697,n739);
nor (n886,n887,n944);
nand (n887,n888,n937);
not (n888,n889);
nor (n889,n890,n928);
xor (n890,n891,n919);
xor (n891,n892,n893);
xor (n892,n380,n393);
xor (n893,n894,n903);
xor (n894,n895,n896);
xor (n895,n366,n372);
and (n896,n897,n900);
nand (n897,n898,n899);
or (n898,n310,n724);
or (n899,n368,n318);
nand (n900,n901,n902);
or (n901,n214,n730);
or (n902,n374,n140);
or (n903,n904,n918);
and (n904,n905,n915);
xor (n905,n906,n911);
nand (n906,n907,n909);
or (n907,n908,n50);
not (n908,n705);
nand (n909,n910,n286);
not (n910,n383);
nor (n911,n75,n912);
nor (n912,n913,n914);
and (n913,n77,n511);
and (n914,n76,n512);
nand (n915,n916,n917);
or (n916,n11,n715);
or (n917,n12,n396);
and (n918,n906,n911);
or (n919,n920,n927);
and (n920,n921,n924);
xor (n921,n922,n923);
xor (n922,n897,n900);
and (n923,n721,n727);
or (n924,n925,n926);
and (n925,n700,n712);
and (n926,n701,n708);
and (n927,n922,n923);
or (n928,n929,n936);
and (n929,n930,n933);
xor (n930,n931,n932);
xor (n931,n905,n915);
xor (n932,n921,n924);
or (n933,n934,n935);
and (n934,n719,n734);
and (n935,n720,n733);
and (n936,n931,n932);
nand (n937,n938,n940);
not (n938,n939);
xor (n939,n930,n933);
not (n940,n941);
or (n941,n942,n943);
and (n942,n698,n737);
and (n943,n699,n718);
nand (n944,n945,n958);
nand (n945,n946,n954);
not (n946,n947);
xor (n947,n948,n951);
xor (n948,n949,n950);
xor (n949,n341,n354);
xor (n950,n363,n378);
or (n951,n952,n953);
and (n952,n894,n903);
and (n953,n895,n896);
not (n954,n955);
or (n955,n956,n957);
and (n956,n891,n919);
and (n957,n892,n893);
nand (n958,n959,n961);
not (n959,n960);
xor (n960,n274,n361);
not (n961,n962);
or (n962,n963,n964);
and (n963,n948,n951);
and (n964,n949,n950);
nand (n965,n966,n958);
nand (n966,n967,n974);
or (n967,n968,n969);
not (n968,n945);
not (n969,n970);
nand (n970,n971,n973);
or (n971,n889,n972);
nand (n972,n939,n941);
nand (n973,n890,n928);
nand (n974,n947,n955);
nand (n975,n962,n960);
not (n976,n977);
nand (n977,n978,n988);
or (n978,n979,n980);
not (n979,n456);
not (n980,n981);
nand (n981,n982,n987);
or (n982,n983,n470);
nor (n983,n984,n986);
and (n984,n985,n434);
and (n985,n272,n402);
nor (n986,n435,n452);
nand (n987,n471,n472);
or (n988,n457,n459);
nor (n989,n990,n994);
and (n990,n991,n993);
not (n991,n992);
nand (n992,n125,n249);
not (n993,n258);
nor (n994,n259,n263);
nand (n995,n120,n2);
xor (n996,n997,n1780);
xor (n997,n998,n2195);
xor (n998,n999,n1775);
xor (n999,n1000,n2188);
xor (n1000,n1001,n1769);
xor (n1001,n1002,n2176);
xor (n1002,n1003,n1763);
xor (n1003,n1004,n2159);
xor (n1004,n1005,n1757);
xor (n1005,n1006,n2137);
xor (n1006,n1007,n1751);
xor (n1007,n1008,n2110);
xor (n1008,n1009,n1745);
xor (n1009,n1010,n2078);
xor (n1010,n1011,n1739);
xor (n1011,n1012,n2041);
xor (n1012,n1013,n1733);
xor (n1013,n1014,n1999);
xor (n1014,n1015,n1727);
xor (n1015,n1016,n1952);
xor (n1016,n1017,n1721);
xor (n1017,n1018,n1900);
xor (n1018,n1019,n1715);
xor (n1019,n1020,n1843);
xor (n1020,n1021,n1709);
xor (n1021,n1022,n1781);
xor (n1022,n1023,n1703);
xor (n1023,n1024,n1700);
xor (n1024,n1025,n114);
xor (n1025,n1026,n1618);
xor (n1026,n1027,n1617);
xor (n1027,n1028,n1524);
xor (n1028,n1029,n1523);
xor (n1029,n1030,n1426);
xor (n1030,n1031,n1425);
xor (n1031,n1032,n1323);
xor (n1032,n1033,n1322);
xor (n1033,n1034,n1045);
xor (n1034,n1035,n1044);
xor (n1035,n1036,n1043);
xor (n1036,n1037,n1042);
xor (n1037,n1038,n1041);
xor (n1038,n1039,n1040);
and (n1039,n41,n231);
and (n1040,n41,n143);
and (n1041,n1039,n1040);
and (n1042,n41,n136);
and (n1043,n1037,n1042);
and (n1044,n41,n20);
or (n1045,n1046,n1047);
and (n1046,n1035,n1044);
and (n1047,n1034,n1048);
or (n1048,n1046,n1049);
and (n1049,n1034,n1050);
or (n1050,n1046,n1051);
and (n1051,n1034,n1052);
or (n1052,n1053,n1237);
and (n1053,n1054,n1236);
xor (n1054,n1036,n1055);
or (n1055,n1056,n1148);
and (n1056,n1057,n1147);
xor (n1057,n1038,n1058);
or (n1058,n1041,n1059);
and (n1059,n1060,n1062);
xor (n1060,n1039,n1061);
and (n1061,n34,n143);
or (n1062,n1063,n1066);
and (n1063,n1064,n1065);
and (n1064,n34,n231);
and (n1065,n67,n143);
and (n1066,n1067,n1068);
xor (n1067,n1064,n1065);
or (n1068,n1069,n1072);
and (n1069,n1070,n1071);
and (n1070,n67,n231);
and (n1071,n83,n143);
and (n1072,n1073,n1074);
xor (n1073,n1070,n1071);
or (n1074,n1075,n1078);
and (n1075,n1076,n1077);
and (n1076,n83,n231);
and (n1077,n98,n143);
and (n1078,n1079,n1080);
xor (n1079,n1076,n1077);
or (n1080,n1081,n1084);
and (n1081,n1082,n1083);
and (n1082,n98,n231);
and (n1083,n161,n143);
and (n1084,n1085,n1086);
xor (n1085,n1082,n1083);
or (n1086,n1087,n1090);
and (n1087,n1088,n1089);
and (n1088,n161,n231);
and (n1089,n186,n143);
and (n1090,n1091,n1092);
xor (n1091,n1088,n1089);
or (n1092,n1093,n1096);
and (n1093,n1094,n1095);
and (n1094,n186,n231);
and (n1095,n227,n143);
and (n1096,n1097,n1098);
xor (n1097,n1094,n1095);
or (n1098,n1099,n1102);
and (n1099,n1100,n1101);
and (n1100,n227,n231);
and (n1101,n282,n143);
and (n1102,n1103,n1104);
xor (n1103,n1100,n1101);
or (n1104,n1105,n1108);
and (n1105,n1106,n1107);
and (n1106,n282,n231);
and (n1107,n294,n143);
and (n1108,n1109,n1110);
xor (n1109,n1106,n1107);
or (n1110,n1111,n1113);
and (n1111,n1112,n575);
and (n1112,n294,n231);
and (n1113,n1114,n1115);
xor (n1114,n1112,n575);
or (n1115,n1116,n1119);
and (n1116,n1117,n1118);
and (n1117,n352,n231);
and (n1118,n391,n143);
and (n1119,n1120,n1121);
xor (n1120,n1117,n1118);
or (n1121,n1122,n1125);
and (n1122,n1123,n1124);
and (n1123,n391,n231);
and (n1124,n512,n143);
and (n1125,n1126,n1127);
xor (n1126,n1123,n1124);
or (n1127,n1128,n1130);
and (n1128,n1129,n808);
and (n1129,n512,n231);
and (n1130,n1131,n1132);
xor (n1131,n1129,n808);
or (n1132,n1133,n1136);
and (n1133,n1134,n1135);
and (n1134,n528,n231);
and (n1135,n522,n143);
and (n1136,n1137,n1138);
xor (n1137,n1134,n1135);
or (n1138,n1139,n1142);
and (n1139,n1140,n1141);
and (n1140,n522,n231);
and (n1141,n503,n143);
and (n1142,n1143,n1144);
xor (n1143,n1140,n1141);
and (n1144,n1145,n1146);
and (n1145,n503,n231);
and (n1146,n497,n143);
and (n1147,n34,n136);
and (n1148,n1149,n1150);
xor (n1149,n1057,n1147);
or (n1150,n1151,n1154);
and (n1151,n1152,n1153);
xor (n1152,n1060,n1062);
and (n1153,n67,n136);
and (n1154,n1155,n1156);
xor (n1155,n1152,n1153);
or (n1156,n1157,n1160);
and (n1157,n1158,n1159);
xor (n1158,n1067,n1068);
and (n1159,n83,n136);
and (n1160,n1161,n1162);
xor (n1161,n1158,n1159);
or (n1162,n1163,n1166);
and (n1163,n1164,n1165);
xor (n1164,n1073,n1074);
and (n1165,n98,n136);
and (n1166,n1167,n1168);
xor (n1167,n1164,n1165);
or (n1168,n1169,n1172);
and (n1169,n1170,n1171);
xor (n1170,n1079,n1080);
and (n1171,n161,n136);
and (n1172,n1173,n1174);
xor (n1173,n1170,n1171);
or (n1174,n1175,n1178);
and (n1175,n1176,n1177);
xor (n1176,n1085,n1086);
and (n1177,n186,n136);
and (n1178,n1179,n1180);
xor (n1179,n1176,n1177);
or (n1180,n1181,n1184);
and (n1181,n1182,n1183);
xor (n1182,n1091,n1092);
and (n1183,n227,n136);
and (n1184,n1185,n1186);
xor (n1185,n1182,n1183);
or (n1186,n1187,n1190);
and (n1187,n1188,n1189);
xor (n1188,n1097,n1098);
and (n1189,n282,n136);
and (n1190,n1191,n1192);
xor (n1191,n1188,n1189);
or (n1192,n1193,n1196);
and (n1193,n1194,n1195);
xor (n1194,n1103,n1104);
and (n1195,n294,n136);
and (n1196,n1197,n1198);
xor (n1197,n1194,n1195);
or (n1198,n1199,n1202);
and (n1199,n1200,n1201);
xor (n1200,n1109,n1110);
and (n1201,n352,n136);
and (n1202,n1203,n1204);
xor (n1203,n1200,n1201);
or (n1204,n1205,n1208);
and (n1205,n1206,n1207);
xor (n1206,n1114,n1115);
and (n1207,n391,n136);
and (n1208,n1209,n1210);
xor (n1209,n1206,n1207);
or (n1210,n1211,n1214);
and (n1211,n1212,n1213);
xor (n1212,n1120,n1121);
and (n1213,n512,n136);
and (n1214,n1215,n1216);
xor (n1215,n1212,n1213);
or (n1216,n1217,n1220);
and (n1217,n1218,n1219);
xor (n1218,n1126,n1127);
and (n1219,n528,n136);
and (n1220,n1221,n1222);
xor (n1221,n1218,n1219);
or (n1222,n1223,n1226);
and (n1223,n1224,n1225);
xor (n1224,n1131,n1132);
and (n1225,n522,n136);
and (n1226,n1227,n1228);
xor (n1227,n1224,n1225);
or (n1228,n1229,n1232);
and (n1229,n1230,n1231);
xor (n1230,n1137,n1138);
and (n1231,n503,n136);
and (n1232,n1233,n1234);
xor (n1233,n1230,n1231);
and (n1234,n1235,n827);
xor (n1235,n1143,n1144);
and (n1236,n34,n20);
and (n1237,n1238,n1239);
xor (n1238,n1054,n1236);
or (n1239,n1240,n1243);
and (n1240,n1241,n1242);
xor (n1241,n1149,n1150);
and (n1242,n67,n20);
and (n1243,n1244,n1245);
xor (n1244,n1241,n1242);
or (n1245,n1246,n1249);
and (n1246,n1247,n1248);
xor (n1247,n1155,n1156);
and (n1248,n83,n20);
and (n1249,n1250,n1251);
xor (n1250,n1247,n1248);
or (n1251,n1252,n1255);
and (n1252,n1253,n1254);
xor (n1253,n1161,n1162);
and (n1254,n98,n20);
and (n1255,n1256,n1257);
xor (n1256,n1253,n1254);
or (n1257,n1258,n1261);
and (n1258,n1259,n1260);
xor (n1259,n1167,n1168);
and (n1260,n161,n20);
and (n1261,n1262,n1263);
xor (n1262,n1259,n1260);
or (n1263,n1264,n1267);
and (n1264,n1265,n1266);
xor (n1265,n1173,n1174);
and (n1266,n186,n20);
and (n1267,n1268,n1269);
xor (n1268,n1265,n1266);
or (n1269,n1270,n1273);
and (n1270,n1271,n1272);
xor (n1271,n1179,n1180);
and (n1272,n227,n20);
and (n1273,n1274,n1275);
xor (n1274,n1271,n1272);
or (n1275,n1276,n1279);
and (n1276,n1277,n1278);
xor (n1277,n1185,n1186);
and (n1278,n282,n20);
and (n1279,n1280,n1281);
xor (n1280,n1277,n1278);
or (n1281,n1282,n1285);
and (n1282,n1283,n1284);
xor (n1283,n1191,n1192);
and (n1284,n294,n20);
and (n1285,n1286,n1287);
xor (n1286,n1283,n1284);
or (n1287,n1288,n1291);
and (n1288,n1289,n1290);
xor (n1289,n1197,n1198);
and (n1290,n352,n20);
and (n1291,n1292,n1293);
xor (n1292,n1289,n1290);
or (n1293,n1294,n1296);
and (n1294,n1295,n516);
xor (n1295,n1203,n1204);
and (n1296,n1297,n1298);
xor (n1297,n1295,n516);
or (n1298,n1299,n1302);
and (n1299,n1300,n1301);
xor (n1300,n1209,n1210);
and (n1301,n512,n20);
and (n1302,n1303,n1304);
xor (n1303,n1300,n1301);
or (n1304,n1305,n1307);
and (n1305,n1306,n642);
xor (n1306,n1215,n1216);
and (n1307,n1308,n1309);
xor (n1308,n1306,n642);
or (n1309,n1310,n1312);
and (n1310,n1311,n757);
xor (n1311,n1221,n1222);
and (n1312,n1313,n1314);
xor (n1313,n1311,n757);
or (n1314,n1315,n1317);
and (n1315,n1316,n800);
xor (n1316,n1227,n1228);
and (n1317,n1318,n1319);
xor (n1318,n1316,n800);
and (n1319,n1320,n1321);
xor (n1320,n1233,n1234);
and (n1321,n497,n20);
and (n1322,n41,n16);
or (n1323,n1324,n1326);
and (n1324,n1325,n1322);
xor (n1325,n1034,n1048);
and (n1326,n1327,n1328);
xor (n1327,n1325,n1322);
or (n1328,n1329,n1331);
and (n1329,n1330,n1322);
xor (n1330,n1034,n1050);
and (n1331,n1332,n1333);
xor (n1332,n1330,n1322);
or (n1333,n1334,n1337);
and (n1334,n1335,n1336);
xor (n1335,n1034,n1052);
and (n1336,n34,n16);
and (n1337,n1338,n1339);
xor (n1338,n1335,n1336);
or (n1339,n1340,n1343);
and (n1340,n1341,n1342);
xor (n1341,n1238,n1239);
and (n1342,n67,n16);
and (n1343,n1344,n1345);
xor (n1344,n1341,n1342);
or (n1345,n1346,n1349);
and (n1346,n1347,n1348);
xor (n1347,n1244,n1245);
and (n1348,n83,n16);
and (n1349,n1350,n1351);
xor (n1350,n1347,n1348);
or (n1351,n1352,n1355);
and (n1352,n1353,n1354);
xor (n1353,n1250,n1251);
and (n1354,n98,n16);
and (n1355,n1356,n1357);
xor (n1356,n1353,n1354);
or (n1357,n1358,n1361);
and (n1358,n1359,n1360);
xor (n1359,n1256,n1257);
and (n1360,n161,n16);
and (n1361,n1362,n1363);
xor (n1362,n1359,n1360);
or (n1363,n1364,n1367);
and (n1364,n1365,n1366);
xor (n1365,n1262,n1263);
and (n1366,n186,n16);
and (n1367,n1368,n1369);
xor (n1368,n1365,n1366);
or (n1369,n1370,n1373);
and (n1370,n1371,n1372);
xor (n1371,n1268,n1269);
and (n1372,n227,n16);
and (n1373,n1374,n1375);
xor (n1374,n1371,n1372);
or (n1375,n1376,n1379);
and (n1376,n1377,n1378);
xor (n1377,n1274,n1275);
and (n1378,n282,n16);
and (n1379,n1380,n1381);
xor (n1380,n1377,n1378);
or (n1381,n1382,n1385);
and (n1382,n1383,n1384);
xor (n1383,n1280,n1281);
and (n1384,n294,n16);
and (n1385,n1386,n1387);
xor (n1386,n1383,n1384);
or (n1387,n1388,n1391);
and (n1388,n1389,n1390);
xor (n1389,n1286,n1287);
and (n1390,n352,n16);
and (n1391,n1392,n1393);
xor (n1392,n1389,n1390);
or (n1393,n1394,n1397);
and (n1394,n1395,n1396);
xor (n1395,n1292,n1293);
and (n1396,n391,n16);
and (n1397,n1398,n1399);
xor (n1398,n1395,n1396);
or (n1399,n1400,n1403);
and (n1400,n1401,n1402);
xor (n1401,n1297,n1298);
and (n1402,n512,n16);
and (n1403,n1404,n1405);
xor (n1404,n1401,n1402);
or (n1405,n1406,n1409);
and (n1406,n1407,n1408);
xor (n1407,n1303,n1304);
and (n1408,n528,n16);
and (n1409,n1410,n1411);
xor (n1410,n1407,n1408);
or (n1411,n1412,n1415);
and (n1412,n1413,n1414);
xor (n1413,n1308,n1309);
and (n1414,n522,n16);
and (n1415,n1416,n1417);
xor (n1416,n1413,n1414);
or (n1417,n1418,n1421);
and (n1418,n1419,n1420);
xor (n1419,n1313,n1314);
and (n1420,n503,n16);
and (n1421,n1422,n1423);
xor (n1422,n1419,n1420);
and (n1423,n1424,n773);
xor (n1424,n1318,n1319);
and (n1425,n41,n26);
or (n1426,n1427,n1429);
and (n1427,n1428,n1425);
xor (n1428,n1327,n1328);
and (n1429,n1430,n1431);
xor (n1430,n1428,n1425);
or (n1431,n1432,n1435);
and (n1432,n1433,n1434);
xor (n1433,n1332,n1333);
and (n1434,n34,n26);
and (n1435,n1436,n1437);
xor (n1436,n1433,n1434);
or (n1437,n1438,n1441);
and (n1438,n1439,n1440);
xor (n1439,n1338,n1339);
and (n1440,n67,n26);
and (n1441,n1442,n1443);
xor (n1442,n1439,n1440);
or (n1443,n1444,n1447);
and (n1444,n1445,n1446);
xor (n1445,n1344,n1345);
and (n1446,n83,n26);
and (n1447,n1448,n1449);
xor (n1448,n1445,n1446);
or (n1449,n1450,n1453);
and (n1450,n1451,n1452);
xor (n1451,n1350,n1351);
and (n1452,n98,n26);
and (n1453,n1454,n1455);
xor (n1454,n1451,n1452);
or (n1455,n1456,n1459);
and (n1456,n1457,n1458);
xor (n1457,n1356,n1357);
and (n1458,n161,n26);
and (n1459,n1460,n1461);
xor (n1460,n1457,n1458);
or (n1461,n1462,n1465);
and (n1462,n1463,n1464);
xor (n1463,n1362,n1363);
and (n1464,n186,n26);
and (n1465,n1466,n1467);
xor (n1466,n1463,n1464);
or (n1467,n1468,n1471);
and (n1468,n1469,n1470);
xor (n1469,n1368,n1369);
and (n1470,n227,n26);
and (n1471,n1472,n1473);
xor (n1472,n1469,n1470);
or (n1473,n1474,n1477);
and (n1474,n1475,n1476);
xor (n1475,n1374,n1375);
and (n1476,n282,n26);
and (n1477,n1478,n1479);
xor (n1478,n1475,n1476);
or (n1479,n1480,n1483);
and (n1480,n1481,n1482);
xor (n1481,n1380,n1381);
and (n1482,n294,n26);
and (n1483,n1484,n1485);
xor (n1484,n1481,n1482);
or (n1485,n1486,n1489);
and (n1486,n1487,n1488);
xor (n1487,n1386,n1387);
and (n1488,n352,n26);
and (n1489,n1490,n1491);
xor (n1490,n1487,n1488);
or (n1491,n1492,n1495);
and (n1492,n1493,n1494);
xor (n1493,n1392,n1393);
and (n1494,n391,n26);
and (n1495,n1496,n1497);
xor (n1496,n1493,n1494);
or (n1497,n1498,n1501);
and (n1498,n1499,n1500);
xor (n1499,n1398,n1399);
and (n1500,n512,n26);
and (n1501,n1502,n1503);
xor (n1502,n1499,n1500);
or (n1503,n1504,n1507);
and (n1504,n1505,n1506);
xor (n1505,n1404,n1405);
and (n1506,n528,n26);
and (n1507,n1508,n1509);
xor (n1508,n1505,n1506);
or (n1509,n1510,n1513);
and (n1510,n1511,n1512);
xor (n1511,n1410,n1411);
and (n1512,n522,n26);
and (n1513,n1514,n1515);
xor (n1514,n1511,n1512);
or (n1515,n1516,n1518);
and (n1516,n1517,n763);
xor (n1517,n1416,n1417);
and (n1518,n1519,n1520);
xor (n1519,n1517,n763);
and (n1520,n1521,n1522);
xor (n1521,n1422,n1423);
and (n1522,n497,n26);
and (n1523,n41,n54);
or (n1524,n1525,n1528);
and (n1525,n1526,n1527);
xor (n1526,n1430,n1431);
and (n1527,n34,n54);
and (n1528,n1529,n1530);
xor (n1529,n1526,n1527);
or (n1530,n1531,n1534);
and (n1531,n1532,n1533);
xor (n1532,n1436,n1437);
and (n1533,n67,n54);
and (n1534,n1535,n1536);
xor (n1535,n1532,n1533);
or (n1536,n1537,n1540);
and (n1537,n1538,n1539);
xor (n1538,n1442,n1443);
and (n1539,n83,n54);
and (n1540,n1541,n1542);
xor (n1541,n1538,n1539);
or (n1542,n1543,n1546);
and (n1543,n1544,n1545);
xor (n1544,n1448,n1449);
and (n1545,n98,n54);
and (n1546,n1547,n1548);
xor (n1547,n1544,n1545);
or (n1548,n1549,n1552);
and (n1549,n1550,n1551);
xor (n1550,n1454,n1455);
and (n1551,n161,n54);
and (n1552,n1553,n1554);
xor (n1553,n1550,n1551);
or (n1554,n1555,n1558);
and (n1555,n1556,n1557);
xor (n1556,n1460,n1461);
and (n1557,n186,n54);
and (n1558,n1559,n1560);
xor (n1559,n1556,n1557);
or (n1560,n1561,n1564);
and (n1561,n1562,n1563);
xor (n1562,n1466,n1467);
and (n1563,n227,n54);
and (n1564,n1565,n1566);
xor (n1565,n1562,n1563);
or (n1566,n1567,n1570);
and (n1567,n1568,n1569);
xor (n1568,n1472,n1473);
and (n1569,n282,n54);
and (n1570,n1571,n1572);
xor (n1571,n1568,n1569);
or (n1572,n1573,n1576);
and (n1573,n1574,n1575);
xor (n1574,n1478,n1479);
and (n1575,n294,n54);
and (n1576,n1577,n1578);
xor (n1577,n1574,n1575);
or (n1578,n1579,n1582);
and (n1579,n1580,n1581);
xor (n1580,n1484,n1485);
and (n1581,n352,n54);
and (n1582,n1583,n1584);
xor (n1583,n1580,n1581);
or (n1584,n1585,n1588);
and (n1585,n1586,n1587);
xor (n1586,n1490,n1491);
and (n1587,n391,n54);
and (n1588,n1589,n1590);
xor (n1589,n1586,n1587);
or (n1590,n1591,n1594);
and (n1591,n1592,n1593);
xor (n1592,n1496,n1497);
and (n1593,n512,n54);
and (n1594,n1595,n1596);
xor (n1595,n1592,n1593);
or (n1596,n1597,n1600);
and (n1597,n1598,n1599);
xor (n1598,n1502,n1503);
and (n1599,n528,n54);
and (n1600,n1601,n1602);
xor (n1601,n1598,n1599);
or (n1602,n1603,n1606);
and (n1603,n1604,n1605);
xor (n1604,n1508,n1509);
and (n1605,n522,n54);
and (n1606,n1607,n1608);
xor (n1607,n1604,n1605);
or (n1608,n1609,n1612);
and (n1609,n1610,n1611);
xor (n1610,n1514,n1515);
and (n1611,n503,n54);
and (n1612,n1613,n1614);
xor (n1613,n1610,n1611);
and (n1614,n1615,n1616);
xor (n1615,n1519,n1520);
not (n1616,n569);
and (n1617,n34,n60);
or (n1618,n1619,n1622);
and (n1619,n1620,n1621);
xor (n1620,n1529,n1530);
and (n1621,n67,n60);
and (n1622,n1623,n1624);
xor (n1623,n1620,n1621);
or (n1624,n1625,n1628);
and (n1625,n1626,n1627);
xor (n1626,n1535,n1536);
and (n1627,n83,n60);
and (n1628,n1629,n1630);
xor (n1629,n1626,n1627);
or (n1630,n1631,n1634);
and (n1631,n1632,n1633);
xor (n1632,n1541,n1542);
and (n1633,n98,n60);
and (n1634,n1635,n1636);
xor (n1635,n1632,n1633);
or (n1636,n1637,n1640);
and (n1637,n1638,n1639);
xor (n1638,n1547,n1548);
and (n1639,n161,n60);
and (n1640,n1641,n1642);
xor (n1641,n1638,n1639);
or (n1642,n1643,n1646);
and (n1643,n1644,n1645);
xor (n1644,n1553,n1554);
and (n1645,n186,n60);
and (n1646,n1647,n1648);
xor (n1647,n1644,n1645);
or (n1648,n1649,n1651);
and (n1649,n1650,n288);
xor (n1650,n1559,n1560);
and (n1651,n1652,n1653);
xor (n1652,n1650,n288);
or (n1653,n1654,n1656);
and (n1654,n1655,n281);
xor (n1655,n1565,n1566);
and (n1656,n1657,n1658);
xor (n1657,n1655,n281);
or (n1658,n1659,n1662);
and (n1659,n1660,n1661);
xor (n1660,n1571,n1572);
and (n1661,n294,n60);
and (n1662,n1663,n1664);
xor (n1663,n1660,n1661);
or (n1664,n1665,n1668);
and (n1665,n1666,n1667);
xor (n1666,n1577,n1578);
and (n1667,n352,n60);
and (n1668,n1669,n1670);
xor (n1669,n1666,n1667);
or (n1670,n1671,n1673);
and (n1671,n1672,n706);
xor (n1672,n1583,n1584);
and (n1673,n1674,n1675);
xor (n1674,n1672,n706);
or (n1675,n1676,n1678);
and (n1676,n1677,n659);
xor (n1677,n1589,n1590);
and (n1678,n1679,n1680);
xor (n1679,n1677,n659);
or (n1680,n1681,n1683);
and (n1681,n1682,n588);
xor (n1682,n1595,n1596);
and (n1683,n1684,n1685);
xor (n1684,n1682,n588);
or (n1685,n1686,n1689);
and (n1686,n1687,n1688);
xor (n1687,n1601,n1602);
and (n1688,n522,n60);
and (n1689,n1690,n1691);
xor (n1690,n1687,n1688);
or (n1691,n1692,n1695);
and (n1692,n1693,n1694);
xor (n1693,n1607,n1608);
and (n1694,n503,n60);
and (n1695,n1696,n1697);
xor (n1696,n1693,n1694);
and (n1697,n1698,n1699);
xor (n1698,n1613,n1614);
and (n1699,n497,n60);
or (n1700,n1701,n1704);
and (n1701,n1702,n1703);
xor (n1702,n1623,n1624);
and (n1703,n83,n77);
and (n1704,n1705,n1706);
xor (n1705,n1702,n1703);
or (n1706,n1707,n1710);
and (n1707,n1708,n1709);
xor (n1708,n1629,n1630);
and (n1709,n98,n77);
and (n1710,n1711,n1712);
xor (n1711,n1708,n1709);
or (n1712,n1713,n1716);
and (n1713,n1714,n1715);
xor (n1714,n1635,n1636);
and (n1715,n161,n77);
and (n1716,n1717,n1718);
xor (n1717,n1714,n1715);
or (n1718,n1719,n1722);
and (n1719,n1720,n1721);
xor (n1720,n1641,n1642);
and (n1721,n186,n77);
and (n1722,n1723,n1724);
xor (n1723,n1720,n1721);
or (n1724,n1725,n1728);
and (n1725,n1726,n1727);
xor (n1726,n1647,n1648);
and (n1727,n227,n77);
and (n1728,n1729,n1730);
xor (n1729,n1726,n1727);
or (n1730,n1731,n1734);
and (n1731,n1732,n1733);
xor (n1732,n1652,n1653);
and (n1733,n282,n77);
and (n1734,n1735,n1736);
xor (n1735,n1732,n1733);
or (n1736,n1737,n1740);
and (n1737,n1738,n1739);
xor (n1738,n1657,n1658);
and (n1739,n294,n77);
and (n1740,n1741,n1742);
xor (n1741,n1738,n1739);
or (n1742,n1743,n1746);
and (n1743,n1744,n1745);
xor (n1744,n1663,n1664);
and (n1745,n352,n77);
and (n1746,n1747,n1748);
xor (n1747,n1744,n1745);
or (n1748,n1749,n1752);
and (n1749,n1750,n1751);
xor (n1750,n1669,n1670);
and (n1751,n391,n77);
and (n1752,n1753,n1754);
xor (n1753,n1750,n1751);
or (n1754,n1755,n1758);
and (n1755,n1756,n1757);
xor (n1756,n1674,n1675);
and (n1757,n512,n77);
and (n1758,n1759,n1760);
xor (n1759,n1756,n1757);
or (n1760,n1761,n1764);
and (n1761,n1762,n1763);
xor (n1762,n1679,n1680);
and (n1763,n528,n77);
and (n1764,n1765,n1766);
xor (n1765,n1762,n1763);
or (n1766,n1767,n1770);
and (n1767,n1768,n1769);
xor (n1768,n1684,n1685);
and (n1769,n522,n77);
and (n1770,n1771,n1772);
xor (n1771,n1768,n1769);
or (n1772,n1773,n1776);
and (n1773,n1774,n1775);
xor (n1774,n1690,n1691);
and (n1775,n503,n77);
and (n1776,n1777,n1778);
xor (n1777,n1774,n1775);
and (n1778,n1779,n1780);
xor (n1779,n1696,n1697);
and (n1780,n497,n77);
or (n1781,n1782,n1784);
and (n1782,n1783,n1709);
xor (n1783,n1705,n1706);
and (n1784,n1785,n1786);
xor (n1785,n1783,n1709);
or (n1786,n1787,n1789);
and (n1787,n1788,n1715);
xor (n1788,n1711,n1712);
and (n1789,n1790,n1791);
xor (n1790,n1788,n1715);
or (n1791,n1792,n1794);
and (n1792,n1793,n1721);
xor (n1793,n1717,n1718);
and (n1794,n1795,n1796);
xor (n1795,n1793,n1721);
or (n1796,n1797,n1799);
and (n1797,n1798,n1727);
xor (n1798,n1723,n1724);
and (n1799,n1800,n1801);
xor (n1800,n1798,n1727);
or (n1801,n1802,n1804);
and (n1802,n1803,n1733);
xor (n1803,n1729,n1730);
and (n1804,n1805,n1806);
xor (n1805,n1803,n1733);
or (n1806,n1807,n1809);
and (n1807,n1808,n1739);
xor (n1808,n1735,n1736);
and (n1809,n1810,n1811);
xor (n1810,n1808,n1739);
or (n1811,n1812,n1814);
and (n1812,n1813,n1745);
xor (n1813,n1741,n1742);
and (n1814,n1815,n1816);
xor (n1815,n1813,n1745);
or (n1816,n1817,n1819);
and (n1817,n1818,n1751);
xor (n1818,n1747,n1748);
and (n1819,n1820,n1821);
xor (n1820,n1818,n1751);
or (n1821,n1822,n1824);
and (n1822,n1823,n1757);
xor (n1823,n1753,n1754);
and (n1824,n1825,n1826);
xor (n1825,n1823,n1757);
or (n1826,n1827,n1829);
and (n1827,n1828,n1763);
xor (n1828,n1759,n1760);
and (n1829,n1830,n1831);
xor (n1830,n1828,n1763);
or (n1831,n1832,n1834);
and (n1832,n1833,n1769);
xor (n1833,n1765,n1766);
and (n1834,n1835,n1836);
xor (n1835,n1833,n1769);
or (n1836,n1837,n1839);
and (n1837,n1838,n1775);
xor (n1838,n1771,n1772);
and (n1839,n1840,n1841);
xor (n1840,n1838,n1775);
and (n1841,n1842,n1780);
xor (n1842,n1777,n1778);
or (n1843,n1844,n1846);
and (n1844,n1845,n1715);
xor (n1845,n1785,n1786);
and (n1846,n1847,n1848);
xor (n1847,n1845,n1715);
or (n1848,n1849,n1851);
and (n1849,n1850,n1721);
xor (n1850,n1790,n1791);
and (n1851,n1852,n1853);
xor (n1852,n1850,n1721);
or (n1853,n1854,n1856);
and (n1854,n1855,n1727);
xor (n1855,n1795,n1796);
and (n1856,n1857,n1858);
xor (n1857,n1855,n1727);
or (n1858,n1859,n1861);
and (n1859,n1860,n1733);
xor (n1860,n1800,n1801);
and (n1861,n1862,n1863);
xor (n1862,n1860,n1733);
or (n1863,n1864,n1866);
and (n1864,n1865,n1739);
xor (n1865,n1805,n1806);
and (n1866,n1867,n1868);
xor (n1867,n1865,n1739);
or (n1868,n1869,n1871);
and (n1869,n1870,n1745);
xor (n1870,n1810,n1811);
and (n1871,n1872,n1873);
xor (n1872,n1870,n1745);
or (n1873,n1874,n1876);
and (n1874,n1875,n1751);
xor (n1875,n1815,n1816);
and (n1876,n1877,n1878);
xor (n1877,n1875,n1751);
or (n1878,n1879,n1881);
and (n1879,n1880,n1757);
xor (n1880,n1820,n1821);
and (n1881,n1882,n1883);
xor (n1882,n1880,n1757);
or (n1883,n1884,n1886);
and (n1884,n1885,n1763);
xor (n1885,n1825,n1826);
and (n1886,n1887,n1888);
xor (n1887,n1885,n1763);
or (n1888,n1889,n1891);
and (n1889,n1890,n1769);
xor (n1890,n1830,n1831);
and (n1891,n1892,n1893);
xor (n1892,n1890,n1769);
or (n1893,n1894,n1896);
and (n1894,n1895,n1775);
xor (n1895,n1835,n1836);
and (n1896,n1897,n1898);
xor (n1897,n1895,n1775);
and (n1898,n1899,n1780);
xor (n1899,n1840,n1841);
or (n1900,n1901,n1903);
and (n1901,n1902,n1721);
xor (n1902,n1847,n1848);
and (n1903,n1904,n1905);
xor (n1904,n1902,n1721);
or (n1905,n1906,n1908);
and (n1906,n1907,n1727);
xor (n1907,n1852,n1853);
and (n1908,n1909,n1910);
xor (n1909,n1907,n1727);
or (n1910,n1911,n1913);
and (n1911,n1912,n1733);
xor (n1912,n1857,n1858);
and (n1913,n1914,n1915);
xor (n1914,n1912,n1733);
or (n1915,n1916,n1918);
and (n1916,n1917,n1739);
xor (n1917,n1862,n1863);
and (n1918,n1919,n1920);
xor (n1919,n1917,n1739);
or (n1920,n1921,n1923);
and (n1921,n1922,n1745);
xor (n1922,n1867,n1868);
and (n1923,n1924,n1925);
xor (n1924,n1922,n1745);
or (n1925,n1926,n1928);
and (n1926,n1927,n1751);
xor (n1927,n1872,n1873);
and (n1928,n1929,n1930);
xor (n1929,n1927,n1751);
or (n1930,n1931,n1933);
and (n1931,n1932,n1757);
xor (n1932,n1877,n1878);
and (n1933,n1934,n1935);
xor (n1934,n1932,n1757);
or (n1935,n1936,n1938);
and (n1936,n1937,n1763);
xor (n1937,n1882,n1883);
and (n1938,n1939,n1940);
xor (n1939,n1937,n1763);
or (n1940,n1941,n1943);
and (n1941,n1942,n1769);
xor (n1942,n1887,n1888);
and (n1943,n1944,n1945);
xor (n1944,n1942,n1769);
or (n1945,n1946,n1948);
and (n1946,n1947,n1775);
xor (n1947,n1892,n1893);
and (n1948,n1949,n1950);
xor (n1949,n1947,n1775);
and (n1950,n1951,n1780);
xor (n1951,n1897,n1898);
or (n1952,n1953,n1955);
and (n1953,n1954,n1727);
xor (n1954,n1904,n1905);
and (n1955,n1956,n1957);
xor (n1956,n1954,n1727);
or (n1957,n1958,n1960);
and (n1958,n1959,n1733);
xor (n1959,n1909,n1910);
and (n1960,n1961,n1962);
xor (n1961,n1959,n1733);
or (n1962,n1963,n1965);
and (n1963,n1964,n1739);
xor (n1964,n1914,n1915);
and (n1965,n1966,n1967);
xor (n1966,n1964,n1739);
or (n1967,n1968,n1970);
and (n1968,n1969,n1745);
xor (n1969,n1919,n1920);
and (n1970,n1971,n1972);
xor (n1971,n1969,n1745);
or (n1972,n1973,n1975);
and (n1973,n1974,n1751);
xor (n1974,n1924,n1925);
and (n1975,n1976,n1977);
xor (n1976,n1974,n1751);
or (n1977,n1978,n1980);
and (n1978,n1979,n1757);
xor (n1979,n1929,n1930);
and (n1980,n1981,n1982);
xor (n1981,n1979,n1757);
or (n1982,n1983,n1985);
and (n1983,n1984,n1763);
xor (n1984,n1934,n1935);
and (n1985,n1986,n1987);
xor (n1986,n1984,n1763);
or (n1987,n1988,n1990);
and (n1988,n1989,n1769);
xor (n1989,n1939,n1940);
and (n1990,n1991,n1992);
xor (n1991,n1989,n1769);
or (n1992,n1993,n1995);
and (n1993,n1994,n1775);
xor (n1994,n1944,n1945);
and (n1995,n1996,n1997);
xor (n1996,n1994,n1775);
and (n1997,n1998,n1780);
xor (n1998,n1949,n1950);
or (n1999,n2000,n2002);
and (n2000,n2001,n1733);
xor (n2001,n1956,n1957);
and (n2002,n2003,n2004);
xor (n2003,n2001,n1733);
or (n2004,n2005,n2007);
and (n2005,n2006,n1739);
xor (n2006,n1961,n1962);
and (n2007,n2008,n2009);
xor (n2008,n2006,n1739);
or (n2009,n2010,n2012);
and (n2010,n2011,n1745);
xor (n2011,n1966,n1967);
and (n2012,n2013,n2014);
xor (n2013,n2011,n1745);
or (n2014,n2015,n2017);
and (n2015,n2016,n1751);
xor (n2016,n1971,n1972);
and (n2017,n2018,n2019);
xor (n2018,n2016,n1751);
or (n2019,n2020,n2022);
and (n2020,n2021,n1757);
xor (n2021,n1976,n1977);
and (n2022,n2023,n2024);
xor (n2023,n2021,n1757);
or (n2024,n2025,n2027);
and (n2025,n2026,n1763);
xor (n2026,n1981,n1982);
and (n2027,n2028,n2029);
xor (n2028,n2026,n1763);
or (n2029,n2030,n2032);
and (n2030,n2031,n1769);
xor (n2031,n1986,n1987);
and (n2032,n2033,n2034);
xor (n2033,n2031,n1769);
or (n2034,n2035,n2037);
and (n2035,n2036,n1775);
xor (n2036,n1991,n1992);
and (n2037,n2038,n2039);
xor (n2038,n2036,n1775);
and (n2039,n2040,n1780);
xor (n2040,n1996,n1997);
or (n2041,n2042,n2044);
and (n2042,n2043,n1739);
xor (n2043,n2003,n2004);
and (n2044,n2045,n2046);
xor (n2045,n2043,n1739);
or (n2046,n2047,n2049);
and (n2047,n2048,n1745);
xor (n2048,n2008,n2009);
and (n2049,n2050,n2051);
xor (n2050,n2048,n1745);
or (n2051,n2052,n2054);
and (n2052,n2053,n1751);
xor (n2053,n2013,n2014);
and (n2054,n2055,n2056);
xor (n2055,n2053,n1751);
or (n2056,n2057,n2059);
and (n2057,n2058,n1757);
xor (n2058,n2018,n2019);
and (n2059,n2060,n2061);
xor (n2060,n2058,n1757);
or (n2061,n2062,n2064);
and (n2062,n2063,n1763);
xor (n2063,n2023,n2024);
and (n2064,n2065,n2066);
xor (n2065,n2063,n1763);
or (n2066,n2067,n2069);
and (n2067,n2068,n1769);
xor (n2068,n2028,n2029);
and (n2069,n2070,n2071);
xor (n2070,n2068,n1769);
or (n2071,n2072,n2074);
and (n2072,n2073,n1775);
xor (n2073,n2033,n2034);
and (n2074,n2075,n2076);
xor (n2075,n2073,n1775);
and (n2076,n2077,n1780);
xor (n2077,n2038,n2039);
or (n2078,n2079,n2081);
and (n2079,n2080,n1745);
xor (n2080,n2045,n2046);
and (n2081,n2082,n2083);
xor (n2082,n2080,n1745);
or (n2083,n2084,n2086);
and (n2084,n2085,n1751);
xor (n2085,n2050,n2051);
and (n2086,n2087,n2088);
xor (n2087,n2085,n1751);
or (n2088,n2089,n2091);
and (n2089,n2090,n1757);
xor (n2090,n2055,n2056);
and (n2091,n2092,n2093);
xor (n2092,n2090,n1757);
or (n2093,n2094,n2096);
and (n2094,n2095,n1763);
xor (n2095,n2060,n2061);
and (n2096,n2097,n2098);
xor (n2097,n2095,n1763);
or (n2098,n2099,n2101);
and (n2099,n2100,n1769);
xor (n2100,n2065,n2066);
and (n2101,n2102,n2103);
xor (n2102,n2100,n1769);
or (n2103,n2104,n2106);
and (n2104,n2105,n1775);
xor (n2105,n2070,n2071);
and (n2106,n2107,n2108);
xor (n2107,n2105,n1775);
and (n2108,n2109,n1780);
xor (n2109,n2075,n2076);
or (n2110,n2111,n2113);
and (n2111,n2112,n1751);
xor (n2112,n2082,n2083);
and (n2113,n2114,n2115);
xor (n2114,n2112,n1751);
or (n2115,n2116,n2118);
and (n2116,n2117,n1757);
xor (n2117,n2087,n2088);
and (n2118,n2119,n2120);
xor (n2119,n2117,n1757);
or (n2120,n2121,n2123);
and (n2121,n2122,n1763);
xor (n2122,n2092,n2093);
and (n2123,n2124,n2125);
xor (n2124,n2122,n1763);
or (n2125,n2126,n2128);
and (n2126,n2127,n1769);
xor (n2127,n2097,n2098);
and (n2128,n2129,n2130);
xor (n2129,n2127,n1769);
or (n2130,n2131,n2133);
and (n2131,n2132,n1775);
xor (n2132,n2102,n2103);
and (n2133,n2134,n2135);
xor (n2134,n2132,n1775);
and (n2135,n2136,n1780);
xor (n2136,n2107,n2108);
or (n2137,n2138,n2140);
and (n2138,n2139,n1757);
xor (n2139,n2114,n2115);
and (n2140,n2141,n2142);
xor (n2141,n2139,n1757);
or (n2142,n2143,n2145);
and (n2143,n2144,n1763);
xor (n2144,n2119,n2120);
and (n2145,n2146,n2147);
xor (n2146,n2144,n1763);
or (n2147,n2148,n2150);
and (n2148,n2149,n1769);
xor (n2149,n2124,n2125);
and (n2150,n2151,n2152);
xor (n2151,n2149,n1769);
or (n2152,n2153,n2155);
and (n2153,n2154,n1775);
xor (n2154,n2129,n2130);
and (n2155,n2156,n2157);
xor (n2156,n2154,n1775);
and (n2157,n2158,n1780);
xor (n2158,n2134,n2135);
or (n2159,n2160,n2162);
and (n2160,n2161,n1763);
xor (n2161,n2141,n2142);
and (n2162,n2163,n2164);
xor (n2163,n2161,n1763);
or (n2164,n2165,n2167);
and (n2165,n2166,n1769);
xor (n2166,n2146,n2147);
and (n2167,n2168,n2169);
xor (n2168,n2166,n1769);
or (n2169,n2170,n2172);
and (n2170,n2171,n1775);
xor (n2171,n2151,n2152);
and (n2172,n2173,n2174);
xor (n2173,n2171,n1775);
and (n2174,n2175,n1780);
xor (n2175,n2156,n2157);
or (n2176,n2177,n2179);
and (n2177,n2178,n1769);
xor (n2178,n2163,n2164);
and (n2179,n2180,n2181);
xor (n2180,n2178,n1769);
or (n2181,n2182,n2184);
and (n2182,n2183,n1775);
xor (n2183,n2168,n2169);
and (n2184,n2185,n2186);
xor (n2185,n2183,n1775);
and (n2186,n2187,n1780);
xor (n2187,n2173,n2174);
or (n2188,n2189,n2191);
and (n2189,n2190,n1775);
xor (n2190,n2180,n2181);
and (n2191,n2192,n2193);
xor (n2192,n2190,n1775);
and (n2193,n2194,n1780);
xor (n2194,n2185,n2186);
and (n2195,n2196,n1780);
xor (n2196,n2192,n2193);
endmodule
