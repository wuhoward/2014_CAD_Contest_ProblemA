module top (out,n5,n20,n23,n24,n32,n33,n35,n36,n46
        ,n55,n59,n69,n70,n72,n73,n80,n86,n98,n99
        ,n101,n102,n105,n111,n123,n124,n133,n139,n168,n209
        ,n256,n311,n346,n376,n677,n1012);
output out;
input n5;
input n20;
input n23;
input n24;
input n32;
input n33;
input n35;
input n36;
input n46;
input n55;
input n59;
input n69;
input n70;
input n72;
input n73;
input n80;
input n86;
input n98;
input n99;
input n101;
input n102;
input n105;
input n111;
input n123;
input n124;
input n133;
input n139;
input n168;
input n209;
input n256;
input n311;
input n346;
input n376;
input n677;
input n1012;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n21;
wire n22;
wire n25;
wire n26;
wire n27;
wire n28;
wire n29;
wire n30;
wire n31;
wire n34;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n54;
wire n56;
wire n57;
wire n58;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n71;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n100;
wire n103;
wire n104;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
xor (out,n0,n1014);
nor (n0,n1,n1013);
not (n1,n2);
nand (n2,n3,n1012);
or (n3,n4,n662);
and (n4,n5,n6);
nand (n6,n7,n661);
or (n7,n8,n268);
not (n8,n9);
nand (n9,n10,n267);
nand (n10,n11,n219);
not (n11,n12);
xor (n12,n13,n177);
xor (n13,n14,n89);
xor (n14,n15,n61);
xor (n15,n16,n49);
nand (n16,n17,n42);
or (n17,n18,n27);
nor (n18,n19,n25);
and (n19,n20,n21);
not (n21,n22);
wire s0n22,s1n22,notn22;
or (n22,s0n22,s1n22);
not(notn22,n5);
and (s0n22,notn22,n23);
and (s1n22,n5,n24);
and (n25,n26,n22);
not (n26,n20);
nand (n27,n28,n39);
nor (n28,n29,n37);
and (n29,n30,n34);
not (n30,n31);
wire s0n31,s1n31,notn31;
or (n31,s0n31,s1n31);
not(notn31,n5);
and (s0n31,notn31,n32);
and (s1n31,n5,n33);
wire s0n34,s1n34,notn34;
or (n34,s0n34,s1n34);
not(notn34,n5);
and (s0n34,notn34,n35);
and (s1n34,n5,n36);
and (n37,n31,n38);
not (n38,n34);
nand (n39,n40,n41);
or (n40,n30,n22);
nand (n41,n22,n30);
nand (n42,n43,n44);
not (n43,n28);
nor (n44,n45,n47);
and (n45,n46,n22);
and (n47,n48,n21);
not (n48,n46);
nor (n49,n50,n56);
nand (n50,n22,n51);
not (n51,n52);
wire s0n52,s1n52,notn52;
or (n52,s0n52,s1n52);
not(notn52,n5);
and (s0n52,notn52,1'b0);
and (s1n52,n5,n54);
and (n54,n55,n24);
nor (n56,n57,n60);
and (n57,n52,n58);
not (n58,n59);
and (n60,n51,n59);
nand (n61,n62,n83);
or (n62,n63,n78);
nand (n63,n64,n75);
not (n64,n65);
nand (n65,n66,n74);
or (n66,n67,n71);
not (n67,n68);
wire s0n68,s1n68,notn68;
or (n68,s0n68,s1n68);
not(notn68,n5);
and (s0n68,notn68,n69);
and (s1n68,n5,n70);
wire s0n71,s1n71,notn71;
or (n71,s0n71,s1n71);
not(notn71,n5);
and (s0n71,notn71,n72);
and (s1n71,n5,n73);
nand (n74,n71,n67);
nand (n75,n76,n77);
or (n76,n67,n34);
nand (n77,n34,n67);
nor (n78,n79,n81);
and (n79,n38,n80);
and (n81,n34,n82);
not (n82,n80);
or (n83,n64,n84);
nor (n84,n85,n87);
and (n85,n38,n86);
and (n87,n34,n88);
not (n88,n86);
xor (n89,n90,n155);
xor (n90,n91,n142);
xor (n91,n92,n115);
nand (n92,n93,n108);
or (n93,n94,n103);
not (n94,n95);
nor (n95,n96,n100);
not (n96,n97);
wire s0n97,s1n97,notn97;
or (n97,s0n97,s1n97);
not(notn97,n5);
and (s0n97,notn97,n98);
and (s1n97,n5,n99);
wire s0n100,s1n100,notn100;
or (n100,s0n100,s1n100);
not(notn100,n5);
and (s0n100,notn100,n101);
and (s1n100,n5,n102);
nor (n103,n104,n106);
and (n104,n96,n105);
and (n106,n97,n107);
not (n107,n105);
or (n108,n109,n114);
nor (n109,n110,n112);
and (n110,n96,n111);
and (n112,n97,n113);
not (n113,n111);
not (n114,n100);
nand (n115,n116,n136);
or (n116,n117,n130);
not (n117,n118);
and (n118,n119,n126);
nand (n119,n120,n125);
or (n120,n121,n71);
not (n121,n122);
wire s0n122,s1n122,notn122;
or (n122,s0n122,s1n122);
not(notn122,n5);
and (s0n122,notn122,n123);
and (s1n122,n5,n124);
nand (n125,n71,n121);
not (n126,n127);
nand (n127,n128,n129);
or (n128,n121,n97);
nand (n129,n97,n121);
nor (n130,n131,n134);
and (n131,n132,n133);
not (n132,n71);
and (n134,n71,n135);
not (n135,n133);
or (n136,n126,n137);
nor (n137,n138,n140);
and (n138,n132,n139);
and (n140,n71,n141);
not (n141,n139);
and (n142,n143,n149);
nand (n143,n144,n148);
or (n144,n94,n145);
nor (n145,n146,n147);
and (n146,n96,n139);
and (n147,n97,n141);
or (n148,n103,n114);
nand (n149,n150,n154);
or (n150,n117,n151);
nor (n151,n152,n153);
and (n152,n132,n86);
and (n153,n71,n88);
or (n154,n130,n126);
or (n155,n156,n176);
and (n156,n157,n170);
xor (n157,n158,n164);
nand (n158,n159,n163);
or (n159,n27,n160);
nor (n160,n161,n162);
and (n161,n21,n59);
and (n162,n22,n58);
or (n163,n28,n18);
nor (n164,n50,n165);
nor (n165,n166,n169);
and (n166,n52,n167);
not (n167,n168);
and (n169,n51,n168);
nand (n170,n171,n172);
or (n171,n78,n64);
or (n172,n63,n173);
nor (n173,n174,n175);
and (n174,n38,n46);
and (n175,n34,n48);
and (n176,n158,n164);
or (n177,n178,n218);
and (n178,n179,n194);
xor (n179,n180,n181);
xor (n180,n143,n149);
and (n181,n182,n188);
nand (n182,n183,n187);
or (n183,n94,n184);
nor (n184,n185,n186);
and (n185,n96,n133);
and (n186,n97,n135);
or (n187,n145,n114);
nand (n188,n189,n193);
or (n189,n117,n190);
nor (n190,n191,n192);
and (n191,n132,n80);
and (n192,n71,n82);
or (n193,n151,n126);
or (n194,n195,n217);
and (n195,n196,n211);
xor (n196,n197,n205);
nand (n197,n198,n203);
or (n198,n199,n27);
not (n199,n200);
nor (n200,n201,n202);
and (n201,n168,n22);
and (n202,n167,n21);
nand (n203,n204,n43);
not (n204,n160);
nor (n205,n50,n206);
nor (n206,n207,n210);
and (n207,n52,n208);
not (n208,n209);
and (n210,n51,n209);
nand (n211,n212,n216);
or (n212,n63,n213);
nor (n213,n214,n215);
and (n214,n38,n20);
and (n215,n34,n26);
or (n216,n64,n173);
and (n217,n197,n205);
and (n218,n180,n181);
not (n219,n220);
or (n220,n221,n266);
and (n221,n222,n225);
xor (n222,n223,n224);
xor (n223,n157,n170);
xor (n224,n179,n194);
or (n225,n226,n265);
and (n226,n227,n242);
xor (n227,n228,n229);
xor (n228,n182,n188);
and (n229,n230,n236);
nand (n230,n231,n235);
or (n231,n94,n232);
nor (n232,n233,n234);
and (n233,n96,n86);
and (n234,n97,n88);
or (n235,n184,n114);
nand (n236,n237,n241);
or (n237,n117,n238);
nor (n238,n239,n240);
and (n239,n132,n46);
and (n240,n71,n48);
or (n241,n126,n190);
or (n242,n243,n264);
and (n243,n244,n258);
xor (n244,n245,n252);
nand (n245,n246,n251);
or (n246,n247,n27);
not (n247,n248);
nor (n248,n249,n250);
and (n249,n209,n22);
and (n250,n208,n21);
nand (n251,n43,n200);
nor (n252,n50,n253);
nor (n253,n254,n257);
and (n254,n52,n255);
not (n255,n256);
and (n257,n51,n256);
nand (n258,n259,n263);
or (n259,n63,n260);
nor (n260,n261,n262);
and (n261,n38,n59);
and (n262,n34,n58);
or (n263,n64,n213);
and (n264,n245,n252);
and (n265,n228,n229);
and (n266,n223,n224);
nand (n267,n12,n220);
not (n268,n269);
nand (n269,n270,n656);
or (n270,n271,n356);
nand (n271,n272,n322);
not (n272,n273);
nor (n273,n274,n275);
xor (n274,n222,n225);
or (n275,n276,n321);
and (n276,n277,n280);
xor (n277,n278,n279);
xor (n278,n196,n211);
xor (n279,n227,n242);
or (n280,n281,n320);
and (n281,n282,n297);
xor (n282,n283,n284);
xor (n283,n230,n236);
and (n284,n285,n291);
nand (n285,n286,n290);
or (n286,n94,n287);
nor (n287,n288,n289);
and (n288,n96,n80);
and (n289,n97,n82);
or (n290,n232,n114);
nand (n291,n292,n296);
or (n292,n117,n293);
nor (n293,n294,n295);
and (n294,n132,n20);
and (n295,n71,n26);
or (n296,n238,n126);
or (n297,n298,n319);
and (n298,n299,n313);
xor (n299,n300,n307);
nand (n300,n301,n306);
or (n301,n302,n27);
not (n302,n303);
nor (n303,n304,n305);
and (n304,n256,n22);
and (n305,n255,n21);
nand (n306,n43,n248);
nor (n307,n50,n308);
nor (n308,n309,n312);
and (n309,n52,n310);
not (n310,n311);
and (n312,n51,n311);
nand (n313,n314,n318);
or (n314,n63,n315);
nor (n315,n316,n317);
and (n316,n38,n168);
and (n317,n34,n167);
or (n318,n64,n260);
and (n319,n300,n307);
and (n320,n283,n284);
and (n321,n278,n279);
nand (n322,n323,n325);
not (n323,n324);
xor (n324,n277,n280);
not (n325,n326);
or (n326,n327,n355);
and (n327,n328,n331);
xor (n328,n329,n330);
xor (n329,n244,n258);
xor (n330,n282,n297);
and (n331,n332,n333);
xor (n332,n285,n291);
or (n333,n334,n354);
and (n334,n335,n348);
xor (n335,n336,n342);
nand (n336,n337,n341);
or (n337,n338,n27);
nor (n338,n339,n340);
and (n339,n311,n21);
and (n340,n310,n22);
nand (n341,n303,n43);
nor (n342,n50,n343);
nor (n343,n344,n347);
and (n344,n52,n345);
not (n345,n346);
and (n347,n51,n346);
nand (n348,n349,n353);
or (n349,n94,n350);
nor (n350,n351,n352);
and (n351,n96,n46);
and (n352,n97,n48);
or (n353,n287,n114);
and (n354,n336,n342);
and (n355,n329,n330);
not (n356,n357);
nand (n357,n358,n511,n655);
nand (n358,n359,n504);
nand (n359,n360,n503);
or (n360,n361,n492);
nor (n361,n362,n491);
and (n362,n363,n463);
not (n363,n364);
nor (n364,n365,n446);
or (n365,n366,n445);
and (n366,n367,n416);
xor (n367,n368,n403);
or (n368,n369,n402);
and (n369,n370,n393);
xor (n370,n371,n383);
nand (n371,n372,n379);
or (n372,n373,n27);
not (n373,n374);
nand (n374,n375,n377);
or (n375,n21,n376);
or (n377,n22,n378);
not (n378,n376);
or (n379,n28,n380);
nor (n380,n381,n382);
and (n381,n346,n21);
and (n382,n345,n22);
nand (n383,n384,n389);
or (n384,n385,n117);
not (n385,n386);
nand (n386,n387,n388);
or (n387,n71,n208);
or (n388,n132,n209);
nand (n389,n127,n390);
nor (n390,n391,n392);
and (n391,n168,n71);
and (n392,n167,n132);
nand (n393,n394,n398);
or (n394,n63,n395);
nor (n395,n396,n397);
and (n396,n38,n311);
and (n397,n34,n310);
or (n398,n64,n399);
nor (n399,n400,n401);
and (n400,n38,n256);
and (n401,n34,n255);
and (n402,n371,n383);
xor (n403,n404,n413);
xor (n404,n405,n407);
and (n405,n406,n376);
not (n406,n50);
nand (n407,n408,n412);
or (n408,n94,n409);
nor (n409,n410,n411);
and (n410,n26,n97);
and (n411,n20,n96);
or (n412,n350,n114);
nand (n413,n414,n415);
or (n414,n27,n380);
or (n415,n28,n338);
xor (n416,n417,n431);
xor (n417,n418,n425);
nand (n418,n419,n421);
or (n419,n117,n420);
not (n420,n390);
or (n421,n126,n422);
nor (n422,n423,n424);
and (n423,n132,n59);
and (n424,n71,n58);
nand (n425,n426,n427);
or (n426,n63,n399);
or (n427,n64,n428);
nor (n428,n429,n430);
and (n429,n38,n209);
and (n430,n34,n208);
and (n431,n432,n437);
nor (n432,n433,n21);
nor (n433,n434,n436);
and (n434,n38,n435);
nand (n435,n31,n376);
and (n436,n30,n378);
nand (n437,n438,n443);
or (n438,n439,n94);
not (n439,n440);
nor (n440,n441,n442);
and (n441,n59,n97);
and (n442,n58,n96);
nand (n443,n444,n100);
not (n444,n409);
and (n445,n368,n403);
xor (n446,n447,n452);
xor (n447,n448,n449);
xor (n448,n335,n348);
or (n449,n450,n451);
and (n450,n417,n431);
and (n451,n418,n425);
xor (n452,n453,n460);
xor (n453,n454,n457);
nand (n454,n455,n456);
or (n455,n63,n428);
or (n456,n64,n315);
nand (n457,n458,n459);
or (n458,n117,n422);
or (n459,n293,n126);
or (n460,n461,n462);
and (n461,n404,n413);
and (n462,n405,n407);
not (n463,n464);
nand (n464,n465,n466);
xor (n465,n367,n416);
or (n466,n467,n490);
and (n467,n468,n489);
xor (n468,n469,n470);
xor (n469,n432,n437);
or (n470,n471,n488);
and (n471,n472,n481);
xor (n472,n473,n474);
and (n473,n43,n376);
nand (n474,n475,n476);
or (n475,n114,n439);
nand (n476,n477,n95);
not (n477,n478);
nor (n478,n479,n480);
and (n479,n168,n96);
and (n480,n167,n97);
nand (n481,n482,n487);
or (n482,n483,n117);
not (n483,n484);
nor (n484,n485,n486);
and (n485,n256,n71);
and (n486,n132,n255);
nand (n487,n127,n386);
and (n488,n473,n474);
xor (n489,n370,n393);
and (n490,n469,n470);
and (n491,n365,n446);
nor (n492,n493,n500);
xor (n493,n494,n497);
xor (n494,n495,n496);
xor (n495,n299,n313);
xor (n496,n332,n333);
or (n497,n498,n499);
and (n498,n453,n460);
and (n499,n454,n457);
or (n500,n501,n502);
and (n501,n447,n452);
and (n502,n448,n449);
nand (n503,n493,n500);
nand (n504,n505,n507);
not (n505,n506);
xor (n506,n328,n331);
not (n507,n508);
or (n508,n509,n510);
and (n509,n494,n497);
and (n510,n495,n496);
nand (n511,n504,n512,n654);
nor (n512,n513,n651);
nor (n513,n514,n649);
and (n514,n515,n644);
or (n515,n516,n643);
and (n516,n517,n559);
xor (n517,n518,n552);
or (n518,n519,n551);
and (n519,n520,n539);
xor (n520,n521,n528);
nand (n521,n522,n527);
or (n522,n523,n117);
not (n523,n524);
nor (n524,n525,n526);
and (n525,n310,n132);
and (n526,n311,n71);
nand (n527,n127,n484);
nand (n528,n529,n534);
or (n529,n530,n64);
not (n530,n531);
nor (n531,n532,n533);
and (n532,n346,n34);
and (n533,n345,n38);
nand (n534,n535,n536);
not (n535,n63);
nand (n536,n537,n538);
or (n537,n38,n376);
or (n538,n34,n378);
xor (n539,n540,n545);
and (n540,n541,n34);
nand (n541,n542,n544);
or (n542,n71,n543);
and (n543,n376,n68);
or (n544,n68,n376);
nand (n545,n546,n550);
or (n546,n94,n547);
nor (n547,n548,n549);
and (n548,n96,n209);
and (n549,n97,n208);
or (n550,n478,n114);
and (n551,n521,n528);
xor (n552,n553,n558);
xor (n553,n554,n557);
nand (n554,n555,n556);
or (n555,n530,n63);
or (n556,n64,n395);
and (n557,n540,n545);
xor (n558,n472,n481);
or (n559,n560,n642);
and (n560,n561,n582);
xor (n561,n562,n581);
or (n562,n563,n580);
and (n563,n564,n573);
xor (n564,n565,n566);
and (n565,n65,n376);
nand (n566,n567,n572);
or (n567,n568,n117);
not (n568,n569);
nor (n569,n570,n571);
and (n570,n346,n71);
and (n571,n345,n132);
nand (n572,n524,n127);
nand (n573,n574,n579);
or (n574,n94,n575);
not (n575,n576);
nor (n576,n577,n578);
and (n577,n255,n96);
and (n578,n256,n97);
or (n579,n547,n114);
and (n580,n565,n566);
xor (n581,n520,n539);
or (n582,n583,n641);
and (n583,n584,n640);
xor (n584,n585,n599);
nor (n585,n586,n594);
not (n586,n587);
nand (n587,n588,n593);
or (n588,n589,n94);
not (n589,n590);
nand (n590,n591,n592);
or (n591,n310,n97);
nand (n592,n97,n310);
nand (n593,n576,n100);
nand (n594,n595,n71);
nand (n595,n596,n598);
or (n596,n97,n597);
and (n597,n376,n122);
or (n598,n122,n376);
nand (n599,n600,n638);
or (n600,n601,n624);
not (n601,n602);
nand (n602,n603,n623);
or (n603,n604,n613);
nor (n604,n605,n612);
nand (n605,n606,n611);
or (n606,n607,n94);
not (n607,n608);
nand (n608,n609,n610);
or (n609,n345,n97);
nand (n610,n97,n345);
nand (n611,n590,n100);
nor (n612,n126,n378);
nand (n613,n614,n621);
nand (n614,n615,n620);
or (n615,n616,n94);
not (n616,n617);
nand (n617,n618,n619);
or (n618,n96,n376);
or (n619,n97,n378);
nand (n620,n608,n100);
nor (n621,n622,n96);
and (n622,n376,n100);
nand (n623,n605,n612);
not (n624,n625);
nand (n625,n626,n634);
not (n626,n627);
nand (n627,n628,n633);
or (n628,n629,n117);
not (n629,n630);
nand (n630,n631,n632);
or (n631,n132,n376);
or (n632,n71,n378);
nand (n633,n127,n569);
nor (n634,n635,n637);
and (n635,n586,n636);
not (n636,n594);
and (n637,n587,n594);
nand (n638,n639,n627);
not (n639,n634);
xor (n640,n564,n573);
and (n641,n585,n599);
and (n642,n562,n581);
and (n643,n518,n552);
or (n644,n645,n646);
xor (n645,n468,n489);
or (n646,n647,n648);
and (n647,n553,n558);
and (n648,n554,n557);
not (n649,n650);
nand (n650,n645,n646);
nand (n651,n652,n363);
not (n652,n653);
nor (n653,n465,n466);
not (n654,n492);
nand (n655,n506,n508);
not (n656,n657);
nand (n657,n658,n660);
or (n658,n273,n659);
nand (n659,n324,n326);
nand (n660,n274,n275);
or (n661,n269,n9);
and (n662,n663,n664);
not (n663,n5);
nand (n664,n665,n1011);
or (n665,n666,n735);
nand (n666,n667,n734);
or (n667,n668,n718);
or (n668,n669,n717);
and (n669,n670,n703);
xor (n670,n671,n686);
not (n671,n672);
nor (n672,n673,n680);
and (n673,n535,n674);
not (n674,n675);
nor (n675,n676,n678);
and (n676,n38,n677);
and (n678,n34,n679);
not (n679,n677);
and (n680,n65,n681);
nand (n681,n682,n685);
or (n682,n34,n683);
not (n683,n684);
and (n684,n55,n677);
or (n685,n38,n684);
xor (n686,n687,n699);
xor (n687,n688,n690);
nand (n688,n689,n681);
or (n689,n535,n65);
nand (n690,n691,n695);
or (n691,n27,n692);
nor (n692,n693,n694);
and (n693,n21,n111);
and (n694,n22,n113);
or (n695,n28,n696);
nor (n696,n697,n698);
and (n697,n21,n677);
and (n698,n22,n679);
nor (n699,n50,n700);
nor (n700,n701,n702);
and (n701,n52,n107);
and (n702,n51,n105);
or (n703,n704,n716);
and (n704,n705,n672);
xor (n705,n706,n712);
nand (n706,n707,n711);
or (n707,n27,n708);
nor (n708,n709,n710);
and (n709,n21,n105);
and (n710,n22,n107);
or (n711,n28,n692);
nor (n712,n50,n713);
nor (n713,n714,n715);
and (n714,n52,n141);
and (n715,n51,n139);
and (n716,n706,n712);
and (n717,n671,n686);
xor (n718,n719,n731);
xor (n719,n720,n727);
nand (n720,n721,n726);
or (n721,n722,n28);
not (n722,n723);
nand (n723,n724,n725);
or (n724,n22,n683);
or (n725,n21,n684);
or (n726,n27,n696);
nand (n727,n728,n729,n406);
or (n728,n52,n111);
not (n729,n730);
and (n730,n111,n52);
or (n731,n732,n733);
and (n732,n687,n699);
and (n733,n688,n690);
nand (n734,n668,n718);
nand (n735,n736,n1005);
or (n736,n737,n852);
not (n737,n738);
nor (n738,n739,n845);
nor (n739,n740,n836);
or (n740,n741,n835);
and (n741,n742,n796);
xor (n742,n743,n760);
xor (n743,n744,n756);
xor (n744,n745,n750);
nand (n745,n746,n747);
or (n746,n118,n127);
nand (n747,n748,n749);
or (n748,n71,n683);
or (n749,n132,n684);
nand (n750,n751,n755);
or (n751,n63,n752);
nor (n752,n753,n754);
and (n753,n38,n111);
and (n754,n34,n113);
or (n755,n64,n675);
nor (n756,n50,n757);
nor (n757,n758,n759);
and (n758,n52,n135);
and (n759,n51,n133);
xor (n760,n761,n776);
xor (n761,n762,n768);
nand (n762,n763,n767);
or (n763,n27,n764);
nor (n764,n765,n766);
and (n765,n21,n139);
and (n766,n22,n141);
or (n767,n28,n708);
nand (n768,n769,n771);
or (n769,n770,n126);
not (n770,n747);
nand (n771,n772,n118);
not (n772,n773);
nor (n773,n774,n775);
and (n774,n132,n677);
and (n775,n71,n679);
or (n776,n777,n795);
and (n777,n778,n789);
xor (n778,n779,n783);
nor (n779,n50,n780);
nor (n780,n781,n782);
and (n781,n52,n88);
and (n782,n51,n86);
nand (n783,n784,n788);
or (n784,n63,n785);
nor (n785,n786,n787);
and (n786,n105,n38);
and (n787,n107,n34);
or (n788,n64,n752);
nand (n789,n790,n794);
or (n790,n27,n791);
nor (n791,n792,n793);
and (n792,n21,n133);
and (n793,n22,n135);
or (n794,n28,n764);
and (n795,n779,n783);
or (n796,n797,n834);
and (n797,n798,n814);
xor (n798,n799,n800);
not (n799,n768);
or (n800,n801,n807);
nand (n801,n802,n806);
or (n802,n27,n803);
nor (n803,n804,n805);
and (n804,n21,n86);
and (n805,n22,n88);
or (n806,n28,n791);
nand (n807,n808,n813);
or (n808,n117,n809);
not (n809,n810);
nand (n810,n811,n812);
or (n811,n71,n113);
or (n812,n132,n111);
or (n813,n126,n773);
or (n814,n815,n833);
and (n815,n816,n827);
xor (n816,n817,n821);
nor (n817,n50,n818);
nor (n818,n819,n820);
and (n819,n52,n82);
and (n820,n51,n80);
nand (n821,n822,n823);
or (n822,n100,n95);
not (n823,n824);
nor (n824,n825,n826);
and (n825,n96,n684);
and (n826,n97,n683);
nand (n827,n828,n829);
or (n828,n785,n64);
or (n829,n63,n830);
nor (n830,n831,n832);
and (n831,n38,n139);
and (n832,n34,n141);
and (n833,n817,n821);
and (n834,n799,n800);
and (n835,n743,n760);
xor (n836,n837,n842);
xor (n837,n838,n841);
or (n838,n839,n840);
and (n839,n744,n756);
and (n840,n745,n750);
xor (n841,n705,n672);
or (n842,n843,n844);
and (n843,n761,n776);
and (n844,n762,n768);
and (n845,n846,n850);
not (n846,n847);
or (n847,n848,n849);
and (n848,n837,n842);
and (n849,n838,n841);
not (n850,n851);
xor (n851,n670,n703);
not (n852,n853);
nand (n853,n854,n992);
or (n854,n855,n975);
not (n855,n856);
and (n856,n857,n956,n969);
nor (n857,n858,n933);
nor (n858,n859,n902);
or (n859,n860,n901);
and (n860,n861,n898);
xor (n861,n862,n881);
xor (n862,n863,n875);
xor (n863,n864,n871);
nand (n864,n865,n867);
or (n865,n866,n27);
not (n866,n44);
nand (n867,n43,n868);
nor (n868,n869,n870);
and (n869,n80,n22);
and (n870,n82,n21);
nor (n871,n50,n872);
nor (n872,n873,n874);
and (n873,n52,n26);
and (n874,n51,n20);
nand (n875,n876,n877);
or (n876,n63,n84);
or (n877,n64,n878);
nor (n878,n879,n880);
and (n879,n38,n133);
and (n880,n34,n135);
xor (n881,n882,n895);
xor (n882,n883,n894);
xor (n883,n884,n890);
nand (n884,n885,n886);
or (n885,n94,n109);
or (n886,n887,n114);
nor (n887,n888,n889);
and (n888,n96,n677);
and (n889,n97,n679);
nand (n890,n891,n892);
or (n891,n117,n137);
or (n892,n893,n126);
xor (n893,n105,n132);
and (n894,n92,n115);
or (n895,n896,n897);
and (n896,n15,n61);
and (n897,n16,n49);
or (n898,n899,n900);
and (n899,n90,n155);
and (n900,n91,n142);
and (n901,n862,n881);
xor (n902,n903,n930);
xor (n903,n904,n917);
xor (n904,n905,n914);
xor (n905,n906,n910);
nand (n906,n907,n909);
or (n907,n908,n27);
not (n908,n868);
or (n909,n28,n803);
nor (n910,n50,n911);
nor (n911,n912,n913);
and (n912,n52,n48);
and (n913,n51,n46);
nand (n914,n915,n916);
or (n915,n63,n878);
or (n916,n64,n830);
xor (n917,n918,n927);
xor (n918,n919,n926);
xor (n919,n920,n923);
nand (n920,n921,n922);
or (n921,n94,n887);
or (n922,n824,n114);
nand (n923,n924,n925);
or (n924,n893,n117);
nand (n925,n127,n810);
and (n926,n884,n890);
or (n927,n928,n929);
and (n928,n863,n875);
and (n929,n864,n871);
or (n930,n931,n932);
and (n931,n882,n895);
and (n932,n883,n894);
not (n933,n934);
nand (n934,n935,n952);
not (n935,n936);
xor (n936,n937,n942);
xor (n937,n938,n939);
xor (n938,n816,n827);
or (n939,n940,n941);
and (n940,n918,n927);
and (n941,n919,n926);
xor (n942,n943,n948);
xor (n943,n944,n945);
and (n944,n920,n923);
or (n945,n946,n947);
and (n946,n905,n914);
and (n947,n906,n910);
nand (n948,n949,n800);
or (n949,n950,n951);
not (n950,n807);
not (n951,n801);
not (n952,n953);
or (n953,n954,n955);
and (n954,n903,n930);
and (n955,n904,n917);
nand (n956,n957,n959);
not (n957,n958);
xor (n958,n742,n796);
not (n959,n960);
or (n960,n961,n968);
and (n961,n962,n965);
xor (n962,n963,n964);
xor (n963,n778,n789);
xor (n964,n798,n814);
or (n965,n966,n967);
and (n966,n943,n948);
and (n967,n944,n945);
and (n968,n963,n964);
not (n969,n970);
nor (n970,n971,n972);
xor (n971,n962,n965);
or (n972,n973,n974);
and (n973,n937,n942);
and (n974,n938,n939);
not (n975,n976);
nand (n976,n977,n987,n991);
nand (n977,n357,n978);
nor (n978,n271,n979);
nand (n979,n10,n980);
nand (n980,n981,n983);
not (n981,n982);
xor (n982,n861,n898);
not (n983,n984);
or (n984,n985,n986);
and (n985,n13,n177);
and (n986,n14,n89);
nand (n987,n988,n980);
nand (n988,n989,n267);
or (n989,n990,n656);
not (n990,n10);
nand (n991,n984,n982);
not (n992,n993);
nand (n993,n994,n1004);
or (n994,n995,n996);
not (n995,n956);
not (n996,n997);
nand (n997,n998,n1003);
or (n998,n999,n970);
nor (n999,n1000,n1002);
and (n1000,n1001,n934);
and (n1001,n859,n902);
nor (n1002,n935,n952);
nand (n1003,n971,n972);
or (n1004,n957,n959);
nor (n1005,n1006,n1010);
and (n1006,n1007,n1009);
not (n1007,n1008);
nand (n1008,n740,n836);
not (n1009,n845);
nor (n1010,n846,n850);
nand (n1011,n735,n666);
nor (n1013,n3,n1012);
xor (n1014,n1012,n1015);
wire s0n1015,s1n1015,notn1015;
or (n1015,s0n1015,s1n1015);
not(notn1015,n5);
and (s0n1015,notn1015,n1016);
and (s1n1015,n5,n2206);
xor (n1016,n1017,n1789);
xor (n1017,n1018,n2204);
xor (n1018,n1019,n1784);
xor (n1019,n1020,n2197);
xor (n1020,n1021,n1778);
xor (n1021,n1022,n2185);
xor (n1022,n1023,n1772);
xor (n1023,n1024,n2168);
xor (n1024,n1025,n1766);
xor (n1025,n1026,n2146);
xor (n1026,n1027,n1760);
xor (n1027,n1028,n2119);
xor (n1028,n1029,n1754);
xor (n1029,n1030,n2087);
xor (n1030,n1031,n1748);
xor (n1031,n1032,n2050);
xor (n1032,n1033,n1742);
xor (n1033,n1034,n2008);
xor (n1034,n1035,n1736);
xor (n1035,n1036,n1961);
xor (n1036,n1037,n1730);
xor (n1037,n1038,n1909);
xor (n1038,n1039,n1724);
xor (n1039,n1040,n1852);
xor (n1040,n1041,n1718);
xor (n1041,n1042,n1790);
xor (n1042,n1043,n1712);
xor (n1043,n1044,n1709);
xor (n1044,n1045,n730);
xor (n1045,n1046,n1627);
xor (n1046,n1047,n1626);
xor (n1047,n1048,n1533);
xor (n1048,n1049,n1532);
xor (n1049,n1050,n1435);
xor (n1050,n1051,n1434);
xor (n1051,n1052,n1067);
xor (n1052,n1053,n1066);
xor (n1053,n1054,n1065);
xor (n1054,n1055,n1064);
xor (n1055,n1056,n1063);
xor (n1056,n1057,n1062);
xor (n1057,n1058,n1061);
xor (n1058,n1059,n1060);
and (n1059,n684,n100);
and (n1060,n684,n97);
and (n1061,n1059,n1060);
and (n1062,n684,n122);
and (n1063,n1057,n1062);
and (n1064,n684,n71);
and (n1065,n1055,n1064);
and (n1066,n684,n68);
or (n1067,n1068,n1069);
and (n1068,n1053,n1066);
and (n1069,n1052,n1070);
or (n1070,n1068,n1071);
and (n1071,n1052,n1072);
or (n1072,n1073,n1346);
and (n1073,n1074,n1345);
xor (n1074,n1054,n1075);
or (n1075,n1076,n1260);
and (n1076,n1077,n1259);
xor (n1077,n1056,n1078);
or (n1078,n1079,n1171);
and (n1079,n1080,n1170);
xor (n1080,n1058,n1081);
or (n1081,n1061,n1082);
and (n1082,n1083,n1085);
xor (n1083,n1059,n1084);
and (n1084,n677,n97);
or (n1085,n1086,n1089);
and (n1086,n1087,n1088);
and (n1087,n677,n100);
and (n1088,n111,n97);
and (n1089,n1090,n1091);
xor (n1090,n1087,n1088);
or (n1091,n1092,n1095);
and (n1092,n1093,n1094);
and (n1093,n111,n100);
and (n1094,n105,n97);
and (n1095,n1096,n1097);
xor (n1096,n1093,n1094);
or (n1097,n1098,n1101);
and (n1098,n1099,n1100);
and (n1099,n105,n100);
and (n1100,n139,n97);
and (n1101,n1102,n1103);
xor (n1102,n1099,n1100);
or (n1103,n1104,n1107);
and (n1104,n1105,n1106);
and (n1105,n139,n100);
and (n1106,n133,n97);
and (n1107,n1108,n1109);
xor (n1108,n1105,n1106);
or (n1109,n1110,n1113);
and (n1110,n1111,n1112);
and (n1111,n133,n100);
and (n1112,n86,n97);
and (n1113,n1114,n1115);
xor (n1114,n1111,n1112);
or (n1115,n1116,n1119);
and (n1116,n1117,n1118);
and (n1117,n86,n100);
and (n1118,n80,n97);
and (n1119,n1120,n1121);
xor (n1120,n1117,n1118);
or (n1121,n1122,n1125);
and (n1122,n1123,n1124);
and (n1123,n80,n100);
and (n1124,n46,n97);
and (n1125,n1126,n1127);
xor (n1126,n1123,n1124);
or (n1127,n1128,n1131);
and (n1128,n1129,n1130);
and (n1129,n46,n100);
and (n1130,n20,n97);
and (n1131,n1132,n1133);
xor (n1132,n1129,n1130);
or (n1133,n1134,n1136);
and (n1134,n1135,n441);
and (n1135,n20,n100);
and (n1136,n1137,n1138);
xor (n1137,n1135,n441);
or (n1138,n1139,n1142);
and (n1139,n1140,n1141);
and (n1140,n59,n100);
and (n1141,n168,n97);
and (n1142,n1143,n1144);
xor (n1143,n1140,n1141);
or (n1144,n1145,n1148);
and (n1145,n1146,n1147);
and (n1146,n168,n100);
and (n1147,n209,n97);
and (n1148,n1149,n1150);
xor (n1149,n1146,n1147);
or (n1150,n1151,n1153);
and (n1151,n1152,n578);
and (n1152,n209,n100);
and (n1153,n1154,n1155);
xor (n1154,n1152,n578);
or (n1155,n1156,n1159);
and (n1156,n1157,n1158);
and (n1157,n256,n100);
and (n1158,n311,n97);
and (n1159,n1160,n1161);
xor (n1160,n1157,n1158);
or (n1161,n1162,n1165);
and (n1162,n1163,n1164);
and (n1163,n311,n100);
and (n1164,n346,n97);
and (n1165,n1166,n1167);
xor (n1166,n1163,n1164);
and (n1167,n1168,n1169);
and (n1168,n346,n100);
and (n1169,n376,n97);
and (n1170,n677,n122);
and (n1171,n1172,n1173);
xor (n1172,n1080,n1170);
or (n1173,n1174,n1177);
and (n1174,n1175,n1176);
xor (n1175,n1083,n1085);
and (n1176,n111,n122);
and (n1177,n1178,n1179);
xor (n1178,n1175,n1176);
or (n1179,n1180,n1183);
and (n1180,n1181,n1182);
xor (n1181,n1090,n1091);
and (n1182,n105,n122);
and (n1183,n1184,n1185);
xor (n1184,n1181,n1182);
or (n1185,n1186,n1189);
and (n1186,n1187,n1188);
xor (n1187,n1096,n1097);
and (n1188,n139,n122);
and (n1189,n1190,n1191);
xor (n1190,n1187,n1188);
or (n1191,n1192,n1195);
and (n1192,n1193,n1194);
xor (n1193,n1102,n1103);
and (n1194,n133,n122);
and (n1195,n1196,n1197);
xor (n1196,n1193,n1194);
or (n1197,n1198,n1201);
and (n1198,n1199,n1200);
xor (n1199,n1108,n1109);
and (n1200,n86,n122);
and (n1201,n1202,n1203);
xor (n1202,n1199,n1200);
or (n1203,n1204,n1207);
and (n1204,n1205,n1206);
xor (n1205,n1114,n1115);
and (n1206,n80,n122);
and (n1207,n1208,n1209);
xor (n1208,n1205,n1206);
or (n1209,n1210,n1213);
and (n1210,n1211,n1212);
xor (n1211,n1120,n1121);
and (n1212,n46,n122);
and (n1213,n1214,n1215);
xor (n1214,n1211,n1212);
or (n1215,n1216,n1219);
and (n1216,n1217,n1218);
xor (n1217,n1126,n1127);
and (n1218,n20,n122);
and (n1219,n1220,n1221);
xor (n1220,n1217,n1218);
or (n1221,n1222,n1225);
and (n1222,n1223,n1224);
xor (n1223,n1132,n1133);
and (n1224,n59,n122);
and (n1225,n1226,n1227);
xor (n1226,n1223,n1224);
or (n1227,n1228,n1231);
and (n1228,n1229,n1230);
xor (n1229,n1137,n1138);
and (n1230,n168,n122);
and (n1231,n1232,n1233);
xor (n1232,n1229,n1230);
or (n1233,n1234,n1237);
and (n1234,n1235,n1236);
xor (n1235,n1143,n1144);
and (n1236,n209,n122);
and (n1237,n1238,n1239);
xor (n1238,n1235,n1236);
or (n1239,n1240,n1243);
and (n1240,n1241,n1242);
xor (n1241,n1149,n1150);
and (n1242,n256,n122);
and (n1243,n1244,n1245);
xor (n1244,n1241,n1242);
or (n1245,n1246,n1249);
and (n1246,n1247,n1248);
xor (n1247,n1154,n1155);
and (n1248,n311,n122);
and (n1249,n1250,n1251);
xor (n1250,n1247,n1248);
or (n1251,n1252,n1255);
and (n1252,n1253,n1254);
xor (n1253,n1160,n1161);
and (n1254,n346,n122);
and (n1255,n1256,n1257);
xor (n1256,n1253,n1254);
and (n1257,n1258,n597);
xor (n1258,n1166,n1167);
and (n1259,n677,n71);
and (n1260,n1261,n1262);
xor (n1261,n1077,n1259);
or (n1262,n1263,n1266);
and (n1263,n1264,n1265);
xor (n1264,n1172,n1173);
and (n1265,n111,n71);
and (n1266,n1267,n1268);
xor (n1267,n1264,n1265);
or (n1268,n1269,n1272);
and (n1269,n1270,n1271);
xor (n1270,n1178,n1179);
and (n1271,n105,n71);
and (n1272,n1273,n1274);
xor (n1273,n1270,n1271);
or (n1274,n1275,n1278);
and (n1275,n1276,n1277);
xor (n1276,n1184,n1185);
and (n1277,n139,n71);
and (n1278,n1279,n1280);
xor (n1279,n1276,n1277);
or (n1280,n1281,n1284);
and (n1281,n1282,n1283);
xor (n1282,n1190,n1191);
and (n1283,n133,n71);
and (n1284,n1285,n1286);
xor (n1285,n1282,n1283);
or (n1286,n1287,n1290);
and (n1287,n1288,n1289);
xor (n1288,n1196,n1197);
and (n1289,n86,n71);
and (n1290,n1291,n1292);
xor (n1291,n1288,n1289);
or (n1292,n1293,n1296);
and (n1293,n1294,n1295);
xor (n1294,n1202,n1203);
and (n1295,n80,n71);
and (n1296,n1297,n1298);
xor (n1297,n1294,n1295);
or (n1298,n1299,n1302);
and (n1299,n1300,n1301);
xor (n1300,n1208,n1209);
and (n1301,n46,n71);
and (n1302,n1303,n1304);
xor (n1303,n1300,n1301);
or (n1304,n1305,n1308);
and (n1305,n1306,n1307);
xor (n1306,n1214,n1215);
and (n1307,n20,n71);
and (n1308,n1309,n1310);
xor (n1309,n1306,n1307);
or (n1310,n1311,n1314);
and (n1311,n1312,n1313);
xor (n1312,n1220,n1221);
and (n1313,n59,n71);
and (n1314,n1315,n1316);
xor (n1315,n1312,n1313);
or (n1316,n1317,n1319);
and (n1317,n1318,n391);
xor (n1318,n1226,n1227);
and (n1319,n1320,n1321);
xor (n1320,n1318,n391);
or (n1321,n1322,n1325);
and (n1322,n1323,n1324);
xor (n1323,n1232,n1233);
and (n1324,n209,n71);
and (n1325,n1326,n1327);
xor (n1326,n1323,n1324);
or (n1327,n1328,n1330);
and (n1328,n1329,n485);
xor (n1329,n1238,n1239);
and (n1330,n1331,n1332);
xor (n1331,n1329,n485);
or (n1332,n1333,n1335);
and (n1333,n1334,n526);
xor (n1334,n1244,n1245);
and (n1335,n1336,n1337);
xor (n1336,n1334,n526);
or (n1337,n1338,n1340);
and (n1338,n1339,n570);
xor (n1339,n1250,n1251);
and (n1340,n1341,n1342);
xor (n1341,n1339,n570);
and (n1342,n1343,n1344);
xor (n1343,n1256,n1257);
and (n1344,n376,n71);
and (n1345,n677,n68);
and (n1346,n1347,n1348);
xor (n1347,n1074,n1345);
or (n1348,n1349,n1352);
and (n1349,n1350,n1351);
xor (n1350,n1261,n1262);
and (n1351,n111,n68);
and (n1352,n1353,n1354);
xor (n1353,n1350,n1351);
or (n1354,n1355,n1358);
and (n1355,n1356,n1357);
xor (n1356,n1267,n1268);
and (n1357,n105,n68);
and (n1358,n1359,n1360);
xor (n1359,n1356,n1357);
or (n1360,n1361,n1364);
and (n1361,n1362,n1363);
xor (n1362,n1273,n1274);
and (n1363,n139,n68);
and (n1364,n1365,n1366);
xor (n1365,n1362,n1363);
or (n1366,n1367,n1370);
and (n1367,n1368,n1369);
xor (n1368,n1279,n1280);
and (n1369,n133,n68);
and (n1370,n1371,n1372);
xor (n1371,n1368,n1369);
or (n1372,n1373,n1376);
and (n1373,n1374,n1375);
xor (n1374,n1285,n1286);
and (n1375,n86,n68);
and (n1376,n1377,n1378);
xor (n1377,n1374,n1375);
or (n1378,n1379,n1382);
and (n1379,n1380,n1381);
xor (n1380,n1291,n1292);
and (n1381,n80,n68);
and (n1382,n1383,n1384);
xor (n1383,n1380,n1381);
or (n1384,n1385,n1388);
and (n1385,n1386,n1387);
xor (n1386,n1297,n1298);
and (n1387,n46,n68);
and (n1388,n1389,n1390);
xor (n1389,n1386,n1387);
or (n1390,n1391,n1394);
and (n1391,n1392,n1393);
xor (n1392,n1303,n1304);
and (n1393,n20,n68);
and (n1394,n1395,n1396);
xor (n1395,n1392,n1393);
or (n1396,n1397,n1400);
and (n1397,n1398,n1399);
xor (n1398,n1309,n1310);
and (n1399,n59,n68);
and (n1400,n1401,n1402);
xor (n1401,n1398,n1399);
or (n1402,n1403,n1406);
and (n1403,n1404,n1405);
xor (n1404,n1315,n1316);
and (n1405,n168,n68);
and (n1406,n1407,n1408);
xor (n1407,n1404,n1405);
or (n1408,n1409,n1412);
and (n1409,n1410,n1411);
xor (n1410,n1320,n1321);
and (n1411,n209,n68);
and (n1412,n1413,n1414);
xor (n1413,n1410,n1411);
or (n1414,n1415,n1418);
and (n1415,n1416,n1417);
xor (n1416,n1326,n1327);
and (n1417,n256,n68);
and (n1418,n1419,n1420);
xor (n1419,n1416,n1417);
or (n1420,n1421,n1424);
and (n1421,n1422,n1423);
xor (n1422,n1331,n1332);
and (n1423,n311,n68);
and (n1424,n1425,n1426);
xor (n1425,n1422,n1423);
or (n1426,n1427,n1430);
and (n1427,n1428,n1429);
xor (n1428,n1336,n1337);
and (n1429,n346,n68);
and (n1430,n1431,n1432);
xor (n1431,n1428,n1429);
and (n1432,n1433,n543);
xor (n1433,n1341,n1342);
and (n1434,n684,n34);
or (n1435,n1436,n1438);
and (n1436,n1437,n1434);
xor (n1437,n1052,n1070);
and (n1438,n1439,n1440);
xor (n1439,n1437,n1434);
or (n1440,n1441,n1444);
and (n1441,n1442,n1443);
xor (n1442,n1052,n1072);
and (n1443,n677,n34);
and (n1444,n1445,n1446);
xor (n1445,n1442,n1443);
or (n1446,n1447,n1450);
and (n1447,n1448,n1449);
xor (n1448,n1347,n1348);
and (n1449,n111,n34);
and (n1450,n1451,n1452);
xor (n1451,n1448,n1449);
or (n1452,n1453,n1456);
and (n1453,n1454,n1455);
xor (n1454,n1353,n1354);
and (n1455,n105,n34);
and (n1456,n1457,n1458);
xor (n1457,n1454,n1455);
or (n1458,n1459,n1462);
and (n1459,n1460,n1461);
xor (n1460,n1359,n1360);
and (n1461,n139,n34);
and (n1462,n1463,n1464);
xor (n1463,n1460,n1461);
or (n1464,n1465,n1468);
and (n1465,n1466,n1467);
xor (n1466,n1365,n1366);
and (n1467,n133,n34);
and (n1468,n1469,n1470);
xor (n1469,n1466,n1467);
or (n1470,n1471,n1474);
and (n1471,n1472,n1473);
xor (n1472,n1371,n1372);
and (n1473,n86,n34);
and (n1474,n1475,n1476);
xor (n1475,n1472,n1473);
or (n1476,n1477,n1480);
and (n1477,n1478,n1479);
xor (n1478,n1377,n1378);
and (n1479,n80,n34);
and (n1480,n1481,n1482);
xor (n1481,n1478,n1479);
or (n1482,n1483,n1486);
and (n1483,n1484,n1485);
xor (n1484,n1383,n1384);
and (n1485,n46,n34);
and (n1486,n1487,n1488);
xor (n1487,n1484,n1485);
or (n1488,n1489,n1492);
and (n1489,n1490,n1491);
xor (n1490,n1389,n1390);
and (n1491,n20,n34);
and (n1492,n1493,n1494);
xor (n1493,n1490,n1491);
or (n1494,n1495,n1498);
and (n1495,n1496,n1497);
xor (n1496,n1395,n1396);
and (n1497,n59,n34);
and (n1498,n1499,n1500);
xor (n1499,n1496,n1497);
or (n1500,n1501,n1504);
and (n1501,n1502,n1503);
xor (n1502,n1401,n1402);
and (n1503,n168,n34);
and (n1504,n1505,n1506);
xor (n1505,n1502,n1503);
or (n1506,n1507,n1510);
and (n1507,n1508,n1509);
xor (n1508,n1407,n1408);
and (n1509,n209,n34);
and (n1510,n1511,n1512);
xor (n1511,n1508,n1509);
or (n1512,n1513,n1516);
and (n1513,n1514,n1515);
xor (n1514,n1413,n1414);
and (n1515,n256,n34);
and (n1516,n1517,n1518);
xor (n1517,n1514,n1515);
or (n1518,n1519,n1522);
and (n1519,n1520,n1521);
xor (n1520,n1419,n1420);
and (n1521,n311,n34);
and (n1522,n1523,n1524);
xor (n1523,n1520,n1521);
or (n1524,n1525,n1527);
and (n1525,n1526,n532);
xor (n1526,n1425,n1426);
and (n1527,n1528,n1529);
xor (n1528,n1526,n532);
and (n1529,n1530,n1531);
xor (n1530,n1431,n1432);
and (n1531,n376,n34);
and (n1532,n684,n31);
or (n1533,n1534,n1537);
and (n1534,n1535,n1536);
xor (n1535,n1439,n1440);
and (n1536,n677,n31);
and (n1537,n1538,n1539);
xor (n1538,n1535,n1536);
or (n1539,n1540,n1543);
and (n1540,n1541,n1542);
xor (n1541,n1445,n1446);
and (n1542,n111,n31);
and (n1543,n1544,n1545);
xor (n1544,n1541,n1542);
or (n1545,n1546,n1549);
and (n1546,n1547,n1548);
xor (n1547,n1451,n1452);
and (n1548,n105,n31);
and (n1549,n1550,n1551);
xor (n1550,n1547,n1548);
or (n1551,n1552,n1555);
and (n1552,n1553,n1554);
xor (n1553,n1457,n1458);
and (n1554,n139,n31);
and (n1555,n1556,n1557);
xor (n1556,n1553,n1554);
or (n1557,n1558,n1561);
and (n1558,n1559,n1560);
xor (n1559,n1463,n1464);
and (n1560,n133,n31);
and (n1561,n1562,n1563);
xor (n1562,n1559,n1560);
or (n1563,n1564,n1567);
and (n1564,n1565,n1566);
xor (n1565,n1469,n1470);
and (n1566,n86,n31);
and (n1567,n1568,n1569);
xor (n1568,n1565,n1566);
or (n1569,n1570,n1573);
and (n1570,n1571,n1572);
xor (n1571,n1475,n1476);
and (n1572,n80,n31);
and (n1573,n1574,n1575);
xor (n1574,n1571,n1572);
or (n1575,n1576,n1579);
and (n1576,n1577,n1578);
xor (n1577,n1481,n1482);
and (n1578,n46,n31);
and (n1579,n1580,n1581);
xor (n1580,n1577,n1578);
or (n1581,n1582,n1585);
and (n1582,n1583,n1584);
xor (n1583,n1487,n1488);
and (n1584,n20,n31);
and (n1585,n1586,n1587);
xor (n1586,n1583,n1584);
or (n1587,n1588,n1591);
and (n1588,n1589,n1590);
xor (n1589,n1493,n1494);
and (n1590,n59,n31);
and (n1591,n1592,n1593);
xor (n1592,n1589,n1590);
or (n1593,n1594,n1597);
and (n1594,n1595,n1596);
xor (n1595,n1499,n1500);
and (n1596,n168,n31);
and (n1597,n1598,n1599);
xor (n1598,n1595,n1596);
or (n1599,n1600,n1603);
and (n1600,n1601,n1602);
xor (n1601,n1505,n1506);
and (n1602,n209,n31);
and (n1603,n1604,n1605);
xor (n1604,n1601,n1602);
or (n1605,n1606,n1609);
and (n1606,n1607,n1608);
xor (n1607,n1511,n1512);
and (n1608,n256,n31);
and (n1609,n1610,n1611);
xor (n1610,n1607,n1608);
or (n1611,n1612,n1615);
and (n1612,n1613,n1614);
xor (n1613,n1517,n1518);
and (n1614,n311,n31);
and (n1615,n1616,n1617);
xor (n1616,n1613,n1614);
or (n1617,n1618,n1621);
and (n1618,n1619,n1620);
xor (n1619,n1523,n1524);
and (n1620,n346,n31);
and (n1621,n1622,n1623);
xor (n1622,n1619,n1620);
and (n1623,n1624,n1625);
xor (n1624,n1528,n1529);
not (n1625,n435);
and (n1626,n677,n22);
or (n1627,n1628,n1631);
and (n1628,n1629,n1630);
xor (n1629,n1538,n1539);
and (n1630,n111,n22);
and (n1631,n1632,n1633);
xor (n1632,n1629,n1630);
or (n1633,n1634,n1637);
and (n1634,n1635,n1636);
xor (n1635,n1544,n1545);
and (n1636,n105,n22);
and (n1637,n1638,n1639);
xor (n1638,n1635,n1636);
or (n1639,n1640,n1643);
and (n1640,n1641,n1642);
xor (n1641,n1550,n1551);
and (n1642,n139,n22);
and (n1643,n1644,n1645);
xor (n1644,n1641,n1642);
or (n1645,n1646,n1649);
and (n1646,n1647,n1648);
xor (n1647,n1556,n1557);
and (n1648,n133,n22);
and (n1649,n1650,n1651);
xor (n1650,n1647,n1648);
or (n1651,n1652,n1655);
and (n1652,n1653,n1654);
xor (n1653,n1562,n1563);
and (n1654,n86,n22);
and (n1655,n1656,n1657);
xor (n1656,n1653,n1654);
or (n1657,n1658,n1660);
and (n1658,n1659,n869);
xor (n1659,n1568,n1569);
and (n1660,n1661,n1662);
xor (n1661,n1659,n869);
or (n1662,n1663,n1665);
and (n1663,n1664,n45);
xor (n1664,n1574,n1575);
and (n1665,n1666,n1667);
xor (n1666,n1664,n45);
or (n1667,n1668,n1671);
and (n1668,n1669,n1670);
xor (n1669,n1580,n1581);
and (n1670,n20,n22);
and (n1671,n1672,n1673);
xor (n1672,n1669,n1670);
or (n1673,n1674,n1677);
and (n1674,n1675,n1676);
xor (n1675,n1586,n1587);
and (n1676,n59,n22);
and (n1677,n1678,n1679);
xor (n1678,n1675,n1676);
or (n1679,n1680,n1682);
and (n1680,n1681,n201);
xor (n1681,n1592,n1593);
and (n1682,n1683,n1684);
xor (n1683,n1681,n201);
or (n1684,n1685,n1687);
and (n1685,n1686,n249);
xor (n1686,n1598,n1599);
and (n1687,n1688,n1689);
xor (n1688,n1686,n249);
or (n1689,n1690,n1692);
and (n1690,n1691,n304);
xor (n1691,n1604,n1605);
and (n1692,n1693,n1694);
xor (n1693,n1691,n304);
or (n1694,n1695,n1698);
and (n1695,n1696,n1697);
xor (n1696,n1610,n1611);
and (n1697,n311,n22);
and (n1698,n1699,n1700);
xor (n1699,n1696,n1697);
or (n1700,n1701,n1704);
and (n1701,n1702,n1703);
xor (n1702,n1616,n1617);
and (n1703,n346,n22);
and (n1704,n1705,n1706);
xor (n1705,n1702,n1703);
and (n1706,n1707,n1708);
xor (n1707,n1622,n1623);
and (n1708,n376,n22);
or (n1709,n1710,n1713);
and (n1710,n1711,n1712);
xor (n1711,n1632,n1633);
and (n1712,n105,n52);
and (n1713,n1714,n1715);
xor (n1714,n1711,n1712);
or (n1715,n1716,n1719);
and (n1716,n1717,n1718);
xor (n1717,n1638,n1639);
and (n1718,n139,n52);
and (n1719,n1720,n1721);
xor (n1720,n1717,n1718);
or (n1721,n1722,n1725);
and (n1722,n1723,n1724);
xor (n1723,n1644,n1645);
and (n1724,n133,n52);
and (n1725,n1726,n1727);
xor (n1726,n1723,n1724);
or (n1727,n1728,n1731);
and (n1728,n1729,n1730);
xor (n1729,n1650,n1651);
and (n1730,n86,n52);
and (n1731,n1732,n1733);
xor (n1732,n1729,n1730);
or (n1733,n1734,n1737);
and (n1734,n1735,n1736);
xor (n1735,n1656,n1657);
and (n1736,n80,n52);
and (n1737,n1738,n1739);
xor (n1738,n1735,n1736);
or (n1739,n1740,n1743);
and (n1740,n1741,n1742);
xor (n1741,n1661,n1662);
and (n1742,n46,n52);
and (n1743,n1744,n1745);
xor (n1744,n1741,n1742);
or (n1745,n1746,n1749);
and (n1746,n1747,n1748);
xor (n1747,n1666,n1667);
and (n1748,n20,n52);
and (n1749,n1750,n1751);
xor (n1750,n1747,n1748);
or (n1751,n1752,n1755);
and (n1752,n1753,n1754);
xor (n1753,n1672,n1673);
and (n1754,n59,n52);
and (n1755,n1756,n1757);
xor (n1756,n1753,n1754);
or (n1757,n1758,n1761);
and (n1758,n1759,n1760);
xor (n1759,n1678,n1679);
and (n1760,n168,n52);
and (n1761,n1762,n1763);
xor (n1762,n1759,n1760);
or (n1763,n1764,n1767);
and (n1764,n1765,n1766);
xor (n1765,n1683,n1684);
and (n1766,n209,n52);
and (n1767,n1768,n1769);
xor (n1768,n1765,n1766);
or (n1769,n1770,n1773);
and (n1770,n1771,n1772);
xor (n1771,n1688,n1689);
and (n1772,n256,n52);
and (n1773,n1774,n1775);
xor (n1774,n1771,n1772);
or (n1775,n1776,n1779);
and (n1776,n1777,n1778);
xor (n1777,n1693,n1694);
and (n1778,n311,n52);
and (n1779,n1780,n1781);
xor (n1780,n1777,n1778);
or (n1781,n1782,n1785);
and (n1782,n1783,n1784);
xor (n1783,n1699,n1700);
and (n1784,n346,n52);
and (n1785,n1786,n1787);
xor (n1786,n1783,n1784);
and (n1787,n1788,n1789);
xor (n1788,n1705,n1706);
and (n1789,n376,n52);
or (n1790,n1791,n1793);
and (n1791,n1792,n1718);
xor (n1792,n1714,n1715);
and (n1793,n1794,n1795);
xor (n1794,n1792,n1718);
or (n1795,n1796,n1798);
and (n1796,n1797,n1724);
xor (n1797,n1720,n1721);
and (n1798,n1799,n1800);
xor (n1799,n1797,n1724);
or (n1800,n1801,n1803);
and (n1801,n1802,n1730);
xor (n1802,n1726,n1727);
and (n1803,n1804,n1805);
xor (n1804,n1802,n1730);
or (n1805,n1806,n1808);
and (n1806,n1807,n1736);
xor (n1807,n1732,n1733);
and (n1808,n1809,n1810);
xor (n1809,n1807,n1736);
or (n1810,n1811,n1813);
and (n1811,n1812,n1742);
xor (n1812,n1738,n1739);
and (n1813,n1814,n1815);
xor (n1814,n1812,n1742);
or (n1815,n1816,n1818);
and (n1816,n1817,n1748);
xor (n1817,n1744,n1745);
and (n1818,n1819,n1820);
xor (n1819,n1817,n1748);
or (n1820,n1821,n1823);
and (n1821,n1822,n1754);
xor (n1822,n1750,n1751);
and (n1823,n1824,n1825);
xor (n1824,n1822,n1754);
or (n1825,n1826,n1828);
and (n1826,n1827,n1760);
xor (n1827,n1756,n1757);
and (n1828,n1829,n1830);
xor (n1829,n1827,n1760);
or (n1830,n1831,n1833);
and (n1831,n1832,n1766);
xor (n1832,n1762,n1763);
and (n1833,n1834,n1835);
xor (n1834,n1832,n1766);
or (n1835,n1836,n1838);
and (n1836,n1837,n1772);
xor (n1837,n1768,n1769);
and (n1838,n1839,n1840);
xor (n1839,n1837,n1772);
or (n1840,n1841,n1843);
and (n1841,n1842,n1778);
xor (n1842,n1774,n1775);
and (n1843,n1844,n1845);
xor (n1844,n1842,n1778);
or (n1845,n1846,n1848);
and (n1846,n1847,n1784);
xor (n1847,n1780,n1781);
and (n1848,n1849,n1850);
xor (n1849,n1847,n1784);
and (n1850,n1851,n1789);
xor (n1851,n1786,n1787);
or (n1852,n1853,n1855);
and (n1853,n1854,n1724);
xor (n1854,n1794,n1795);
and (n1855,n1856,n1857);
xor (n1856,n1854,n1724);
or (n1857,n1858,n1860);
and (n1858,n1859,n1730);
xor (n1859,n1799,n1800);
and (n1860,n1861,n1862);
xor (n1861,n1859,n1730);
or (n1862,n1863,n1865);
and (n1863,n1864,n1736);
xor (n1864,n1804,n1805);
and (n1865,n1866,n1867);
xor (n1866,n1864,n1736);
or (n1867,n1868,n1870);
and (n1868,n1869,n1742);
xor (n1869,n1809,n1810);
and (n1870,n1871,n1872);
xor (n1871,n1869,n1742);
or (n1872,n1873,n1875);
and (n1873,n1874,n1748);
xor (n1874,n1814,n1815);
and (n1875,n1876,n1877);
xor (n1876,n1874,n1748);
or (n1877,n1878,n1880);
and (n1878,n1879,n1754);
xor (n1879,n1819,n1820);
and (n1880,n1881,n1882);
xor (n1881,n1879,n1754);
or (n1882,n1883,n1885);
and (n1883,n1884,n1760);
xor (n1884,n1824,n1825);
and (n1885,n1886,n1887);
xor (n1886,n1884,n1760);
or (n1887,n1888,n1890);
and (n1888,n1889,n1766);
xor (n1889,n1829,n1830);
and (n1890,n1891,n1892);
xor (n1891,n1889,n1766);
or (n1892,n1893,n1895);
and (n1893,n1894,n1772);
xor (n1894,n1834,n1835);
and (n1895,n1896,n1897);
xor (n1896,n1894,n1772);
or (n1897,n1898,n1900);
and (n1898,n1899,n1778);
xor (n1899,n1839,n1840);
and (n1900,n1901,n1902);
xor (n1901,n1899,n1778);
or (n1902,n1903,n1905);
and (n1903,n1904,n1784);
xor (n1904,n1844,n1845);
and (n1905,n1906,n1907);
xor (n1906,n1904,n1784);
and (n1907,n1908,n1789);
xor (n1908,n1849,n1850);
or (n1909,n1910,n1912);
and (n1910,n1911,n1730);
xor (n1911,n1856,n1857);
and (n1912,n1913,n1914);
xor (n1913,n1911,n1730);
or (n1914,n1915,n1917);
and (n1915,n1916,n1736);
xor (n1916,n1861,n1862);
and (n1917,n1918,n1919);
xor (n1918,n1916,n1736);
or (n1919,n1920,n1922);
and (n1920,n1921,n1742);
xor (n1921,n1866,n1867);
and (n1922,n1923,n1924);
xor (n1923,n1921,n1742);
or (n1924,n1925,n1927);
and (n1925,n1926,n1748);
xor (n1926,n1871,n1872);
and (n1927,n1928,n1929);
xor (n1928,n1926,n1748);
or (n1929,n1930,n1932);
and (n1930,n1931,n1754);
xor (n1931,n1876,n1877);
and (n1932,n1933,n1934);
xor (n1933,n1931,n1754);
or (n1934,n1935,n1937);
and (n1935,n1936,n1760);
xor (n1936,n1881,n1882);
and (n1937,n1938,n1939);
xor (n1938,n1936,n1760);
or (n1939,n1940,n1942);
and (n1940,n1941,n1766);
xor (n1941,n1886,n1887);
and (n1942,n1943,n1944);
xor (n1943,n1941,n1766);
or (n1944,n1945,n1947);
and (n1945,n1946,n1772);
xor (n1946,n1891,n1892);
and (n1947,n1948,n1949);
xor (n1948,n1946,n1772);
or (n1949,n1950,n1952);
and (n1950,n1951,n1778);
xor (n1951,n1896,n1897);
and (n1952,n1953,n1954);
xor (n1953,n1951,n1778);
or (n1954,n1955,n1957);
and (n1955,n1956,n1784);
xor (n1956,n1901,n1902);
and (n1957,n1958,n1959);
xor (n1958,n1956,n1784);
and (n1959,n1960,n1789);
xor (n1960,n1906,n1907);
or (n1961,n1962,n1964);
and (n1962,n1963,n1736);
xor (n1963,n1913,n1914);
and (n1964,n1965,n1966);
xor (n1965,n1963,n1736);
or (n1966,n1967,n1969);
and (n1967,n1968,n1742);
xor (n1968,n1918,n1919);
and (n1969,n1970,n1971);
xor (n1970,n1968,n1742);
or (n1971,n1972,n1974);
and (n1972,n1973,n1748);
xor (n1973,n1923,n1924);
and (n1974,n1975,n1976);
xor (n1975,n1973,n1748);
or (n1976,n1977,n1979);
and (n1977,n1978,n1754);
xor (n1978,n1928,n1929);
and (n1979,n1980,n1981);
xor (n1980,n1978,n1754);
or (n1981,n1982,n1984);
and (n1982,n1983,n1760);
xor (n1983,n1933,n1934);
and (n1984,n1985,n1986);
xor (n1985,n1983,n1760);
or (n1986,n1987,n1989);
and (n1987,n1988,n1766);
xor (n1988,n1938,n1939);
and (n1989,n1990,n1991);
xor (n1990,n1988,n1766);
or (n1991,n1992,n1994);
and (n1992,n1993,n1772);
xor (n1993,n1943,n1944);
and (n1994,n1995,n1996);
xor (n1995,n1993,n1772);
or (n1996,n1997,n1999);
and (n1997,n1998,n1778);
xor (n1998,n1948,n1949);
and (n1999,n2000,n2001);
xor (n2000,n1998,n1778);
or (n2001,n2002,n2004);
and (n2002,n2003,n1784);
xor (n2003,n1953,n1954);
and (n2004,n2005,n2006);
xor (n2005,n2003,n1784);
and (n2006,n2007,n1789);
xor (n2007,n1958,n1959);
or (n2008,n2009,n2011);
and (n2009,n2010,n1742);
xor (n2010,n1965,n1966);
and (n2011,n2012,n2013);
xor (n2012,n2010,n1742);
or (n2013,n2014,n2016);
and (n2014,n2015,n1748);
xor (n2015,n1970,n1971);
and (n2016,n2017,n2018);
xor (n2017,n2015,n1748);
or (n2018,n2019,n2021);
and (n2019,n2020,n1754);
xor (n2020,n1975,n1976);
and (n2021,n2022,n2023);
xor (n2022,n2020,n1754);
or (n2023,n2024,n2026);
and (n2024,n2025,n1760);
xor (n2025,n1980,n1981);
and (n2026,n2027,n2028);
xor (n2027,n2025,n1760);
or (n2028,n2029,n2031);
and (n2029,n2030,n1766);
xor (n2030,n1985,n1986);
and (n2031,n2032,n2033);
xor (n2032,n2030,n1766);
or (n2033,n2034,n2036);
and (n2034,n2035,n1772);
xor (n2035,n1990,n1991);
and (n2036,n2037,n2038);
xor (n2037,n2035,n1772);
or (n2038,n2039,n2041);
and (n2039,n2040,n1778);
xor (n2040,n1995,n1996);
and (n2041,n2042,n2043);
xor (n2042,n2040,n1778);
or (n2043,n2044,n2046);
and (n2044,n2045,n1784);
xor (n2045,n2000,n2001);
and (n2046,n2047,n2048);
xor (n2047,n2045,n1784);
and (n2048,n2049,n1789);
xor (n2049,n2005,n2006);
or (n2050,n2051,n2053);
and (n2051,n2052,n1748);
xor (n2052,n2012,n2013);
and (n2053,n2054,n2055);
xor (n2054,n2052,n1748);
or (n2055,n2056,n2058);
and (n2056,n2057,n1754);
xor (n2057,n2017,n2018);
and (n2058,n2059,n2060);
xor (n2059,n2057,n1754);
or (n2060,n2061,n2063);
and (n2061,n2062,n1760);
xor (n2062,n2022,n2023);
and (n2063,n2064,n2065);
xor (n2064,n2062,n1760);
or (n2065,n2066,n2068);
and (n2066,n2067,n1766);
xor (n2067,n2027,n2028);
and (n2068,n2069,n2070);
xor (n2069,n2067,n1766);
or (n2070,n2071,n2073);
and (n2071,n2072,n1772);
xor (n2072,n2032,n2033);
and (n2073,n2074,n2075);
xor (n2074,n2072,n1772);
or (n2075,n2076,n2078);
and (n2076,n2077,n1778);
xor (n2077,n2037,n2038);
and (n2078,n2079,n2080);
xor (n2079,n2077,n1778);
or (n2080,n2081,n2083);
and (n2081,n2082,n1784);
xor (n2082,n2042,n2043);
and (n2083,n2084,n2085);
xor (n2084,n2082,n1784);
and (n2085,n2086,n1789);
xor (n2086,n2047,n2048);
or (n2087,n2088,n2090);
and (n2088,n2089,n1754);
xor (n2089,n2054,n2055);
and (n2090,n2091,n2092);
xor (n2091,n2089,n1754);
or (n2092,n2093,n2095);
and (n2093,n2094,n1760);
xor (n2094,n2059,n2060);
and (n2095,n2096,n2097);
xor (n2096,n2094,n1760);
or (n2097,n2098,n2100);
and (n2098,n2099,n1766);
xor (n2099,n2064,n2065);
and (n2100,n2101,n2102);
xor (n2101,n2099,n1766);
or (n2102,n2103,n2105);
and (n2103,n2104,n1772);
xor (n2104,n2069,n2070);
and (n2105,n2106,n2107);
xor (n2106,n2104,n1772);
or (n2107,n2108,n2110);
and (n2108,n2109,n1778);
xor (n2109,n2074,n2075);
and (n2110,n2111,n2112);
xor (n2111,n2109,n1778);
or (n2112,n2113,n2115);
and (n2113,n2114,n1784);
xor (n2114,n2079,n2080);
and (n2115,n2116,n2117);
xor (n2116,n2114,n1784);
and (n2117,n2118,n1789);
xor (n2118,n2084,n2085);
or (n2119,n2120,n2122);
and (n2120,n2121,n1760);
xor (n2121,n2091,n2092);
and (n2122,n2123,n2124);
xor (n2123,n2121,n1760);
or (n2124,n2125,n2127);
and (n2125,n2126,n1766);
xor (n2126,n2096,n2097);
and (n2127,n2128,n2129);
xor (n2128,n2126,n1766);
or (n2129,n2130,n2132);
and (n2130,n2131,n1772);
xor (n2131,n2101,n2102);
and (n2132,n2133,n2134);
xor (n2133,n2131,n1772);
or (n2134,n2135,n2137);
and (n2135,n2136,n1778);
xor (n2136,n2106,n2107);
and (n2137,n2138,n2139);
xor (n2138,n2136,n1778);
or (n2139,n2140,n2142);
and (n2140,n2141,n1784);
xor (n2141,n2111,n2112);
and (n2142,n2143,n2144);
xor (n2143,n2141,n1784);
and (n2144,n2145,n1789);
xor (n2145,n2116,n2117);
or (n2146,n2147,n2149);
and (n2147,n2148,n1766);
xor (n2148,n2123,n2124);
and (n2149,n2150,n2151);
xor (n2150,n2148,n1766);
or (n2151,n2152,n2154);
and (n2152,n2153,n1772);
xor (n2153,n2128,n2129);
and (n2154,n2155,n2156);
xor (n2155,n2153,n1772);
or (n2156,n2157,n2159);
and (n2157,n2158,n1778);
xor (n2158,n2133,n2134);
and (n2159,n2160,n2161);
xor (n2160,n2158,n1778);
or (n2161,n2162,n2164);
and (n2162,n2163,n1784);
xor (n2163,n2138,n2139);
and (n2164,n2165,n2166);
xor (n2165,n2163,n1784);
and (n2166,n2167,n1789);
xor (n2167,n2143,n2144);
or (n2168,n2169,n2171);
and (n2169,n2170,n1772);
xor (n2170,n2150,n2151);
and (n2171,n2172,n2173);
xor (n2172,n2170,n1772);
or (n2173,n2174,n2176);
and (n2174,n2175,n1778);
xor (n2175,n2155,n2156);
and (n2176,n2177,n2178);
xor (n2177,n2175,n1778);
or (n2178,n2179,n2181);
and (n2179,n2180,n1784);
xor (n2180,n2160,n2161);
and (n2181,n2182,n2183);
xor (n2182,n2180,n1784);
and (n2183,n2184,n1789);
xor (n2184,n2165,n2166);
or (n2185,n2186,n2188);
and (n2186,n2187,n1778);
xor (n2187,n2172,n2173);
and (n2188,n2189,n2190);
xor (n2189,n2187,n1778);
or (n2190,n2191,n2193);
and (n2191,n2192,n1784);
xor (n2192,n2177,n2178);
and (n2193,n2194,n2195);
xor (n2194,n2192,n1784);
and (n2195,n2196,n1789);
xor (n2196,n2182,n2183);
or (n2197,n2198,n2200);
and (n2198,n2199,n1784);
xor (n2199,n2189,n2190);
and (n2200,n2201,n2202);
xor (n2201,n2199,n1784);
and (n2202,n2203,n1789);
xor (n2203,n2194,n2195);
and (n2204,n2205,n1789);
xor (n2205,n2201,n2202);
xor (n2206,n2086,n1789);
endmodule
