module top (out,n23,n24,n28,n30,n37,n44,n51,n58,n65
        ,n72,n79,n86,n93,n99,n101,n168,n235,n302,n369
        ,n436,n503,n570,n635,n694,n768,n769,n773,n775,n782
        ,n789,n796,n803,n810,n817,n824,n831,n838,n844,n846
        ,n913,n980,n1047,n1114,n1181,n1248,n1315,n1380,n1439,n1491);
output out;
input n23;
input n24;
input n28;
input n30;
input n37;
input n44;
input n51;
input n58;
input n65;
input n72;
input n79;
input n86;
input n93;
input n99;
input n101;
input n168;
input n235;
input n302;
input n369;
input n436;
input n503;
input n570;
input n635;
input n694;
input n768;
input n769;
input n773;
input n775;
input n782;
input n789;
input n796;
input n803;
input n810;
input n817;
input n824;
input n831;
input n838;
input n844;
input n846;
input n913;
input n980;
input n1047;
input n1114;
input n1181;
input n1248;
input n1315;
input n1380;
input n1439;
input n1491;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n25;
wire n26;
wire n27;
wire n29;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n100;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n770;
wire n771;
wire n772;
wire n774;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n845;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
xor (out,n0,n1492);
wire s0n0,s1n0,notn0;
or (n0,s0n0,s1n0);
not(notn0,n1491);
and (s0n0,notn0,n1);
and (s1n0,n1491,n746);
xor (n1,n2,n695);
xor (n2,n3,n693);
xor (n3,n4,n636);
xor (n4,n5,n634);
xor (n5,n6,n571);
xor (n6,n7,n569);
or (n7,n8,n504);
and (n8,n9,n502);
or (n9,n10,n437);
and (n10,n11,n435);
or (n11,n12,n370);
and (n12,n13,n368);
or (n13,n14,n303);
and (n14,n15,n301);
or (n15,n16,n236);
and (n16,n17,n234);
or (n17,n18,n169);
and (n18,n19,n167);
or (n19,n20,n102);
and (n20,n21,n100);
and (n21,n22,n25);
and (n22,n23,n24);
or (n25,n26,n31);
and (n26,n27,n29);
and (n27,n23,n28);
and (n29,n30,n24);
and (n31,n32,n33);
xor (n32,n27,n29);
or (n33,n34,n38);
and (n34,n35,n36);
and (n35,n30,n28);
and (n36,n37,n24);
and (n38,n39,n40);
xor (n39,n35,n36);
or (n40,n41,n45);
and (n41,n42,n43);
and (n42,n37,n28);
and (n43,n44,n24);
and (n45,n46,n47);
xor (n46,n42,n43);
or (n47,n48,n52);
and (n48,n49,n50);
and (n49,n44,n28);
and (n50,n51,n24);
and (n52,n53,n54);
xor (n53,n49,n50);
or (n54,n55,n59);
and (n55,n56,n57);
and (n56,n51,n28);
and (n57,n58,n24);
and (n59,n60,n61);
xor (n60,n56,n57);
or (n61,n62,n66);
and (n62,n63,n64);
and (n63,n58,n28);
and (n64,n65,n24);
and (n66,n67,n68);
xor (n67,n63,n64);
or (n68,n69,n73);
and (n69,n70,n71);
and (n70,n65,n28);
and (n71,n72,n24);
and (n73,n74,n75);
xor (n74,n70,n71);
or (n75,n76,n80);
and (n76,n77,n78);
and (n77,n72,n28);
and (n78,n79,n24);
and (n80,n81,n82);
xor (n81,n77,n78);
or (n82,n83,n87);
and (n83,n84,n85);
and (n84,n79,n28);
and (n85,n86,n24);
and (n87,n88,n89);
xor (n88,n84,n85);
or (n89,n90,n94);
and (n90,n91,n92);
and (n91,n86,n28);
and (n92,n93,n24);
and (n94,n95,n96);
xor (n95,n91,n92);
and (n96,n97,n98);
and (n97,n93,n28);
and (n98,n99,n24);
and (n100,n23,n101);
and (n102,n103,n104);
xor (n103,n21,n100);
or (n104,n105,n108);
and (n105,n106,n107);
xor (n106,n22,n25);
and (n107,n30,n101);
and (n108,n109,n110);
xor (n109,n106,n107);
or (n110,n111,n114);
and (n111,n112,n113);
xor (n112,n32,n33);
and (n113,n37,n101);
and (n114,n115,n116);
xor (n115,n112,n113);
or (n116,n117,n120);
and (n117,n118,n119);
xor (n118,n39,n40);
and (n119,n44,n101);
and (n120,n121,n122);
xor (n121,n118,n119);
or (n122,n123,n126);
and (n123,n124,n125);
xor (n124,n46,n47);
and (n125,n51,n101);
and (n126,n127,n128);
xor (n127,n124,n125);
or (n128,n129,n132);
and (n129,n130,n131);
xor (n130,n53,n54);
and (n131,n58,n101);
and (n132,n133,n134);
xor (n133,n130,n131);
or (n134,n135,n138);
and (n135,n136,n137);
xor (n136,n60,n61);
and (n137,n65,n101);
and (n138,n139,n140);
xor (n139,n136,n137);
or (n140,n141,n144);
and (n141,n142,n143);
xor (n142,n67,n68);
and (n143,n72,n101);
and (n144,n145,n146);
xor (n145,n142,n143);
or (n146,n147,n150);
and (n147,n148,n149);
xor (n148,n74,n75);
and (n149,n79,n101);
and (n150,n151,n152);
xor (n151,n148,n149);
or (n152,n153,n156);
and (n153,n154,n155);
xor (n154,n81,n82);
and (n155,n86,n101);
and (n156,n157,n158);
xor (n157,n154,n155);
or (n158,n159,n162);
and (n159,n160,n161);
xor (n160,n88,n89);
and (n161,n93,n101);
and (n162,n163,n164);
xor (n163,n160,n161);
and (n164,n165,n166);
xor (n165,n95,n96);
and (n166,n99,n101);
and (n167,n23,n168);
and (n169,n170,n171);
xor (n170,n19,n167);
or (n171,n172,n175);
and (n172,n173,n174);
xor (n173,n103,n104);
and (n174,n30,n168);
and (n175,n176,n177);
xor (n176,n173,n174);
or (n177,n178,n181);
and (n178,n179,n180);
xor (n179,n109,n110);
and (n180,n37,n168);
and (n181,n182,n183);
xor (n182,n179,n180);
or (n183,n184,n187);
and (n184,n185,n186);
xor (n185,n115,n116);
and (n186,n44,n168);
and (n187,n188,n189);
xor (n188,n185,n186);
or (n189,n190,n193);
and (n190,n191,n192);
xor (n191,n121,n122);
and (n192,n51,n168);
and (n193,n194,n195);
xor (n194,n191,n192);
or (n195,n196,n199);
and (n196,n197,n198);
xor (n197,n127,n128);
and (n198,n58,n168);
and (n199,n200,n201);
xor (n200,n197,n198);
or (n201,n202,n205);
and (n202,n203,n204);
xor (n203,n133,n134);
and (n204,n65,n168);
and (n205,n206,n207);
xor (n206,n203,n204);
or (n207,n208,n211);
and (n208,n209,n210);
xor (n209,n139,n140);
and (n210,n72,n168);
and (n211,n212,n213);
xor (n212,n209,n210);
or (n213,n214,n217);
and (n214,n215,n216);
xor (n215,n145,n146);
and (n216,n79,n168);
and (n217,n218,n219);
xor (n218,n215,n216);
or (n219,n220,n223);
and (n220,n221,n222);
xor (n221,n151,n152);
and (n222,n86,n168);
and (n223,n224,n225);
xor (n224,n221,n222);
or (n225,n226,n229);
and (n226,n227,n228);
xor (n227,n157,n158);
and (n228,n93,n168);
and (n229,n230,n231);
xor (n230,n227,n228);
and (n231,n232,n233);
xor (n232,n163,n164);
and (n233,n99,n168);
and (n234,n23,n235);
and (n236,n237,n238);
xor (n237,n17,n234);
or (n238,n239,n242);
and (n239,n240,n241);
xor (n240,n170,n171);
and (n241,n30,n235);
and (n242,n243,n244);
xor (n243,n240,n241);
or (n244,n245,n248);
and (n245,n246,n247);
xor (n246,n176,n177);
and (n247,n37,n235);
and (n248,n249,n250);
xor (n249,n246,n247);
or (n250,n251,n254);
and (n251,n252,n253);
xor (n252,n182,n183);
and (n253,n44,n235);
and (n254,n255,n256);
xor (n255,n252,n253);
or (n256,n257,n260);
and (n257,n258,n259);
xor (n258,n188,n189);
and (n259,n51,n235);
and (n260,n261,n262);
xor (n261,n258,n259);
or (n262,n263,n266);
and (n263,n264,n265);
xor (n264,n194,n195);
and (n265,n58,n235);
and (n266,n267,n268);
xor (n267,n264,n265);
or (n268,n269,n272);
and (n269,n270,n271);
xor (n270,n200,n201);
and (n271,n65,n235);
and (n272,n273,n274);
xor (n273,n270,n271);
or (n274,n275,n278);
and (n275,n276,n277);
xor (n276,n206,n207);
and (n277,n72,n235);
and (n278,n279,n280);
xor (n279,n276,n277);
or (n280,n281,n284);
and (n281,n282,n283);
xor (n282,n212,n213);
and (n283,n79,n235);
and (n284,n285,n286);
xor (n285,n282,n283);
or (n286,n287,n290);
and (n287,n288,n289);
xor (n288,n218,n219);
and (n289,n86,n235);
and (n290,n291,n292);
xor (n291,n288,n289);
or (n292,n293,n296);
and (n293,n294,n295);
xor (n294,n224,n225);
and (n295,n93,n235);
and (n296,n297,n298);
xor (n297,n294,n295);
and (n298,n299,n300);
xor (n299,n230,n231);
and (n300,n99,n235);
and (n301,n23,n302);
and (n303,n304,n305);
xor (n304,n15,n301);
or (n305,n306,n309);
and (n306,n307,n308);
xor (n307,n237,n238);
and (n308,n30,n302);
and (n309,n310,n311);
xor (n310,n307,n308);
or (n311,n312,n315);
and (n312,n313,n314);
xor (n313,n243,n244);
and (n314,n37,n302);
and (n315,n316,n317);
xor (n316,n313,n314);
or (n317,n318,n321);
and (n318,n319,n320);
xor (n319,n249,n250);
and (n320,n44,n302);
and (n321,n322,n323);
xor (n322,n319,n320);
or (n323,n324,n327);
and (n324,n325,n326);
xor (n325,n255,n256);
and (n326,n51,n302);
and (n327,n328,n329);
xor (n328,n325,n326);
or (n329,n330,n333);
and (n330,n331,n332);
xor (n331,n261,n262);
and (n332,n58,n302);
and (n333,n334,n335);
xor (n334,n331,n332);
or (n335,n336,n339);
and (n336,n337,n338);
xor (n337,n267,n268);
and (n338,n65,n302);
and (n339,n340,n341);
xor (n340,n337,n338);
or (n341,n342,n345);
and (n342,n343,n344);
xor (n343,n273,n274);
and (n344,n72,n302);
and (n345,n346,n347);
xor (n346,n343,n344);
or (n347,n348,n351);
and (n348,n349,n350);
xor (n349,n279,n280);
and (n350,n79,n302);
and (n351,n352,n353);
xor (n352,n349,n350);
or (n353,n354,n357);
and (n354,n355,n356);
xor (n355,n285,n286);
and (n356,n86,n302);
and (n357,n358,n359);
xor (n358,n355,n356);
or (n359,n360,n363);
and (n360,n361,n362);
xor (n361,n291,n292);
and (n362,n93,n302);
and (n363,n364,n365);
xor (n364,n361,n362);
and (n365,n366,n367);
xor (n366,n297,n298);
and (n367,n99,n302);
and (n368,n23,n369);
and (n370,n371,n372);
xor (n371,n13,n368);
or (n372,n373,n376);
and (n373,n374,n375);
xor (n374,n304,n305);
and (n375,n30,n369);
and (n376,n377,n378);
xor (n377,n374,n375);
or (n378,n379,n382);
and (n379,n380,n381);
xor (n380,n310,n311);
and (n381,n37,n369);
and (n382,n383,n384);
xor (n383,n380,n381);
or (n384,n385,n388);
and (n385,n386,n387);
xor (n386,n316,n317);
and (n387,n44,n369);
and (n388,n389,n390);
xor (n389,n386,n387);
or (n390,n391,n394);
and (n391,n392,n393);
xor (n392,n322,n323);
and (n393,n51,n369);
and (n394,n395,n396);
xor (n395,n392,n393);
or (n396,n397,n400);
and (n397,n398,n399);
xor (n398,n328,n329);
and (n399,n58,n369);
and (n400,n401,n402);
xor (n401,n398,n399);
or (n402,n403,n406);
and (n403,n404,n405);
xor (n404,n334,n335);
and (n405,n65,n369);
and (n406,n407,n408);
xor (n407,n404,n405);
or (n408,n409,n412);
and (n409,n410,n411);
xor (n410,n340,n341);
and (n411,n72,n369);
and (n412,n413,n414);
xor (n413,n410,n411);
or (n414,n415,n418);
and (n415,n416,n417);
xor (n416,n346,n347);
and (n417,n79,n369);
and (n418,n419,n420);
xor (n419,n416,n417);
or (n420,n421,n424);
and (n421,n422,n423);
xor (n422,n352,n353);
and (n423,n86,n369);
and (n424,n425,n426);
xor (n425,n422,n423);
or (n426,n427,n430);
and (n427,n428,n429);
xor (n428,n358,n359);
and (n429,n93,n369);
and (n430,n431,n432);
xor (n431,n428,n429);
and (n432,n433,n434);
xor (n433,n364,n365);
and (n434,n99,n369);
and (n435,n23,n436);
and (n437,n438,n439);
xor (n438,n11,n435);
or (n439,n440,n443);
and (n440,n441,n442);
xor (n441,n371,n372);
and (n442,n30,n436);
and (n443,n444,n445);
xor (n444,n441,n442);
or (n445,n446,n449);
and (n446,n447,n448);
xor (n447,n377,n378);
and (n448,n37,n436);
and (n449,n450,n451);
xor (n450,n447,n448);
or (n451,n452,n455);
and (n452,n453,n454);
xor (n453,n383,n384);
and (n454,n44,n436);
and (n455,n456,n457);
xor (n456,n453,n454);
or (n457,n458,n461);
and (n458,n459,n460);
xor (n459,n389,n390);
and (n460,n51,n436);
and (n461,n462,n463);
xor (n462,n459,n460);
or (n463,n464,n467);
and (n464,n465,n466);
xor (n465,n395,n396);
and (n466,n58,n436);
and (n467,n468,n469);
xor (n468,n465,n466);
or (n469,n470,n473);
and (n470,n471,n472);
xor (n471,n401,n402);
and (n472,n65,n436);
and (n473,n474,n475);
xor (n474,n471,n472);
or (n475,n476,n479);
and (n476,n477,n478);
xor (n477,n407,n408);
and (n478,n72,n436);
and (n479,n480,n481);
xor (n480,n477,n478);
or (n481,n482,n485);
and (n482,n483,n484);
xor (n483,n413,n414);
and (n484,n79,n436);
and (n485,n486,n487);
xor (n486,n483,n484);
or (n487,n488,n491);
and (n488,n489,n490);
xor (n489,n419,n420);
and (n490,n86,n436);
and (n491,n492,n493);
xor (n492,n489,n490);
or (n493,n494,n497);
and (n494,n495,n496);
xor (n495,n425,n426);
and (n496,n93,n436);
and (n497,n498,n499);
xor (n498,n495,n496);
and (n499,n500,n501);
xor (n500,n431,n432);
and (n501,n99,n436);
and (n502,n23,n503);
and (n504,n505,n506);
xor (n505,n9,n502);
or (n506,n507,n510);
and (n507,n508,n509);
xor (n508,n438,n439);
and (n509,n30,n503);
and (n510,n511,n512);
xor (n511,n508,n509);
or (n512,n513,n516);
and (n513,n514,n515);
xor (n514,n444,n445);
and (n515,n37,n503);
and (n516,n517,n518);
xor (n517,n514,n515);
or (n518,n519,n522);
and (n519,n520,n521);
xor (n520,n450,n451);
and (n521,n44,n503);
and (n522,n523,n524);
xor (n523,n520,n521);
or (n524,n525,n528);
and (n525,n526,n527);
xor (n526,n456,n457);
and (n527,n51,n503);
and (n528,n529,n530);
xor (n529,n526,n527);
or (n530,n531,n534);
and (n531,n532,n533);
xor (n532,n462,n463);
and (n533,n58,n503);
and (n534,n535,n536);
xor (n535,n532,n533);
or (n536,n537,n540);
and (n537,n538,n539);
xor (n538,n468,n469);
and (n539,n65,n503);
and (n540,n541,n542);
xor (n541,n538,n539);
or (n542,n543,n546);
and (n543,n544,n545);
xor (n544,n474,n475);
and (n545,n72,n503);
and (n546,n547,n548);
xor (n547,n544,n545);
or (n548,n549,n552);
and (n549,n550,n551);
xor (n550,n480,n481);
and (n551,n79,n503);
and (n552,n553,n554);
xor (n553,n550,n551);
or (n554,n555,n558);
and (n555,n556,n557);
xor (n556,n486,n487);
and (n557,n86,n503);
and (n558,n559,n560);
xor (n559,n556,n557);
or (n560,n561,n564);
and (n561,n562,n563);
xor (n562,n492,n493);
and (n563,n93,n503);
and (n564,n565,n566);
xor (n565,n562,n563);
and (n566,n567,n568);
xor (n567,n498,n499);
and (n568,n99,n503);
and (n569,n23,n570);
or (n571,n572,n575);
and (n572,n573,n574);
xor (n573,n505,n506);
and (n574,n30,n570);
and (n575,n576,n577);
xor (n576,n573,n574);
or (n577,n578,n581);
and (n578,n579,n580);
xor (n579,n511,n512);
and (n580,n37,n570);
and (n581,n582,n583);
xor (n582,n579,n580);
or (n583,n584,n587);
and (n584,n585,n586);
xor (n585,n517,n518);
and (n586,n44,n570);
and (n587,n588,n589);
xor (n588,n585,n586);
or (n589,n590,n593);
and (n590,n591,n592);
xor (n591,n523,n524);
and (n592,n51,n570);
and (n593,n594,n595);
xor (n594,n591,n592);
or (n595,n596,n599);
and (n596,n597,n598);
xor (n597,n529,n530);
and (n598,n58,n570);
and (n599,n600,n601);
xor (n600,n597,n598);
or (n601,n602,n605);
and (n602,n603,n604);
xor (n603,n535,n536);
and (n604,n65,n570);
and (n605,n606,n607);
xor (n606,n603,n604);
or (n607,n608,n611);
and (n608,n609,n610);
xor (n609,n541,n542);
and (n610,n72,n570);
and (n611,n612,n613);
xor (n612,n609,n610);
or (n613,n614,n617);
and (n614,n615,n616);
xor (n615,n547,n548);
and (n616,n79,n570);
and (n617,n618,n619);
xor (n618,n615,n616);
or (n619,n620,n623);
and (n620,n621,n622);
xor (n621,n553,n554);
and (n622,n86,n570);
and (n623,n624,n625);
xor (n624,n621,n622);
or (n625,n626,n629);
and (n626,n627,n628);
xor (n627,n559,n560);
and (n628,n93,n570);
and (n629,n630,n631);
xor (n630,n627,n628);
and (n631,n632,n633);
xor (n632,n565,n566);
and (n633,n99,n570);
and (n634,n30,n635);
or (n636,n637,n640);
and (n637,n638,n639);
xor (n638,n576,n577);
and (n639,n37,n635);
and (n640,n641,n642);
xor (n641,n638,n639);
or (n642,n643,n646);
and (n643,n644,n645);
xor (n644,n582,n583);
and (n645,n44,n635);
and (n646,n647,n648);
xor (n647,n644,n645);
or (n648,n649,n652);
and (n649,n650,n651);
xor (n650,n588,n589);
and (n651,n51,n635);
and (n652,n653,n654);
xor (n653,n650,n651);
or (n654,n655,n658);
and (n655,n656,n657);
xor (n656,n594,n595);
and (n657,n58,n635);
and (n658,n659,n660);
xor (n659,n656,n657);
or (n660,n661,n664);
and (n661,n662,n663);
xor (n662,n600,n601);
and (n663,n65,n635);
and (n664,n665,n666);
xor (n665,n662,n663);
or (n666,n667,n670);
and (n667,n668,n669);
xor (n668,n606,n607);
and (n669,n72,n635);
and (n670,n671,n672);
xor (n671,n668,n669);
or (n672,n673,n676);
and (n673,n674,n675);
xor (n674,n612,n613);
and (n675,n79,n635);
and (n676,n677,n678);
xor (n677,n674,n675);
or (n678,n679,n682);
and (n679,n680,n681);
xor (n680,n618,n619);
and (n681,n86,n635);
and (n682,n683,n684);
xor (n683,n680,n681);
or (n684,n685,n688);
and (n685,n686,n687);
xor (n686,n624,n625);
and (n687,n93,n635);
and (n688,n689,n690);
xor (n689,n686,n687);
and (n690,n691,n692);
xor (n691,n630,n631);
and (n692,n99,n635);
and (n693,n37,n694);
or (n695,n696,n699);
and (n696,n697,n698);
xor (n697,n641,n642);
and (n698,n44,n694);
and (n699,n700,n701);
xor (n700,n697,n698);
or (n701,n702,n705);
and (n702,n703,n704);
xor (n703,n647,n648);
and (n704,n51,n694);
and (n705,n706,n707);
xor (n706,n703,n704);
or (n707,n708,n711);
and (n708,n709,n710);
xor (n709,n653,n654);
and (n710,n58,n694);
and (n711,n712,n713);
xor (n712,n709,n710);
or (n713,n714,n717);
and (n714,n715,n716);
xor (n715,n659,n660);
and (n716,n65,n694);
and (n717,n718,n719);
xor (n718,n715,n716);
or (n719,n720,n723);
and (n720,n721,n722);
xor (n721,n665,n666);
and (n722,n72,n694);
and (n723,n724,n725);
xor (n724,n721,n722);
or (n725,n726,n729);
and (n726,n727,n728);
xor (n727,n671,n672);
and (n728,n79,n694);
and (n729,n730,n731);
xor (n730,n727,n728);
or (n731,n732,n735);
and (n732,n733,n734);
xor (n733,n677,n678);
and (n734,n86,n694);
and (n735,n736,n737);
xor (n736,n733,n734);
or (n737,n738,n741);
and (n738,n739,n740);
xor (n739,n683,n684);
and (n740,n93,n694);
and (n741,n742,n743);
xor (n742,n739,n740);
and (n743,n744,n745);
xor (n744,n689,n690);
and (n745,n99,n694);
xor (n746,n747,n1440);
xor (n747,n748,n1438);
xor (n748,n749,n1381);
xor (n749,n750,n1379);
xor (n750,n751,n1316);
xor (n751,n752,n1314);
or (n752,n753,n1249);
and (n753,n754,n1247);
or (n754,n755,n1182);
and (n755,n756,n1180);
or (n756,n757,n1115);
and (n757,n758,n1113);
or (n758,n759,n1048);
and (n759,n760,n1046);
or (n760,n761,n981);
and (n761,n762,n979);
or (n762,n763,n914);
and (n763,n764,n912);
or (n764,n765,n847);
and (n765,n766,n845);
and (n766,n767,n770);
and (n767,n768,n769);
or (n770,n771,n776);
and (n771,n772,n774);
and (n772,n768,n773);
and (n774,n775,n769);
and (n776,n777,n778);
xor (n777,n772,n774);
or (n778,n779,n783);
and (n779,n780,n781);
and (n780,n775,n773);
and (n781,n782,n769);
and (n783,n784,n785);
xor (n784,n780,n781);
or (n785,n786,n790);
and (n786,n787,n788);
and (n787,n782,n773);
and (n788,n789,n769);
and (n790,n791,n792);
xor (n791,n787,n788);
or (n792,n793,n797);
and (n793,n794,n795);
and (n794,n789,n773);
and (n795,n796,n769);
and (n797,n798,n799);
xor (n798,n794,n795);
or (n799,n800,n804);
and (n800,n801,n802);
and (n801,n796,n773);
and (n802,n803,n769);
and (n804,n805,n806);
xor (n805,n801,n802);
or (n806,n807,n811);
and (n807,n808,n809);
and (n808,n803,n773);
and (n809,n810,n769);
and (n811,n812,n813);
xor (n812,n808,n809);
or (n813,n814,n818);
and (n814,n815,n816);
and (n815,n810,n773);
and (n816,n817,n769);
and (n818,n819,n820);
xor (n819,n815,n816);
or (n820,n821,n825);
and (n821,n822,n823);
and (n822,n817,n773);
and (n823,n824,n769);
and (n825,n826,n827);
xor (n826,n822,n823);
or (n827,n828,n832);
and (n828,n829,n830);
and (n829,n824,n773);
and (n830,n831,n769);
and (n832,n833,n834);
xor (n833,n829,n830);
or (n834,n835,n839);
and (n835,n836,n837);
and (n836,n831,n773);
and (n837,n838,n769);
and (n839,n840,n841);
xor (n840,n836,n837);
and (n841,n842,n843);
and (n842,n838,n773);
and (n843,n844,n769);
and (n845,n768,n846);
and (n847,n848,n849);
xor (n848,n766,n845);
or (n849,n850,n853);
and (n850,n851,n852);
xor (n851,n767,n770);
and (n852,n775,n846);
and (n853,n854,n855);
xor (n854,n851,n852);
or (n855,n856,n859);
and (n856,n857,n858);
xor (n857,n777,n778);
and (n858,n782,n846);
and (n859,n860,n861);
xor (n860,n857,n858);
or (n861,n862,n865);
and (n862,n863,n864);
xor (n863,n784,n785);
and (n864,n789,n846);
and (n865,n866,n867);
xor (n866,n863,n864);
or (n867,n868,n871);
and (n868,n869,n870);
xor (n869,n791,n792);
and (n870,n796,n846);
and (n871,n872,n873);
xor (n872,n869,n870);
or (n873,n874,n877);
and (n874,n875,n876);
xor (n875,n798,n799);
and (n876,n803,n846);
and (n877,n878,n879);
xor (n878,n875,n876);
or (n879,n880,n883);
and (n880,n881,n882);
xor (n881,n805,n806);
and (n882,n810,n846);
and (n883,n884,n885);
xor (n884,n881,n882);
or (n885,n886,n889);
and (n886,n887,n888);
xor (n887,n812,n813);
and (n888,n817,n846);
and (n889,n890,n891);
xor (n890,n887,n888);
or (n891,n892,n895);
and (n892,n893,n894);
xor (n893,n819,n820);
and (n894,n824,n846);
and (n895,n896,n897);
xor (n896,n893,n894);
or (n897,n898,n901);
and (n898,n899,n900);
xor (n899,n826,n827);
and (n900,n831,n846);
and (n901,n902,n903);
xor (n902,n899,n900);
or (n903,n904,n907);
and (n904,n905,n906);
xor (n905,n833,n834);
and (n906,n838,n846);
and (n907,n908,n909);
xor (n908,n905,n906);
and (n909,n910,n911);
xor (n910,n840,n841);
and (n911,n844,n846);
and (n912,n768,n913);
and (n914,n915,n916);
xor (n915,n764,n912);
or (n916,n917,n920);
and (n917,n918,n919);
xor (n918,n848,n849);
and (n919,n775,n913);
and (n920,n921,n922);
xor (n921,n918,n919);
or (n922,n923,n926);
and (n923,n924,n925);
xor (n924,n854,n855);
and (n925,n782,n913);
and (n926,n927,n928);
xor (n927,n924,n925);
or (n928,n929,n932);
and (n929,n930,n931);
xor (n930,n860,n861);
and (n931,n789,n913);
and (n932,n933,n934);
xor (n933,n930,n931);
or (n934,n935,n938);
and (n935,n936,n937);
xor (n936,n866,n867);
and (n937,n796,n913);
and (n938,n939,n940);
xor (n939,n936,n937);
or (n940,n941,n944);
and (n941,n942,n943);
xor (n942,n872,n873);
and (n943,n803,n913);
and (n944,n945,n946);
xor (n945,n942,n943);
or (n946,n947,n950);
and (n947,n948,n949);
xor (n948,n878,n879);
and (n949,n810,n913);
and (n950,n951,n952);
xor (n951,n948,n949);
or (n952,n953,n956);
and (n953,n954,n955);
xor (n954,n884,n885);
and (n955,n817,n913);
and (n956,n957,n958);
xor (n957,n954,n955);
or (n958,n959,n962);
and (n959,n960,n961);
xor (n960,n890,n891);
and (n961,n824,n913);
and (n962,n963,n964);
xor (n963,n960,n961);
or (n964,n965,n968);
and (n965,n966,n967);
xor (n966,n896,n897);
and (n967,n831,n913);
and (n968,n969,n970);
xor (n969,n966,n967);
or (n970,n971,n974);
and (n971,n972,n973);
xor (n972,n902,n903);
and (n973,n838,n913);
and (n974,n975,n976);
xor (n975,n972,n973);
and (n976,n977,n978);
xor (n977,n908,n909);
and (n978,n844,n913);
and (n979,n768,n980);
and (n981,n982,n983);
xor (n982,n762,n979);
or (n983,n984,n987);
and (n984,n985,n986);
xor (n985,n915,n916);
and (n986,n775,n980);
and (n987,n988,n989);
xor (n988,n985,n986);
or (n989,n990,n993);
and (n990,n991,n992);
xor (n991,n921,n922);
and (n992,n782,n980);
and (n993,n994,n995);
xor (n994,n991,n992);
or (n995,n996,n999);
and (n996,n997,n998);
xor (n997,n927,n928);
and (n998,n789,n980);
and (n999,n1000,n1001);
xor (n1000,n997,n998);
or (n1001,n1002,n1005);
and (n1002,n1003,n1004);
xor (n1003,n933,n934);
and (n1004,n796,n980);
and (n1005,n1006,n1007);
xor (n1006,n1003,n1004);
or (n1007,n1008,n1011);
and (n1008,n1009,n1010);
xor (n1009,n939,n940);
and (n1010,n803,n980);
and (n1011,n1012,n1013);
xor (n1012,n1009,n1010);
or (n1013,n1014,n1017);
and (n1014,n1015,n1016);
xor (n1015,n945,n946);
and (n1016,n810,n980);
and (n1017,n1018,n1019);
xor (n1018,n1015,n1016);
or (n1019,n1020,n1023);
and (n1020,n1021,n1022);
xor (n1021,n951,n952);
and (n1022,n817,n980);
and (n1023,n1024,n1025);
xor (n1024,n1021,n1022);
or (n1025,n1026,n1029);
and (n1026,n1027,n1028);
xor (n1027,n957,n958);
and (n1028,n824,n980);
and (n1029,n1030,n1031);
xor (n1030,n1027,n1028);
or (n1031,n1032,n1035);
and (n1032,n1033,n1034);
xor (n1033,n963,n964);
and (n1034,n831,n980);
and (n1035,n1036,n1037);
xor (n1036,n1033,n1034);
or (n1037,n1038,n1041);
and (n1038,n1039,n1040);
xor (n1039,n969,n970);
and (n1040,n838,n980);
and (n1041,n1042,n1043);
xor (n1042,n1039,n1040);
and (n1043,n1044,n1045);
xor (n1044,n975,n976);
and (n1045,n844,n980);
and (n1046,n768,n1047);
and (n1048,n1049,n1050);
xor (n1049,n760,n1046);
or (n1050,n1051,n1054);
and (n1051,n1052,n1053);
xor (n1052,n982,n983);
and (n1053,n775,n1047);
and (n1054,n1055,n1056);
xor (n1055,n1052,n1053);
or (n1056,n1057,n1060);
and (n1057,n1058,n1059);
xor (n1058,n988,n989);
and (n1059,n782,n1047);
and (n1060,n1061,n1062);
xor (n1061,n1058,n1059);
or (n1062,n1063,n1066);
and (n1063,n1064,n1065);
xor (n1064,n994,n995);
and (n1065,n789,n1047);
and (n1066,n1067,n1068);
xor (n1067,n1064,n1065);
or (n1068,n1069,n1072);
and (n1069,n1070,n1071);
xor (n1070,n1000,n1001);
and (n1071,n796,n1047);
and (n1072,n1073,n1074);
xor (n1073,n1070,n1071);
or (n1074,n1075,n1078);
and (n1075,n1076,n1077);
xor (n1076,n1006,n1007);
and (n1077,n803,n1047);
and (n1078,n1079,n1080);
xor (n1079,n1076,n1077);
or (n1080,n1081,n1084);
and (n1081,n1082,n1083);
xor (n1082,n1012,n1013);
and (n1083,n810,n1047);
and (n1084,n1085,n1086);
xor (n1085,n1082,n1083);
or (n1086,n1087,n1090);
and (n1087,n1088,n1089);
xor (n1088,n1018,n1019);
and (n1089,n817,n1047);
and (n1090,n1091,n1092);
xor (n1091,n1088,n1089);
or (n1092,n1093,n1096);
and (n1093,n1094,n1095);
xor (n1094,n1024,n1025);
and (n1095,n824,n1047);
and (n1096,n1097,n1098);
xor (n1097,n1094,n1095);
or (n1098,n1099,n1102);
and (n1099,n1100,n1101);
xor (n1100,n1030,n1031);
and (n1101,n831,n1047);
and (n1102,n1103,n1104);
xor (n1103,n1100,n1101);
or (n1104,n1105,n1108);
and (n1105,n1106,n1107);
xor (n1106,n1036,n1037);
and (n1107,n838,n1047);
and (n1108,n1109,n1110);
xor (n1109,n1106,n1107);
and (n1110,n1111,n1112);
xor (n1111,n1042,n1043);
and (n1112,n844,n1047);
and (n1113,n768,n1114);
and (n1115,n1116,n1117);
xor (n1116,n758,n1113);
or (n1117,n1118,n1121);
and (n1118,n1119,n1120);
xor (n1119,n1049,n1050);
and (n1120,n775,n1114);
and (n1121,n1122,n1123);
xor (n1122,n1119,n1120);
or (n1123,n1124,n1127);
and (n1124,n1125,n1126);
xor (n1125,n1055,n1056);
and (n1126,n782,n1114);
and (n1127,n1128,n1129);
xor (n1128,n1125,n1126);
or (n1129,n1130,n1133);
and (n1130,n1131,n1132);
xor (n1131,n1061,n1062);
and (n1132,n789,n1114);
and (n1133,n1134,n1135);
xor (n1134,n1131,n1132);
or (n1135,n1136,n1139);
and (n1136,n1137,n1138);
xor (n1137,n1067,n1068);
and (n1138,n796,n1114);
and (n1139,n1140,n1141);
xor (n1140,n1137,n1138);
or (n1141,n1142,n1145);
and (n1142,n1143,n1144);
xor (n1143,n1073,n1074);
and (n1144,n803,n1114);
and (n1145,n1146,n1147);
xor (n1146,n1143,n1144);
or (n1147,n1148,n1151);
and (n1148,n1149,n1150);
xor (n1149,n1079,n1080);
and (n1150,n810,n1114);
and (n1151,n1152,n1153);
xor (n1152,n1149,n1150);
or (n1153,n1154,n1157);
and (n1154,n1155,n1156);
xor (n1155,n1085,n1086);
and (n1156,n817,n1114);
and (n1157,n1158,n1159);
xor (n1158,n1155,n1156);
or (n1159,n1160,n1163);
and (n1160,n1161,n1162);
xor (n1161,n1091,n1092);
and (n1162,n824,n1114);
and (n1163,n1164,n1165);
xor (n1164,n1161,n1162);
or (n1165,n1166,n1169);
and (n1166,n1167,n1168);
xor (n1167,n1097,n1098);
and (n1168,n831,n1114);
and (n1169,n1170,n1171);
xor (n1170,n1167,n1168);
or (n1171,n1172,n1175);
and (n1172,n1173,n1174);
xor (n1173,n1103,n1104);
and (n1174,n838,n1114);
and (n1175,n1176,n1177);
xor (n1176,n1173,n1174);
and (n1177,n1178,n1179);
xor (n1178,n1109,n1110);
and (n1179,n844,n1114);
and (n1180,n768,n1181);
and (n1182,n1183,n1184);
xor (n1183,n756,n1180);
or (n1184,n1185,n1188);
and (n1185,n1186,n1187);
xor (n1186,n1116,n1117);
and (n1187,n775,n1181);
and (n1188,n1189,n1190);
xor (n1189,n1186,n1187);
or (n1190,n1191,n1194);
and (n1191,n1192,n1193);
xor (n1192,n1122,n1123);
and (n1193,n782,n1181);
and (n1194,n1195,n1196);
xor (n1195,n1192,n1193);
or (n1196,n1197,n1200);
and (n1197,n1198,n1199);
xor (n1198,n1128,n1129);
and (n1199,n789,n1181);
and (n1200,n1201,n1202);
xor (n1201,n1198,n1199);
or (n1202,n1203,n1206);
and (n1203,n1204,n1205);
xor (n1204,n1134,n1135);
and (n1205,n796,n1181);
and (n1206,n1207,n1208);
xor (n1207,n1204,n1205);
or (n1208,n1209,n1212);
and (n1209,n1210,n1211);
xor (n1210,n1140,n1141);
and (n1211,n803,n1181);
and (n1212,n1213,n1214);
xor (n1213,n1210,n1211);
or (n1214,n1215,n1218);
and (n1215,n1216,n1217);
xor (n1216,n1146,n1147);
and (n1217,n810,n1181);
and (n1218,n1219,n1220);
xor (n1219,n1216,n1217);
or (n1220,n1221,n1224);
and (n1221,n1222,n1223);
xor (n1222,n1152,n1153);
and (n1223,n817,n1181);
and (n1224,n1225,n1226);
xor (n1225,n1222,n1223);
or (n1226,n1227,n1230);
and (n1227,n1228,n1229);
xor (n1228,n1158,n1159);
and (n1229,n824,n1181);
and (n1230,n1231,n1232);
xor (n1231,n1228,n1229);
or (n1232,n1233,n1236);
and (n1233,n1234,n1235);
xor (n1234,n1164,n1165);
and (n1235,n831,n1181);
and (n1236,n1237,n1238);
xor (n1237,n1234,n1235);
or (n1238,n1239,n1242);
and (n1239,n1240,n1241);
xor (n1240,n1170,n1171);
and (n1241,n838,n1181);
and (n1242,n1243,n1244);
xor (n1243,n1240,n1241);
and (n1244,n1245,n1246);
xor (n1245,n1176,n1177);
and (n1246,n844,n1181);
and (n1247,n768,n1248);
and (n1249,n1250,n1251);
xor (n1250,n754,n1247);
or (n1251,n1252,n1255);
and (n1252,n1253,n1254);
xor (n1253,n1183,n1184);
and (n1254,n775,n1248);
and (n1255,n1256,n1257);
xor (n1256,n1253,n1254);
or (n1257,n1258,n1261);
and (n1258,n1259,n1260);
xor (n1259,n1189,n1190);
and (n1260,n782,n1248);
and (n1261,n1262,n1263);
xor (n1262,n1259,n1260);
or (n1263,n1264,n1267);
and (n1264,n1265,n1266);
xor (n1265,n1195,n1196);
and (n1266,n789,n1248);
and (n1267,n1268,n1269);
xor (n1268,n1265,n1266);
or (n1269,n1270,n1273);
and (n1270,n1271,n1272);
xor (n1271,n1201,n1202);
and (n1272,n796,n1248);
and (n1273,n1274,n1275);
xor (n1274,n1271,n1272);
or (n1275,n1276,n1279);
and (n1276,n1277,n1278);
xor (n1277,n1207,n1208);
and (n1278,n803,n1248);
and (n1279,n1280,n1281);
xor (n1280,n1277,n1278);
or (n1281,n1282,n1285);
and (n1282,n1283,n1284);
xor (n1283,n1213,n1214);
and (n1284,n810,n1248);
and (n1285,n1286,n1287);
xor (n1286,n1283,n1284);
or (n1287,n1288,n1291);
and (n1288,n1289,n1290);
xor (n1289,n1219,n1220);
and (n1290,n817,n1248);
and (n1291,n1292,n1293);
xor (n1292,n1289,n1290);
or (n1293,n1294,n1297);
and (n1294,n1295,n1296);
xor (n1295,n1225,n1226);
and (n1296,n824,n1248);
and (n1297,n1298,n1299);
xor (n1298,n1295,n1296);
or (n1299,n1300,n1303);
and (n1300,n1301,n1302);
xor (n1301,n1231,n1232);
and (n1302,n831,n1248);
and (n1303,n1304,n1305);
xor (n1304,n1301,n1302);
or (n1305,n1306,n1309);
and (n1306,n1307,n1308);
xor (n1307,n1237,n1238);
and (n1308,n838,n1248);
and (n1309,n1310,n1311);
xor (n1310,n1307,n1308);
and (n1311,n1312,n1313);
xor (n1312,n1243,n1244);
and (n1313,n844,n1248);
and (n1314,n768,n1315);
or (n1316,n1317,n1320);
and (n1317,n1318,n1319);
xor (n1318,n1250,n1251);
and (n1319,n775,n1315);
and (n1320,n1321,n1322);
xor (n1321,n1318,n1319);
or (n1322,n1323,n1326);
and (n1323,n1324,n1325);
xor (n1324,n1256,n1257);
and (n1325,n782,n1315);
and (n1326,n1327,n1328);
xor (n1327,n1324,n1325);
or (n1328,n1329,n1332);
and (n1329,n1330,n1331);
xor (n1330,n1262,n1263);
and (n1331,n789,n1315);
and (n1332,n1333,n1334);
xor (n1333,n1330,n1331);
or (n1334,n1335,n1338);
and (n1335,n1336,n1337);
xor (n1336,n1268,n1269);
and (n1337,n796,n1315);
and (n1338,n1339,n1340);
xor (n1339,n1336,n1337);
or (n1340,n1341,n1344);
and (n1341,n1342,n1343);
xor (n1342,n1274,n1275);
and (n1343,n803,n1315);
and (n1344,n1345,n1346);
xor (n1345,n1342,n1343);
or (n1346,n1347,n1350);
and (n1347,n1348,n1349);
xor (n1348,n1280,n1281);
and (n1349,n810,n1315);
and (n1350,n1351,n1352);
xor (n1351,n1348,n1349);
or (n1352,n1353,n1356);
and (n1353,n1354,n1355);
xor (n1354,n1286,n1287);
and (n1355,n817,n1315);
and (n1356,n1357,n1358);
xor (n1357,n1354,n1355);
or (n1358,n1359,n1362);
and (n1359,n1360,n1361);
xor (n1360,n1292,n1293);
and (n1361,n824,n1315);
and (n1362,n1363,n1364);
xor (n1363,n1360,n1361);
or (n1364,n1365,n1368);
and (n1365,n1366,n1367);
xor (n1366,n1298,n1299);
and (n1367,n831,n1315);
and (n1368,n1369,n1370);
xor (n1369,n1366,n1367);
or (n1370,n1371,n1374);
and (n1371,n1372,n1373);
xor (n1372,n1304,n1305);
and (n1373,n838,n1315);
and (n1374,n1375,n1376);
xor (n1375,n1372,n1373);
and (n1376,n1377,n1378);
xor (n1377,n1310,n1311);
and (n1378,n844,n1315);
and (n1379,n775,n1380);
or (n1381,n1382,n1385);
and (n1382,n1383,n1384);
xor (n1383,n1321,n1322);
and (n1384,n782,n1380);
and (n1385,n1386,n1387);
xor (n1386,n1383,n1384);
or (n1387,n1388,n1391);
and (n1388,n1389,n1390);
xor (n1389,n1327,n1328);
and (n1390,n789,n1380);
and (n1391,n1392,n1393);
xor (n1392,n1389,n1390);
or (n1393,n1394,n1397);
and (n1394,n1395,n1396);
xor (n1395,n1333,n1334);
and (n1396,n796,n1380);
and (n1397,n1398,n1399);
xor (n1398,n1395,n1396);
or (n1399,n1400,n1403);
and (n1400,n1401,n1402);
xor (n1401,n1339,n1340);
and (n1402,n803,n1380);
and (n1403,n1404,n1405);
xor (n1404,n1401,n1402);
or (n1405,n1406,n1409);
and (n1406,n1407,n1408);
xor (n1407,n1345,n1346);
and (n1408,n810,n1380);
and (n1409,n1410,n1411);
xor (n1410,n1407,n1408);
or (n1411,n1412,n1415);
and (n1412,n1413,n1414);
xor (n1413,n1351,n1352);
and (n1414,n817,n1380);
and (n1415,n1416,n1417);
xor (n1416,n1413,n1414);
or (n1417,n1418,n1421);
and (n1418,n1419,n1420);
xor (n1419,n1357,n1358);
and (n1420,n824,n1380);
and (n1421,n1422,n1423);
xor (n1422,n1419,n1420);
or (n1423,n1424,n1427);
and (n1424,n1425,n1426);
xor (n1425,n1363,n1364);
and (n1426,n831,n1380);
and (n1427,n1428,n1429);
xor (n1428,n1425,n1426);
or (n1429,n1430,n1433);
and (n1430,n1431,n1432);
xor (n1431,n1369,n1370);
and (n1432,n838,n1380);
and (n1433,n1434,n1435);
xor (n1434,n1431,n1432);
and (n1435,n1436,n1437);
xor (n1436,n1375,n1376);
and (n1437,n844,n1380);
and (n1438,n782,n1439);
or (n1440,n1441,n1444);
and (n1441,n1442,n1443);
xor (n1442,n1386,n1387);
and (n1443,n789,n1439);
and (n1444,n1445,n1446);
xor (n1445,n1442,n1443);
or (n1446,n1447,n1450);
and (n1447,n1448,n1449);
xor (n1448,n1392,n1393);
and (n1449,n796,n1439);
and (n1450,n1451,n1452);
xor (n1451,n1448,n1449);
or (n1452,n1453,n1456);
and (n1453,n1454,n1455);
xor (n1454,n1398,n1399);
and (n1455,n803,n1439);
and (n1456,n1457,n1458);
xor (n1457,n1454,n1455);
or (n1458,n1459,n1462);
and (n1459,n1460,n1461);
xor (n1460,n1404,n1405);
and (n1461,n810,n1439);
and (n1462,n1463,n1464);
xor (n1463,n1460,n1461);
or (n1464,n1465,n1468);
and (n1465,n1466,n1467);
xor (n1466,n1410,n1411);
and (n1467,n817,n1439);
and (n1468,n1469,n1470);
xor (n1469,n1466,n1467);
or (n1470,n1471,n1474);
and (n1471,n1472,n1473);
xor (n1472,n1416,n1417);
and (n1473,n824,n1439);
and (n1474,n1475,n1476);
xor (n1475,n1472,n1473);
or (n1476,n1477,n1480);
and (n1477,n1478,n1479);
xor (n1478,n1422,n1423);
and (n1479,n831,n1439);
and (n1480,n1481,n1482);
xor (n1481,n1478,n1479);
or (n1482,n1483,n1486);
and (n1483,n1484,n1485);
xor (n1484,n1428,n1429);
and (n1485,n838,n1439);
and (n1486,n1487,n1488);
xor (n1487,n1484,n1485);
and (n1488,n1489,n1490);
xor (n1489,n1434,n1435);
and (n1490,n844,n1439);
xor (n1492,n1493,n2186);
xor (n1493,n1494,n2184);
xor (n1494,n1495,n2127);
xor (n1495,n1496,n2125);
xor (n1496,n1497,n2062);
xor (n1497,n1498,n2060);
or (n1498,n1499,n1995);
and (n1499,n1500,n1993);
or (n1500,n1501,n1928);
and (n1501,n1502,n1926);
or (n1502,n1503,n1861);
and (n1503,n1504,n1859);
or (n1504,n1505,n1794);
and (n1505,n1506,n1792);
or (n1506,n1507,n1727);
and (n1507,n1508,n1725);
or (n1508,n1509,n1660);
and (n1509,n1510,n1658);
or (n1510,n1511,n1593);
and (n1511,n1512,n1591);
and (n1512,n1513,n1516);
and (n1513,n1514,n1515);
wire s0n1514,s1n1514,notn1514;
or (n1514,s0n1514,s1n1514);
not(notn1514,n1491);
and (s0n1514,notn1514,n23);
and (s1n1514,n1491,n768);
wire s0n1515,s1n1515,notn1515;
or (n1515,s0n1515,s1n1515);
not(notn1515,n1491);
and (s0n1515,notn1515,n24);
and (s1n1515,n1491,n769);
or (n1516,n1517,n1522);
and (n1517,n1518,n1520);
and (n1518,n1514,n1519);
wire s0n1519,s1n1519,notn1519;
or (n1519,s0n1519,s1n1519);
not(notn1519,n1491);
and (s0n1519,notn1519,n28);
and (s1n1519,n1491,n773);
and (n1520,n1521,n1515);
wire s0n1521,s1n1521,notn1521;
or (n1521,s0n1521,s1n1521);
not(notn1521,n1491);
and (s0n1521,notn1521,n30);
and (s1n1521,n1491,n775);
and (n1522,n1523,n1524);
xor (n1523,n1518,n1520);
or (n1524,n1525,n1529);
and (n1525,n1526,n1527);
and (n1526,n1521,n1519);
and (n1527,n1528,n1515);
wire s0n1528,s1n1528,notn1528;
or (n1528,s0n1528,s1n1528);
not(notn1528,n1491);
and (s0n1528,notn1528,n37);
and (s1n1528,n1491,n782);
and (n1529,n1530,n1531);
xor (n1530,n1526,n1527);
or (n1531,n1532,n1536);
and (n1532,n1533,n1534);
and (n1533,n1528,n1519);
and (n1534,n1535,n1515);
wire s0n1535,s1n1535,notn1535;
or (n1535,s0n1535,s1n1535);
not(notn1535,n1491);
and (s0n1535,notn1535,n44);
and (s1n1535,n1491,n789);
and (n1536,n1537,n1538);
xor (n1537,n1533,n1534);
or (n1538,n1539,n1543);
and (n1539,n1540,n1541);
and (n1540,n1535,n1519);
and (n1541,n1542,n1515);
wire s0n1542,s1n1542,notn1542;
or (n1542,s0n1542,s1n1542);
not(notn1542,n1491);
and (s0n1542,notn1542,n51);
and (s1n1542,n1491,n796);
and (n1543,n1544,n1545);
xor (n1544,n1540,n1541);
or (n1545,n1546,n1550);
and (n1546,n1547,n1548);
and (n1547,n1542,n1519);
and (n1548,n1549,n1515);
wire s0n1549,s1n1549,notn1549;
or (n1549,s0n1549,s1n1549);
not(notn1549,n1491);
and (s0n1549,notn1549,n58);
and (s1n1549,n1491,n803);
and (n1550,n1551,n1552);
xor (n1551,n1547,n1548);
or (n1552,n1553,n1557);
and (n1553,n1554,n1555);
and (n1554,n1549,n1519);
and (n1555,n1556,n1515);
wire s0n1556,s1n1556,notn1556;
or (n1556,s0n1556,s1n1556);
not(notn1556,n1491);
and (s0n1556,notn1556,n65);
and (s1n1556,n1491,n810);
and (n1557,n1558,n1559);
xor (n1558,n1554,n1555);
or (n1559,n1560,n1564);
and (n1560,n1561,n1562);
and (n1561,n1556,n1519);
and (n1562,n1563,n1515);
wire s0n1563,s1n1563,notn1563;
or (n1563,s0n1563,s1n1563);
not(notn1563,n1491);
and (s0n1563,notn1563,n72);
and (s1n1563,n1491,n817);
and (n1564,n1565,n1566);
xor (n1565,n1561,n1562);
or (n1566,n1567,n1571);
and (n1567,n1568,n1569);
and (n1568,n1563,n1519);
and (n1569,n1570,n1515);
wire s0n1570,s1n1570,notn1570;
or (n1570,s0n1570,s1n1570);
not(notn1570,n1491);
and (s0n1570,notn1570,n79);
and (s1n1570,n1491,n824);
and (n1571,n1572,n1573);
xor (n1572,n1568,n1569);
or (n1573,n1574,n1578);
and (n1574,n1575,n1576);
and (n1575,n1570,n1519);
and (n1576,n1577,n1515);
wire s0n1577,s1n1577,notn1577;
or (n1577,s0n1577,s1n1577);
not(notn1577,n1491);
and (s0n1577,notn1577,n86);
and (s1n1577,n1491,n831);
and (n1578,n1579,n1580);
xor (n1579,n1575,n1576);
or (n1580,n1581,n1585);
and (n1581,n1582,n1583);
and (n1582,n1577,n1519);
and (n1583,n1584,n1515);
wire s0n1584,s1n1584,notn1584;
or (n1584,s0n1584,s1n1584);
not(notn1584,n1491);
and (s0n1584,notn1584,n93);
and (s1n1584,n1491,n838);
and (n1585,n1586,n1587);
xor (n1586,n1582,n1583);
and (n1587,n1588,n1589);
and (n1588,n1584,n1519);
and (n1589,n1590,n1515);
wire s0n1590,s1n1590,notn1590;
or (n1590,s0n1590,s1n1590);
not(notn1590,n1491);
and (s0n1590,notn1590,n99);
and (s1n1590,n1491,n844);
and (n1591,n1514,n1592);
wire s0n1592,s1n1592,notn1592;
or (n1592,s0n1592,s1n1592);
not(notn1592,n1491);
and (s0n1592,notn1592,n101);
and (s1n1592,n1491,n846);
and (n1593,n1594,n1595);
xor (n1594,n1512,n1591);
or (n1595,n1596,n1599);
and (n1596,n1597,n1598);
xor (n1597,n1513,n1516);
and (n1598,n1521,n1592);
and (n1599,n1600,n1601);
xor (n1600,n1597,n1598);
or (n1601,n1602,n1605);
and (n1602,n1603,n1604);
xor (n1603,n1523,n1524);
and (n1604,n1528,n1592);
and (n1605,n1606,n1607);
xor (n1606,n1603,n1604);
or (n1607,n1608,n1611);
and (n1608,n1609,n1610);
xor (n1609,n1530,n1531);
and (n1610,n1535,n1592);
and (n1611,n1612,n1613);
xor (n1612,n1609,n1610);
or (n1613,n1614,n1617);
and (n1614,n1615,n1616);
xor (n1615,n1537,n1538);
and (n1616,n1542,n1592);
and (n1617,n1618,n1619);
xor (n1618,n1615,n1616);
or (n1619,n1620,n1623);
and (n1620,n1621,n1622);
xor (n1621,n1544,n1545);
and (n1622,n1549,n1592);
and (n1623,n1624,n1625);
xor (n1624,n1621,n1622);
or (n1625,n1626,n1629);
and (n1626,n1627,n1628);
xor (n1627,n1551,n1552);
and (n1628,n1556,n1592);
and (n1629,n1630,n1631);
xor (n1630,n1627,n1628);
or (n1631,n1632,n1635);
and (n1632,n1633,n1634);
xor (n1633,n1558,n1559);
and (n1634,n1563,n1592);
and (n1635,n1636,n1637);
xor (n1636,n1633,n1634);
or (n1637,n1638,n1641);
and (n1638,n1639,n1640);
xor (n1639,n1565,n1566);
and (n1640,n1570,n1592);
and (n1641,n1642,n1643);
xor (n1642,n1639,n1640);
or (n1643,n1644,n1647);
and (n1644,n1645,n1646);
xor (n1645,n1572,n1573);
and (n1646,n1577,n1592);
and (n1647,n1648,n1649);
xor (n1648,n1645,n1646);
or (n1649,n1650,n1653);
and (n1650,n1651,n1652);
xor (n1651,n1579,n1580);
and (n1652,n1584,n1592);
and (n1653,n1654,n1655);
xor (n1654,n1651,n1652);
and (n1655,n1656,n1657);
xor (n1656,n1586,n1587);
and (n1657,n1590,n1592);
and (n1658,n1514,n1659);
wire s0n1659,s1n1659,notn1659;
or (n1659,s0n1659,s1n1659);
not(notn1659,n1491);
and (s0n1659,notn1659,n168);
and (s1n1659,n1491,n913);
and (n1660,n1661,n1662);
xor (n1661,n1510,n1658);
or (n1662,n1663,n1666);
and (n1663,n1664,n1665);
xor (n1664,n1594,n1595);
and (n1665,n1521,n1659);
and (n1666,n1667,n1668);
xor (n1667,n1664,n1665);
or (n1668,n1669,n1672);
and (n1669,n1670,n1671);
xor (n1670,n1600,n1601);
and (n1671,n1528,n1659);
and (n1672,n1673,n1674);
xor (n1673,n1670,n1671);
or (n1674,n1675,n1678);
and (n1675,n1676,n1677);
xor (n1676,n1606,n1607);
and (n1677,n1535,n1659);
and (n1678,n1679,n1680);
xor (n1679,n1676,n1677);
or (n1680,n1681,n1684);
and (n1681,n1682,n1683);
xor (n1682,n1612,n1613);
and (n1683,n1542,n1659);
and (n1684,n1685,n1686);
xor (n1685,n1682,n1683);
or (n1686,n1687,n1690);
and (n1687,n1688,n1689);
xor (n1688,n1618,n1619);
and (n1689,n1549,n1659);
and (n1690,n1691,n1692);
xor (n1691,n1688,n1689);
or (n1692,n1693,n1696);
and (n1693,n1694,n1695);
xor (n1694,n1624,n1625);
and (n1695,n1556,n1659);
and (n1696,n1697,n1698);
xor (n1697,n1694,n1695);
or (n1698,n1699,n1702);
and (n1699,n1700,n1701);
xor (n1700,n1630,n1631);
and (n1701,n1563,n1659);
and (n1702,n1703,n1704);
xor (n1703,n1700,n1701);
or (n1704,n1705,n1708);
and (n1705,n1706,n1707);
xor (n1706,n1636,n1637);
and (n1707,n1570,n1659);
and (n1708,n1709,n1710);
xor (n1709,n1706,n1707);
or (n1710,n1711,n1714);
and (n1711,n1712,n1713);
xor (n1712,n1642,n1643);
and (n1713,n1577,n1659);
and (n1714,n1715,n1716);
xor (n1715,n1712,n1713);
or (n1716,n1717,n1720);
and (n1717,n1718,n1719);
xor (n1718,n1648,n1649);
and (n1719,n1584,n1659);
and (n1720,n1721,n1722);
xor (n1721,n1718,n1719);
and (n1722,n1723,n1724);
xor (n1723,n1654,n1655);
and (n1724,n1590,n1659);
and (n1725,n1514,n1726);
wire s0n1726,s1n1726,notn1726;
or (n1726,s0n1726,s1n1726);
not(notn1726,n1491);
and (s0n1726,notn1726,n235);
and (s1n1726,n1491,n980);
and (n1727,n1728,n1729);
xor (n1728,n1508,n1725);
or (n1729,n1730,n1733);
and (n1730,n1731,n1732);
xor (n1731,n1661,n1662);
and (n1732,n1521,n1726);
and (n1733,n1734,n1735);
xor (n1734,n1731,n1732);
or (n1735,n1736,n1739);
and (n1736,n1737,n1738);
xor (n1737,n1667,n1668);
and (n1738,n1528,n1726);
and (n1739,n1740,n1741);
xor (n1740,n1737,n1738);
or (n1741,n1742,n1745);
and (n1742,n1743,n1744);
xor (n1743,n1673,n1674);
and (n1744,n1535,n1726);
and (n1745,n1746,n1747);
xor (n1746,n1743,n1744);
or (n1747,n1748,n1751);
and (n1748,n1749,n1750);
xor (n1749,n1679,n1680);
and (n1750,n1542,n1726);
and (n1751,n1752,n1753);
xor (n1752,n1749,n1750);
or (n1753,n1754,n1757);
and (n1754,n1755,n1756);
xor (n1755,n1685,n1686);
and (n1756,n1549,n1726);
and (n1757,n1758,n1759);
xor (n1758,n1755,n1756);
or (n1759,n1760,n1763);
and (n1760,n1761,n1762);
xor (n1761,n1691,n1692);
and (n1762,n1556,n1726);
and (n1763,n1764,n1765);
xor (n1764,n1761,n1762);
or (n1765,n1766,n1769);
and (n1766,n1767,n1768);
xor (n1767,n1697,n1698);
and (n1768,n1563,n1726);
and (n1769,n1770,n1771);
xor (n1770,n1767,n1768);
or (n1771,n1772,n1775);
and (n1772,n1773,n1774);
xor (n1773,n1703,n1704);
and (n1774,n1570,n1726);
and (n1775,n1776,n1777);
xor (n1776,n1773,n1774);
or (n1777,n1778,n1781);
and (n1778,n1779,n1780);
xor (n1779,n1709,n1710);
and (n1780,n1577,n1726);
and (n1781,n1782,n1783);
xor (n1782,n1779,n1780);
or (n1783,n1784,n1787);
and (n1784,n1785,n1786);
xor (n1785,n1715,n1716);
and (n1786,n1584,n1726);
and (n1787,n1788,n1789);
xor (n1788,n1785,n1786);
and (n1789,n1790,n1791);
xor (n1790,n1721,n1722);
and (n1791,n1590,n1726);
and (n1792,n1514,n1793);
wire s0n1793,s1n1793,notn1793;
or (n1793,s0n1793,s1n1793);
not(notn1793,n1491);
and (s0n1793,notn1793,n302);
and (s1n1793,n1491,n1047);
and (n1794,n1795,n1796);
xor (n1795,n1506,n1792);
or (n1796,n1797,n1800);
and (n1797,n1798,n1799);
xor (n1798,n1728,n1729);
and (n1799,n1521,n1793);
and (n1800,n1801,n1802);
xor (n1801,n1798,n1799);
or (n1802,n1803,n1806);
and (n1803,n1804,n1805);
xor (n1804,n1734,n1735);
and (n1805,n1528,n1793);
and (n1806,n1807,n1808);
xor (n1807,n1804,n1805);
or (n1808,n1809,n1812);
and (n1809,n1810,n1811);
xor (n1810,n1740,n1741);
and (n1811,n1535,n1793);
and (n1812,n1813,n1814);
xor (n1813,n1810,n1811);
or (n1814,n1815,n1818);
and (n1815,n1816,n1817);
xor (n1816,n1746,n1747);
and (n1817,n1542,n1793);
and (n1818,n1819,n1820);
xor (n1819,n1816,n1817);
or (n1820,n1821,n1824);
and (n1821,n1822,n1823);
xor (n1822,n1752,n1753);
and (n1823,n1549,n1793);
and (n1824,n1825,n1826);
xor (n1825,n1822,n1823);
or (n1826,n1827,n1830);
and (n1827,n1828,n1829);
xor (n1828,n1758,n1759);
and (n1829,n1556,n1793);
and (n1830,n1831,n1832);
xor (n1831,n1828,n1829);
or (n1832,n1833,n1836);
and (n1833,n1834,n1835);
xor (n1834,n1764,n1765);
and (n1835,n1563,n1793);
and (n1836,n1837,n1838);
xor (n1837,n1834,n1835);
or (n1838,n1839,n1842);
and (n1839,n1840,n1841);
xor (n1840,n1770,n1771);
and (n1841,n1570,n1793);
and (n1842,n1843,n1844);
xor (n1843,n1840,n1841);
or (n1844,n1845,n1848);
and (n1845,n1846,n1847);
xor (n1846,n1776,n1777);
and (n1847,n1577,n1793);
and (n1848,n1849,n1850);
xor (n1849,n1846,n1847);
or (n1850,n1851,n1854);
and (n1851,n1852,n1853);
xor (n1852,n1782,n1783);
and (n1853,n1584,n1793);
and (n1854,n1855,n1856);
xor (n1855,n1852,n1853);
and (n1856,n1857,n1858);
xor (n1857,n1788,n1789);
and (n1858,n1590,n1793);
and (n1859,n1514,n1860);
wire s0n1860,s1n1860,notn1860;
or (n1860,s0n1860,s1n1860);
not(notn1860,n1491);
and (s0n1860,notn1860,n369);
and (s1n1860,n1491,n1114);
and (n1861,n1862,n1863);
xor (n1862,n1504,n1859);
or (n1863,n1864,n1867);
and (n1864,n1865,n1866);
xor (n1865,n1795,n1796);
and (n1866,n1521,n1860);
and (n1867,n1868,n1869);
xor (n1868,n1865,n1866);
or (n1869,n1870,n1873);
and (n1870,n1871,n1872);
xor (n1871,n1801,n1802);
and (n1872,n1528,n1860);
and (n1873,n1874,n1875);
xor (n1874,n1871,n1872);
or (n1875,n1876,n1879);
and (n1876,n1877,n1878);
xor (n1877,n1807,n1808);
and (n1878,n1535,n1860);
and (n1879,n1880,n1881);
xor (n1880,n1877,n1878);
or (n1881,n1882,n1885);
and (n1882,n1883,n1884);
xor (n1883,n1813,n1814);
and (n1884,n1542,n1860);
and (n1885,n1886,n1887);
xor (n1886,n1883,n1884);
or (n1887,n1888,n1891);
and (n1888,n1889,n1890);
xor (n1889,n1819,n1820);
and (n1890,n1549,n1860);
and (n1891,n1892,n1893);
xor (n1892,n1889,n1890);
or (n1893,n1894,n1897);
and (n1894,n1895,n1896);
xor (n1895,n1825,n1826);
and (n1896,n1556,n1860);
and (n1897,n1898,n1899);
xor (n1898,n1895,n1896);
or (n1899,n1900,n1903);
and (n1900,n1901,n1902);
xor (n1901,n1831,n1832);
and (n1902,n1563,n1860);
and (n1903,n1904,n1905);
xor (n1904,n1901,n1902);
or (n1905,n1906,n1909);
and (n1906,n1907,n1908);
xor (n1907,n1837,n1838);
and (n1908,n1570,n1860);
and (n1909,n1910,n1911);
xor (n1910,n1907,n1908);
or (n1911,n1912,n1915);
and (n1912,n1913,n1914);
xor (n1913,n1843,n1844);
and (n1914,n1577,n1860);
and (n1915,n1916,n1917);
xor (n1916,n1913,n1914);
or (n1917,n1918,n1921);
and (n1918,n1919,n1920);
xor (n1919,n1849,n1850);
and (n1920,n1584,n1860);
and (n1921,n1922,n1923);
xor (n1922,n1919,n1920);
and (n1923,n1924,n1925);
xor (n1924,n1855,n1856);
and (n1925,n1590,n1860);
and (n1926,n1514,n1927);
wire s0n1927,s1n1927,notn1927;
or (n1927,s0n1927,s1n1927);
not(notn1927,n1491);
and (s0n1927,notn1927,n436);
and (s1n1927,n1491,n1181);
and (n1928,n1929,n1930);
xor (n1929,n1502,n1926);
or (n1930,n1931,n1934);
and (n1931,n1932,n1933);
xor (n1932,n1862,n1863);
and (n1933,n1521,n1927);
and (n1934,n1935,n1936);
xor (n1935,n1932,n1933);
or (n1936,n1937,n1940);
and (n1937,n1938,n1939);
xor (n1938,n1868,n1869);
and (n1939,n1528,n1927);
and (n1940,n1941,n1942);
xor (n1941,n1938,n1939);
or (n1942,n1943,n1946);
and (n1943,n1944,n1945);
xor (n1944,n1874,n1875);
and (n1945,n1535,n1927);
and (n1946,n1947,n1948);
xor (n1947,n1944,n1945);
or (n1948,n1949,n1952);
and (n1949,n1950,n1951);
xor (n1950,n1880,n1881);
and (n1951,n1542,n1927);
and (n1952,n1953,n1954);
xor (n1953,n1950,n1951);
or (n1954,n1955,n1958);
and (n1955,n1956,n1957);
xor (n1956,n1886,n1887);
and (n1957,n1549,n1927);
and (n1958,n1959,n1960);
xor (n1959,n1956,n1957);
or (n1960,n1961,n1964);
and (n1961,n1962,n1963);
xor (n1962,n1892,n1893);
and (n1963,n1556,n1927);
and (n1964,n1965,n1966);
xor (n1965,n1962,n1963);
or (n1966,n1967,n1970);
and (n1967,n1968,n1969);
xor (n1968,n1898,n1899);
and (n1969,n1563,n1927);
and (n1970,n1971,n1972);
xor (n1971,n1968,n1969);
or (n1972,n1973,n1976);
and (n1973,n1974,n1975);
xor (n1974,n1904,n1905);
and (n1975,n1570,n1927);
and (n1976,n1977,n1978);
xor (n1977,n1974,n1975);
or (n1978,n1979,n1982);
and (n1979,n1980,n1981);
xor (n1980,n1910,n1911);
and (n1981,n1577,n1927);
and (n1982,n1983,n1984);
xor (n1983,n1980,n1981);
or (n1984,n1985,n1988);
and (n1985,n1986,n1987);
xor (n1986,n1916,n1917);
and (n1987,n1584,n1927);
and (n1988,n1989,n1990);
xor (n1989,n1986,n1987);
and (n1990,n1991,n1992);
xor (n1991,n1922,n1923);
and (n1992,n1590,n1927);
and (n1993,n1514,n1994);
wire s0n1994,s1n1994,notn1994;
or (n1994,s0n1994,s1n1994);
not(notn1994,n1491);
and (s0n1994,notn1994,n503);
and (s1n1994,n1491,n1248);
and (n1995,n1996,n1997);
xor (n1996,n1500,n1993);
or (n1997,n1998,n2001);
and (n1998,n1999,n2000);
xor (n1999,n1929,n1930);
and (n2000,n1521,n1994);
and (n2001,n2002,n2003);
xor (n2002,n1999,n2000);
or (n2003,n2004,n2007);
and (n2004,n2005,n2006);
xor (n2005,n1935,n1936);
and (n2006,n1528,n1994);
and (n2007,n2008,n2009);
xor (n2008,n2005,n2006);
or (n2009,n2010,n2013);
and (n2010,n2011,n2012);
xor (n2011,n1941,n1942);
and (n2012,n1535,n1994);
and (n2013,n2014,n2015);
xor (n2014,n2011,n2012);
or (n2015,n2016,n2019);
and (n2016,n2017,n2018);
xor (n2017,n1947,n1948);
and (n2018,n1542,n1994);
and (n2019,n2020,n2021);
xor (n2020,n2017,n2018);
or (n2021,n2022,n2025);
and (n2022,n2023,n2024);
xor (n2023,n1953,n1954);
and (n2024,n1549,n1994);
and (n2025,n2026,n2027);
xor (n2026,n2023,n2024);
or (n2027,n2028,n2031);
and (n2028,n2029,n2030);
xor (n2029,n1959,n1960);
and (n2030,n1556,n1994);
and (n2031,n2032,n2033);
xor (n2032,n2029,n2030);
or (n2033,n2034,n2037);
and (n2034,n2035,n2036);
xor (n2035,n1965,n1966);
and (n2036,n1563,n1994);
and (n2037,n2038,n2039);
xor (n2038,n2035,n2036);
or (n2039,n2040,n2043);
and (n2040,n2041,n2042);
xor (n2041,n1971,n1972);
and (n2042,n1570,n1994);
and (n2043,n2044,n2045);
xor (n2044,n2041,n2042);
or (n2045,n2046,n2049);
and (n2046,n2047,n2048);
xor (n2047,n1977,n1978);
and (n2048,n1577,n1994);
and (n2049,n2050,n2051);
xor (n2050,n2047,n2048);
or (n2051,n2052,n2055);
and (n2052,n2053,n2054);
xor (n2053,n1983,n1984);
and (n2054,n1584,n1994);
and (n2055,n2056,n2057);
xor (n2056,n2053,n2054);
and (n2057,n2058,n2059);
xor (n2058,n1989,n1990);
and (n2059,n1590,n1994);
and (n2060,n1514,n2061);
wire s0n2061,s1n2061,notn2061;
or (n2061,s0n2061,s1n2061);
not(notn2061,n1491);
and (s0n2061,notn2061,n570);
and (s1n2061,n1491,n1315);
or (n2062,n2063,n2066);
and (n2063,n2064,n2065);
xor (n2064,n1996,n1997);
and (n2065,n1521,n2061);
and (n2066,n2067,n2068);
xor (n2067,n2064,n2065);
or (n2068,n2069,n2072);
and (n2069,n2070,n2071);
xor (n2070,n2002,n2003);
and (n2071,n1528,n2061);
and (n2072,n2073,n2074);
xor (n2073,n2070,n2071);
or (n2074,n2075,n2078);
and (n2075,n2076,n2077);
xor (n2076,n2008,n2009);
and (n2077,n1535,n2061);
and (n2078,n2079,n2080);
xor (n2079,n2076,n2077);
or (n2080,n2081,n2084);
and (n2081,n2082,n2083);
xor (n2082,n2014,n2015);
and (n2083,n1542,n2061);
and (n2084,n2085,n2086);
xor (n2085,n2082,n2083);
or (n2086,n2087,n2090);
and (n2087,n2088,n2089);
xor (n2088,n2020,n2021);
and (n2089,n1549,n2061);
and (n2090,n2091,n2092);
xor (n2091,n2088,n2089);
or (n2092,n2093,n2096);
and (n2093,n2094,n2095);
xor (n2094,n2026,n2027);
and (n2095,n1556,n2061);
and (n2096,n2097,n2098);
xor (n2097,n2094,n2095);
or (n2098,n2099,n2102);
and (n2099,n2100,n2101);
xor (n2100,n2032,n2033);
and (n2101,n1563,n2061);
and (n2102,n2103,n2104);
xor (n2103,n2100,n2101);
or (n2104,n2105,n2108);
and (n2105,n2106,n2107);
xor (n2106,n2038,n2039);
and (n2107,n1570,n2061);
and (n2108,n2109,n2110);
xor (n2109,n2106,n2107);
or (n2110,n2111,n2114);
and (n2111,n2112,n2113);
xor (n2112,n2044,n2045);
and (n2113,n1577,n2061);
and (n2114,n2115,n2116);
xor (n2115,n2112,n2113);
or (n2116,n2117,n2120);
and (n2117,n2118,n2119);
xor (n2118,n2050,n2051);
and (n2119,n1584,n2061);
and (n2120,n2121,n2122);
xor (n2121,n2118,n2119);
and (n2122,n2123,n2124);
xor (n2123,n2056,n2057);
and (n2124,n1590,n2061);
and (n2125,n1521,n2126);
wire s0n2126,s1n2126,notn2126;
or (n2126,s0n2126,s1n2126);
not(notn2126,n1491);
and (s0n2126,notn2126,n635);
and (s1n2126,n1491,n1380);
or (n2127,n2128,n2131);
and (n2128,n2129,n2130);
xor (n2129,n2067,n2068);
and (n2130,n1528,n2126);
and (n2131,n2132,n2133);
xor (n2132,n2129,n2130);
or (n2133,n2134,n2137);
and (n2134,n2135,n2136);
xor (n2135,n2073,n2074);
and (n2136,n1535,n2126);
and (n2137,n2138,n2139);
xor (n2138,n2135,n2136);
or (n2139,n2140,n2143);
and (n2140,n2141,n2142);
xor (n2141,n2079,n2080);
and (n2142,n1542,n2126);
and (n2143,n2144,n2145);
xor (n2144,n2141,n2142);
or (n2145,n2146,n2149);
and (n2146,n2147,n2148);
xor (n2147,n2085,n2086);
and (n2148,n1549,n2126);
and (n2149,n2150,n2151);
xor (n2150,n2147,n2148);
or (n2151,n2152,n2155);
and (n2152,n2153,n2154);
xor (n2153,n2091,n2092);
and (n2154,n1556,n2126);
and (n2155,n2156,n2157);
xor (n2156,n2153,n2154);
or (n2157,n2158,n2161);
and (n2158,n2159,n2160);
xor (n2159,n2097,n2098);
and (n2160,n1563,n2126);
and (n2161,n2162,n2163);
xor (n2162,n2159,n2160);
or (n2163,n2164,n2167);
and (n2164,n2165,n2166);
xor (n2165,n2103,n2104);
and (n2166,n1570,n2126);
and (n2167,n2168,n2169);
xor (n2168,n2165,n2166);
or (n2169,n2170,n2173);
and (n2170,n2171,n2172);
xor (n2171,n2109,n2110);
and (n2172,n1577,n2126);
and (n2173,n2174,n2175);
xor (n2174,n2171,n2172);
or (n2175,n2176,n2179);
and (n2176,n2177,n2178);
xor (n2177,n2115,n2116);
and (n2178,n1584,n2126);
and (n2179,n2180,n2181);
xor (n2180,n2177,n2178);
and (n2181,n2182,n2183);
xor (n2182,n2121,n2122);
and (n2183,n1590,n2126);
and (n2184,n1528,n2185);
wire s0n2185,s1n2185,notn2185;
or (n2185,s0n2185,s1n2185);
not(notn2185,n1491);
and (s0n2185,notn2185,n694);
and (s1n2185,n1491,n1439);
or (n2186,n2187,n2190);
and (n2187,n2188,n2189);
xor (n2188,n2132,n2133);
and (n2189,n1535,n2185);
and (n2190,n2191,n2192);
xor (n2191,n2188,n2189);
or (n2192,n2193,n2196);
and (n2193,n2194,n2195);
xor (n2194,n2138,n2139);
and (n2195,n1542,n2185);
and (n2196,n2197,n2198);
xor (n2197,n2194,n2195);
or (n2198,n2199,n2202);
and (n2199,n2200,n2201);
xor (n2200,n2144,n2145);
and (n2201,n1549,n2185);
and (n2202,n2203,n2204);
xor (n2203,n2200,n2201);
or (n2204,n2205,n2208);
and (n2205,n2206,n2207);
xor (n2206,n2150,n2151);
and (n2207,n1556,n2185);
and (n2208,n2209,n2210);
xor (n2209,n2206,n2207);
or (n2210,n2211,n2214);
and (n2211,n2212,n2213);
xor (n2212,n2156,n2157);
and (n2213,n1563,n2185);
and (n2214,n2215,n2216);
xor (n2215,n2212,n2213);
or (n2216,n2217,n2220);
and (n2217,n2218,n2219);
xor (n2218,n2162,n2163);
and (n2219,n1570,n2185);
and (n2220,n2221,n2222);
xor (n2221,n2218,n2219);
or (n2222,n2223,n2226);
and (n2223,n2224,n2225);
xor (n2224,n2168,n2169);
and (n2225,n1577,n2185);
and (n2226,n2227,n2228);
xor (n2227,n2224,n2225);
or (n2228,n2229,n2232);
and (n2229,n2230,n2231);
xor (n2230,n2174,n2175);
and (n2231,n1584,n2185);
and (n2232,n2233,n2234);
xor (n2233,n2230,n2231);
and (n2234,n2235,n2236);
xor (n2235,n2180,n2181);
and (n2236,n1590,n2185);
endmodule
