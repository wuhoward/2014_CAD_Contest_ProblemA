module top (out,n23,n24,n28,n30,n37,n44,n51,n58,n65
        ,n72,n79,n86,n93,n99,n101,n166,n225,n278,n325
        ,n366,n401,n430,n453,n470,n502,n503,n507,n509,n516
        ,n523,n530,n537,n544,n551,n558,n565,n572,n578,n580
        ,n645,n704,n757,n804,n845,n880,n909,n932,n949,n959);
output out;
input n23;
input n24;
input n28;
input n30;
input n37;
input n44;
input n51;
input n58;
input n65;
input n72;
input n79;
input n86;
input n93;
input n99;
input n101;
input n166;
input n225;
input n278;
input n325;
input n366;
input n401;
input n430;
input n453;
input n470;
input n502;
input n503;
input n507;
input n509;
input n516;
input n523;
input n530;
input n537;
input n544;
input n551;
input n558;
input n565;
input n572;
input n578;
input n580;
input n645;
input n704;
input n757;
input n804;
input n845;
input n880;
input n909;
input n932;
input n949;
input n959;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n25;
wire n26;
wire n27;
wire n29;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n100;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n504;
wire n505;
wire n506;
wire n508;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n579;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
xor (out,n0,n960);
wire s0n0,s1n0,notn0;
or (n0,s0n0,s1n0);
not(notn0,n959);
and (s0n0,notn0,n1);
and (s1n0,n959,n480);
xor (n1,n2,n471);
xor (n2,n3,n469);
xor (n3,n4,n454);
xor (n4,n5,n452);
xor (n5,n6,n431);
xor (n6,n7,n429);
xor (n7,n8,n402);
xor (n8,n9,n400);
xor (n9,n10,n367);
xor (n10,n11,n365);
xor (n11,n12,n326);
xor (n12,n13,n324);
xor (n13,n14,n279);
xor (n14,n15,n277);
xor (n15,n16,n226);
xor (n16,n17,n224);
xor (n17,n18,n167);
xor (n18,n19,n165);
xor (n19,n20,n102);
xor (n20,n21,n100);
and (n21,n22,n25);
and (n22,n23,n24);
or (n25,n26,n31);
and (n26,n27,n29);
and (n27,n23,n28);
and (n29,n30,n24);
and (n31,n32,n33);
xor (n32,n27,n29);
or (n33,n34,n38);
and (n34,n35,n36);
and (n35,n30,n28);
and (n36,n37,n24);
and (n38,n39,n40);
xor (n39,n35,n36);
or (n40,n41,n45);
and (n41,n42,n43);
and (n42,n37,n28);
and (n43,n44,n24);
and (n45,n46,n47);
xor (n46,n42,n43);
or (n47,n48,n52);
and (n48,n49,n50);
and (n49,n44,n28);
and (n50,n51,n24);
and (n52,n53,n54);
xor (n53,n49,n50);
or (n54,n55,n59);
and (n55,n56,n57);
and (n56,n51,n28);
and (n57,n58,n24);
and (n59,n60,n61);
xor (n60,n56,n57);
or (n61,n62,n66);
and (n62,n63,n64);
and (n63,n58,n28);
and (n64,n65,n24);
and (n66,n67,n68);
xor (n67,n63,n64);
or (n68,n69,n73);
and (n69,n70,n71);
and (n70,n65,n28);
and (n71,n72,n24);
and (n73,n74,n75);
xor (n74,n70,n71);
or (n75,n76,n80);
and (n76,n77,n78);
and (n77,n72,n28);
and (n78,n79,n24);
and (n80,n81,n82);
xor (n81,n77,n78);
or (n82,n83,n87);
and (n83,n84,n85);
and (n84,n79,n28);
and (n85,n86,n24);
and (n87,n88,n89);
xor (n88,n84,n85);
or (n89,n90,n94);
and (n90,n91,n92);
and (n91,n86,n28);
and (n92,n93,n24);
and (n94,n95,n96);
xor (n95,n91,n92);
and (n96,n97,n98);
and (n97,n93,n28);
and (n98,n99,n24);
and (n100,n23,n101);
or (n102,n103,n106);
and (n103,n104,n105);
xor (n104,n22,n25);
and (n105,n30,n101);
and (n106,n107,n108);
xor (n107,n104,n105);
or (n108,n109,n112);
and (n109,n110,n111);
xor (n110,n32,n33);
and (n111,n37,n101);
and (n112,n113,n114);
xor (n113,n110,n111);
or (n114,n115,n118);
and (n115,n116,n117);
xor (n116,n39,n40);
and (n117,n44,n101);
and (n118,n119,n120);
xor (n119,n116,n117);
or (n120,n121,n124);
and (n121,n122,n123);
xor (n122,n46,n47);
and (n123,n51,n101);
and (n124,n125,n126);
xor (n125,n122,n123);
or (n126,n127,n130);
and (n127,n128,n129);
xor (n128,n53,n54);
and (n129,n58,n101);
and (n130,n131,n132);
xor (n131,n128,n129);
or (n132,n133,n136);
and (n133,n134,n135);
xor (n134,n60,n61);
and (n135,n65,n101);
and (n136,n137,n138);
xor (n137,n134,n135);
or (n138,n139,n142);
and (n139,n140,n141);
xor (n140,n67,n68);
and (n141,n72,n101);
and (n142,n143,n144);
xor (n143,n140,n141);
or (n144,n145,n148);
and (n145,n146,n147);
xor (n146,n74,n75);
and (n147,n79,n101);
and (n148,n149,n150);
xor (n149,n146,n147);
or (n150,n151,n154);
and (n151,n152,n153);
xor (n152,n81,n82);
and (n153,n86,n101);
and (n154,n155,n156);
xor (n155,n152,n153);
or (n156,n157,n160);
and (n157,n158,n159);
xor (n158,n88,n89);
and (n159,n93,n101);
and (n160,n161,n162);
xor (n161,n158,n159);
and (n162,n163,n164);
xor (n163,n95,n96);
and (n164,n99,n101);
and (n165,n30,n166);
or (n167,n168,n171);
and (n168,n169,n170);
xor (n169,n107,n108);
and (n170,n37,n166);
and (n171,n172,n173);
xor (n172,n169,n170);
or (n173,n174,n177);
and (n174,n175,n176);
xor (n175,n113,n114);
and (n176,n44,n166);
and (n177,n178,n179);
xor (n178,n175,n176);
or (n179,n180,n183);
and (n180,n181,n182);
xor (n181,n119,n120);
and (n182,n51,n166);
and (n183,n184,n185);
xor (n184,n181,n182);
or (n185,n186,n189);
and (n186,n187,n188);
xor (n187,n125,n126);
and (n188,n58,n166);
and (n189,n190,n191);
xor (n190,n187,n188);
or (n191,n192,n195);
and (n192,n193,n194);
xor (n193,n131,n132);
and (n194,n65,n166);
and (n195,n196,n197);
xor (n196,n193,n194);
or (n197,n198,n201);
and (n198,n199,n200);
xor (n199,n137,n138);
and (n200,n72,n166);
and (n201,n202,n203);
xor (n202,n199,n200);
or (n203,n204,n207);
and (n204,n205,n206);
xor (n205,n143,n144);
and (n206,n79,n166);
and (n207,n208,n209);
xor (n208,n205,n206);
or (n209,n210,n213);
and (n210,n211,n212);
xor (n211,n149,n150);
and (n212,n86,n166);
and (n213,n214,n215);
xor (n214,n211,n212);
or (n215,n216,n219);
and (n216,n217,n218);
xor (n217,n155,n156);
and (n218,n93,n166);
and (n219,n220,n221);
xor (n220,n217,n218);
and (n221,n222,n223);
xor (n222,n161,n162);
and (n223,n99,n166);
and (n224,n37,n225);
or (n226,n227,n230);
and (n227,n228,n229);
xor (n228,n172,n173);
and (n229,n44,n225);
and (n230,n231,n232);
xor (n231,n228,n229);
or (n232,n233,n236);
and (n233,n234,n235);
xor (n234,n178,n179);
and (n235,n51,n225);
and (n236,n237,n238);
xor (n237,n234,n235);
or (n238,n239,n242);
and (n239,n240,n241);
xor (n240,n184,n185);
and (n241,n58,n225);
and (n242,n243,n244);
xor (n243,n240,n241);
or (n244,n245,n248);
and (n245,n246,n247);
xor (n246,n190,n191);
and (n247,n65,n225);
and (n248,n249,n250);
xor (n249,n246,n247);
or (n250,n251,n254);
and (n251,n252,n253);
xor (n252,n196,n197);
and (n253,n72,n225);
and (n254,n255,n256);
xor (n255,n252,n253);
or (n256,n257,n260);
and (n257,n258,n259);
xor (n258,n202,n203);
and (n259,n79,n225);
and (n260,n261,n262);
xor (n261,n258,n259);
or (n262,n263,n266);
and (n263,n264,n265);
xor (n264,n208,n209);
and (n265,n86,n225);
and (n266,n267,n268);
xor (n267,n264,n265);
or (n268,n269,n272);
and (n269,n270,n271);
xor (n270,n214,n215);
and (n271,n93,n225);
and (n272,n273,n274);
xor (n273,n270,n271);
and (n274,n275,n276);
xor (n275,n220,n221);
and (n276,n99,n225);
and (n277,n44,n278);
or (n279,n280,n283);
and (n280,n281,n282);
xor (n281,n231,n232);
and (n282,n51,n278);
and (n283,n284,n285);
xor (n284,n281,n282);
or (n285,n286,n289);
and (n286,n287,n288);
xor (n287,n237,n238);
and (n288,n58,n278);
and (n289,n290,n291);
xor (n290,n287,n288);
or (n291,n292,n295);
and (n292,n293,n294);
xor (n293,n243,n244);
and (n294,n65,n278);
and (n295,n296,n297);
xor (n296,n293,n294);
or (n297,n298,n301);
and (n298,n299,n300);
xor (n299,n249,n250);
and (n300,n72,n278);
and (n301,n302,n303);
xor (n302,n299,n300);
or (n303,n304,n307);
and (n304,n305,n306);
xor (n305,n255,n256);
and (n306,n79,n278);
and (n307,n308,n309);
xor (n308,n305,n306);
or (n309,n310,n313);
and (n310,n311,n312);
xor (n311,n261,n262);
and (n312,n86,n278);
and (n313,n314,n315);
xor (n314,n311,n312);
or (n315,n316,n319);
and (n316,n317,n318);
xor (n317,n267,n268);
and (n318,n93,n278);
and (n319,n320,n321);
xor (n320,n317,n318);
and (n321,n322,n323);
xor (n322,n273,n274);
and (n323,n99,n278);
and (n324,n51,n325);
or (n326,n327,n330);
and (n327,n328,n329);
xor (n328,n284,n285);
and (n329,n58,n325);
and (n330,n331,n332);
xor (n331,n328,n329);
or (n332,n333,n336);
and (n333,n334,n335);
xor (n334,n290,n291);
and (n335,n65,n325);
and (n336,n337,n338);
xor (n337,n334,n335);
or (n338,n339,n342);
and (n339,n340,n341);
xor (n340,n296,n297);
and (n341,n72,n325);
and (n342,n343,n344);
xor (n343,n340,n341);
or (n344,n345,n348);
and (n345,n346,n347);
xor (n346,n302,n303);
and (n347,n79,n325);
and (n348,n349,n350);
xor (n349,n346,n347);
or (n350,n351,n354);
and (n351,n352,n353);
xor (n352,n308,n309);
and (n353,n86,n325);
and (n354,n355,n356);
xor (n355,n352,n353);
or (n356,n357,n360);
and (n357,n358,n359);
xor (n358,n314,n315);
and (n359,n93,n325);
and (n360,n361,n362);
xor (n361,n358,n359);
and (n362,n363,n364);
xor (n363,n320,n321);
and (n364,n99,n325);
and (n365,n58,n366);
or (n367,n368,n371);
and (n368,n369,n370);
xor (n369,n331,n332);
and (n370,n65,n366);
and (n371,n372,n373);
xor (n372,n369,n370);
or (n373,n374,n377);
and (n374,n375,n376);
xor (n375,n337,n338);
and (n376,n72,n366);
and (n377,n378,n379);
xor (n378,n375,n376);
or (n379,n380,n383);
and (n380,n381,n382);
xor (n381,n343,n344);
and (n382,n79,n366);
and (n383,n384,n385);
xor (n384,n381,n382);
or (n385,n386,n389);
and (n386,n387,n388);
xor (n387,n349,n350);
and (n388,n86,n366);
and (n389,n390,n391);
xor (n390,n387,n388);
or (n391,n392,n395);
and (n392,n393,n394);
xor (n393,n355,n356);
and (n394,n93,n366);
and (n395,n396,n397);
xor (n396,n393,n394);
and (n397,n398,n399);
xor (n398,n361,n362);
and (n399,n99,n366);
and (n400,n65,n401);
or (n402,n403,n406);
and (n403,n404,n405);
xor (n404,n372,n373);
and (n405,n72,n401);
and (n406,n407,n408);
xor (n407,n404,n405);
or (n408,n409,n412);
and (n409,n410,n411);
xor (n410,n378,n379);
and (n411,n79,n401);
and (n412,n413,n414);
xor (n413,n410,n411);
or (n414,n415,n418);
and (n415,n416,n417);
xor (n416,n384,n385);
and (n417,n86,n401);
and (n418,n419,n420);
xor (n419,n416,n417);
or (n420,n421,n424);
and (n421,n422,n423);
xor (n422,n390,n391);
and (n423,n93,n401);
and (n424,n425,n426);
xor (n425,n422,n423);
and (n426,n427,n428);
xor (n427,n396,n397);
and (n428,n99,n401);
and (n429,n72,n430);
or (n431,n432,n435);
and (n432,n433,n434);
xor (n433,n407,n408);
and (n434,n79,n430);
and (n435,n436,n437);
xor (n436,n433,n434);
or (n437,n438,n441);
and (n438,n439,n440);
xor (n439,n413,n414);
and (n440,n86,n430);
and (n441,n442,n443);
xor (n442,n439,n440);
or (n443,n444,n447);
and (n444,n445,n446);
xor (n445,n419,n420);
and (n446,n93,n430);
and (n447,n448,n449);
xor (n448,n445,n446);
and (n449,n450,n451);
xor (n450,n425,n426);
and (n451,n99,n430);
and (n452,n79,n453);
or (n454,n455,n458);
and (n455,n456,n457);
xor (n456,n436,n437);
and (n457,n86,n453);
and (n458,n459,n460);
xor (n459,n456,n457);
or (n460,n461,n464);
and (n461,n462,n463);
xor (n462,n442,n443);
and (n463,n93,n453);
and (n464,n465,n466);
xor (n465,n462,n463);
and (n466,n467,n468);
xor (n467,n448,n449);
and (n468,n99,n453);
and (n469,n86,n470);
or (n471,n472,n475);
and (n472,n473,n474);
xor (n473,n459,n460);
and (n474,n93,n470);
and (n475,n476,n477);
xor (n476,n473,n474);
and (n477,n478,n479);
xor (n478,n465,n466);
and (n479,n99,n470);
xor (n480,n481,n950);
xor (n481,n482,n948);
xor (n482,n483,n933);
xor (n483,n484,n931);
xor (n484,n485,n910);
xor (n485,n486,n908);
xor (n486,n487,n881);
xor (n487,n488,n879);
xor (n488,n489,n846);
xor (n489,n490,n844);
xor (n490,n491,n805);
xor (n491,n492,n803);
xor (n492,n493,n758);
xor (n493,n494,n756);
xor (n494,n495,n705);
xor (n495,n496,n703);
xor (n496,n497,n646);
xor (n497,n498,n644);
xor (n498,n499,n581);
xor (n499,n500,n579);
and (n500,n501,n504);
and (n501,n502,n503);
or (n504,n505,n510);
and (n505,n506,n508);
and (n506,n502,n507);
and (n508,n509,n503);
and (n510,n511,n512);
xor (n511,n506,n508);
or (n512,n513,n517);
and (n513,n514,n515);
and (n514,n509,n507);
and (n515,n516,n503);
and (n517,n518,n519);
xor (n518,n514,n515);
or (n519,n520,n524);
and (n520,n521,n522);
and (n521,n516,n507);
and (n522,n523,n503);
and (n524,n525,n526);
xor (n525,n521,n522);
or (n526,n527,n531);
and (n527,n528,n529);
and (n528,n523,n507);
and (n529,n530,n503);
and (n531,n532,n533);
xor (n532,n528,n529);
or (n533,n534,n538);
and (n534,n535,n536);
and (n535,n530,n507);
and (n536,n537,n503);
and (n538,n539,n540);
xor (n539,n535,n536);
or (n540,n541,n545);
and (n541,n542,n543);
and (n542,n537,n507);
and (n543,n544,n503);
and (n545,n546,n547);
xor (n546,n542,n543);
or (n547,n548,n552);
and (n548,n549,n550);
and (n549,n544,n507);
and (n550,n551,n503);
and (n552,n553,n554);
xor (n553,n549,n550);
or (n554,n555,n559);
and (n555,n556,n557);
and (n556,n551,n507);
and (n557,n558,n503);
and (n559,n560,n561);
xor (n560,n556,n557);
or (n561,n562,n566);
and (n562,n563,n564);
and (n563,n558,n507);
and (n564,n565,n503);
and (n566,n567,n568);
xor (n567,n563,n564);
or (n568,n569,n573);
and (n569,n570,n571);
and (n570,n565,n507);
and (n571,n572,n503);
and (n573,n574,n575);
xor (n574,n570,n571);
and (n575,n576,n577);
and (n576,n572,n507);
and (n577,n578,n503);
and (n579,n502,n580);
or (n581,n582,n585);
and (n582,n583,n584);
xor (n583,n501,n504);
and (n584,n509,n580);
and (n585,n586,n587);
xor (n586,n583,n584);
or (n587,n588,n591);
and (n588,n589,n590);
xor (n589,n511,n512);
and (n590,n516,n580);
and (n591,n592,n593);
xor (n592,n589,n590);
or (n593,n594,n597);
and (n594,n595,n596);
xor (n595,n518,n519);
and (n596,n523,n580);
and (n597,n598,n599);
xor (n598,n595,n596);
or (n599,n600,n603);
and (n600,n601,n602);
xor (n601,n525,n526);
and (n602,n530,n580);
and (n603,n604,n605);
xor (n604,n601,n602);
or (n605,n606,n609);
and (n606,n607,n608);
xor (n607,n532,n533);
and (n608,n537,n580);
and (n609,n610,n611);
xor (n610,n607,n608);
or (n611,n612,n615);
and (n612,n613,n614);
xor (n613,n539,n540);
and (n614,n544,n580);
and (n615,n616,n617);
xor (n616,n613,n614);
or (n617,n618,n621);
and (n618,n619,n620);
xor (n619,n546,n547);
and (n620,n551,n580);
and (n621,n622,n623);
xor (n622,n619,n620);
or (n623,n624,n627);
and (n624,n625,n626);
xor (n625,n553,n554);
and (n626,n558,n580);
and (n627,n628,n629);
xor (n628,n625,n626);
or (n629,n630,n633);
and (n630,n631,n632);
xor (n631,n560,n561);
and (n632,n565,n580);
and (n633,n634,n635);
xor (n634,n631,n632);
or (n635,n636,n639);
and (n636,n637,n638);
xor (n637,n567,n568);
and (n638,n572,n580);
and (n639,n640,n641);
xor (n640,n637,n638);
and (n641,n642,n643);
xor (n642,n574,n575);
and (n643,n578,n580);
and (n644,n509,n645);
or (n646,n647,n650);
and (n647,n648,n649);
xor (n648,n586,n587);
and (n649,n516,n645);
and (n650,n651,n652);
xor (n651,n648,n649);
or (n652,n653,n656);
and (n653,n654,n655);
xor (n654,n592,n593);
and (n655,n523,n645);
and (n656,n657,n658);
xor (n657,n654,n655);
or (n658,n659,n662);
and (n659,n660,n661);
xor (n660,n598,n599);
and (n661,n530,n645);
and (n662,n663,n664);
xor (n663,n660,n661);
or (n664,n665,n668);
and (n665,n666,n667);
xor (n666,n604,n605);
and (n667,n537,n645);
and (n668,n669,n670);
xor (n669,n666,n667);
or (n670,n671,n674);
and (n671,n672,n673);
xor (n672,n610,n611);
and (n673,n544,n645);
and (n674,n675,n676);
xor (n675,n672,n673);
or (n676,n677,n680);
and (n677,n678,n679);
xor (n678,n616,n617);
and (n679,n551,n645);
and (n680,n681,n682);
xor (n681,n678,n679);
or (n682,n683,n686);
and (n683,n684,n685);
xor (n684,n622,n623);
and (n685,n558,n645);
and (n686,n687,n688);
xor (n687,n684,n685);
or (n688,n689,n692);
and (n689,n690,n691);
xor (n690,n628,n629);
and (n691,n565,n645);
and (n692,n693,n694);
xor (n693,n690,n691);
or (n694,n695,n698);
and (n695,n696,n697);
xor (n696,n634,n635);
and (n697,n572,n645);
and (n698,n699,n700);
xor (n699,n696,n697);
and (n700,n701,n702);
xor (n701,n640,n641);
and (n702,n578,n645);
and (n703,n516,n704);
or (n705,n706,n709);
and (n706,n707,n708);
xor (n707,n651,n652);
and (n708,n523,n704);
and (n709,n710,n711);
xor (n710,n707,n708);
or (n711,n712,n715);
and (n712,n713,n714);
xor (n713,n657,n658);
and (n714,n530,n704);
and (n715,n716,n717);
xor (n716,n713,n714);
or (n717,n718,n721);
and (n718,n719,n720);
xor (n719,n663,n664);
and (n720,n537,n704);
and (n721,n722,n723);
xor (n722,n719,n720);
or (n723,n724,n727);
and (n724,n725,n726);
xor (n725,n669,n670);
and (n726,n544,n704);
and (n727,n728,n729);
xor (n728,n725,n726);
or (n729,n730,n733);
and (n730,n731,n732);
xor (n731,n675,n676);
and (n732,n551,n704);
and (n733,n734,n735);
xor (n734,n731,n732);
or (n735,n736,n739);
and (n736,n737,n738);
xor (n737,n681,n682);
and (n738,n558,n704);
and (n739,n740,n741);
xor (n740,n737,n738);
or (n741,n742,n745);
and (n742,n743,n744);
xor (n743,n687,n688);
and (n744,n565,n704);
and (n745,n746,n747);
xor (n746,n743,n744);
or (n747,n748,n751);
and (n748,n749,n750);
xor (n749,n693,n694);
and (n750,n572,n704);
and (n751,n752,n753);
xor (n752,n749,n750);
and (n753,n754,n755);
xor (n754,n699,n700);
and (n755,n578,n704);
and (n756,n523,n757);
or (n758,n759,n762);
and (n759,n760,n761);
xor (n760,n710,n711);
and (n761,n530,n757);
and (n762,n763,n764);
xor (n763,n760,n761);
or (n764,n765,n768);
and (n765,n766,n767);
xor (n766,n716,n717);
and (n767,n537,n757);
and (n768,n769,n770);
xor (n769,n766,n767);
or (n770,n771,n774);
and (n771,n772,n773);
xor (n772,n722,n723);
and (n773,n544,n757);
and (n774,n775,n776);
xor (n775,n772,n773);
or (n776,n777,n780);
and (n777,n778,n779);
xor (n778,n728,n729);
and (n779,n551,n757);
and (n780,n781,n782);
xor (n781,n778,n779);
or (n782,n783,n786);
and (n783,n784,n785);
xor (n784,n734,n735);
and (n785,n558,n757);
and (n786,n787,n788);
xor (n787,n784,n785);
or (n788,n789,n792);
and (n789,n790,n791);
xor (n790,n740,n741);
and (n791,n565,n757);
and (n792,n793,n794);
xor (n793,n790,n791);
or (n794,n795,n798);
and (n795,n796,n797);
xor (n796,n746,n747);
and (n797,n572,n757);
and (n798,n799,n800);
xor (n799,n796,n797);
and (n800,n801,n802);
xor (n801,n752,n753);
and (n802,n578,n757);
and (n803,n530,n804);
or (n805,n806,n809);
and (n806,n807,n808);
xor (n807,n763,n764);
and (n808,n537,n804);
and (n809,n810,n811);
xor (n810,n807,n808);
or (n811,n812,n815);
and (n812,n813,n814);
xor (n813,n769,n770);
and (n814,n544,n804);
and (n815,n816,n817);
xor (n816,n813,n814);
or (n817,n818,n821);
and (n818,n819,n820);
xor (n819,n775,n776);
and (n820,n551,n804);
and (n821,n822,n823);
xor (n822,n819,n820);
or (n823,n824,n827);
and (n824,n825,n826);
xor (n825,n781,n782);
and (n826,n558,n804);
and (n827,n828,n829);
xor (n828,n825,n826);
or (n829,n830,n833);
and (n830,n831,n832);
xor (n831,n787,n788);
and (n832,n565,n804);
and (n833,n834,n835);
xor (n834,n831,n832);
or (n835,n836,n839);
and (n836,n837,n838);
xor (n837,n793,n794);
and (n838,n572,n804);
and (n839,n840,n841);
xor (n840,n837,n838);
and (n841,n842,n843);
xor (n842,n799,n800);
and (n843,n578,n804);
and (n844,n537,n845);
or (n846,n847,n850);
and (n847,n848,n849);
xor (n848,n810,n811);
and (n849,n544,n845);
and (n850,n851,n852);
xor (n851,n848,n849);
or (n852,n853,n856);
and (n853,n854,n855);
xor (n854,n816,n817);
and (n855,n551,n845);
and (n856,n857,n858);
xor (n857,n854,n855);
or (n858,n859,n862);
and (n859,n860,n861);
xor (n860,n822,n823);
and (n861,n558,n845);
and (n862,n863,n864);
xor (n863,n860,n861);
or (n864,n865,n868);
and (n865,n866,n867);
xor (n866,n828,n829);
and (n867,n565,n845);
and (n868,n869,n870);
xor (n869,n866,n867);
or (n870,n871,n874);
and (n871,n872,n873);
xor (n872,n834,n835);
and (n873,n572,n845);
and (n874,n875,n876);
xor (n875,n872,n873);
and (n876,n877,n878);
xor (n877,n840,n841);
and (n878,n578,n845);
and (n879,n544,n880);
or (n881,n882,n885);
and (n882,n883,n884);
xor (n883,n851,n852);
and (n884,n551,n880);
and (n885,n886,n887);
xor (n886,n883,n884);
or (n887,n888,n891);
and (n888,n889,n890);
xor (n889,n857,n858);
and (n890,n558,n880);
and (n891,n892,n893);
xor (n892,n889,n890);
or (n893,n894,n897);
and (n894,n895,n896);
xor (n895,n863,n864);
and (n896,n565,n880);
and (n897,n898,n899);
xor (n898,n895,n896);
or (n899,n900,n903);
and (n900,n901,n902);
xor (n901,n869,n870);
and (n902,n572,n880);
and (n903,n904,n905);
xor (n904,n901,n902);
and (n905,n906,n907);
xor (n906,n875,n876);
and (n907,n578,n880);
and (n908,n551,n909);
or (n910,n911,n914);
and (n911,n912,n913);
xor (n912,n886,n887);
and (n913,n558,n909);
and (n914,n915,n916);
xor (n915,n912,n913);
or (n916,n917,n920);
and (n917,n918,n919);
xor (n918,n892,n893);
and (n919,n565,n909);
and (n920,n921,n922);
xor (n921,n918,n919);
or (n922,n923,n926);
and (n923,n924,n925);
xor (n924,n898,n899);
and (n925,n572,n909);
and (n926,n927,n928);
xor (n927,n924,n925);
and (n928,n929,n930);
xor (n929,n904,n905);
and (n930,n578,n909);
and (n931,n558,n932);
or (n933,n934,n937);
and (n934,n935,n936);
xor (n935,n915,n916);
and (n936,n565,n932);
and (n937,n938,n939);
xor (n938,n935,n936);
or (n939,n940,n943);
and (n940,n941,n942);
xor (n941,n921,n922);
and (n942,n572,n932);
and (n943,n944,n945);
xor (n944,n941,n942);
and (n945,n946,n947);
xor (n946,n927,n928);
and (n947,n578,n932);
and (n948,n565,n949);
or (n950,n951,n954);
and (n951,n952,n953);
xor (n952,n938,n939);
and (n953,n572,n949);
and (n954,n955,n956);
xor (n955,n952,n953);
and (n956,n957,n958);
xor (n957,n944,n945);
and (n958,n578,n949);
xor (n960,n961,n1430);
xor (n961,n962,n1428);
xor (n962,n963,n1413);
xor (n963,n964,n1411);
xor (n964,n965,n1390);
xor (n965,n966,n1388);
xor (n966,n967,n1361);
xor (n967,n968,n1359);
xor (n968,n969,n1326);
xor (n969,n970,n1324);
xor (n970,n971,n1285);
xor (n971,n972,n1283);
xor (n972,n973,n1238);
xor (n973,n974,n1236);
xor (n974,n975,n1185);
xor (n975,n976,n1183);
xor (n976,n977,n1126);
xor (n977,n978,n1124);
xor (n978,n979,n1061);
xor (n979,n980,n1059);
and (n980,n981,n984);
and (n981,n982,n983);
wire s0n982,s1n982,notn982;
or (n982,s0n982,s1n982);
not(notn982,n959);
and (s0n982,notn982,n23);
and (s1n982,n959,n502);
wire s0n983,s1n983,notn983;
or (n983,s0n983,s1n983);
not(notn983,n959);
and (s0n983,notn983,n24);
and (s1n983,n959,n503);
or (n984,n985,n990);
and (n985,n986,n988);
and (n986,n982,n987);
wire s0n987,s1n987,notn987;
or (n987,s0n987,s1n987);
not(notn987,n959);
and (s0n987,notn987,n28);
and (s1n987,n959,n507);
and (n988,n989,n983);
wire s0n989,s1n989,notn989;
or (n989,s0n989,s1n989);
not(notn989,n959);
and (s0n989,notn989,n30);
and (s1n989,n959,n509);
and (n990,n991,n992);
xor (n991,n986,n988);
or (n992,n993,n997);
and (n993,n994,n995);
and (n994,n989,n987);
and (n995,n996,n983);
wire s0n996,s1n996,notn996;
or (n996,s0n996,s1n996);
not(notn996,n959);
and (s0n996,notn996,n37);
and (s1n996,n959,n516);
and (n997,n998,n999);
xor (n998,n994,n995);
or (n999,n1000,n1004);
and (n1000,n1001,n1002);
and (n1001,n996,n987);
and (n1002,n1003,n983);
wire s0n1003,s1n1003,notn1003;
or (n1003,s0n1003,s1n1003);
not(notn1003,n959);
and (s0n1003,notn1003,n44);
and (s1n1003,n959,n523);
and (n1004,n1005,n1006);
xor (n1005,n1001,n1002);
or (n1006,n1007,n1011);
and (n1007,n1008,n1009);
and (n1008,n1003,n987);
and (n1009,n1010,n983);
wire s0n1010,s1n1010,notn1010;
or (n1010,s0n1010,s1n1010);
not(notn1010,n959);
and (s0n1010,notn1010,n51);
and (s1n1010,n959,n530);
and (n1011,n1012,n1013);
xor (n1012,n1008,n1009);
or (n1013,n1014,n1018);
and (n1014,n1015,n1016);
and (n1015,n1010,n987);
and (n1016,n1017,n983);
wire s0n1017,s1n1017,notn1017;
or (n1017,s0n1017,s1n1017);
not(notn1017,n959);
and (s0n1017,notn1017,n58);
and (s1n1017,n959,n537);
and (n1018,n1019,n1020);
xor (n1019,n1015,n1016);
or (n1020,n1021,n1025);
and (n1021,n1022,n1023);
and (n1022,n1017,n987);
and (n1023,n1024,n983);
wire s0n1024,s1n1024,notn1024;
or (n1024,s0n1024,s1n1024);
not(notn1024,n959);
and (s0n1024,notn1024,n65);
and (s1n1024,n959,n544);
and (n1025,n1026,n1027);
xor (n1026,n1022,n1023);
or (n1027,n1028,n1032);
and (n1028,n1029,n1030);
and (n1029,n1024,n987);
and (n1030,n1031,n983);
wire s0n1031,s1n1031,notn1031;
or (n1031,s0n1031,s1n1031);
not(notn1031,n959);
and (s0n1031,notn1031,n72);
and (s1n1031,n959,n551);
and (n1032,n1033,n1034);
xor (n1033,n1029,n1030);
or (n1034,n1035,n1039);
and (n1035,n1036,n1037);
and (n1036,n1031,n987);
and (n1037,n1038,n983);
wire s0n1038,s1n1038,notn1038;
or (n1038,s0n1038,s1n1038);
not(notn1038,n959);
and (s0n1038,notn1038,n79);
and (s1n1038,n959,n558);
and (n1039,n1040,n1041);
xor (n1040,n1036,n1037);
or (n1041,n1042,n1046);
and (n1042,n1043,n1044);
and (n1043,n1038,n987);
and (n1044,n1045,n983);
wire s0n1045,s1n1045,notn1045;
or (n1045,s0n1045,s1n1045);
not(notn1045,n959);
and (s0n1045,notn1045,n86);
and (s1n1045,n959,n565);
and (n1046,n1047,n1048);
xor (n1047,n1043,n1044);
or (n1048,n1049,n1053);
and (n1049,n1050,n1051);
and (n1050,n1045,n987);
and (n1051,n1052,n983);
wire s0n1052,s1n1052,notn1052;
or (n1052,s0n1052,s1n1052);
not(notn1052,n959);
and (s0n1052,notn1052,n93);
and (s1n1052,n959,n572);
and (n1053,n1054,n1055);
xor (n1054,n1050,n1051);
and (n1055,n1056,n1057);
and (n1056,n1052,n987);
and (n1057,n1058,n983);
wire s0n1058,s1n1058,notn1058;
or (n1058,s0n1058,s1n1058);
not(notn1058,n959);
and (s0n1058,notn1058,n99);
and (s1n1058,n959,n578);
and (n1059,n982,n1060);
wire s0n1060,s1n1060,notn1060;
or (n1060,s0n1060,s1n1060);
not(notn1060,n959);
and (s0n1060,notn1060,n101);
and (s1n1060,n959,n580);
or (n1061,n1062,n1065);
and (n1062,n1063,n1064);
xor (n1063,n981,n984);
and (n1064,n989,n1060);
and (n1065,n1066,n1067);
xor (n1066,n1063,n1064);
or (n1067,n1068,n1071);
and (n1068,n1069,n1070);
xor (n1069,n991,n992);
and (n1070,n996,n1060);
and (n1071,n1072,n1073);
xor (n1072,n1069,n1070);
or (n1073,n1074,n1077);
and (n1074,n1075,n1076);
xor (n1075,n998,n999);
and (n1076,n1003,n1060);
and (n1077,n1078,n1079);
xor (n1078,n1075,n1076);
or (n1079,n1080,n1083);
and (n1080,n1081,n1082);
xor (n1081,n1005,n1006);
and (n1082,n1010,n1060);
and (n1083,n1084,n1085);
xor (n1084,n1081,n1082);
or (n1085,n1086,n1089);
and (n1086,n1087,n1088);
xor (n1087,n1012,n1013);
and (n1088,n1017,n1060);
and (n1089,n1090,n1091);
xor (n1090,n1087,n1088);
or (n1091,n1092,n1095);
and (n1092,n1093,n1094);
xor (n1093,n1019,n1020);
and (n1094,n1024,n1060);
and (n1095,n1096,n1097);
xor (n1096,n1093,n1094);
or (n1097,n1098,n1101);
and (n1098,n1099,n1100);
xor (n1099,n1026,n1027);
and (n1100,n1031,n1060);
and (n1101,n1102,n1103);
xor (n1102,n1099,n1100);
or (n1103,n1104,n1107);
and (n1104,n1105,n1106);
xor (n1105,n1033,n1034);
and (n1106,n1038,n1060);
and (n1107,n1108,n1109);
xor (n1108,n1105,n1106);
or (n1109,n1110,n1113);
and (n1110,n1111,n1112);
xor (n1111,n1040,n1041);
and (n1112,n1045,n1060);
and (n1113,n1114,n1115);
xor (n1114,n1111,n1112);
or (n1115,n1116,n1119);
and (n1116,n1117,n1118);
xor (n1117,n1047,n1048);
and (n1118,n1052,n1060);
and (n1119,n1120,n1121);
xor (n1120,n1117,n1118);
and (n1121,n1122,n1123);
xor (n1122,n1054,n1055);
and (n1123,n1058,n1060);
and (n1124,n989,n1125);
wire s0n1125,s1n1125,notn1125;
or (n1125,s0n1125,s1n1125);
not(notn1125,n959);
and (s0n1125,notn1125,n166);
and (s1n1125,n959,n645);
or (n1126,n1127,n1130);
and (n1127,n1128,n1129);
xor (n1128,n1066,n1067);
and (n1129,n996,n1125);
and (n1130,n1131,n1132);
xor (n1131,n1128,n1129);
or (n1132,n1133,n1136);
and (n1133,n1134,n1135);
xor (n1134,n1072,n1073);
and (n1135,n1003,n1125);
and (n1136,n1137,n1138);
xor (n1137,n1134,n1135);
or (n1138,n1139,n1142);
and (n1139,n1140,n1141);
xor (n1140,n1078,n1079);
and (n1141,n1010,n1125);
and (n1142,n1143,n1144);
xor (n1143,n1140,n1141);
or (n1144,n1145,n1148);
and (n1145,n1146,n1147);
xor (n1146,n1084,n1085);
and (n1147,n1017,n1125);
and (n1148,n1149,n1150);
xor (n1149,n1146,n1147);
or (n1150,n1151,n1154);
and (n1151,n1152,n1153);
xor (n1152,n1090,n1091);
and (n1153,n1024,n1125);
and (n1154,n1155,n1156);
xor (n1155,n1152,n1153);
or (n1156,n1157,n1160);
and (n1157,n1158,n1159);
xor (n1158,n1096,n1097);
and (n1159,n1031,n1125);
and (n1160,n1161,n1162);
xor (n1161,n1158,n1159);
or (n1162,n1163,n1166);
and (n1163,n1164,n1165);
xor (n1164,n1102,n1103);
and (n1165,n1038,n1125);
and (n1166,n1167,n1168);
xor (n1167,n1164,n1165);
or (n1168,n1169,n1172);
and (n1169,n1170,n1171);
xor (n1170,n1108,n1109);
and (n1171,n1045,n1125);
and (n1172,n1173,n1174);
xor (n1173,n1170,n1171);
or (n1174,n1175,n1178);
and (n1175,n1176,n1177);
xor (n1176,n1114,n1115);
and (n1177,n1052,n1125);
and (n1178,n1179,n1180);
xor (n1179,n1176,n1177);
and (n1180,n1181,n1182);
xor (n1181,n1120,n1121);
and (n1182,n1058,n1125);
and (n1183,n996,n1184);
wire s0n1184,s1n1184,notn1184;
or (n1184,s0n1184,s1n1184);
not(notn1184,n959);
and (s0n1184,notn1184,n225);
and (s1n1184,n959,n704);
or (n1185,n1186,n1189);
and (n1186,n1187,n1188);
xor (n1187,n1131,n1132);
and (n1188,n1003,n1184);
and (n1189,n1190,n1191);
xor (n1190,n1187,n1188);
or (n1191,n1192,n1195);
and (n1192,n1193,n1194);
xor (n1193,n1137,n1138);
and (n1194,n1010,n1184);
and (n1195,n1196,n1197);
xor (n1196,n1193,n1194);
or (n1197,n1198,n1201);
and (n1198,n1199,n1200);
xor (n1199,n1143,n1144);
and (n1200,n1017,n1184);
and (n1201,n1202,n1203);
xor (n1202,n1199,n1200);
or (n1203,n1204,n1207);
and (n1204,n1205,n1206);
xor (n1205,n1149,n1150);
and (n1206,n1024,n1184);
and (n1207,n1208,n1209);
xor (n1208,n1205,n1206);
or (n1209,n1210,n1213);
and (n1210,n1211,n1212);
xor (n1211,n1155,n1156);
and (n1212,n1031,n1184);
and (n1213,n1214,n1215);
xor (n1214,n1211,n1212);
or (n1215,n1216,n1219);
and (n1216,n1217,n1218);
xor (n1217,n1161,n1162);
and (n1218,n1038,n1184);
and (n1219,n1220,n1221);
xor (n1220,n1217,n1218);
or (n1221,n1222,n1225);
and (n1222,n1223,n1224);
xor (n1223,n1167,n1168);
and (n1224,n1045,n1184);
and (n1225,n1226,n1227);
xor (n1226,n1223,n1224);
or (n1227,n1228,n1231);
and (n1228,n1229,n1230);
xor (n1229,n1173,n1174);
and (n1230,n1052,n1184);
and (n1231,n1232,n1233);
xor (n1232,n1229,n1230);
and (n1233,n1234,n1235);
xor (n1234,n1179,n1180);
and (n1235,n1058,n1184);
and (n1236,n1003,n1237);
wire s0n1237,s1n1237,notn1237;
or (n1237,s0n1237,s1n1237);
not(notn1237,n959);
and (s0n1237,notn1237,n278);
and (s1n1237,n959,n757);
or (n1238,n1239,n1242);
and (n1239,n1240,n1241);
xor (n1240,n1190,n1191);
and (n1241,n1010,n1237);
and (n1242,n1243,n1244);
xor (n1243,n1240,n1241);
or (n1244,n1245,n1248);
and (n1245,n1246,n1247);
xor (n1246,n1196,n1197);
and (n1247,n1017,n1237);
and (n1248,n1249,n1250);
xor (n1249,n1246,n1247);
or (n1250,n1251,n1254);
and (n1251,n1252,n1253);
xor (n1252,n1202,n1203);
and (n1253,n1024,n1237);
and (n1254,n1255,n1256);
xor (n1255,n1252,n1253);
or (n1256,n1257,n1260);
and (n1257,n1258,n1259);
xor (n1258,n1208,n1209);
and (n1259,n1031,n1237);
and (n1260,n1261,n1262);
xor (n1261,n1258,n1259);
or (n1262,n1263,n1266);
and (n1263,n1264,n1265);
xor (n1264,n1214,n1215);
and (n1265,n1038,n1237);
and (n1266,n1267,n1268);
xor (n1267,n1264,n1265);
or (n1268,n1269,n1272);
and (n1269,n1270,n1271);
xor (n1270,n1220,n1221);
and (n1271,n1045,n1237);
and (n1272,n1273,n1274);
xor (n1273,n1270,n1271);
or (n1274,n1275,n1278);
and (n1275,n1276,n1277);
xor (n1276,n1226,n1227);
and (n1277,n1052,n1237);
and (n1278,n1279,n1280);
xor (n1279,n1276,n1277);
and (n1280,n1281,n1282);
xor (n1281,n1232,n1233);
and (n1282,n1058,n1237);
and (n1283,n1010,n1284);
wire s0n1284,s1n1284,notn1284;
or (n1284,s0n1284,s1n1284);
not(notn1284,n959);
and (s0n1284,notn1284,n325);
and (s1n1284,n959,n804);
or (n1285,n1286,n1289);
and (n1286,n1287,n1288);
xor (n1287,n1243,n1244);
and (n1288,n1017,n1284);
and (n1289,n1290,n1291);
xor (n1290,n1287,n1288);
or (n1291,n1292,n1295);
and (n1292,n1293,n1294);
xor (n1293,n1249,n1250);
and (n1294,n1024,n1284);
and (n1295,n1296,n1297);
xor (n1296,n1293,n1294);
or (n1297,n1298,n1301);
and (n1298,n1299,n1300);
xor (n1299,n1255,n1256);
and (n1300,n1031,n1284);
and (n1301,n1302,n1303);
xor (n1302,n1299,n1300);
or (n1303,n1304,n1307);
and (n1304,n1305,n1306);
xor (n1305,n1261,n1262);
and (n1306,n1038,n1284);
and (n1307,n1308,n1309);
xor (n1308,n1305,n1306);
or (n1309,n1310,n1313);
and (n1310,n1311,n1312);
xor (n1311,n1267,n1268);
and (n1312,n1045,n1284);
and (n1313,n1314,n1315);
xor (n1314,n1311,n1312);
or (n1315,n1316,n1319);
and (n1316,n1317,n1318);
xor (n1317,n1273,n1274);
and (n1318,n1052,n1284);
and (n1319,n1320,n1321);
xor (n1320,n1317,n1318);
and (n1321,n1322,n1323);
xor (n1322,n1279,n1280);
and (n1323,n1058,n1284);
and (n1324,n1017,n1325);
wire s0n1325,s1n1325,notn1325;
or (n1325,s0n1325,s1n1325);
not(notn1325,n959);
and (s0n1325,notn1325,n366);
and (s1n1325,n959,n845);
or (n1326,n1327,n1330);
and (n1327,n1328,n1329);
xor (n1328,n1290,n1291);
and (n1329,n1024,n1325);
and (n1330,n1331,n1332);
xor (n1331,n1328,n1329);
or (n1332,n1333,n1336);
and (n1333,n1334,n1335);
xor (n1334,n1296,n1297);
and (n1335,n1031,n1325);
and (n1336,n1337,n1338);
xor (n1337,n1334,n1335);
or (n1338,n1339,n1342);
and (n1339,n1340,n1341);
xor (n1340,n1302,n1303);
and (n1341,n1038,n1325);
and (n1342,n1343,n1344);
xor (n1343,n1340,n1341);
or (n1344,n1345,n1348);
and (n1345,n1346,n1347);
xor (n1346,n1308,n1309);
and (n1347,n1045,n1325);
and (n1348,n1349,n1350);
xor (n1349,n1346,n1347);
or (n1350,n1351,n1354);
and (n1351,n1352,n1353);
xor (n1352,n1314,n1315);
and (n1353,n1052,n1325);
and (n1354,n1355,n1356);
xor (n1355,n1352,n1353);
and (n1356,n1357,n1358);
xor (n1357,n1320,n1321);
and (n1358,n1058,n1325);
and (n1359,n1024,n1360);
wire s0n1360,s1n1360,notn1360;
or (n1360,s0n1360,s1n1360);
not(notn1360,n959);
and (s0n1360,notn1360,n401);
and (s1n1360,n959,n880);
or (n1361,n1362,n1365);
and (n1362,n1363,n1364);
xor (n1363,n1331,n1332);
and (n1364,n1031,n1360);
and (n1365,n1366,n1367);
xor (n1366,n1363,n1364);
or (n1367,n1368,n1371);
and (n1368,n1369,n1370);
xor (n1369,n1337,n1338);
and (n1370,n1038,n1360);
and (n1371,n1372,n1373);
xor (n1372,n1369,n1370);
or (n1373,n1374,n1377);
and (n1374,n1375,n1376);
xor (n1375,n1343,n1344);
and (n1376,n1045,n1360);
and (n1377,n1378,n1379);
xor (n1378,n1375,n1376);
or (n1379,n1380,n1383);
and (n1380,n1381,n1382);
xor (n1381,n1349,n1350);
and (n1382,n1052,n1360);
and (n1383,n1384,n1385);
xor (n1384,n1381,n1382);
and (n1385,n1386,n1387);
xor (n1386,n1355,n1356);
and (n1387,n1058,n1360);
and (n1388,n1031,n1389);
wire s0n1389,s1n1389,notn1389;
or (n1389,s0n1389,s1n1389);
not(notn1389,n959);
and (s0n1389,notn1389,n430);
and (s1n1389,n959,n909);
or (n1390,n1391,n1394);
and (n1391,n1392,n1393);
xor (n1392,n1366,n1367);
and (n1393,n1038,n1389);
and (n1394,n1395,n1396);
xor (n1395,n1392,n1393);
or (n1396,n1397,n1400);
and (n1397,n1398,n1399);
xor (n1398,n1372,n1373);
and (n1399,n1045,n1389);
and (n1400,n1401,n1402);
xor (n1401,n1398,n1399);
or (n1402,n1403,n1406);
and (n1403,n1404,n1405);
xor (n1404,n1378,n1379);
and (n1405,n1052,n1389);
and (n1406,n1407,n1408);
xor (n1407,n1404,n1405);
and (n1408,n1409,n1410);
xor (n1409,n1384,n1385);
and (n1410,n1058,n1389);
and (n1411,n1038,n1412);
wire s0n1412,s1n1412,notn1412;
or (n1412,s0n1412,s1n1412);
not(notn1412,n959);
and (s0n1412,notn1412,n453);
and (s1n1412,n959,n932);
or (n1413,n1414,n1417);
and (n1414,n1415,n1416);
xor (n1415,n1395,n1396);
and (n1416,n1045,n1412);
and (n1417,n1418,n1419);
xor (n1418,n1415,n1416);
or (n1419,n1420,n1423);
and (n1420,n1421,n1422);
xor (n1421,n1401,n1402);
and (n1422,n1052,n1412);
and (n1423,n1424,n1425);
xor (n1424,n1421,n1422);
and (n1425,n1426,n1427);
xor (n1426,n1407,n1408);
and (n1427,n1058,n1412);
and (n1428,n1045,n1429);
wire s0n1429,s1n1429,notn1429;
or (n1429,s0n1429,s1n1429);
not(notn1429,n959);
and (s0n1429,notn1429,n470);
and (s1n1429,n959,n949);
or (n1430,n1431,n1434);
and (n1431,n1432,n1433);
xor (n1432,n1418,n1419);
and (n1433,n1052,n1429);
and (n1434,n1435,n1436);
xor (n1435,n1432,n1433);
and (n1436,n1437,n1438);
xor (n1437,n1424,n1425);
and (n1438,n1058,n1429);
endmodule
