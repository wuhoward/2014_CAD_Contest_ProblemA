module top (out,n2,n4,n5,n25,n27,n33,n35,n45,n53
        ,n54,n60,n61,n69,n81,n86,n90,n96,n105,n106
        ,n108,n113,n114,n118,n125,n133,n139,n148,n159,n165
        ,n174,n182,n184,n189,n195,n209,n220,n227);
output out;
input n2;
input n4;
input n5;
input n25;
input n27;
input n33;
input n35;
input n45;
input n53;
input n54;
input n60;
input n61;
input n69;
input n81;
input n86;
input n90;
input n96;
input n105;
input n106;
input n108;
input n113;
input n114;
input n118;
input n125;
input n133;
input n139;
input n148;
input n159;
input n165;
input n174;
input n182;
input n184;
input n189;
input n195;
input n209;
input n220;
input n227;
wire n0;
wire n1;
wire n3;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n24;
wire n26;
wire n28;
wire n29;
wire n30;
wire n31;
wire n32;
wire n34;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n82;
wire n83;
wire n84;
wire n85;
wire n87;
wire n88;
wire n89;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n107;
wire n109;
wire n110;
wire n111;
wire n112;
wire n115;
wire n116;
wire n117;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n183;
wire n185;
wire n186;
wire n187;
wire n188;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
xnor (out,n0,n1016);
nor (n0,n1,n6);
and (n1,n2,n3);
nor (n3,n4,n5);
and (n6,n7,n1013);
nand (n7,n8,n1012);
or (n8,n9,n501);
not (n9,n10);
nand (n10,n11,n500);
not (n11,n12);
nor (n12,n13,n441);
xor (n13,n14,n371);
xor (n14,n15,n229);
xor (n15,n16,n151);
xor (n16,n17,n99);
xor (n17,n18,n75);
xor (n18,n19,n47);
nand (n19,n20,n41);
or (n20,n21,n29);
not (n21,n22);
nor (n22,n23,n28);
and (n23,n24,n26);
not (n24,n25);
not (n26,n27);
and (n28,n25,n27);
not (n29,n30);
nor (n30,n31,n37);
nand (n31,n32,n36);
or (n32,n33,n34);
not (n34,n35);
nand (n36,n33,n34);
nor (n37,n38,n40);
and (n38,n39,n27);
not (n39,n33);
and (n40,n33,n26);
nand (n41,n31,n42);
nand (n42,n43,n46);
or (n43,n44,n27);
not (n44,n45);
or (n46,n26,n45);
nand (n47,n48,n64);
or (n48,n49,n56);
not (n49,n50);
nand (n50,n51,n55);
or (n51,n52,n54);
not (n52,n53);
nand (n55,n54,n52);
not (n56,n57);
nand (n57,n58,n62);
or (n58,n59,n61);
not (n59,n60);
or (n62,n63,n60);
not (n63,n61);
nand (n64,n65,n71);
not (n65,n66);
nor (n66,n67,n70);
and (n67,n61,n68);
not (n68,n69);
and (n70,n63,n69);
and (n71,n49,n72);
nand (n72,n73,n74);
nand (n73,n61,n52);
nand (n74,n53,n63);
nand (n75,n76,n93);
or (n76,n77,n88);
nand (n77,n78,n83);
nor (n78,n79,n82);
and (n79,n80,n61);
not (n80,n81);
and (n82,n81,n63);
nor (n83,n84,n87);
and (n84,n80,n85);
not (n85,n86);
and (n87,n81,n86);
nor (n88,n89,n91);
and (n89,n90,n85);
and (n91,n86,n92);
not (n92,n90);
or (n93,n94,n78);
nor (n94,n95,n97);
and (n95,n96,n85);
and (n97,n86,n98);
not (n98,n96);
xor (n99,n100,n127);
xor (n100,n101,n109);
and (n101,n102,n108);
nand (n102,n103,n107);
or (n103,n104,n106);
not (n104,n105);
nand (n107,n106,n104);
nand (n109,n110,n121);
or (n110,n111,n115);
nand (n111,n112,n114);
not (n112,n113);
nor (n115,n116,n119);
and (n116,n117,n118);
not (n117,n114);
and (n119,n114,n120);
not (n120,n118);
nand (n121,n122,n113);
nor (n122,n123,n126);
and (n123,n124,n117);
not (n124,n125);
and (n126,n125,n114);
nand (n127,n128,n141);
or (n128,n129,n135);
not (n129,n130);
nor (n130,n131,n134);
and (n131,n132,n34);
not (n132,n133);
and (n134,n133,n35);
not (n135,n136);
nand (n136,n137,n140);
or (n137,n138,n114);
not (n138,n139);
nand (n140,n114,n138);
or (n141,n142,n146);
nand (n142,n135,n143);
nand (n143,n144,n145);
or (n144,n138,n35);
nand (n145,n138,n35);
nor (n146,n147,n149);
and (n147,n34,n148);
and (n149,n35,n150);
not (n150,n148);
xor (n151,n152,n203);
xor (n152,n153,n176);
nand (n153,n154,n170);
or (n154,n155,n161);
not (n155,n156);
nor (n156,n157,n160);
and (n157,n158,n104);
not (n158,n159);
and (n160,n159,n105);
nand (n161,n162,n167);
not (n162,n163);
nand (n163,n164,n166);
or (n164,n85,n165);
nand (n166,n165,n85);
nand (n167,n168,n169);
or (n168,n165,n104);
nand (n169,n104,n165);
nand (n170,n163,n171);
nor (n171,n172,n175);
and (n172,n173,n104);
not (n173,n174);
and (n175,n174,n105);
nand (n176,n177,n191);
or (n177,n178,n186);
not (n178,n179);
nor (n179,n180,n185);
and (n180,n181,n183);
not (n181,n182);
not (n183,n184);
and (n185,n182,n184);
not (n186,n187);
nand (n187,n188,n190);
or (n188,n26,n189);
nand (n190,n189,n26);
nand (n191,n192,n198);
not (n192,n193);
nor (n193,n194,n196);
and (n194,n183,n195);
and (n196,n184,n197);
not (n197,n195);
not (n198,n199);
nand (n199,n200,n186);
nand (n200,n201,n202);
or (n201,n189,n183);
nand (n202,n183,n189);
nand (n203,n204,n222);
or (n204,n205,n216);
not (n205,n206);
nor (n206,n207,n211);
nand (n207,n208,n210);
or (n208,n183,n209);
nand (n210,n183,n209);
nor (n211,n212,n214);
and (n212,n213,n209);
not (n213,n54);
and (n214,n54,n215);
not (n215,n209);
not (n216,n217);
nor (n217,n218,n221);
and (n218,n219,n213);
not (n219,n220);
and (n221,n220,n54);
or (n222,n223,n224);
not (n223,n207);
nor (n224,n225,n228);
and (n225,n226,n54);
not (n226,n227);
and (n228,n227,n213);
or (n229,n230,n370);
and (n230,n231,n309);
xor (n231,n232,n272);
or (n232,n233,n271);
and (n233,n234,n254);
xor (n234,n235,n245);
nand (n235,n236,n241);
or (n236,n237,n238);
not (n237,n71);
nor (n238,n239,n240);
and (n239,n63,n90);
and (n240,n61,n92);
or (n241,n49,n242);
nor (n242,n243,n244);
and (n243,n63,n96);
and (n244,n61,n98);
nand (n245,n246,n250);
or (n246,n77,n247);
nor (n247,n248,n249);
and (n248,n85,n159);
and (n249,n86,n158);
or (n250,n78,n251);
nor (n251,n252,n253);
and (n252,n85,n174);
and (n253,n86,n173);
and (n254,n255,n261);
nor (n255,n256,n85);
nor (n256,n257,n259);
and (n257,n258,n63);
nand (n258,n108,n81);
and (n259,n260,n80);
not (n260,n108);
nand (n261,n262,n267);
or (n262,n111,n263);
not (n263,n264);
nor (n264,n265,n266);
and (n265,n44,n117);
and (n266,n45,n114);
or (n267,n268,n112);
nor (n268,n269,n270);
and (n269,n117,n148);
and (n270,n114,n150);
and (n271,n235,n245);
xor (n272,n273,n291);
xor (n273,n274,n277);
nand (n274,n275,n276);
or (n275,n77,n251);
or (n276,n78,n88);
xor (n277,n278,n284);
nor (n278,n279,n104);
nor (n279,n280,n282);
and (n280,n281,n85);
nand (n281,n108,n165);
and (n282,n260,n283);
not (n283,n165);
nand (n284,n285,n290);
or (n285,n111,n286);
not (n286,n287);
nor (n287,n288,n289);
and (n288,n133,n114);
and (n289,n132,n117);
or (n290,n115,n112);
or (n291,n292,n308);
and (n292,n293,n298);
xor (n293,n294,n295);
nor (n294,n162,n260);
nand (n295,n296,n297);
or (n296,n112,n286);
or (n297,n268,n111);
nand (n298,n299,n303);
or (n299,n142,n300);
nor (n300,n301,n302);
and (n301,n25,n34);
and (n302,n24,n35);
or (n303,n135,n304);
not (n304,n305);
nor (n305,n306,n307);
and (n306,n45,n35);
and (n307,n44,n34);
and (n308,n294,n295);
or (n309,n310,n369);
and (n310,n311,n368);
xor (n311,n312,n342);
or (n312,n313,n341);
and (n313,n314,n332);
xor (n314,n315,n322);
nand (n315,n316,n320);
or (n316,n142,n317);
nor (n317,n318,n319);
and (n318,n182,n34);
and (n319,n181,n35);
nand (n320,n321,n136);
not (n321,n300);
nand (n322,n323,n328);
or (n323,n324,n186);
not (n324,n325);
nor (n325,n326,n327);
and (n326,n220,n184);
and (n327,n219,n183);
or (n328,n199,n329);
nor (n329,n330,n331);
and (n330,n59,n184);
and (n331,n60,n183);
nand (n332,n333,n337);
or (n333,n205,n334);
nor (n334,n335,n336);
and (n335,n213,n96);
and (n336,n98,n54);
or (n337,n223,n338);
nor (n338,n339,n340);
and (n339,n213,n69);
and (n340,n54,n68);
and (n341,n315,n322);
or (n342,n343,n367);
and (n343,n344,n361);
xor (n344,n345,n355);
nand (n345,n346,n350);
or (n346,n347,n29);
nor (n347,n348,n349);
and (n348,n26,n227);
and (n349,n27,n226);
nand (n350,n351,n31);
not (n351,n352);
nor (n352,n353,n354);
and (n353,n26,n195);
and (n354,n27,n197);
nand (n355,n356,n360);
or (n356,n237,n357);
nor (n357,n358,n359);
and (n358,n63,n174);
and (n359,n61,n173);
or (n360,n49,n238);
nand (n361,n362,n366);
or (n362,n77,n363);
nor (n363,n364,n365);
and (n364,n260,n86);
and (n365,n108,n85);
or (n366,n247,n78);
and (n367,n345,n355);
xor (n368,n293,n298);
and (n369,n312,n342);
and (n370,n232,n272);
xor (n371,n372,n422);
xor (n372,n373,n376);
or (n373,n374,n375);
and (n374,n273,n291);
and (n375,n274,n277);
xor (n376,n377,n401);
xor (n377,n378,n379);
and (n378,n278,n284);
or (n379,n380,n400);
and (n380,n381,n393);
xor (n381,n382,n386);
nand (n382,n383,n384);
or (n383,n304,n142);
nand (n384,n385,n136);
not (n385,n146);
nand (n386,n387,n392);
or (n387,n388,n161);
not (n388,n389);
nand (n389,n390,n391);
or (n390,n104,n108);
or (n391,n260,n105);
nand (n392,n163,n156);
nand (n393,n394,n399);
or (n394,n199,n395);
not (n395,n396);
nor (n396,n397,n398);
and (n397,n227,n184);
and (n398,n226,n183);
or (n399,n186,n193);
and (n400,n382,n386);
or (n401,n402,n421);
and (n402,n403,n418);
xor (n403,n404,n411);
nand (n404,n405,n410);
or (n405,n406,n205);
not (n406,n407);
nor (n407,n408,n409);
and (n408,n59,n213);
and (n409,n60,n54);
nand (n410,n207,n217);
nand (n411,n412,n414);
or (n412,n21,n413);
not (n413,n31);
or (n414,n29,n415);
nor (n415,n416,n417);
and (n416,n26,n182);
and (n417,n27,n181);
nand (n418,n419,n420);
or (n419,n237,n242);
or (n420,n49,n66);
and (n421,n404,n411);
or (n422,n423,n440);
and (n423,n424,n439);
xor (n424,n425,n438);
or (n425,n426,n437);
and (n426,n427,n434);
xor (n427,n428,n431);
nand (n428,n429,n430);
or (n429,n324,n199);
nand (n430,n187,n396);
nand (n431,n432,n433);
or (n432,n205,n338);
nand (n433,n207,n407);
nand (n434,n435,n436);
or (n435,n29,n352);
or (n436,n413,n415);
and (n437,n428,n431);
xor (n438,n403,n418);
xor (n439,n381,n393);
and (n440,n425,n438);
or (n441,n442,n499);
and (n442,n443,n498);
xor (n443,n444,n445);
xor (n444,n424,n439);
or (n445,n446,n497);
and (n446,n447,n450);
xor (n447,n448,n449);
xor (n448,n427,n434);
xor (n449,n234,n254);
or (n450,n451,n496);
and (n451,n452,n471);
xor (n452,n453,n454);
xor (n453,n255,n261);
or (n454,n455,n470);
and (n455,n456,n463);
xor (n456,n457,n458);
nor (n457,n78,n260);
nand (n458,n459,n461);
or (n459,n142,n460);
xor (n460,n195,n34);
nand (n461,n462,n136);
not (n462,n317);
nand (n463,n464,n469);
or (n464,n199,n465);
not (n465,n466);
nor (n466,n467,n468);
and (n467,n68,n183);
and (n468,n69,n184);
or (n469,n186,n329);
and (n470,n457,n458);
or (n471,n472,n495);
and (n472,n473,n489);
xor (n473,n474,n482);
nand (n474,n475,n480);
or (n475,n476,n205);
not (n476,n477);
nand (n477,n478,n479);
or (n478,n54,n92);
or (n479,n90,n213);
nand (n480,n481,n207);
not (n481,n334);
nand (n482,n483,n488);
or (n483,n111,n484);
not (n484,n485);
nor (n485,n486,n487);
and (n486,n24,n117);
and (n487,n25,n114);
nand (n488,n264,n113);
nand (n489,n490,n494);
or (n490,n237,n491);
nor (n491,n492,n493);
and (n492,n63,n159);
and (n493,n61,n158);
or (n494,n49,n357);
and (n495,n474,n482);
and (n496,n453,n454);
and (n497,n448,n449);
xor (n498,n231,n309);
and (n499,n444,n445);
nand (n500,n13,n441);
not (n501,n502);
nand (n502,n503,n718);
nor (n503,n504,n717);
and (n504,n505,n569);
nand (n505,n506,n508);
not (n506,n507);
xor (n507,n443,n498);
not (n508,n509);
or (n509,n510,n568);
and (n510,n511,n514);
xor (n511,n512,n513);
xor (n512,n311,n368);
xor (n513,n447,n450);
or (n514,n515,n567);
and (n515,n516,n519);
xor (n516,n517,n518);
xor (n517,n344,n361);
xor (n518,n314,n332);
or (n519,n520,n566);
and (n520,n521,n542);
xor (n521,n522,n528);
nand (n522,n523,n527);
or (n523,n29,n524);
nor (n524,n525,n526);
and (n525,n26,n220);
and (n526,n27,n219);
or (n527,n413,n347);
and (n528,n529,n535);
nand (n529,n530,n531);
or (n530,n460,n135);
or (n531,n142,n532);
nor (n532,n533,n534);
and (n533,n227,n34);
and (n534,n226,n35);
not (n535,n536);
nand (n536,n537,n61);
nand (n537,n538,n539);
or (n538,n108,n53);
nand (n539,n540,n213);
not (n540,n541);
and (n541,n108,n53);
or (n542,n543,n565);
and (n543,n544,n559);
xor (n544,n545,n552);
nand (n545,n546,n551);
or (n546,n547,n199);
not (n547,n548);
nand (n548,n549,n550);
or (n549,n184,n98);
or (n550,n183,n96);
nand (n551,n187,n466);
nand (n552,n553,n558);
or (n553,n554,n205);
not (n554,n555);
nand (n555,n556,n557);
or (n556,n54,n173);
or (n557,n213,n174);
nand (n558,n207,n477);
nand (n559,n560,n561);
or (n560,n112,n484);
or (n561,n562,n111);
nor (n562,n563,n564);
and (n563,n117,n182);
and (n564,n114,n181);
and (n565,n545,n552);
and (n566,n522,n528);
and (n567,n517,n518);
and (n568,n512,n513);
nand (n569,n570,n716);
or (n570,n571,n708);
not (n571,n572);
nand (n572,n573,n707);
or (n573,n574,n657);
nor (n574,n575,n605);
xor (n575,n576,n604);
xor (n576,n577,n578);
xor (n577,n452,n471);
or (n578,n579,n603);
and (n579,n580,n583);
xor (n580,n581,n582);
xor (n581,n473,n489);
xor (n582,n456,n463);
or (n583,n584,n602);
and (n584,n585,n598);
xor (n585,n586,n592);
nand (n586,n587,n591);
or (n587,n237,n588);
nor (n588,n589,n590);
and (n589,n260,n61);
and (n590,n108,n63);
or (n591,n49,n491);
nand (n592,n593,n597);
or (n593,n29,n594);
nor (n594,n595,n596);
and (n595,n26,n60);
and (n596,n27,n59);
or (n597,n413,n524);
nand (n598,n599,n601);
or (n599,n535,n600);
not (n600,n529);
or (n601,n529,n536);
and (n602,n586,n592);
and (n603,n581,n582);
xor (n604,n516,n519);
or (n605,n606,n656);
and (n606,n607,n655);
xor (n607,n608,n609);
xor (n608,n521,n542);
or (n609,n610,n654);
and (n610,n611,n653);
xor (n611,n612,n630);
or (n612,n613,n629);
and (n613,n614,n623);
xor (n614,n615,n616);
nor (n615,n49,n260);
nand (n616,n617,n621);
or (n617,n618,n142);
nor (n618,n619,n620);
and (n619,n34,n220);
and (n620,n35,n219);
nand (n621,n622,n136);
not (n622,n532);
nand (n623,n624,n625);
or (n624,n547,n186);
or (n625,n199,n626);
nor (n626,n627,n628);
and (n627,n183,n90);
and (n628,n184,n92);
and (n629,n615,n616);
or (n630,n631,n652);
and (n631,n632,n646);
xor (n632,n633,n640);
nand (n633,n634,n639);
or (n634,n635,n205);
not (n635,n636);
nand (n636,n637,n638);
or (n637,n54,n158);
or (n638,n213,n159);
nand (n639,n207,n555);
nand (n640,n641,n645);
or (n641,n642,n111);
nor (n642,n643,n644);
and (n643,n117,n195);
and (n644,n114,n197);
or (n645,n562,n112);
nand (n646,n647,n651);
or (n647,n29,n648);
nor (n648,n649,n650);
and (n649,n26,n69);
and (n650,n27,n68);
or (n651,n413,n594);
and (n652,n633,n640);
xor (n653,n544,n559);
and (n654,n612,n630);
xor (n655,n580,n583);
and (n656,n608,n609);
nand (n657,n658,n706);
or (n658,n659,n705);
and (n659,n660,n663);
xor (n660,n661,n662);
xor (n661,n585,n598);
xor (n662,n611,n653);
or (n663,n664,n704);
and (n664,n665,n703);
xor (n665,n666,n679);
and (n666,n667,n673);
and (n667,n668,n54);
nand (n668,n669,n670);
or (n669,n108,n209);
nand (n670,n671,n183);
not (n671,n672);
and (n672,n108,n209);
nand (n673,n674,n678);
or (n674,n142,n675);
nor (n675,n676,n677);
and (n676,n34,n60);
and (n677,n35,n59);
or (n678,n135,n618);
or (n679,n680,n702);
and (n680,n681,n696);
xor (n681,n682,n689);
nand (n682,n683,n687);
or (n683,n684,n199);
nor (n684,n685,n686);
and (n685,n183,n174);
and (n686,n184,n173);
nand (n687,n688,n187);
not (n688,n626);
nand (n689,n690,n691);
or (n690,n635,n223);
nand (n691,n692,n206);
not (n692,n693);
nor (n693,n694,n695);
and (n694,n260,n54);
and (n695,n213,n108);
nand (n696,n697,n701);
or (n697,n111,n698);
nor (n698,n699,n700);
and (n699,n117,n227);
and (n700,n114,n226);
or (n701,n642,n112);
and (n702,n682,n689);
xor (n703,n614,n623);
and (n704,n666,n679);
and (n705,n661,n662);
xor (n706,n607,n655);
nand (n707,n575,n605);
not (n708,n709);
nand (n709,n710,n712);
not (n710,n711);
xor (n711,n511,n514);
not (n712,n713);
or (n713,n714,n715);
and (n714,n576,n604);
and (n715,n577,n578);
nand (n716,n711,n713);
nor (n717,n506,n508);
nand (n718,n719,n505,n1008);
nand (n719,n720,n1007);
or (n720,n721,n758);
not (n721,n722);
or (n722,n723,n724);
xor (n723,n660,n663);
or (n724,n725,n757);
and (n725,n726,n756);
xor (n726,n727,n728);
xor (n727,n632,n646);
or (n728,n729,n755);
and (n729,n730,n738);
xor (n730,n731,n737);
nand (n731,n732,n736);
or (n732,n29,n733);
nor (n733,n734,n735);
and (n734,n26,n96);
and (n735,n27,n98);
or (n736,n413,n648);
xor (n737,n667,n673);
or (n738,n739,n754);
and (n739,n740,n748);
xor (n740,n741,n742);
nor (n741,n223,n260);
nand (n742,n743,n747);
or (n743,n744,n111);
nor (n744,n745,n746);
and (n745,n219,n114);
and (n746,n220,n117);
or (n747,n698,n112);
nand (n748,n749,n753);
or (n749,n199,n750);
nor (n750,n751,n752);
and (n751,n183,n159);
and (n752,n184,n158);
or (n753,n186,n684);
and (n754,n741,n742);
and (n755,n731,n737);
xor (n756,n665,n703);
and (n757,n727,n728);
not (n758,n759);
or (n759,n760,n1006);
and (n760,n761,n801);
xor (n761,n762,n800);
or (n762,n763,n799);
and (n763,n764,n798);
xor (n764,n765,n766);
xor (n765,n681,n696);
or (n766,n767,n797);
and (n767,n768,n783);
xor (n768,n769,n777);
nand (n769,n770,n775);
or (n770,n771,n142);
not (n771,n772);
nand (n772,n773,n774);
or (n773,n35,n68);
or (n774,n34,n69);
nand (n775,n776,n136);
not (n776,n675);
nand (n777,n778,n782);
or (n778,n29,n779);
nor (n779,n780,n781);
and (n780,n26,n90);
and (n781,n27,n92);
or (n782,n413,n733);
and (n783,n784,n790);
nor (n784,n785,n183);
nor (n785,n786,n788);
and (n786,n260,n787);
not (n787,n189);
nor (n788,n789,n27);
and (n789,n108,n189);
nand (n790,n791,n796);
or (n791,n111,n792);
not (n792,n793);
nor (n793,n794,n795);
and (n794,n59,n117);
and (n795,n60,n114);
or (n796,n744,n112);
and (n797,n769,n777);
xor (n798,n730,n738);
and (n799,n765,n766);
xor (n800,n726,n756);
nand (n801,n802,n1003,n1005);
nand (n802,n803,n838,n998);
nand (n803,n804,n806);
not (n804,n805);
xor (n805,n764,n798);
not (n806,n807);
or (n807,n808,n837);
and (n808,n809,n836);
xor (n809,n810,n835);
or (n810,n811,n834);
and (n811,n812,n828);
xor (n812,n813,n821);
nand (n813,n814,n819);
or (n814,n815,n199);
not (n815,n816);
nand (n816,n817,n818);
or (n817,n183,n108);
or (n818,n260,n184);
nand (n819,n820,n187);
not (n820,n750);
nand (n821,n822,n827);
or (n822,n823,n142);
not (n823,n824);
nand (n824,n825,n826);
or (n825,n35,n98);
or (n826,n34,n96);
nand (n827,n136,n772);
nand (n828,n829,n833);
or (n829,n29,n830);
nor (n830,n831,n832);
and (n831,n26,n174);
and (n832,n27,n173);
or (n833,n413,n779);
and (n834,n813,n821);
xor (n835,n740,n748);
xor (n836,n768,n783);
and (n837,n810,n835);
nand (n838,n839,n997);
or (n839,n840,n890);
not (n840,n841);
nand (n841,n842,n866);
not (n842,n843);
xor (n843,n844,n865);
xor (n844,n845,n846);
xor (n845,n784,n790);
or (n846,n847,n864);
and (n847,n848,n857);
xor (n848,n849,n850);
and (n849,n187,n108);
nand (n850,n851,n856);
or (n851,n111,n852);
not (n852,n853);
nor (n853,n854,n855);
and (n854,n68,n117);
and (n855,n69,n114);
nand (n856,n793,n113);
nand (n857,n858,n863);
or (n858,n859,n142);
not (n859,n860);
nor (n860,n861,n862);
and (n861,n92,n34);
and (n862,n90,n35);
nand (n863,n136,n824);
and (n864,n849,n850);
xor (n865,n812,n828);
not (n866,n867);
or (n867,n868,n889);
and (n868,n869,n888);
xor (n869,n870,n876);
nand (n870,n871,n875);
or (n871,n29,n872);
nor (n872,n873,n874);
and (n873,n158,n27);
and (n874,n159,n26);
or (n875,n413,n830);
and (n876,n877,n882);
and (n877,n878,n27);
nand (n878,n879,n881);
or (n879,n880,n35);
and (n880,n108,n33);
or (n881,n108,n33);
nand (n882,n883,n884);
or (n883,n112,n852);
or (n884,n885,n111);
nor (n885,n886,n887);
and (n886,n117,n96);
and (n887,n114,n98);
xor (n888,n848,n857);
and (n889,n870,n876);
not (n890,n891);
nand (n891,n892,n996);
or (n892,n893,n916);
not (n893,n894);
nand (n894,n895,n897);
not (n895,n896);
xor (n896,n869,n888);
not (n897,n898);
or (n898,n899,n915);
and (n899,n900,n914);
xor (n900,n901,n908);
nand (n901,n902,n907);
or (n902,n903,n142);
not (n903,n904);
nor (n904,n905,n906);
and (n905,n173,n34);
and (n906,n174,n35);
nand (n907,n860,n136);
nand (n908,n909,n910);
or (n909,n413,n872);
nand (n910,n30,n911);
nand (n911,n912,n913);
or (n912,n108,n26);
or (n913,n260,n27);
xor (n914,n877,n882);
and (n915,n901,n908);
not (n916,n917);
or (n917,n918,n995);
and (n918,n919,n940);
xor (n919,n920,n939);
or (n920,n921,n938);
and (n921,n922,n931);
xor (n922,n923,n924);
and (n923,n31,n108);
nand (n924,n925,n930);
or (n925,n926,n142);
not (n926,n927);
nor (n927,n928,n929);
and (n928,n158,n34);
and (n929,n159,n35);
nand (n930,n904,n136);
nand (n931,n932,n937);
or (n932,n111,n933);
not (n933,n934);
nor (n934,n935,n936);
and (n935,n92,n117);
and (n936,n90,n114);
or (n937,n885,n112);
and (n938,n923,n924);
xor (n939,n900,n914);
nand (n940,n941,n994);
or (n941,n942,n958);
nor (n942,n943,n944);
xor (n943,n922,n931);
nor (n944,n945,n953);
not (n945,n946);
nand (n946,n947,n948);
or (n947,n112,n933);
nand (n948,n949,n952);
nand (n949,n950,n951);
or (n950,n174,n117);
nand (n951,n117,n174);
not (n952,n111);
nand (n953,n954,n35);
nand (n954,n955,n957);
or (n955,n956,n114);
and (n956,n108,n139);
or (n957,n108,n139);
nor (n958,n959,n993);
and (n959,n960,n972);
nand (n960,n961,n968);
not (n961,n962);
nand (n962,n963,n967);
or (n963,n142,n964);
nor (n964,n965,n966);
and (n965,n35,n260);
and (n966,n108,n34);
or (n967,n135,n926);
nor (n968,n969,n970);
and (n969,n953,n946);
and (n970,n971,n945);
not (n971,n953);
or (n972,n973,n992);
and (n973,n974,n983);
xor (n974,n975,n976);
nor (n975,n135,n260);
nand (n976,n977,n982);
or (n977,n111,n978);
not (n978,n979);
nand (n979,n980,n981);
or (n980,n158,n114);
nand (n981,n114,n158);
nand (n982,n949,n113);
nor (n983,n984,n990);
nor (n984,n985,n986);
and (n985,n979,n113);
nor (n986,n987,n111);
nor (n987,n988,n989);
and (n988,n260,n114);
and (n989,n108,n117);
or (n990,n991,n117);
and (n991,n108,n113);
and (n992,n975,n976);
nor (n993,n961,n968);
nand (n994,n943,n944);
and (n995,n920,n939);
nand (n996,n896,n898);
nand (n997,n843,n867);
or (n998,n999,n1002);
or (n999,n1000,n1001);
and (n1000,n844,n865);
and (n1001,n845,n846);
xor (n1002,n809,n836);
nand (n1003,n803,n1004);
and (n1004,n1002,n999);
nand (n1005,n807,n805);
and (n1006,n762,n800);
nand (n1007,n723,n724);
nor (n1008,n708,n1009);
nand (n1009,n1010,n1011);
not (n1010,n574);
or (n1011,n658,n706);
or (n1012,n502,n10);
not (n1013,n1014);
nand (n1014,n1015,n4);
not (n1015,n5);
wire s0n1016,s1n1016,notn1016;
or (n1016,s0n1016,s1n1016);
not(notn1016,n5);
and (s0n1016,notn1016,n1017);
and (s1n1016,n5,1'b0);
wire s0n1017,s1n1017,notn1017;
or (n1017,s0n1017,s1n1017);
not(notn1017,n4);
and (s0n1017,notn1017,n2);
and (s1n1017,n4,n1018);
xor (n1018,n1019,n1718);
xor (n1019,n1020,n1715);
xor (n1020,n1021,n160);
xor (n1021,n1022,n1706);
xor (n1022,n1023,n1705);
xor (n1023,n1024,n1690);
xor (n1024,n1025,n1689);
xor (n1025,n1026,n1668);
xor (n1026,n1027,n1667);
xor (n1027,n1028,n1640);
xor (n1028,n1029,n1639);
xor (n1029,n1030,n1607);
xor (n1030,n1031,n1606);
xor (n1031,n1032,n1568);
xor (n1032,n1033,n221);
xor (n1033,n1034,n1524);
xor (n1034,n1035,n1523);
xor (n1035,n1036,n1475);
xor (n1036,n1037,n1474);
xor (n1037,n1038,n1418);
xor (n1038,n1039,n1417);
xor (n1039,n1040,n1354);
xor (n1040,n1041,n28);
xor (n1041,n1042,n1286);
xor (n1042,n1043,n1285);
xor (n1043,n1044,n1214);
xor (n1044,n1045,n1213);
xor (n1045,n1046,n1133);
xor (n1046,n1047,n1132);
xor (n1047,n1048,n1051);
xor (n1048,n1049,n1050);
and (n1049,n125,n113);
and (n1050,n118,n114);
or (n1051,n1052,n1054);
and (n1052,n1053,n288);
and (n1053,n118,n113);
and (n1054,n1055,n1056);
xor (n1055,n1053,n288);
or (n1056,n1057,n1060);
and (n1057,n1058,n1059);
and (n1058,n133,n113);
and (n1059,n148,n114);
and (n1060,n1061,n1062);
xor (n1061,n1058,n1059);
or (n1062,n1063,n1065);
and (n1063,n1064,n266);
and (n1064,n148,n113);
and (n1065,n1066,n1067);
xor (n1066,n1064,n266);
or (n1067,n1068,n1070);
and (n1068,n1069,n487);
and (n1069,n45,n113);
and (n1070,n1071,n1072);
xor (n1071,n1069,n487);
or (n1072,n1073,n1076);
and (n1073,n1074,n1075);
and (n1074,n25,n113);
and (n1075,n182,n114);
and (n1076,n1077,n1078);
xor (n1077,n1074,n1075);
or (n1078,n1079,n1082);
and (n1079,n1080,n1081);
and (n1080,n182,n113);
and (n1081,n195,n114);
and (n1082,n1083,n1084);
xor (n1083,n1080,n1081);
or (n1084,n1085,n1088);
and (n1085,n1086,n1087);
and (n1086,n195,n113);
and (n1087,n227,n114);
and (n1088,n1089,n1090);
xor (n1089,n1086,n1087);
or (n1090,n1091,n1094);
and (n1091,n1092,n1093);
and (n1092,n227,n113);
and (n1093,n220,n114);
and (n1094,n1095,n1096);
xor (n1095,n1092,n1093);
or (n1096,n1097,n1099);
and (n1097,n1098,n795);
and (n1098,n220,n113);
and (n1099,n1100,n1101);
xor (n1100,n1098,n795);
or (n1101,n1102,n1104);
and (n1102,n1103,n855);
and (n1103,n60,n113);
and (n1104,n1105,n1106);
xor (n1105,n1103,n855);
or (n1106,n1107,n1110);
and (n1107,n1108,n1109);
and (n1108,n69,n113);
and (n1109,n96,n114);
and (n1110,n1111,n1112);
xor (n1111,n1108,n1109);
or (n1112,n1113,n1115);
and (n1113,n1114,n936);
and (n1114,n96,n113);
and (n1115,n1116,n1117);
xor (n1116,n1114,n936);
or (n1117,n1118,n1121);
and (n1118,n1119,n1120);
and (n1119,n90,n113);
and (n1120,n174,n114);
and (n1121,n1122,n1123);
xor (n1122,n1119,n1120);
or (n1123,n1124,n1127);
and (n1124,n1125,n1126);
and (n1125,n174,n113);
and (n1126,n159,n114);
and (n1127,n1128,n1129);
xor (n1128,n1125,n1126);
and (n1129,n1130,n1131);
and (n1130,n159,n113);
and (n1131,n108,n114);
and (n1132,n133,n139);
or (n1133,n1134,n1137);
and (n1134,n1135,n1136);
xor (n1135,n1055,n1056);
and (n1136,n148,n139);
and (n1137,n1138,n1139);
xor (n1138,n1135,n1136);
or (n1139,n1140,n1143);
and (n1140,n1141,n1142);
xor (n1141,n1061,n1062);
and (n1142,n45,n139);
and (n1143,n1144,n1145);
xor (n1144,n1141,n1142);
or (n1145,n1146,n1149);
and (n1146,n1147,n1148);
xor (n1147,n1066,n1067);
and (n1148,n25,n139);
and (n1149,n1150,n1151);
xor (n1150,n1147,n1148);
or (n1151,n1152,n1155);
and (n1152,n1153,n1154);
xor (n1153,n1071,n1072);
and (n1154,n182,n139);
and (n1155,n1156,n1157);
xor (n1156,n1153,n1154);
or (n1157,n1158,n1161);
and (n1158,n1159,n1160);
xor (n1159,n1077,n1078);
and (n1160,n195,n139);
and (n1161,n1162,n1163);
xor (n1162,n1159,n1160);
or (n1163,n1164,n1167);
and (n1164,n1165,n1166);
xor (n1165,n1083,n1084);
and (n1166,n227,n139);
and (n1167,n1168,n1169);
xor (n1168,n1165,n1166);
or (n1169,n1170,n1173);
and (n1170,n1171,n1172);
xor (n1171,n1089,n1090);
and (n1172,n220,n139);
and (n1173,n1174,n1175);
xor (n1174,n1171,n1172);
or (n1175,n1176,n1179);
and (n1176,n1177,n1178);
xor (n1177,n1095,n1096);
and (n1178,n60,n139);
and (n1179,n1180,n1181);
xor (n1180,n1177,n1178);
or (n1181,n1182,n1185);
and (n1182,n1183,n1184);
xor (n1183,n1100,n1101);
and (n1184,n69,n139);
and (n1185,n1186,n1187);
xor (n1186,n1183,n1184);
or (n1187,n1188,n1191);
and (n1188,n1189,n1190);
xor (n1189,n1105,n1106);
and (n1190,n96,n139);
and (n1191,n1192,n1193);
xor (n1192,n1189,n1190);
or (n1193,n1194,n1197);
and (n1194,n1195,n1196);
xor (n1195,n1111,n1112);
and (n1196,n90,n139);
and (n1197,n1198,n1199);
xor (n1198,n1195,n1196);
or (n1199,n1200,n1203);
and (n1200,n1201,n1202);
xor (n1201,n1116,n1117);
and (n1202,n174,n139);
and (n1203,n1204,n1205);
xor (n1204,n1201,n1202);
or (n1205,n1206,n1209);
and (n1206,n1207,n1208);
xor (n1207,n1122,n1123);
and (n1208,n159,n139);
and (n1209,n1210,n1211);
xor (n1210,n1207,n1208);
and (n1211,n1212,n956);
xor (n1212,n1128,n1129);
and (n1213,n148,n35);
or (n1214,n1215,n1217);
and (n1215,n1216,n306);
xor (n1216,n1138,n1139);
and (n1217,n1218,n1219);
xor (n1218,n1216,n306);
or (n1219,n1220,n1223);
and (n1220,n1221,n1222);
xor (n1221,n1144,n1145);
and (n1222,n25,n35);
and (n1223,n1224,n1225);
xor (n1224,n1221,n1222);
or (n1225,n1226,n1229);
and (n1226,n1227,n1228);
xor (n1227,n1150,n1151);
and (n1228,n182,n35);
and (n1229,n1230,n1231);
xor (n1230,n1227,n1228);
or (n1231,n1232,n1235);
and (n1232,n1233,n1234);
xor (n1233,n1156,n1157);
and (n1234,n195,n35);
and (n1235,n1236,n1237);
xor (n1236,n1233,n1234);
or (n1237,n1238,n1241);
and (n1238,n1239,n1240);
xor (n1239,n1162,n1163);
and (n1240,n227,n35);
and (n1241,n1242,n1243);
xor (n1242,n1239,n1240);
or (n1243,n1244,n1247);
and (n1244,n1245,n1246);
xor (n1245,n1168,n1169);
and (n1246,n220,n35);
and (n1247,n1248,n1249);
xor (n1248,n1245,n1246);
or (n1249,n1250,n1253);
and (n1250,n1251,n1252);
xor (n1251,n1174,n1175);
and (n1252,n60,n35);
and (n1253,n1254,n1255);
xor (n1254,n1251,n1252);
or (n1255,n1256,n1259);
and (n1256,n1257,n1258);
xor (n1257,n1180,n1181);
and (n1258,n69,n35);
and (n1259,n1260,n1261);
xor (n1260,n1257,n1258);
or (n1261,n1262,n1265);
and (n1262,n1263,n1264);
xor (n1263,n1186,n1187);
and (n1264,n96,n35);
and (n1265,n1266,n1267);
xor (n1266,n1263,n1264);
or (n1267,n1268,n1270);
and (n1268,n1269,n862);
xor (n1269,n1192,n1193);
and (n1270,n1271,n1272);
xor (n1271,n1269,n862);
or (n1272,n1273,n1275);
and (n1273,n1274,n906);
xor (n1274,n1198,n1199);
and (n1275,n1276,n1277);
xor (n1276,n1274,n906);
or (n1277,n1278,n1280);
and (n1278,n1279,n929);
xor (n1279,n1204,n1205);
and (n1280,n1281,n1282);
xor (n1281,n1279,n929);
and (n1282,n1283,n1284);
xor (n1283,n1210,n1211);
and (n1284,n108,n35);
and (n1285,n45,n33);
or (n1286,n1287,n1290);
and (n1287,n1288,n1289);
xor (n1288,n1218,n1219);
and (n1289,n25,n33);
and (n1290,n1291,n1292);
xor (n1291,n1288,n1289);
or (n1292,n1293,n1296);
and (n1293,n1294,n1295);
xor (n1294,n1224,n1225);
and (n1295,n182,n33);
and (n1296,n1297,n1298);
xor (n1297,n1294,n1295);
or (n1298,n1299,n1302);
and (n1299,n1300,n1301);
xor (n1300,n1230,n1231);
and (n1301,n195,n33);
and (n1302,n1303,n1304);
xor (n1303,n1300,n1301);
or (n1304,n1305,n1308);
and (n1305,n1306,n1307);
xor (n1306,n1236,n1237);
and (n1307,n227,n33);
and (n1308,n1309,n1310);
xor (n1309,n1306,n1307);
or (n1310,n1311,n1314);
and (n1311,n1312,n1313);
xor (n1312,n1242,n1243);
and (n1313,n220,n33);
and (n1314,n1315,n1316);
xor (n1315,n1312,n1313);
or (n1316,n1317,n1320);
and (n1317,n1318,n1319);
xor (n1318,n1248,n1249);
and (n1319,n60,n33);
and (n1320,n1321,n1322);
xor (n1321,n1318,n1319);
or (n1322,n1323,n1326);
and (n1323,n1324,n1325);
xor (n1324,n1254,n1255);
and (n1325,n69,n33);
and (n1326,n1327,n1328);
xor (n1327,n1324,n1325);
or (n1328,n1329,n1332);
and (n1329,n1330,n1331);
xor (n1330,n1260,n1261);
and (n1331,n96,n33);
and (n1332,n1333,n1334);
xor (n1333,n1330,n1331);
or (n1334,n1335,n1338);
and (n1335,n1336,n1337);
xor (n1336,n1266,n1267);
and (n1337,n90,n33);
and (n1338,n1339,n1340);
xor (n1339,n1336,n1337);
or (n1340,n1341,n1344);
and (n1341,n1342,n1343);
xor (n1342,n1271,n1272);
and (n1343,n174,n33);
and (n1344,n1345,n1346);
xor (n1345,n1342,n1343);
or (n1346,n1347,n1350);
and (n1347,n1348,n1349);
xor (n1348,n1276,n1277);
and (n1349,n159,n33);
and (n1350,n1351,n1352);
xor (n1351,n1348,n1349);
and (n1352,n1353,n880);
xor (n1353,n1281,n1282);
or (n1354,n1355,n1358);
and (n1355,n1356,n1357);
xor (n1356,n1291,n1292);
and (n1357,n182,n27);
and (n1358,n1359,n1360);
xor (n1359,n1356,n1357);
or (n1360,n1361,n1364);
and (n1361,n1362,n1363);
xor (n1362,n1297,n1298);
and (n1363,n195,n27);
and (n1364,n1365,n1366);
xor (n1365,n1362,n1363);
or (n1366,n1367,n1370);
and (n1367,n1368,n1369);
xor (n1368,n1303,n1304);
and (n1369,n227,n27);
and (n1370,n1371,n1372);
xor (n1371,n1368,n1369);
or (n1372,n1373,n1376);
and (n1373,n1374,n1375);
xor (n1374,n1309,n1310);
and (n1375,n220,n27);
and (n1376,n1377,n1378);
xor (n1377,n1374,n1375);
or (n1378,n1379,n1382);
and (n1379,n1380,n1381);
xor (n1380,n1315,n1316);
and (n1381,n60,n27);
and (n1382,n1383,n1384);
xor (n1383,n1380,n1381);
or (n1384,n1385,n1388);
and (n1385,n1386,n1387);
xor (n1386,n1321,n1322);
and (n1387,n69,n27);
and (n1388,n1389,n1390);
xor (n1389,n1386,n1387);
or (n1390,n1391,n1394);
and (n1391,n1392,n1393);
xor (n1392,n1327,n1328);
and (n1393,n96,n27);
and (n1394,n1395,n1396);
xor (n1395,n1392,n1393);
or (n1396,n1397,n1400);
and (n1397,n1398,n1399);
xor (n1398,n1333,n1334);
and (n1399,n90,n27);
and (n1400,n1401,n1402);
xor (n1401,n1398,n1399);
or (n1402,n1403,n1406);
and (n1403,n1404,n1405);
xor (n1404,n1339,n1340);
and (n1405,n174,n27);
and (n1406,n1407,n1408);
xor (n1407,n1404,n1405);
or (n1408,n1409,n1412);
and (n1409,n1410,n1411);
xor (n1410,n1345,n1346);
and (n1411,n159,n27);
and (n1412,n1413,n1414);
xor (n1413,n1410,n1411);
and (n1414,n1415,n1416);
xor (n1415,n1351,n1352);
and (n1416,n108,n27);
and (n1417,n182,n189);
or (n1418,n1419,n1422);
and (n1419,n1420,n1421);
xor (n1420,n1359,n1360);
and (n1421,n195,n189);
and (n1422,n1423,n1424);
xor (n1423,n1420,n1421);
or (n1424,n1425,n1428);
and (n1425,n1426,n1427);
xor (n1426,n1365,n1366);
and (n1427,n227,n189);
and (n1428,n1429,n1430);
xor (n1429,n1426,n1427);
or (n1430,n1431,n1434);
and (n1431,n1432,n1433);
xor (n1432,n1371,n1372);
and (n1433,n220,n189);
and (n1434,n1435,n1436);
xor (n1435,n1432,n1433);
or (n1436,n1437,n1440);
and (n1437,n1438,n1439);
xor (n1438,n1377,n1378);
and (n1439,n60,n189);
and (n1440,n1441,n1442);
xor (n1441,n1438,n1439);
or (n1442,n1443,n1446);
and (n1443,n1444,n1445);
xor (n1444,n1383,n1384);
and (n1445,n69,n189);
and (n1446,n1447,n1448);
xor (n1447,n1444,n1445);
or (n1448,n1449,n1452);
and (n1449,n1450,n1451);
xor (n1450,n1389,n1390);
and (n1451,n96,n189);
and (n1452,n1453,n1454);
xor (n1453,n1450,n1451);
or (n1454,n1455,n1458);
and (n1455,n1456,n1457);
xor (n1456,n1395,n1396);
and (n1457,n90,n189);
and (n1458,n1459,n1460);
xor (n1459,n1456,n1457);
or (n1460,n1461,n1464);
and (n1461,n1462,n1463);
xor (n1462,n1401,n1402);
and (n1463,n174,n189);
and (n1464,n1465,n1466);
xor (n1465,n1462,n1463);
or (n1466,n1467,n1470);
and (n1467,n1468,n1469);
xor (n1468,n1407,n1408);
and (n1469,n159,n189);
and (n1470,n1471,n1472);
xor (n1471,n1468,n1469);
and (n1472,n1473,n789);
xor (n1473,n1413,n1414);
and (n1474,n195,n184);
or (n1475,n1476,n1478);
and (n1476,n1477,n397);
xor (n1477,n1423,n1424);
and (n1478,n1479,n1480);
xor (n1479,n1477,n397);
or (n1480,n1481,n1483);
and (n1481,n1482,n326);
xor (n1482,n1429,n1430);
and (n1483,n1484,n1485);
xor (n1484,n1482,n326);
or (n1485,n1486,n1489);
and (n1486,n1487,n1488);
xor (n1487,n1435,n1436);
and (n1488,n60,n184);
and (n1489,n1490,n1491);
xor (n1490,n1487,n1488);
or (n1491,n1492,n1494);
and (n1492,n1493,n468);
xor (n1493,n1441,n1442);
and (n1494,n1495,n1496);
xor (n1495,n1493,n468);
or (n1496,n1497,n1500);
and (n1497,n1498,n1499);
xor (n1498,n1447,n1448);
and (n1499,n96,n184);
and (n1500,n1501,n1502);
xor (n1501,n1498,n1499);
or (n1502,n1503,n1506);
and (n1503,n1504,n1505);
xor (n1504,n1453,n1454);
and (n1505,n90,n184);
and (n1506,n1507,n1508);
xor (n1507,n1504,n1505);
or (n1508,n1509,n1512);
and (n1509,n1510,n1511);
xor (n1510,n1459,n1460);
and (n1511,n174,n184);
and (n1512,n1513,n1514);
xor (n1513,n1510,n1511);
or (n1514,n1515,n1518);
and (n1515,n1516,n1517);
xor (n1516,n1465,n1466);
and (n1517,n159,n184);
and (n1518,n1519,n1520);
xor (n1519,n1516,n1517);
and (n1520,n1521,n1522);
xor (n1521,n1471,n1472);
and (n1522,n108,n184);
and (n1523,n227,n209);
or (n1524,n1525,n1528);
and (n1525,n1526,n1527);
xor (n1526,n1479,n1480);
and (n1527,n220,n209);
and (n1528,n1529,n1530);
xor (n1529,n1526,n1527);
or (n1530,n1531,n1534);
and (n1531,n1532,n1533);
xor (n1532,n1484,n1485);
and (n1533,n60,n209);
and (n1534,n1535,n1536);
xor (n1535,n1532,n1533);
or (n1536,n1537,n1540);
and (n1537,n1538,n1539);
xor (n1538,n1490,n1491);
and (n1539,n69,n209);
and (n1540,n1541,n1542);
xor (n1541,n1538,n1539);
or (n1542,n1543,n1546);
and (n1543,n1544,n1545);
xor (n1544,n1495,n1496);
and (n1545,n96,n209);
and (n1546,n1547,n1548);
xor (n1547,n1544,n1545);
or (n1548,n1549,n1552);
and (n1549,n1550,n1551);
xor (n1550,n1501,n1502);
and (n1551,n90,n209);
and (n1552,n1553,n1554);
xor (n1553,n1550,n1551);
or (n1554,n1555,n1558);
and (n1555,n1556,n1557);
xor (n1556,n1507,n1508);
and (n1557,n174,n209);
and (n1558,n1559,n1560);
xor (n1559,n1556,n1557);
or (n1560,n1561,n1564);
and (n1561,n1562,n1563);
xor (n1562,n1513,n1514);
and (n1563,n159,n209);
and (n1564,n1565,n1566);
xor (n1565,n1562,n1563);
and (n1566,n1567,n672);
xor (n1567,n1519,n1520);
or (n1568,n1569,n1571);
and (n1569,n1570,n409);
xor (n1570,n1529,n1530);
and (n1571,n1572,n1573);
xor (n1572,n1570,n409);
or (n1573,n1574,n1577);
and (n1574,n1575,n1576);
xor (n1575,n1535,n1536);
and (n1576,n69,n54);
and (n1577,n1578,n1579);
xor (n1578,n1575,n1576);
or (n1579,n1580,n1583);
and (n1580,n1581,n1582);
xor (n1581,n1541,n1542);
and (n1582,n96,n54);
and (n1583,n1584,n1585);
xor (n1584,n1581,n1582);
or (n1585,n1586,n1589);
and (n1586,n1587,n1588);
xor (n1587,n1547,n1548);
and (n1588,n90,n54);
and (n1589,n1590,n1591);
xor (n1590,n1587,n1588);
or (n1591,n1592,n1595);
and (n1592,n1593,n1594);
xor (n1593,n1553,n1554);
and (n1594,n174,n54);
and (n1595,n1596,n1597);
xor (n1596,n1593,n1594);
or (n1597,n1598,n1601);
and (n1598,n1599,n1600);
xor (n1599,n1559,n1560);
and (n1600,n159,n54);
and (n1601,n1602,n1603);
xor (n1602,n1599,n1600);
and (n1603,n1604,n1605);
xor (n1604,n1565,n1566);
and (n1605,n108,n54);
and (n1606,n60,n53);
or (n1607,n1608,n1611);
and (n1608,n1609,n1610);
xor (n1609,n1572,n1573);
and (n1610,n69,n53);
and (n1611,n1612,n1613);
xor (n1612,n1609,n1610);
or (n1613,n1614,n1617);
and (n1614,n1615,n1616);
xor (n1615,n1578,n1579);
and (n1616,n96,n53);
and (n1617,n1618,n1619);
xor (n1618,n1615,n1616);
or (n1619,n1620,n1623);
and (n1620,n1621,n1622);
xor (n1621,n1584,n1585);
and (n1622,n90,n53);
and (n1623,n1624,n1625);
xor (n1624,n1621,n1622);
or (n1625,n1626,n1629);
and (n1626,n1627,n1628);
xor (n1627,n1590,n1591);
and (n1628,n174,n53);
and (n1629,n1630,n1631);
xor (n1630,n1627,n1628);
or (n1631,n1632,n1635);
and (n1632,n1633,n1634);
xor (n1633,n1596,n1597);
and (n1634,n159,n53);
and (n1635,n1636,n1637);
xor (n1636,n1633,n1634);
and (n1637,n1638,n541);
xor (n1638,n1602,n1603);
and (n1639,n69,n61);
or (n1640,n1641,n1644);
and (n1641,n1642,n1643);
xor (n1642,n1612,n1613);
and (n1643,n96,n61);
and (n1644,n1645,n1646);
xor (n1645,n1642,n1643);
or (n1646,n1647,n1650);
and (n1647,n1648,n1649);
xor (n1648,n1618,n1619);
and (n1649,n90,n61);
and (n1650,n1651,n1652);
xor (n1651,n1648,n1649);
or (n1652,n1653,n1656);
and (n1653,n1654,n1655);
xor (n1654,n1624,n1625);
and (n1655,n174,n61);
and (n1656,n1657,n1658);
xor (n1657,n1654,n1655);
or (n1658,n1659,n1662);
and (n1659,n1660,n1661);
xor (n1660,n1630,n1631);
and (n1661,n159,n61);
and (n1662,n1663,n1664);
xor (n1663,n1660,n1661);
and (n1664,n1665,n1666);
xor (n1665,n1636,n1637);
and (n1666,n108,n61);
and (n1667,n96,n81);
or (n1668,n1669,n1672);
and (n1669,n1670,n1671);
xor (n1670,n1645,n1646);
and (n1671,n90,n81);
and (n1672,n1673,n1674);
xor (n1673,n1670,n1671);
or (n1674,n1675,n1678);
and (n1675,n1676,n1677);
xor (n1676,n1651,n1652);
and (n1677,n174,n81);
and (n1678,n1679,n1680);
xor (n1679,n1676,n1677);
or (n1680,n1681,n1684);
and (n1681,n1682,n1683);
xor (n1682,n1657,n1658);
and (n1683,n159,n81);
and (n1684,n1685,n1686);
xor (n1685,n1682,n1683);
and (n1686,n1687,n1688);
xor (n1687,n1663,n1664);
not (n1688,n258);
and (n1689,n90,n86);
or (n1690,n1691,n1694);
and (n1691,n1692,n1693);
xor (n1692,n1673,n1674);
and (n1693,n174,n86);
and (n1694,n1695,n1696);
xor (n1695,n1692,n1693);
or (n1696,n1697,n1700);
and (n1697,n1698,n1699);
xor (n1698,n1679,n1680);
and (n1699,n159,n86);
and (n1700,n1701,n1702);
xor (n1701,n1698,n1699);
and (n1702,n1703,n1704);
xor (n1703,n1685,n1686);
and (n1704,n108,n86);
and (n1705,n174,n165);
or (n1706,n1707,n1710);
and (n1707,n1708,n1709);
xor (n1708,n1695,n1696);
and (n1709,n159,n165);
and (n1710,n1711,n1712);
xor (n1711,n1708,n1709);
and (n1712,n1713,n1714);
xor (n1713,n1701,n1702);
not (n1714,n281);
and (n1715,n1716,n1717);
xor (n1716,n1711,n1712);
and (n1717,n108,n105);
and (n1718,n108,n106);
endmodule
