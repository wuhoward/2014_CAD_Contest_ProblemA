module top (out,n20,n25,n26,n27,n29,n30,n41,n44,n47
        ,n50,n53,n56,n59,n62,n65,n68,n71,n74,n77
        ,n80,n83,n86,n89,n92,n95,n98,n101,n104,n107
        ,n110,n113,n116,n118,n121,n124,n132,n158,n163,n166
        ,n169,n172,n175,n178,n181,n184,n187,n190,n193,n196
        ,n199,n202,n205,n208,n211,n214,n217,n220,n223,n226
        ,n229,n232,n235,n243,n400,n414);
output out;
input n20;
input n25;
input n26;
input n27;
input n29;
input n30;
input n41;
input n44;
input n47;
input n50;
input n53;
input n56;
input n59;
input n62;
input n65;
input n68;
input n71;
input n74;
input n77;
input n80;
input n83;
input n86;
input n89;
input n92;
input n95;
input n98;
input n101;
input n104;
input n107;
input n110;
input n113;
input n116;
input n118;
input n121;
input n124;
input n132;
input n158;
input n163;
input n166;
input n169;
input n172;
input n175;
input n178;
input n181;
input n184;
input n187;
input n190;
input n193;
input n196;
input n199;
input n202;
input n205;
input n208;
input n211;
input n214;
input n217;
input n220;
input n223;
input n226;
input n229;
input n232;
input n235;
input n243;
input n400;
input n414;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n21;
wire n22;
wire n23;
wire n24;
wire n28;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n42;
wire n43;
wire n45;
wire n46;
wire n48;
wire n49;
wire n51;
wire n52;
wire n54;
wire n55;
wire n57;
wire n58;
wire n60;
wire n61;
wire n63;
wire n64;
wire n66;
wire n67;
wire n69;
wire n70;
wire n72;
wire n73;
wire n75;
wire n76;
wire n78;
wire n79;
wire n81;
wire n82;
wire n84;
wire n85;
wire n87;
wire n88;
wire n90;
wire n91;
wire n93;
wire n94;
wire n96;
wire n97;
wire n99;
wire n100;
wire n102;
wire n103;
wire n105;
wire n106;
wire n108;
wire n109;
wire n111;
wire n112;
wire n114;
wire n115;
wire n117;
wire n119;
wire n120;
wire n122;
wire n123;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n159;
wire n160;
wire n161;
wire n162;
wire n164;
wire n165;
wire n167;
wire n168;
wire n170;
wire n171;
wire n173;
wire n174;
wire n176;
wire n177;
wire n179;
wire n180;
wire n182;
wire n183;
wire n185;
wire n186;
wire n188;
wire n189;
wire n191;
wire n192;
wire n194;
wire n195;
wire n197;
wire n198;
wire n200;
wire n201;
wire n203;
wire n204;
wire n206;
wire n207;
wire n209;
wire n210;
wire n212;
wire n213;
wire n215;
wire n216;
wire n218;
wire n219;
wire n221;
wire n222;
wire n224;
wire n225;
wire n227;
wire n228;
wire n230;
wire n231;
wire n233;
wire n234;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2988;
wire n2989;
wire n2990;
wire n2991;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2996;
wire n2997;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3003;
wire n3004;
wire n3005;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3010;
wire n3011;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3038;
wire n3039;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
wire n3056;
wire n3057;
wire n3058;
wire n3059;
wire n3060;
wire n3061;
wire n3062;
wire n3063;
wire n3064;
wire n3065;
wire n3066;
wire n3067;
wire n3068;
wire n3069;
wire n3070;
wire n3071;
wire n3072;
wire n3073;
wire n3074;
wire n3075;
wire n3076;
wire n3077;
wire n3078;
wire n3079;
wire n3080;
wire n3081;
wire n3082;
wire n3083;
wire n3084;
wire n3085;
wire n3086;
wire n3087;
wire n3088;
wire n3089;
wire n3090;
wire n3091;
wire n3092;
wire n3093;
wire n3094;
wire n3095;
wire n3096;
wire n3097;
wire n3098;
wire n3099;
wire n3100;
wire n3101;
wire n3102;
wire n3103;
wire n3104;
wire n3105;
wire n3106;
wire n3107;
wire n3108;
wire n3109;
wire n3110;
wire n3111;
wire n3112;
wire n3113;
wire n3114;
wire n3115;
wire n3116;
wire n3117;
wire n3118;
wire n3119;
wire n3120;
wire n3121;
wire n3122;
wire n3123;
wire n3124;
wire n3125;
wire n3126;
wire n3127;
wire n3128;
wire n3129;
wire n3130;
wire n3131;
wire n3132;
wire n3133;
wire n3134;
wire n3135;
wire n3136;
wire n3137;
wire n3138;
wire n3139;
wire n3140;
wire n3141;
wire n3142;
wire n3143;
wire n3144;
wire n3145;
wire n3146;
wire n3147;
wire n3148;
wire n3149;
wire n3150;
wire n3151;
wire n3152;
wire n3153;
wire n3154;
wire n3155;
wire n3156;
wire n3157;
wire n3158;
wire n3159;
wire n3160;
wire n3161;
wire n3162;
wire n3163;
wire n3164;
wire n3165;
wire n3166;
wire n3167;
wire n3168;
wire n3169;
wire n3170;
wire n3171;
wire n3172;
wire n3173;
wire n3174;
wire n3175;
wire n3176;
wire n3177;
wire n3178;
wire n3179;
wire n3180;
wire n3181;
wire n3182;
wire n3183;
wire n3184;
wire n3185;
wire n3186;
wire n3187;
wire n3188;
wire n3189;
wire n3190;
wire n3191;
wire n3192;
wire n3193;
wire n3194;
wire n3195;
wire n3196;
wire n3197;
wire n3198;
wire n3199;
wire n3200;
wire n3201;
wire n3202;
wire n3203;
wire n3204;
wire n3205;
wire n3206;
wire n3207;
wire n3208;
wire n3209;
wire n3210;
wire n3211;
wire n3212;
wire n3213;
wire n3214;
wire n3215;
wire n3216;
wire n3217;
wire n3218;
wire n3219;
wire n3220;
wire n3221;
wire n3222;
wire n3223;
wire n3224;
wire n3225;
wire n3226;
wire n3227;
wire n3228;
wire n3229;
wire n3230;
wire n3231;
wire n3232;
wire n3233;
wire n3234;
wire n3235;
wire n3236;
wire n3237;
wire n3238;
wire n3239;
wire n3240;
wire n3241;
wire n3242;
wire n3243;
wire n3244;
wire n3245;
wire n3246;
wire n3247;
wire n3248;
wire n3249;
wire n3250;
wire n3251;
wire n3252;
wire n3253;
wire n3254;
wire n3255;
wire n3256;
wire n3257;
wire n3258;
wire n3259;
wire n3260;
wire n3261;
wire n3262;
wire n3263;
wire n3264;
wire n3265;
wire n3266;
wire n3267;
wire n3268;
wire n3269;
wire n3270;
wire n3271;
wire n3272;
wire n3273;
wire n3274;
wire n3275;
wire n3276;
wire n3277;
wire n3278;
wire n3279;
wire n3280;
wire n3281;
wire n3282;
wire n3283;
wire n3284;
wire n3285;
wire n3286;
wire n3287;
wire n3288;
wire n3289;
wire n3290;
wire n3291;
wire n3292;
wire n3293;
wire n3294;
wire n3295;
wire n3296;
wire n3297;
wire n3298;
wire n3299;
wire n3300;
wire n3301;
wire n3302;
wire n3303;
wire n3304;
wire n3305;
wire n3306;
wire n3307;
wire n3308;
wire n3309;
wire n3310;
wire n3311;
wire n3312;
wire n3313;
wire n3314;
wire n3315;
wire n3316;
wire n3317;
wire n3318;
wire n3319;
wire n3320;
wire n3321;
wire n3322;
wire n3323;
wire n3324;
wire n3325;
wire n3326;
wire n3327;
wire n3328;
wire n3329;
wire n3330;
wire n3331;
wire n3332;
wire n3333;
wire n3334;
wire n3335;
wire n3336;
wire n3337;
wire n3338;
wire n3339;
wire n3340;
wire n3341;
wire n3342;
wire n3343;
wire n3344;
wire n3345;
wire n3346;
wire n3347;
wire n3348;
wire n3349;
wire n3350;
wire n3351;
wire n3352;
wire n3353;
wire n3354;
wire n3355;
wire n3356;
wire n3357;
wire n3358;
wire n3359;
wire n3360;
wire n3361;
wire n3362;
wire n3363;
wire n3364;
wire n3365;
wire n3366;
wire n3367;
wire n3368;
wire n3369;
wire n3370;
wire n3371;
wire n3372;
wire n3373;
wire n3374;
wire n3375;
wire n3376;
wire n3377;
wire n3378;
wire n3379;
wire n3380;
wire n3381;
wire n3382;
wire n3383;
wire n3384;
wire n3385;
wire n3386;
wire n3387;
wire n3388;
wire n3389;
wire n3390;
wire n3391;
wire n3392;
wire n3393;
wire n3394;
wire n3395;
wire n3396;
wire n3397;
wire n3398;
wire n3399;
wire n3400;
wire n3401;
wire n3402;
wire n3403;
wire n3404;
wire n3405;
wire n3406;
wire n3407;
wire n3408;
wire n3409;
wire n3410;
wire n3411;
wire n3412;
wire n3413;
wire n3414;
wire n3415;
wire n3416;
wire n3417;
wire n3418;
wire n3419;
wire n3420;
wire n3421;
wire n3422;
wire n3423;
wire n3424;
wire n3425;
wire n3426;
wire n3427;
wire n3428;
wire n3429;
wire n3430;
wire n3431;
wire n3432;
wire n3433;
wire n3434;
wire n3435;
wire n3436;
wire n3437;
wire n3438;
wire n3439;
wire n3440;
wire n3441;
wire n3442;
wire n3443;
wire n3444;
wire n3445;
wire n3446;
wire n3447;
wire n3448;
wire n3449;
wire n3450;
wire n3451;
wire n3452;
wire n3453;
wire n3454;
wire n3455;
wire n3456;
wire n3457;
wire n3458;
wire n3459;
wire n3460;
wire n3461;
wire n3462;
wire n3463;
wire n3464;
wire n3465;
wire n3466;
wire n3467;
wire n3468;
wire n3469;
wire n3470;
wire n3471;
wire n3472;
wire n3473;
wire n3474;
wire n3475;
wire n3476;
wire n3477;
wire n3478;
wire n3479;
wire n3480;
wire n3481;
wire n3482;
wire n3483;
wire n3484;
wire n3485;
wire n3486;
wire n3487;
wire n3488;
wire n3489;
wire n3490;
wire n3491;
wire n3492;
wire n3493;
wire n3494;
wire n3495;
wire n3496;
wire n3497;
wire n3498;
wire n3499;
wire n3500;
wire n3501;
wire n3502;
wire n3503;
wire n3504;
wire n3505;
wire n3506;
wire n3507;
wire n3508;
wire n3509;
wire n3510;
wire n3511;
wire n3512;
wire n3513;
wire n3514;
wire n3515;
wire n3516;
wire n3517;
wire n3518;
wire n3519;
wire n3520;
wire n3521;
wire n3522;
wire n3523;
wire n3524;
wire n3525;
wire n3526;
wire n3527;
wire n3528;
wire n3529;
wire n3530;
wire n3531;
wire n3532;
wire n3533;
wire n3534;
wire n3535;
wire n3536;
wire n3537;
wire n3538;
wire n3539;
wire n3540;
wire n3541;
wire n3542;
wire n3543;
wire n3544;
wire n3545;
wire n3546;
wire n3547;
wire n3548;
wire n3549;
wire n3550;
wire n3551;
wire n3552;
wire n3553;
wire n3554;
wire n3555;
wire n3556;
wire n3557;
wire n3558;
wire n3559;
wire n3560;
wire n3561;
wire n3562;
wire n3563;
wire n3564;
wire n3565;
wire n3566;
wire n3567;
wire n3568;
wire n3569;
wire n3570;
wire n3571;
wire n3572;
wire n3573;
wire n3574;
wire n3575;
wire n3576;
wire n3577;
wire n3578;
wire n3579;
wire n3580;
wire n3581;
wire n3582;
wire n3583;
wire n3584;
wire n3585;
wire n3586;
wire n3587;
wire n3588;
wire n3589;
wire n3590;
wire n3591;
wire n3592;
wire n3593;
wire n3594;
wire n3595;
wire n3596;
wire n3597;
wire n3598;
wire n3599;
wire n3600;
wire n3601;
wire n3602;
wire n3603;
wire n3604;
wire n3605;
wire n3606;
wire n3607;
wire n3608;
wire n3609;
wire n3610;
wire n3611;
wire n3612;
wire n3613;
wire n3614;
wire n3615;
wire n3616;
wire n3617;
wire n3618;
wire n3619;
wire n3620;
wire n3621;
wire n3622;
wire n3623;
wire n3624;
wire n3625;
wire n3626;
wire n3627;
wire n3628;
wire n3629;
wire n3630;
wire n3631;
wire n3632;
wire n3633;
wire n3634;
wire n3635;
wire n3636;
wire n3637;
wire n3638;
wire n3639;
wire n3640;
wire n3641;
wire n3642;
wire n3643;
wire n3644;
wire n3645;
wire n3646;
wire n3647;
wire n3648;
wire n3649;
wire n3650;
wire n3651;
wire n3652;
wire n3653;
wire n3654;
wire n3655;
wire n3656;
wire n3657;
wire n3658;
wire n3659;
wire n3660;
wire n3661;
wire n3662;
wire n3663;
wire n3664;
wire n3665;
wire n3666;
wire n3667;
wire n3668;
wire n3669;
wire n3670;
wire n3671;
wire n3672;
wire n3673;
wire n3674;
wire n3675;
wire n3676;
wire n3677;
wire n3678;
wire n3679;
wire n3680;
wire n3681;
wire n3682;
wire n3683;
wire n3684;
wire n3685;
wire n3686;
wire n3687;
wire n3688;
wire n3689;
wire n3690;
wire n3691;
wire n3692;
wire n3693;
wire n3694;
wire n3695;
wire n3696;
wire n3697;
wire n3698;
wire n3699;
wire n3700;
wire n3701;
wire n3702;
wire n3703;
wire n3704;
wire n3705;
wire n3706;
wire n3707;
wire n3708;
wire n3709;
wire n3710;
wire n3711;
wire n3712;
wire n3713;
wire n3714;
wire n3715;
wire n3716;
wire n3717;
wire n3718;
wire n3719;
wire n3720;
wire n3721;
wire n3722;
wire n3723;
wire n3724;
wire n3725;
wire n3726;
wire n3727;
wire n3728;
wire n3729;
wire n3730;
wire n3731;
wire n3732;
wire n3733;
wire n3734;
wire n3735;
wire n3736;
wire n3737;
wire n3738;
wire n3739;
wire n3740;
wire n3741;
wire n3742;
wire n3743;
wire n3744;
wire n3745;
wire n3746;
wire n3747;
wire n3748;
wire n3749;
wire n3750;
wire n3751;
wire n3752;
wire n3753;
wire n3754;
wire n3755;
wire n3756;
wire n3757;
wire n3758;
wire n3759;
wire n3760;
wire n3761;
wire n3762;
wire n3763;
wire n3764;
wire n3765;
wire n3766;
wire n3767;
wire n3768;
wire n3769;
wire n3770;
wire n3771;
wire n3772;
wire n3773;
wire n3774;
wire n3775;
wire n3776;
wire n3777;
wire n3778;
wire n3779;
wire n3780;
wire n3781;
wire n3782;
wire n3783;
wire n3784;
wire n3785;
wire n3786;
wire n3787;
wire n3788;
wire n3789;
wire n3790;
wire n3791;
wire n3792;
wire n3793;
wire n3794;
wire n3795;
wire n3796;
wire n3797;
wire n3798;
wire n3799;
wire n3800;
wire n3801;
wire n3802;
wire n3803;
wire n3804;
wire n3805;
wire n3806;
wire n3807;
wire n3808;
wire n3809;
wire n3810;
wire n3811;
wire n3812;
wire n3813;
wire n3814;
wire n3815;
wire n3816;
wire n3817;
wire n3818;
wire n3819;
wire n3820;
wire n3821;
wire n3822;
wire n3823;
wire n3824;
wire n3825;
wire n3826;
wire n3827;
wire n3828;
wire n3829;
wire n3830;
wire n3831;
wire n3832;
wire n3833;
wire n3834;
wire n3835;
wire n3836;
wire n3837;
wire n3838;
wire n3839;
wire n3840;
wire n3841;
wire n3842;
wire n3843;
wire n3844;
wire n3845;
wire n3846;
wire n3847;
wire n3848;
wire n3849;
wire n3850;
wire n3851;
wire n3852;
wire n3853;
wire n3854;
wire n3855;
wire n3856;
wire n3857;
wire n3858;
wire n3859;
wire n3860;
wire n3861;
wire n3862;
wire n3863;
wire n3864;
wire n3865;
wire n3866;
wire n3867;
wire n3868;
wire n3869;
wire n3870;
wire n3871;
wire n3872;
wire n3873;
wire n3874;
wire n3875;
wire n3876;
wire n3877;
wire n3878;
wire n3879;
wire n3880;
wire n3881;
wire n3882;
wire n3883;
wire n3884;
wire n3885;
wire n3886;
wire n3887;
wire n3888;
wire n3889;
wire n3890;
wire n3891;
wire n3892;
wire n3893;
wire n3894;
wire n3895;
wire n3896;
wire n3897;
wire n3898;
wire n3899;
wire n3900;
wire n3901;
wire n3902;
wire n3903;
wire n3904;
wire n3905;
wire n3906;
wire n3907;
wire n3908;
wire n3909;
wire n3910;
wire n3911;
wire n3912;
wire n3913;
wire n3914;
wire n3915;
wire n3916;
wire n3917;
wire n3918;
wire n3919;
wire n3920;
wire n3921;
wire n3922;
wire n3923;
wire n3924;
wire n3925;
wire n3926;
wire n3927;
wire n3928;
wire n3929;
wire n3930;
wire n3931;
wire n3932;
wire n3933;
wire n3934;
wire n3935;
wire n3936;
wire n3937;
wire n3938;
wire n3939;
wire n3940;
wire n3941;
wire n3942;
wire n3943;
wire n3944;
wire n3945;
wire n3946;
wire n3947;
wire n3948;
wire n3949;
wire n3950;
wire n3951;
wire n3952;
wire n3953;
wire n3954;
wire n3955;
wire n3956;
wire n3957;
wire n3958;
wire n3959;
wire n3960;
wire n3961;
wire n3962;
wire n3963;
wire n3964;
wire n3965;
wire n3966;
wire n3967;
wire n3968;
wire n3969;
wire n3970;
wire n3971;
wire n3972;
wire n3973;
wire n3974;
wire n3975;
wire n3976;
wire n3977;
wire n3978;
wire n3979;
wire n3980;
wire n3981;
wire n3982;
wire n3983;
wire n3984;
wire n3985;
wire n3986;
wire n3987;
wire n3988;
wire n3989;
wire n3990;
wire n3991;
wire n3992;
wire n3993;
wire n3994;
wire n3995;
wire n3996;
wire n3997;
wire n3998;
wire n3999;
wire n4000;
wire n4001;
wire n4002;
wire n4003;
wire n4004;
wire n4005;
wire n4006;
wire n4007;
wire n4008;
wire n4009;
wire n4010;
wire n4011;
wire n4012;
wire n4013;
wire n4014;
wire n4015;
wire n4016;
wire n4017;
wire n4018;
wire n4019;
wire n4020;
wire n4021;
wire n4022;
wire n4023;
wire n4024;
wire n4025;
wire n4026;
wire n4027;
wire n4028;
wire n4029;
wire n4030;
wire n4031;
wire n4032;
wire n4033;
wire n4034;
wire n4035;
wire n4036;
wire n4037;
wire n4038;
wire n4039;
wire n4040;
wire n4041;
wire n4042;
wire n4043;
wire n4044;
wire n4045;
wire n4046;
wire n4047;
wire n4048;
wire n4049;
wire n4050;
wire n4051;
wire n4052;
wire n4053;
wire n4054;
wire n4055;
wire n4056;
wire n4057;
wire n4058;
wire n4059;
wire n4060;
wire n4061;
wire n4062;
wire n4063;
wire n4064;
wire n4065;
wire n4066;
wire n4067;
wire n4068;
wire n4069;
wire n4070;
wire n4071;
wire n4072;
wire n4073;
wire n4074;
wire n4075;
wire n4076;
wire n4077;
wire n4078;
wire n4079;
wire n4080;
wire n4081;
wire n4082;
wire n4083;
wire n4084;
wire n4085;
wire n4086;
wire n4087;
wire n4088;
wire n4089;
wire n4090;
wire n4091;
wire n4092;
wire n4093;
wire n4094;
wire n4095;
wire n4096;
wire n4097;
wire n4098;
wire n4099;
wire n4100;
wire n4101;
wire n4102;
wire n4103;
wire n4104;
wire n4105;
wire n4106;
wire n4107;
wire n4108;
wire n4109;
wire n4110;
wire n4111;
wire n4112;
wire n4113;
wire n4114;
wire n4115;
wire n4116;
wire n4117;
wire n4118;
wire n4119;
wire n4120;
wire n4121;
wire n4122;
wire n4123;
wire n4124;
wire n4125;
wire n4126;
wire n4127;
wire n4128;
wire n4129;
wire n4130;
wire n4131;
wire n4132;
wire n4133;
wire n4134;
wire n4135;
wire n4136;
wire n4137;
wire n4138;
wire n4139;
wire n4140;
wire n4141;
wire n4142;
wire n4143;
wire n4144;
wire n4145;
wire n4146;
wire n4147;
wire n4148;
wire n4149;
wire n4150;
wire n4151;
wire n4152;
wire n4153;
wire n4154;
wire n4155;
wire n4156;
wire n4157;
wire n4158;
wire n4159;
wire n4160;
wire n4161;
wire n4162;
wire n4163;
wire n4164;
wire n4165;
wire n4166;
wire n4167;
wire n4168;
wire n4169;
wire n4170;
wire n4171;
wire n4172;
wire n4173;
wire n4174;
wire n4175;
wire n4176;
wire n4177;
wire n4178;
wire n4179;
wire n4180;
wire n4181;
wire n4182;
wire n4183;
wire n4184;
wire n4185;
wire n4186;
wire n4187;
wire n4188;
wire n4189;
wire n4190;
wire n4191;
wire n4192;
wire n4193;
wire n4194;
wire n4195;
wire n4196;
wire n4197;
wire n4198;
wire n4199;
wire n4200;
wire n4201;
wire n4202;
wire n4203;
wire n4204;
wire n4205;
wire n4206;
wire n4207;
wire n4208;
wire n4209;
wire n4210;
wire n4211;
wire n4212;
wire n4213;
wire n4214;
wire n4215;
wire n4216;
wire n4217;
wire n4218;
wire n4219;
wire n4220;
wire n4221;
wire n4222;
wire n4223;
wire n4224;
wire n4225;
wire n4226;
wire n4227;
wire n4228;
wire n4229;
wire n4230;
wire n4231;
wire n4232;
wire n4233;
wire n4234;
wire n4235;
wire n4236;
wire n4237;
wire n4238;
wire n4239;
wire n4240;
wire n4241;
wire n4242;
wire n4243;
wire n4244;
wire n4245;
wire n4246;
wire n4247;
wire n4248;
wire n4249;
wire n4250;
wire n4251;
wire n4252;
wire n4253;
wire n4254;
wire n4255;
wire n4256;
wire n4257;
wire n4258;
wire n4259;
wire n4260;
wire n4261;
wire n4262;
wire n4263;
wire n4264;
wire n4265;
wire n4266;
wire n4267;
wire n4268;
wire n4269;
wire n4270;
wire n4271;
wire n4272;
wire n4273;
wire n4274;
wire n4275;
wire n4276;
wire n4277;
wire n4278;
wire n4279;
wire n4280;
wire n4281;
wire n4282;
wire n4283;
wire n4284;
wire n4285;
wire n4286;
wire n4287;
wire n4288;
wire n4289;
wire n4290;
wire n4291;
wire n4292;
wire n4293;
wire n4294;
wire n4295;
wire n4296;
wire n4297;
wire n4298;
wire n4299;
wire n4300;
wire n4301;
wire n4302;
wire n4303;
wire n4304;
wire n4305;
wire n4306;
wire n4307;
wire n4308;
wire n4309;
wire n4310;
wire n4311;
wire n4312;
wire n4313;
wire n4314;
wire n4315;
wire n4316;
wire n4317;
wire n4318;
wire n4319;
wire n4320;
wire n4321;
wire n4322;
wire n4323;
wire n4324;
wire n4325;
wire n4326;
wire n4327;
wire n4328;
wire n4329;
wire n4330;
wire n4331;
wire n4332;
wire n4333;
wire n4334;
wire n4335;
wire n4336;
wire n4337;
wire n4338;
wire n4339;
wire n4340;
wire n4341;
wire n4342;
wire n4343;
wire n4344;
wire n4345;
wire n4346;
wire n4347;
wire n4348;
wire n4349;
wire n4350;
wire n4351;
wire n4352;
wire n4353;
wire n4354;
wire n4355;
wire n4356;
wire n4357;
wire n4358;
wire n4359;
wire n4360;
wire n4361;
wire n4362;
wire n4363;
wire n4364;
wire n4365;
wire n4366;
wire n4367;
wire n4368;
wire n4369;
wire n4370;
wire n4371;
wire n4372;
wire n4373;
wire n4374;
wire n4375;
wire n4376;
wire n4377;
wire n4378;
wire n4379;
wire n4380;
wire n4381;
wire n4382;
wire n4383;
wire n4384;
wire n4385;
wire n4386;
wire n4387;
wire n4388;
wire n4389;
wire n4390;
wire n4391;
wire n4392;
wire n4393;
wire n4394;
wire n4395;
wire n4396;
wire n4397;
wire n4398;
wire n4399;
wire n4400;
wire n4401;
wire n4402;
wire n4403;
wire n4404;
wire n4405;
wire n4406;
wire n4407;
wire n4408;
wire n4409;
wire n4410;
wire n4411;
wire n4412;
wire n4413;
wire n4414;
wire n4415;
wire n4416;
wire n4417;
wire n4418;
wire n4419;
wire n4420;
wire n4421;
wire n4422;
wire n4423;
wire n4424;
wire n4425;
wire n4426;
wire n4427;
wire n4428;
wire n4429;
wire n4430;
wire n4431;
wire n4432;
wire n4433;
wire n4434;
wire n4435;
wire n4436;
wire n4437;
wire n4438;
wire n4439;
wire n4440;
wire n4441;
wire n4442;
wire n4443;
wire n4444;
wire n4445;
wire n4446;
wire n4447;
wire n4448;
wire n4449;
wire n4450;
wire n4451;
wire n4452;
wire n4453;
wire n4454;
wire n4455;
wire n4456;
wire n4457;
wire n4458;
wire n4459;
wire n4460;
wire n4461;
wire n4462;
wire n4463;
wire n4464;
wire n4465;
wire n4466;
wire n4467;
wire n4468;
wire n4469;
wire n4470;
wire n4471;
wire n4472;
wire n4473;
wire n4474;
wire n4475;
wire n4476;
wire n4477;
wire n4478;
wire n4479;
wire n4480;
wire n4481;
wire n4482;
wire n4483;
wire n4484;
wire n4485;
wire n4486;
wire n4487;
wire n4488;
wire n4489;
wire n4490;
wire n4491;
wire n4492;
wire n4493;
wire n4494;
wire n4495;
wire n4496;
wire n4497;
wire n4498;
wire n4499;
wire n4500;
wire n4501;
wire n4502;
wire n4503;
wire n4504;
wire n4505;
wire n4506;
wire n4507;
wire n4508;
wire n4509;
wire n4510;
wire n4511;
wire n4512;
wire n4513;
wire n4514;
wire n4515;
wire n4516;
wire n4517;
wire n4518;
wire n4519;
wire n4520;
wire n4521;
wire n4522;
wire n4523;
wire n4524;
wire n4525;
wire n4526;
wire n4527;
wire n4528;
wire n4529;
wire n4530;
wire n4531;
wire n4532;
wire n4533;
wire n4534;
wire n4535;
wire n4536;
wire n4537;
wire n4538;
wire n4539;
wire n4540;
wire n4541;
wire n4542;
wire n4543;
wire n4544;
wire n4545;
wire n4546;
wire n4547;
wire n4548;
wire n4549;
wire n4550;
wire n4551;
wire n4552;
wire n4553;
wire n4554;
wire n4555;
wire n4556;
wire n4557;
wire n4558;
wire n4559;
wire n4560;
wire n4561;
wire n4562;
wire n4563;
wire n4564;
wire n4565;
wire n4566;
wire n4567;
wire n4568;
wire n4569;
wire n4570;
wire n4571;
wire n4572;
wire n4573;
wire n4574;
wire n4575;
wire n4576;
wire n4577;
wire n4578;
wire n4579;
wire n4580;
wire n4581;
wire n4582;
wire n4583;
wire n4584;
wire n4585;
wire n4586;
wire n4587;
wire n4588;
wire n4589;
wire n4590;
wire n4591;
wire n4592;
wire n4593;
wire n4594;
wire n4595;
wire n4596;
wire n4597;
wire n4598;
wire n4599;
wire n4600;
wire n4601;
wire n4602;
wire n4603;
wire n4604;
wire n4605;
wire n4606;
wire n4607;
wire n4608;
wire n4609;
wire n4610;
wire n4611;
wire n4612;
wire n4613;
wire n4614;
wire n4615;
wire n4616;
wire n4617;
wire n4618;
wire n4619;
wire n4620;
wire n4621;
wire n4622;
wire n4623;
wire n4624;
wire n4625;
wire n4626;
wire n4627;
wire n4628;
wire n4629;
wire n4630;
wire n4631;
wire n4632;
wire n4633;
wire n4634;
wire n4635;
wire n4636;
wire n4637;
wire n4638;
wire n4639;
wire n4640;
wire n4641;
wire n4642;
wire n4643;
wire n4644;
wire n4645;
wire n4646;
wire n4647;
wire n4648;
wire n4649;
wire n4650;
wire n4651;
wire n4652;
wire n4653;
wire n4654;
wire n4655;
wire n4656;
wire n4657;
wire n4658;
wire n4659;
wire n4660;
wire n4661;
wire n4662;
wire n4663;
wire n4664;
wire n4665;
wire n4666;
wire n4667;
wire n4668;
wire n4669;
wire n4670;
wire n4671;
wire n4672;
wire n4673;
wire n4674;
wire n4675;
wire n4676;
wire n4677;
wire n4678;
wire n4679;
wire n4680;
wire n4681;
wire n4682;
wire n4683;
wire n4684;
wire n4685;
wire n4686;
wire n4687;
wire n4688;
wire n4689;
wire n4690;
wire n4691;
wire n4692;
wire n4693;
wire n4694;
wire n4695;
wire n4696;
wire n4697;
wire n4698;
wire n4699;
wire n4700;
wire n4701;
wire n4702;
wire n4703;
wire n4704;
wire n4705;
wire n4706;
wire n4707;
wire n4708;
wire n4709;
wire n4710;
wire n4711;
wire n4712;
wire n4713;
wire n4714;
wire n4715;
wire n4716;
wire n4717;
wire n4718;
wire n4719;
wire n4720;
wire n4721;
wire n4722;
wire n4723;
wire n4724;
wire n4725;
wire n4726;
wire n4727;
wire n4728;
wire n4729;
wire n4730;
wire n4731;
wire n4732;
wire n4733;
wire n4734;
wire n4735;
wire n4736;
wire n4737;
wire n4738;
wire n4739;
wire n4740;
wire n4741;
wire n4742;
wire n4743;
wire n4744;
wire n4745;
wire n4746;
wire n4747;
wire n4748;
wire n4749;
wire n4750;
wire n4751;
wire n4752;
wire n4753;
wire n4754;
wire n4755;
wire n4756;
wire n4757;
wire n4758;
wire n4759;
wire n4760;
wire n4761;
wire n4762;
wire n4763;
wire n4764;
wire n4765;
wire n4766;
wire n4767;
wire n4768;
wire n4769;
wire n4770;
wire n4771;
wire n4772;
wire n4773;
wire n4774;
wire n4775;
wire n4776;
wire n4777;
wire n4778;
wire n4779;
wire n4780;
wire n4781;
wire n4782;
wire n4783;
wire n4784;
wire n4785;
wire n4786;
wire n4787;
wire n4788;
wire n4789;
wire n4790;
wire n4791;
wire n4792;
wire n4793;
wire n4794;
wire n4795;
wire n4796;
wire n4797;
wire n4798;
wire n4799;
wire n4800;
wire n4801;
wire n4802;
wire n4803;
wire n4804;
wire n4805;
wire n4806;
wire n4807;
wire n4808;
wire n4809;
wire n4810;
wire n4811;
wire n4812;
wire n4813;
wire n4814;
wire n4815;
wire n4816;
wire n4817;
wire n4818;
wire n4819;
wire n4820;
wire n4821;
wire n4822;
wire n4823;
wire n4824;
wire n4825;
wire n4826;
wire n4827;
wire n4828;
wire n4829;
wire n4830;
wire n4831;
wire n4832;
wire n4833;
wire n4834;
wire n4835;
wire n4836;
wire n4837;
wire n4838;
wire n4839;
wire n4840;
wire n4841;
wire n4842;
wire n4843;
wire n4844;
wire n4845;
wire n4846;
wire n4847;
wire n4848;
wire n4849;
wire n4850;
wire n4851;
wire n4852;
wire n4853;
wire n4854;
wire n4855;
wire n4856;
wire n4857;
wire n4858;
wire n4859;
wire n4860;
wire n4861;
wire n4862;
wire n4863;
wire n4864;
wire n4865;
wire n4866;
wire n4867;
wire n4868;
wire n4869;
wire n4870;
wire n4871;
wire n4872;
wire n4873;
wire n4874;
wire n4875;
wire n4876;
wire n4877;
wire n4878;
wire n4879;
wire n4880;
wire n4881;
wire n4882;
wire n4883;
wire n4884;
wire n4885;
wire n4886;
wire n4887;
wire n4888;
wire n4889;
wire n4890;
wire n4891;
wire n4892;
wire n4893;
wire n4894;
wire n4895;
wire n4896;
wire n4897;
wire n4898;
wire n4899;
wire n4900;
wire n4901;
wire n4902;
wire n4903;
wire n4904;
wire n4905;
wire n4906;
wire n4907;
wire n4908;
wire n4909;
wire n4910;
wire n4911;
wire n4912;
wire n4913;
wire n4914;
wire n4915;
wire n4916;
wire n4917;
wire n4918;
wire n4919;
wire n4920;
wire n4921;
wire n4922;
wire n4923;
wire n4924;
wire n4925;
wire n4926;
wire n4927;
wire n4928;
wire n4929;
wire n4930;
wire n4931;
wire n4932;
wire n4933;
wire n4934;
wire n4935;
wire n4936;
wire n4937;
wire n4938;
wire n4939;
wire n4940;
wire n4941;
wire n4942;
wire n4943;
wire n4944;
wire n4945;
wire n4946;
wire n4947;
wire n4948;
wire n4949;
wire n4950;
wire n4951;
wire n4952;
wire n4953;
wire n4954;
wire n4955;
wire n4956;
wire n4957;
wire n4958;
wire n4959;
wire n4960;
wire n4961;
wire n4962;
wire n4963;
wire n4964;
wire n4965;
wire n4966;
wire n4967;
wire n4968;
wire n4969;
wire n4970;
wire n4971;
wire n4972;
wire n4973;
wire n4974;
wire n4975;
wire n4976;
wire n4977;
wire n4978;
wire n4979;
wire n4980;
wire n4981;
wire n4982;
wire n4983;
wire n4984;
wire n4985;
wire n4986;
wire n4987;
wire n4988;
wire n4989;
wire n4990;
wire n4991;
wire n4992;
wire n4993;
wire n4994;
wire n4995;
wire n4996;
wire n4997;
wire n4998;
wire n4999;
wire n5000;
wire n5001;
wire n5002;
wire n5003;
wire n5004;
wire n5005;
wire n5006;
wire n5007;
wire n5008;
wire n5009;
wire n5010;
wire n5011;
wire n5012;
wire n5013;
wire n5014;
wire n5015;
wire n5016;
wire n5017;
wire n5018;
wire n5019;
wire n5020;
wire n5021;
wire n5022;
wire n5023;
wire n5024;
wire n5025;
wire n5026;
wire n5027;
wire n5028;
wire n5029;
wire n5030;
wire n5031;
wire n5032;
wire n5033;
wire n5034;
wire n5035;
wire n5036;
wire n5037;
wire n5038;
wire n5039;
wire n5040;
wire n5041;
wire n5042;
wire n5043;
wire n5044;
wire n5045;
wire n5046;
wire n5047;
wire n5048;
wire n5049;
wire n5050;
wire n5051;
wire n5052;
wire n5053;
wire n5054;
wire n5055;
wire n5056;
wire n5057;
wire n5058;
wire n5059;
wire n5060;
wire n5061;
wire n5062;
wire n5063;
wire n5064;
wire n5065;
wire n5066;
wire n5067;
wire n5068;
wire n5069;
wire n5070;
wire n5071;
wire n5072;
wire n5073;
wire n5074;
wire n5075;
wire n5076;
wire n5077;
wire n5078;
wire n5079;
wire n5080;
wire n5081;
wire n5082;
wire n5083;
wire n5084;
wire n5085;
wire n5086;
wire n5087;
wire n5088;
wire n5089;
wire n5090;
wire n5091;
wire n5092;
wire n5093;
wire n5094;
wire n5095;
wire n5096;
wire n5097;
wire n5098;
wire n5099;
wire n5100;
wire n5101;
wire n5102;
wire n5103;
wire n5104;
wire n5105;
wire n5106;
wire n5107;
wire n5108;
wire n5109;
wire n5110;
wire n5111;
wire n5112;
wire n5113;
wire n5114;
wire n5115;
wire n5116;
wire n5117;
wire n5118;
wire n5119;
wire n5120;
wire n5121;
wire n5122;
wire n5123;
wire n5124;
wire n5125;
wire n5126;
wire n5127;
wire n5128;
wire n5129;
wire n5130;
wire n5131;
wire n5132;
wire n5133;
wire n5134;
wire n5135;
wire n5136;
wire n5137;
wire n5138;
wire n5139;
wire n5140;
wire n5141;
wire n5142;
wire n5143;
wire n5144;
wire n5145;
wire n5146;
wire n5147;
wire n5148;
wire n5149;
wire n5150;
xor (out,n0,n2895);
nand (n0,n1,n2894);
or (n1,n2,n1280);
not (n2,n3);
nor (n3,n4,n1279);
and (n4,n5,n1156);
xor (n5,n6,n1040);
xor (n6,n7,n884);
xor (n7,n8,n586);
xor (n8,n9,n485);
xor (n9,n10,n392);
xor (n10,n11,n285);
xor (n11,n12,n249);
xor (n12,n13,n133);
nor (n13,n14,n130);
nor (n14,n15,n128);
and (n15,n16,n122);
not (n16,n17);
wire s0n17,s1n17,notn17;
or (n17,s0n17,s1n17);
not(notn17,n119);
and (s0n17,notn17,n18);
and (s1n17,n119,n37);
wire s0n18,s1n18,notn18;
or (n18,s0n18,s1n18);
not(notn18,n21);
and (s0n18,notn18,1'b0);
and (s1n18,n21,n20);
or (n21,n22,n33);
or (n22,n23,n31);
nor (n23,n24,n26,n27,n28,n30);
not (n24,n25);
not (n28,n29);
nor (n31,n25,n32,n27,n28,n30);
not (n32,n26);
or (n33,n34,n36);
and (n34,n24,n26,n27,n28,n35);
not (n35,n30);
nor (n36,n24,n32,n27,n28,n30);
xor (n37,n38,n39);
not (n38,n20);
and (n39,n40,n42);
not (n40,n41);
and (n42,n43,n45);
not (n43,n44);
and (n45,n46,n48);
not (n46,n47);
and (n48,n49,n51);
not (n49,n50);
and (n51,n52,n54);
not (n52,n53);
and (n54,n55,n57);
not (n55,n56);
and (n57,n58,n60);
not (n58,n59);
and (n60,n61,n63);
not (n61,n62);
and (n63,n64,n66);
not (n64,n65);
and (n66,n67,n69);
not (n67,n68);
and (n69,n70,n72);
not (n70,n71);
and (n72,n73,n75);
not (n73,n74);
and (n75,n76,n78);
not (n76,n77);
and (n78,n79,n81);
not (n79,n80);
and (n81,n82,n84);
not (n82,n83);
and (n84,n85,n87);
not (n85,n86);
and (n87,n88,n90);
not (n88,n89);
and (n90,n91,n93);
not (n91,n92);
and (n93,n94,n96);
not (n94,n95);
and (n96,n97,n99);
not (n97,n98);
and (n99,n100,n102);
not (n100,n101);
and (n102,n103,n105);
not (n103,n104);
and (n105,n106,n108);
not (n106,n107);
and (n108,n109,n111);
not (n109,n110);
and (n111,n112,n114);
not (n112,n113);
and (n114,n115,n117);
not (n115,n116);
not (n117,n118);
and (n119,n120,n121);
or (n120,n23,n34);
wire s0n122,s1n122,notn122;
or (n122,s0n122,s1n122);
not(notn122,n119);
and (s0n122,notn122,n123);
and (s1n122,n119,n125);
wire s0n123,s1n123,notn123;
or (n123,s0n123,s1n123);
not(notn123,n21);
and (s0n123,notn123,1'b0);
and (s1n123,n21,n124);
xor (n125,n126,n127);
not (n126,n124);
and (n127,n38,n39);
and (n128,n17,n129);
not (n129,n122);
not (n130,n131);
wire s0n131,s1n131,notn131;
or (n131,s0n131,s1n131);
not(notn131,n21);
and (s0n131,notn131,1'b0);
and (s1n131,n21,n132);
nand (n133,n134,n238);
or (n134,n135,n154);
nand (n135,n136,n147);
nor (n136,n137,n145);
and (n137,n138,n142);
not (n138,n139);
wire s0n139,s1n139,notn139;
or (n139,s0n139,s1n139);
not(notn139,n119);
and (s0n139,notn139,n140);
and (s1n139,n119,n141);
wire s0n140,s1n140,notn140;
or (n140,s0n140,s1n140);
not(notn140,n21);
and (s0n140,notn140,1'b0);
and (s1n140,n21,n116);
xor (n141,n115,n117);
wire s0n142,s1n142,notn142;
or (n142,s0n142,s1n142);
not(notn142,n119);
and (s0n142,notn142,n143);
and (s1n142,n119,n144);
wire s0n143,s1n143,notn143;
or (n143,s0n143,s1n143);
not(notn143,n21);
and (s0n143,notn143,1'b0);
and (s1n143,n21,n113);
xor (n144,n112,n114);
and (n145,n139,n146);
not (n146,n142);
nand (n147,n148,n153);
or (n148,n149,n142);
not (n149,n150);
wire s0n150,s1n150,notn150;
or (n150,s0n150,s1n150);
not(notn150,n119);
and (s0n150,notn150,n151);
and (s1n150,n119,n152);
wire s0n151,s1n151,notn151;
or (n151,s0n151,s1n151);
not(notn151,n21);
and (s0n151,notn151,1'b0);
and (s1n151,n21,n110);
xor (n152,n109,n111);
nand (n153,n149,n142);
nor (n154,n155,n236);
and (n155,n156,n149);
wire s0n156,s1n156,notn156;
or (n156,s0n156,s1n156);
not(notn156,n234);
and (s0n156,notn156,n157);
and (s1n156,n234,n159);
wire s0n157,s1n157,notn157;
or (n157,s0n157,s1n157);
not(notn157,n21);
and (s0n157,notn157,1'b0);
and (s1n157,n21,n158);
xor (n159,n160,n161);
not (n160,n158);
and (n161,n162,n164);
not (n162,n163);
and (n164,n165,n167);
not (n165,n166);
and (n167,n168,n170);
not (n168,n169);
and (n170,n171,n173);
not (n171,n172);
and (n173,n174,n176);
not (n174,n175);
and (n176,n177,n179);
not (n177,n178);
and (n179,n180,n182);
not (n180,n181);
and (n182,n183,n185);
not (n183,n184);
and (n185,n186,n188);
not (n186,n187);
and (n188,n189,n191);
not (n189,n190);
and (n191,n192,n194);
not (n192,n193);
and (n194,n195,n197);
not (n195,n196);
and (n197,n198,n200);
not (n198,n199);
and (n200,n201,n203);
not (n201,n202);
and (n203,n204,n206);
not (n204,n205);
and (n206,n207,n209);
not (n207,n208);
and (n209,n210,n212);
not (n210,n211);
and (n212,n213,n215);
not (n213,n214);
and (n215,n216,n218);
not (n216,n217);
and (n218,n219,n221);
not (n219,n220);
and (n221,n222,n224);
not (n222,n223);
and (n224,n225,n227);
not (n225,n226);
and (n227,n228,n230);
not (n228,n229);
and (n230,n231,n233);
not (n231,n232);
not (n233,n132);
and (n234,n120,n235);
and (n236,n237,n150);
not (n237,n156);
or (n238,n239,n136);
nor (n239,n240,n247);
and (n240,n241,n149);
wire s0n241,s1n241,notn241;
or (n241,s0n241,s1n241);
not(notn241,n234);
and (s0n241,notn241,n242);
and (s1n241,n234,n244);
wire s0n242,s1n242,notn242;
or (n242,s0n242,s1n242);
not(notn242,n21);
and (s0n242,notn242,1'b0);
and (s1n242,n21,n243);
xor (n244,n245,n246);
not (n245,n243);
and (n246,n160,n161);
and (n247,n248,n150);
not (n248,n241);
nand (n249,n250,n277);
or (n250,n251,n270);
nand (n251,n252,n263);
or (n252,n253,n260);
and (n253,n254,n257);
wire s0n254,s1n254,notn254;
or (n254,s0n254,s1n254);
not(notn254,n119);
and (s0n254,notn254,n255);
and (s1n254,n119,n256);
wire s0n255,s1n255,notn255;
or (n255,s0n255,s1n255);
not(notn255,n21);
and (s0n255,notn255,1'b0);
and (s1n255,n21,n104);
xor (n256,n103,n105);
wire s0n257,s1n257,notn257;
or (n257,s0n257,s1n257);
not(notn257,n119);
and (s0n257,notn257,n258);
and (s1n257,n119,n259);
wire s0n258,s1n258,notn258;
or (n258,s0n258,s1n258);
not(notn258,n21);
and (s0n258,notn258,1'b0);
and (s1n258,n21,n101);
xor (n259,n100,n102);
and (n260,n261,n262);
not (n261,n254);
not (n262,n257);
nor (n263,n264,n268);
and (n264,n265,n257);
wire s0n265,s1n265,notn265;
or (n265,s0n265,s1n265);
not(notn265,n119);
and (s0n265,notn265,n266);
and (s1n265,n119,n267);
wire s0n266,s1n266,notn266;
or (n266,s0n266,s1n266);
not(notn266,n21);
and (s0n266,notn266,1'b0);
and (s1n266,n21,n98);
xor (n267,n97,n99);
and (n268,n269,n262);
not (n269,n265);
nor (n270,n271,n275);
and (n271,n272,n269);
wire s0n272,s1n272,notn272;
or (n272,s0n272,s1n272);
not(notn272,n234);
and (s0n272,notn272,n273);
and (s1n272,n234,n274);
wire s0n273,s1n273,notn273;
or (n273,s0n273,s1n273);
not(notn273,n21);
and (s0n273,notn273,1'b0);
and (s1n273,n21,n172);
xor (n274,n171,n173);
and (n275,n276,n265);
not (n276,n272);
or (n277,n278,n252);
nor (n278,n279,n283);
and (n279,n280,n269);
wire s0n280,s1n280,notn280;
or (n280,s0n280,s1n280);
not(notn280,n234);
and (s0n280,notn280,n281);
and (s1n280,n234,n282);
wire s0n281,s1n281,notn281;
or (n281,s0n281,s1n281);
not(notn281,n21);
and (s0n281,notn281,1'b0);
and (s1n281,n21,n169);
xor (n282,n168,n170);
and (n283,n284,n265);
not (n284,n280);
or (n285,n286,n391);
and (n286,n287,n357);
xor (n287,n288,n324);
nand (n288,n289,n316);
or (n289,n290,n309);
nand (n290,n291,n302);
nor (n291,n292,n300);
and (n292,n293,n297);
not (n293,n294);
wire s0n294,s1n294,notn294;
or (n294,s0n294,s1n294);
not(notn294,n119);
and (s0n294,notn294,n295);
and (s1n294,n119,n296);
wire s0n295,s1n295,notn295;
or (n295,s0n295,s1n295);
not(notn295,n21);
and (s0n295,notn295,1'b0);
and (s1n295,n21,n62);
xor (n296,n61,n63);
wire s0n297,s1n297,notn297;
or (n297,s0n297,s1n297);
not(notn297,n119);
and (s0n297,notn297,n298);
and (s1n297,n119,n299);
wire s0n298,s1n298,notn298;
or (n298,s0n298,s1n298);
not(notn298,n21);
and (s0n298,notn298,1'b0);
and (s1n298,n21,n59);
xor (n299,n58,n60);
and (n300,n294,n301);
not (n301,n297);
nand (n302,n303,n307);
or (n303,n301,n304);
wire s0n304,s1n304,notn304;
or (n304,s0n304,s1n304);
not(notn304,n119);
and (s0n304,notn304,n305);
and (s1n304,n119,n306);
wire s0n305,s1n305,notn305;
or (n305,s0n305,s1n305);
not(notn305,n21);
and (s0n305,notn305,1'b0);
and (s1n305,n21,n56);
xor (n306,n55,n57);
or (n307,n297,n308);
not (n308,n304);
nor (n309,n310,n314);
and (n310,n308,n311);
wire s0n311,s1n311,notn311;
or (n311,s0n311,s1n311);
not(notn311,n234);
and (s0n311,notn311,n312);
and (s1n311,n234,n313);
wire s0n312,s1n312,notn312;
or (n312,s0n312,s1n312);
not(notn312,n21);
and (s0n312,notn312,1'b0);
and (s1n312,n21,n217);
xor (n313,n216,n218);
and (n314,n315,n304);
not (n315,n311);
or (n316,n291,n317);
nor (n317,n318,n322);
and (n318,n308,n319);
wire s0n319,s1n319,notn319;
or (n319,s0n319,s1n319);
not(notn319,n234);
and (s0n319,notn319,n320);
and (s1n319,n234,n321);
wire s0n320,s1n320,notn320;
or (n320,s0n320,s1n320);
not(notn320,n21);
and (s0n320,notn320,1'b0);
and (s1n320,n21,n214);
xor (n321,n213,n215);
and (n322,n323,n304);
not (n323,n319);
nand (n324,n325,n349);
or (n325,n326,n342);
or (n326,n327,n335);
not (n327,n328);
and (n328,n329,n334);
nand (n329,n330,n304);
not (n330,n331);
wire s0n331,s1n331,notn331;
or (n331,s0n331,s1n331);
not(notn331,n119);
and (s0n331,notn331,n332);
and (s1n331,n119,n333);
wire s0n332,s1n332,notn332;
or (n332,s0n332,s1n332);
not(notn332,n21);
and (s0n332,notn332,1'b0);
and (s1n332,n21,n53);
xor (n333,n52,n54);
nand (n334,n331,n308);
nor (n335,n336,n341);
and (n336,n331,n337);
not (n337,n338);
wire s0n338,s1n338,notn338;
or (n338,s0n338,s1n338);
not(notn338,n119);
and (s0n338,notn338,n339);
and (s1n338,n119,n340);
wire s0n339,s1n339,notn339;
or (n339,s0n339,s1n339);
not(notn339,n21);
and (s0n339,notn339,1'b0);
and (s1n339,n21,n50);
xor (n340,n49,n51);
and (n341,n330,n338);
nor (n342,n343,n347);
and (n343,n337,n344);
wire s0n344,s1n344,notn344;
or (n344,s0n344,s1n344);
not(notn344,n234);
and (s0n344,notn344,n345);
and (s1n344,n234,n346);
wire s0n345,s1n345,notn345;
or (n345,s0n345,s1n345);
not(notn345,n21);
and (s0n345,notn345,1'b0);
and (s1n345,n21,n223);
xor (n346,n222,n224);
and (n347,n348,n338);
not (n348,n344);
or (n349,n328,n350);
nor (n350,n351,n355);
and (n351,n337,n352);
wire s0n352,s1n352,notn352;
or (n352,s0n352,s1n352);
not(notn352,n234);
and (s0n352,notn352,n353);
and (s1n352,n234,n354);
wire s0n353,s1n353,notn353;
or (n353,s0n353,s1n353);
not(notn353,n21);
and (s0n353,notn353,1'b0);
and (s1n353,n21,n220);
xor (n354,n219,n221);
and (n355,n356,n338);
not (n356,n352);
nand (n357,n358,n383);
or (n358,n359,n376);
nand (n359,n360,n373);
or (n360,n361,n370);
not (n361,n362);
nand (n362,n363,n366);
wire s0n363,s1n363,notn363;
or (n363,s0n363,s1n363);
not(notn363,n119);
and (s0n363,notn363,n364);
and (s1n363,n119,n365);
wire s0n364,s1n364,notn364;
or (n364,s0n364,s1n364);
not(notn364,n21);
and (s0n364,notn364,1'b0);
and (s1n364,n21,n47);
xor (n365,n46,n48);
not (n366,n367);
wire s0n367,s1n367,notn367;
or (n367,s0n367,s1n367);
not(notn367,n119);
and (s0n367,notn367,n368);
and (s1n367,n119,n369);
wire s0n368,s1n368,notn368;
or (n368,s0n368,s1n368);
not(notn368,n21);
and (s0n368,notn368,1'b0);
and (s1n368,n21,n44);
xor (n369,n43,n45);
not (n370,n371);
nand (n371,n372,n367);
not (n372,n363);
and (n373,n374,n375);
nand (n374,n372,n338);
nand (n375,n363,n337);
nor (n376,n377,n381);
and (n377,n378,n366);
wire s0n378,s1n378,notn378;
or (n378,s0n378,s1n378);
not(notn378,n234);
and (s0n378,notn378,n379);
and (s1n378,n234,n380);
wire s0n379,s1n379,notn379;
or (n379,s0n379,s1n379);
not(notn379,n21);
and (s0n379,notn379,1'b0);
and (s1n379,n21,n229);
xor (n380,n228,n230);
and (n381,n382,n367);
not (n382,n378);
or (n383,n373,n384);
nor (n384,n385,n389);
and (n385,n386,n366);
wire s0n386,s1n386,notn386;
or (n386,s0n386,s1n386);
not(notn386,n234);
and (s0n386,notn386,n387);
and (s1n386,n234,n388);
wire s0n387,s1n387,notn387;
or (n387,s0n387,s1n387);
not(notn387,n21);
and (s0n387,notn387,1'b0);
and (s1n387,n21,n226);
xor (n388,n225,n227);
and (n389,n390,n367);
not (n390,n386);
and (n391,n288,n324);
xor (n392,n393,n456);
xor (n393,n394,n420);
nand (n394,n395,n409);
or (n395,n396,n406);
nor (n396,n397,n404);
and (n397,n398,n138);
wire s0n398,s1n398,notn398;
or (n398,s0n398,s1n398);
not(notn398,n234);
and (s0n398,notn398,n399);
and (s1n398,n234,n401);
wire s0n399,s1n399,notn399;
or (n399,s0n399,s1n399);
not(notn399,n21);
and (s0n399,notn399,1'b0);
and (s1n399,n21,n400);
xor (n401,n402,n403);
not (n402,n400);
and (n403,n245,n246);
and (n404,n405,n139);
not (n405,n398);
nand (n406,n139,n407);
not (n407,n408);
wire s0n408,s1n408,notn408;
or (n408,s0n408,s1n408);
not(notn408,n21);
and (s0n408,notn408,1'b0);
and (s1n408,n21,n118);
or (n409,n410,n407);
nor (n410,n411,n418);
and (n411,n412,n138);
wire s0n412,s1n412,notn412;
or (n412,s0n412,s1n412);
not(notn412,n234);
and (s0n412,notn412,n413);
and (s1n412,n234,n415);
wire s0n413,s1n413,notn413;
or (n413,s0n413,s1n413);
not(notn413,n21);
and (s0n413,notn413,1'b0);
and (s1n413,n21,n414);
xor (n415,n416,n417);
not (n416,n414);
and (n417,n402,n403);
and (n418,n419,n139);
not (n419,n412);
nand (n420,n421,n448);
or (n421,n422,n441);
nand (n422,n423,n434);
or (n423,n424,n431);
and (n424,n425,n428);
wire s0n425,s1n425,notn425;
or (n425,s0n425,s1n425);
not(notn425,n119);
and (s0n425,notn425,n426);
and (s1n425,n119,n427);
wire s0n426,s1n426,notn426;
or (n426,s0n426,s1n426);
not(notn426,n21);
and (s0n426,notn426,1'b0);
and (s1n426,n21,n89);
xor (n427,n88,n90);
wire s0n428,s1n428,notn428;
or (n428,s0n428,s1n428);
not(notn428,n119);
and (s0n428,notn428,n429);
and (s1n428,n119,n430);
wire s0n429,s1n429,notn429;
or (n429,s0n429,s1n429);
not(notn429,n21);
and (s0n429,notn429,1'b0);
and (s1n429,n21,n92);
xor (n430,n91,n93);
and (n431,n432,n433);
not (n432,n425);
not (n433,n428);
nand (n434,n435,n439);
or (n435,n432,n436);
wire s0n436,s1n436,notn436;
or (n436,s0n436,s1n436);
not(notn436,n119);
and (s0n436,notn436,n437);
and (s1n436,n119,n438);
wire s0n437,s1n437,notn437;
or (n437,s0n437,s1n437);
not(notn437,n21);
and (s0n437,notn437,1'b0);
and (s1n437,n21,n86);
xor (n438,n85,n87);
or (n439,n440,n425);
not (n440,n436);
nor (n441,n442,n446);
and (n442,n443,n440);
wire s0n443,s1n443,notn443;
or (n443,s0n443,s1n443);
not(notn443,n234);
and (s0n443,notn443,n444);
and (s1n443,n234,n445);
wire s0n444,s1n444,notn444;
or (n444,s0n444,s1n444);
not(notn444,n21);
and (s0n444,notn444,1'b0);
and (s1n444,n21,n184);
xor (n445,n183,n185);
and (n446,n447,n436);
not (n447,n443);
or (n448,n423,n449);
nor (n449,n450,n454);
and (n450,n440,n451);
wire s0n451,s1n451,notn451;
or (n451,s0n451,s1n451);
not(notn451,n234);
and (s0n451,notn451,n452);
and (s1n451,n234,n453);
wire s0n452,s1n452,notn452;
or (n452,s0n452,s1n452);
not(notn452,n21);
and (s0n452,notn452,1'b0);
and (s1n452,n21,n181);
xor (n453,n180,n182);
and (n454,n455,n436);
not (n455,n451);
nand (n456,n457,n477);
or (n457,n458,n470);
nand (n458,n459,n466);
not (n459,n460);
nand (n460,n461,n465);
or (n461,n149,n462);
wire s0n462,s1n462,notn462;
or (n462,s0n462,s1n462);
not(notn462,n119);
and (s0n462,notn462,n463);
and (s1n462,n119,n464);
wire s0n463,s1n463,notn463;
or (n463,s0n463,s1n463);
not(notn463,n21);
and (s0n463,notn463,1'b0);
and (s1n463,n21,n107);
xor (n464,n106,n108);
nand (n465,n462,n149);
nor (n466,n467,n469);
and (n467,n261,n468);
not (n468,n462);
and (n469,n254,n462);
nor (n470,n471,n475);
and (n471,n472,n261);
wire s0n472,s1n472,notn472;
or (n472,s0n472,s1n472);
not(notn472,n234);
and (s0n472,notn472,n473);
and (s1n472,n234,n474);
wire s0n473,s1n473,notn473;
or (n473,s0n473,s1n473);
not(notn473,n21);
and (s0n473,notn473,1'b0);
and (s1n473,n21,n166);
xor (n474,n165,n167);
and (n475,n476,n254);
not (n476,n472);
or (n477,n478,n459);
nor (n478,n479,n483);
and (n479,n480,n261);
wire s0n480,s1n480,notn480;
or (n480,s0n480,s1n480);
not(notn480,n234);
and (s0n480,notn480,n481);
and (s1n480,n234,n482);
wire s0n481,s1n481,notn481;
or (n481,s0n481,s1n481);
not(notn481,n21);
and (s0n481,notn481,1'b0);
and (s1n481,n21,n163);
xor (n482,n162,n164);
and (n483,n484,n254);
not (n484,n480);
or (n485,n486,n585);
and (n486,n487,n525);
xor (n487,n488,n489);
xor (n488,n287,n357);
or (n489,n490,n524);
and (n490,n491,n508);
xor (n491,n492,n498);
nand (n492,n493,n497);
or (n493,n326,n494);
nor (n494,n495,n496);
and (n495,n386,n337);
and (n496,n390,n338);
or (n497,n328,n342);
nand (n498,n499,n507);
or (n499,n359,n500);
nor (n500,n501,n505);
and (n501,n502,n366);
wire s0n502,s1n502,notn502;
or (n502,s0n502,s1n502);
not(notn502,n234);
and (s0n502,notn502,n503);
and (s1n502,n234,n504);
wire s0n503,s1n503,notn503;
or (n503,s0n503,s1n503);
not(notn503,n21);
and (s0n503,notn503,1'b0);
and (s1n503,n21,n232);
xor (n504,n231,n233);
and (n505,n506,n367);
not (n506,n502);
or (n507,n376,n373);
and (n508,n509,n515);
nor (n509,n510,n366);
nor (n510,n511,n514);
and (n511,n512,n337);
not (n512,n513);
and (n513,n131,n363);
and (n514,n372,n130);
nand (n515,n516,n520);
or (n516,n135,n517);
nor (n517,n518,n519);
and (n518,n280,n149);
and (n519,n284,n150);
or (n520,n136,n521);
nor (n521,n522,n523);
and (n522,n472,n149);
and (n523,n476,n150);
and (n524,n492,n498);
xor (n525,n526,n560);
xor (n526,n527,n547);
nand (n527,n528,n543);
or (n528,n529,n540);
nand (n529,n530,n537);
nor (n530,n531,n535);
and (n531,n366,n532);
wire s0n532,s1n532,notn532;
or (n532,s0n532,s1n532);
not(notn532,n119);
and (s0n532,notn532,n533);
and (s1n532,n119,n534);
wire s0n533,s1n533,notn533;
or (n533,s0n533,s1n533);
not(notn533,n21);
and (s0n533,notn533,1'b0);
and (s1n533,n21,n41);
xor (n534,n40,n42);
and (n535,n367,n536);
not (n536,n532);
nand (n537,n538,n539);
or (n538,n536,n17);
or (n539,n532,n16);
nor (n540,n541,n542);
and (n541,n17,n130);
and (n542,n16,n131);
or (n543,n530,n544);
nor (n544,n545,n546);
and (n545,n16,n502);
and (n546,n506,n17);
xor (n547,n548,n554);
nor (n548,n549,n16);
nor (n549,n550,n553);
and (n550,n366,n551);
not (n551,n552);
and (n552,n131,n532);
and (n553,n536,n130);
nand (n554,n555,n559);
or (n555,n135,n556);
nor (n556,n557,n558);
and (n557,n480,n149);
and (n558,n484,n150);
or (n559,n154,n136);
or (n560,n561,n584);
and (n561,n562,n567);
xor (n562,n563,n564);
nor (n563,n530,n130);
nand (n564,n565,n566);
or (n565,n135,n521);
or (n566,n556,n136);
nand (n567,n568,n576);
or (n568,n251,n569);
nor (n569,n570,n574);
and (n570,n571,n269);
wire s0n571,s1n571,notn571;
or (n571,s0n571,s1n571);
not(notn571,n234);
and (s0n571,notn571,n572);
and (s1n571,n234,n573);
wire s0n572,s1n572,notn572;
or (n572,s0n572,s1n572);
not(notn572,n21);
and (s0n572,notn572,1'b0);
and (s1n572,n21,n178);
xor (n573,n177,n179);
and (n574,n575,n265);
not (n575,n571);
or (n576,n577,n252);
nor (n577,n578,n582);
and (n578,n579,n269);
wire s0n579,s1n579,notn579;
or (n579,s0n579,s1n579);
not(notn579,n234);
and (s0n579,notn579,n580);
and (s1n579,n234,n581);
wire s0n580,s1n580,notn580;
or (n580,s0n580,s1n580);
not(notn580,n21);
and (s0n580,notn580,1'b0);
and (s1n580,n21,n175);
xor (n581,n174,n176);
and (n582,n583,n265);
not (n583,n579);
and (n584,n563,n564);
and (n585,n488,n489);
or (n586,n587,n883);
and (n587,n588,n842);
xor (n588,n589,n754);
or (n589,n590,n753);
and (n590,n591,n728);
xor (n591,n592,n673);
or (n592,n593,n672);
and (n593,n594,n639);
xor (n594,n595,n601);
nand (n595,n596,n600);
or (n596,n251,n597);
nor (n597,n598,n599);
and (n598,n451,n269);
and (n599,n455,n265);
or (n600,n569,n252);
nand (n601,n602,n630);
or (n602,n603,n623);
not (n603,n604);
nor (n604,n605,n615);
nand (n605,n606,n614);
or (n606,n607,n611);
not (n607,n608);
wire s0n608,s1n608,notn608;
or (n608,s0n608,s1n608);
not(notn608,n119);
and (s0n608,notn608,n609);
and (s1n608,n119,n610);
wire s0n609,s1n609,notn609;
or (n609,s0n609,s1n609);
not(notn609,n21);
and (s0n609,notn609,1'b0);
and (s1n609,n21,n80);
xor (n610,n79,n81);
wire s0n611,s1n611,notn611;
or (n611,s0n611,s1n611);
not(notn611,n119);
and (s0n611,notn611,n612);
and (s1n611,n119,n613);
wire s0n612,s1n612,notn612;
or (n612,s0n612,s1n612);
not(notn612,n21);
and (s0n612,notn612,1'b0);
and (s1n612,n21,n77);
xor (n613,n76,n78);
nand (n614,n607,n611);
nor (n615,n616,n621);
and (n616,n617,n611);
not (n617,n618);
wire s0n618,s1n618,notn618;
or (n618,s0n618,s1n618);
not(notn618,n119);
and (s0n618,notn618,n619);
and (s1n618,n119,n620);
wire s0n619,s1n619,notn619;
or (n619,s0n619,s1n619);
not(notn619,n21);
and (s0n619,notn619,1'b0);
and (s1n619,n21,n74);
xor (n620,n73,n75);
and (n621,n622,n618);
not (n622,n611);
nor (n623,n624,n628);
and (n624,n617,n625);
wire s0n625,s1n625,notn625;
or (n625,s0n625,s1n625);
not(notn625,n234);
and (s0n625,notn625,n626);
and (s1n625,n234,n627);
wire s0n626,s1n626,notn626;
or (n626,s0n626,s1n626);
not(notn626,n21);
and (s0n626,notn626,1'b0);
and (s1n626,n21,n205);
xor (n627,n204,n206);
and (n628,n618,n629);
not (n629,n625);
or (n630,n631,n632);
not (n631,n605);
nor (n632,n633,n637);
and (n633,n617,n634);
wire s0n634,s1n634,notn634;
or (n634,s0n634,s1n634);
not(notn634,n234);
and (s0n634,notn634,n635);
and (s1n634,n234,n636);
wire s0n635,s1n635,notn635;
or (n635,s0n635,s1n635);
not(notn635,n21);
and (s0n635,notn635,1'b0);
and (s1n635,n21,n202);
xor (n636,n201,n203);
and (n637,n618,n638);
not (n638,n634);
nand (n639,n640,n664);
or (n640,n641,n657);
not (n641,n642);
and (n642,n643,n650);
nor (n643,n644,n649);
and (n644,n618,n645);
not (n645,n646);
wire s0n646,s1n646,notn646;
or (n646,s0n646,s1n646);
not(notn646,n119);
and (s0n646,notn646,n647);
and (s1n646,n119,n648);
wire s0n647,s1n647,notn647;
or (n647,s0n647,s1n647);
not(notn647,n21);
and (s0n647,notn647,1'b0);
and (s1n647,n21,n71);
xor (n648,n70,n72);
and (n649,n617,n646);
nand (n650,n651,n655);
or (n651,n645,n652);
wire s0n652,s1n652,notn652;
or (n652,s0n652,s1n652);
not(notn652,n119);
and (s0n652,notn652,n653);
and (s1n652,n119,n654);
wire s0n653,s1n653,notn653;
or (n653,s0n653,s1n653);
not(notn653,n21);
and (s0n653,notn653,1'b0);
and (s1n653,n21,n68);
xor (n654,n67,n69);
or (n655,n656,n646);
not (n656,n652);
nor (n657,n658,n662);
and (n658,n656,n659);
wire s0n659,s1n659,notn659;
or (n659,s0n659,s1n659);
not(notn659,n234);
and (s0n659,notn659,n660);
and (s1n659,n234,n661);
wire s0n660,s1n660,notn660;
or (n660,s0n660,s1n660);
not(notn660,n21);
and (s0n660,notn660,1'b0);
and (s1n660,n21,n211);
xor (n661,n210,n212);
and (n662,n652,n663);
not (n663,n659);
or (n664,n665,n643);
nor (n665,n666,n670);
and (n666,n656,n667);
wire s0n667,s1n667,notn667;
or (n667,s0n667,s1n667);
not(notn667,n234);
and (s0n667,notn667,n668);
and (s1n667,n234,n669);
wire s0n668,s1n668,notn668;
or (n668,s0n668,s1n668);
not(notn668,n21);
and (s0n668,notn668,1'b0);
and (s1n668,n21,n208);
xor (n669,n207,n209);
and (n670,n652,n671);
not (n671,n667);
and (n672,n595,n601);
or (n673,n674,n727);
and (n674,n675,n710);
xor (n675,n676,n701);
nand (n676,n677,n697);
or (n677,n678,n690);
nand (n678,n679,n686);
nor (n679,n680,n684);
and (n680,n681,n428);
wire s0n681,s1n681,notn681;
or (n681,s0n681,s1n681);
not(notn681,n119);
and (s0n681,notn681,n682);
and (s1n681,n119,n683);
wire s0n682,s1n682,notn682;
or (n682,s0n682,s1n682);
not(notn682,n21);
and (s0n682,notn682,1'b0);
and (s1n682,n21,n95);
xor (n683,n94,n96);
and (n684,n685,n433);
not (n685,n681);
not (n686,n687);
nor (n687,n688,n689);
and (n688,n265,n681);
and (n689,n269,n685);
nor (n690,n691,n695);
and (n691,n433,n692);
wire s0n692,s1n692,notn692;
or (n692,s0n692,s1n692);
not(notn692,n234);
and (s0n692,notn692,n693);
and (s1n692,n234,n694);
wire s0n693,s1n693,notn693;
or (n693,s0n693,s1n693);
not(notn693,n21);
and (s0n693,notn693,1'b0);
and (s1n693,n21,n187);
xor (n694,n186,n188);
and (n695,n428,n696);
not (n696,n692);
or (n697,n698,n686);
nor (n698,n699,n700);
and (n699,n443,n433);
and (n700,n447,n428);
nand (n701,n702,n706);
or (n702,n703,n406);
nor (n703,n704,n705);
and (n704,n480,n138);
and (n705,n484,n139);
or (n706,n707,n407);
nor (n707,n708,n709);
and (n708,n156,n138);
and (n709,n237,n139);
nand (n710,n711,n719);
or (n711,n422,n712);
nor (n712,n713,n717);
and (n713,n440,n714);
wire s0n714,s1n714,notn714;
or (n714,s0n714,s1n714);
not(notn714,n234);
and (s0n714,notn714,n715);
and (s1n714,n234,n716);
wire s0n715,s1n715,notn715;
or (n715,s0n715,s1n715);
not(notn715,n21);
and (s0n715,notn715,1'b0);
and (s1n715,n21,n193);
xor (n716,n192,n194);
and (n717,n436,n718);
not (n718,n714);
or (n719,n423,n720);
nor (n720,n721,n725);
and (n721,n440,n722);
wire s0n722,s1n722,notn722;
or (n722,s0n722,s1n722);
not(notn722,n234);
and (s0n722,notn722,n723);
and (s1n722,n234,n724);
wire s0n723,s1n723,notn723;
or (n723,s0n723,s1n723);
not(notn723,n21);
and (s0n723,notn723,1'b0);
and (s1n723,n21,n190);
xor (n724,n189,n191);
and (n725,n436,n726);
not (n726,n722);
and (n727,n676,n701);
or (n728,n729,n752);
and (n729,n730,n746);
xor (n730,n731,n740);
nand (n731,n732,n736);
or (n732,n290,n733);
nor (n733,n734,n735);
and (n734,n308,n344);
and (n735,n304,n348);
or (n736,n291,n737);
nor (n737,n738,n739);
and (n738,n308,n352);
and (n739,n356,n304);
nand (n740,n741,n745);
or (n741,n326,n742);
nor (n742,n743,n744);
and (n743,n378,n337);
and (n744,n382,n338);
or (n745,n328,n494);
nand (n746,n747,n751);
or (n747,n359,n748);
nor (n748,n749,n750);
and (n749,n367,n130);
and (n750,n366,n131);
or (n751,n373,n500);
and (n752,n731,n740);
and (n753,n592,n673);
or (n754,n755,n841);
and (n755,n756,n840);
xor (n756,n757,n820);
or (n757,n758,n819);
and (n758,n759,n798);
xor (n759,n760,n769);
nand (n760,n761,n765);
or (n761,n458,n762);
nor (n762,n763,n764);
and (n763,n579,n261);
and (n764,n583,n254);
or (n765,n766,n459);
nor (n766,n767,n768);
and (n767,n272,n261);
and (n768,n276,n254);
nand (n769,n770,n789);
or (n770,n771,n782);
or (n771,n772,n779);
nor (n772,n773,n777);
and (n773,n607,n774);
wire s0n774,s1n774,notn774;
or (n774,s0n774,s1n774);
not(notn774,n119);
and (s0n774,notn774,n775);
and (s1n774,n119,n776);
wire s0n775,s1n775,notn775;
or (n775,s0n775,s1n775);
not(notn775,n21);
and (s0n775,notn775,1'b0);
and (s1n775,n21,n83);
xor (n776,n82,n84);
and (n777,n778,n608);
not (n778,n774);
nor (n779,n780,n781);
and (n780,n774,n436);
and (n781,n778,n440);
nor (n782,n783,n787);
and (n783,n607,n784);
wire s0n784,s1n784,notn784;
or (n784,s0n784,s1n784);
not(notn784,n234);
and (s0n784,notn784,n785);
and (s1n784,n234,n786);
wire s0n785,s1n785,notn785;
or (n785,s0n785,s1n785);
not(notn785,n21);
and (s0n785,notn785,1'b0);
and (s1n785,n21,n199);
xor (n786,n198,n200);
and (n787,n608,n788);
not (n788,n784);
or (n789,n790,n791);
not (n790,n779);
nor (n791,n792,n796);
and (n792,n607,n793);
wire s0n793,s1n793,notn793;
or (n793,s0n793,s1n793);
not(notn793,n234);
and (s0n793,notn793,n794);
and (s1n793,n234,n795);
wire s0n794,s1n794,notn794;
or (n794,s0n794,s1n794);
not(notn794,n21);
and (s0n794,notn794,1'b0);
and (s1n794,n21,n196);
xor (n795,n195,n197);
and (n796,n608,n797);
not (n797,n793);
nand (n798,n799,n814);
or (n799,n800,n811);
or (n800,n801,n808);
nor (n801,n802,n806);
and (n802,n803,n652);
wire s0n803,s1n803,notn803;
or (n803,s0n803,s1n803);
not(notn803,n119);
and (s0n803,notn803,n804);
and (s1n803,n119,n805);
wire s0n804,s1n804,notn804;
or (n804,s0n804,s1n804);
not(notn804,n21);
and (s0n804,notn804,1'b0);
and (s1n804,n21,n65);
xor (n805,n64,n66);
and (n806,n807,n656);
not (n807,n803);
nor (n808,n809,n810);
and (n809,n803,n293);
and (n810,n807,n294);
nor (n811,n812,n813);
and (n812,n293,n311);
and (n813,n294,n315);
or (n814,n815,n816);
not (n815,n801);
nor (n816,n817,n818);
and (n817,n293,n319);
and (n818,n294,n323);
and (n819,n760,n769);
xor (n820,n821,n834);
xor (n821,n822,n828);
nand (n822,n823,n824);
or (n823,n707,n406);
or (n824,n825,n407);
nor (n825,n826,n827);
and (n826,n241,n138);
and (n827,n248,n139);
nand (n828,n829,n830);
or (n829,n422,n720);
or (n830,n423,n831);
nor (n831,n832,n833);
and (n832,n440,n692);
and (n833,n436,n696);
nand (n834,n835,n836);
or (n835,n458,n766);
or (n836,n837,n459);
nor (n837,n838,n839);
and (n838,n280,n261);
and (n839,n284,n254);
xor (n840,n562,n567);
and (n841,n757,n820);
xor (n842,n843,n869);
xor (n843,n844,n866);
or (n844,n845,n865);
and (n845,n846,n859);
xor (n846,n847,n853);
nand (n847,n848,n849);
or (n848,n603,n632);
or (n849,n631,n850);
nor (n850,n851,n852);
and (n851,n617,n784);
and (n852,n618,n788);
nand (n853,n854,n855);
or (n854,n641,n665);
or (n855,n643,n856);
nor (n856,n857,n858);
and (n857,n656,n625);
and (n858,n652,n629);
nand (n859,n860,n861);
or (n860,n678,n698);
or (n861,n862,n686);
nor (n862,n863,n864);
and (n863,n451,n433);
and (n864,n455,n428);
and (n865,n847,n853);
or (n866,n867,n868);
and (n867,n821,n834);
and (n868,n822,n828);
xor (n869,n870,n880);
xor (n870,n871,n877);
nand (n871,n872,n873);
or (n872,n678,n862);
or (n873,n874,n686);
nor (n874,n875,n876);
and (n875,n571,n433);
and (n876,n575,n428);
nand (n877,n878,n879);
or (n878,n825,n406);
or (n879,n396,n407);
nand (n880,n881,n882);
or (n881,n422,n831);
or (n882,n423,n441);
and (n883,n589,n754);
xor (n884,n885,n1027);
xor (n885,n886,n942);
xor (n886,n887,n917);
xor (n887,n888,n914);
xor (n888,n889,n908);
xor (n889,n890,n899);
nand (n890,n891,n895);
or (n891,n771,n892);
nor (n892,n893,n894);
and (n893,n607,n722);
and (n894,n608,n726);
or (n895,n790,n896);
nor (n896,n897,n898);
and (n897,n607,n692);
and (n898,n608,n696);
nand (n899,n900,n904);
or (n900,n800,n901);
nor (n901,n902,n903);
and (n902,n293,n667);
and (n903,n294,n671);
or (n904,n815,n905);
nor (n905,n906,n907);
and (n906,n293,n625);
and (n907,n294,n629);
nand (n908,n909,n910);
or (n909,n290,n317);
or (n910,n291,n911);
nor (n911,n912,n913);
and (n912,n308,n659);
and (n913,n663,n304);
or (n914,n915,n916);
and (n915,n526,n560);
and (n916,n527,n547);
xor (n917,n918,n939);
xor (n918,n919,n920);
and (n919,n548,n554);
or (n920,n921,n938);
and (n921,n922,n932);
xor (n922,n923,n926);
nand (n923,n924,n925);
or (n924,n251,n577);
or (n925,n270,n252);
nand (n926,n927,n928);
or (n927,n603,n850);
or (n928,n631,n929);
nor (n929,n930,n931);
and (n930,n617,n793);
and (n931,n618,n797);
nand (n932,n933,n934);
or (n933,n641,n856);
or (n934,n643,n935);
nor (n935,n936,n937);
and (n936,n656,n634);
and (n937,n652,n638);
and (n938,n923,n926);
or (n939,n940,n941);
and (n940,n870,n880);
and (n941,n871,n877);
xor (n942,n943,n982);
xor (n943,n944,n947);
or (n944,n945,n946);
and (n945,n843,n869);
and (n946,n844,n866);
or (n947,n948,n981);
and (n948,n949,n968);
xor (n949,n950,n967);
xor (n950,n951,n961);
xor (n951,n952,n955);
nand (n952,n953,n954);
or (n953,n458,n837);
or (n954,n470,n459);
nand (n955,n956,n960);
or (n956,n771,n957);
nor (n957,n958,n959);
and (n958,n607,n714);
and (n959,n608,n718);
or (n960,n790,n892);
nand (n961,n962,n966);
or (n962,n800,n963);
nor (n963,n964,n965);
and (n964,n293,n659);
and (n965,n294,n663);
or (n966,n815,n901);
xor (n967,n922,n932);
or (n968,n969,n980);
and (n969,n970,n977);
xor (n970,n971,n974);
nand (n971,n972,n973);
or (n972,n771,n791);
or (n973,n790,n957);
nand (n974,n975,n976);
or (n975,n800,n816);
or (n976,n815,n963);
nand (n977,n978,n979);
or (n978,n290,n737);
or (n979,n291,n309);
and (n980,n971,n974);
and (n981,n950,n967);
xor (n982,n983,n1007);
xor (n983,n984,n987);
or (n984,n985,n986);
and (n985,n951,n961);
and (n986,n952,n955);
xor (n987,n988,n1001);
xor (n988,n989,n995);
nand (n989,n990,n991);
or (n990,n603,n929);
or (n991,n631,n992);
nor (n992,n993,n994);
and (n993,n617,n714);
and (n994,n618,n718);
nand (n995,n996,n997);
or (n996,n641,n935);
or (n997,n643,n998);
nor (n998,n999,n1000);
and (n999,n656,n784);
and (n1000,n652,n788);
nand (n1001,n1002,n1003);
or (n1002,n678,n874);
or (n1003,n1004,n686);
nor (n1004,n1005,n1006);
and (n1005,n433,n579);
and (n1006,n583,n428);
xor (n1007,n1008,n1021);
xor (n1008,n1009,n1015);
nand (n1009,n1010,n1011);
or (n1010,n326,n350);
or (n1011,n328,n1012);
nor (n1012,n1013,n1014);
and (n1013,n337,n311);
and (n1014,n315,n338);
nand (n1015,n1016,n1017);
or (n1016,n359,n384);
or (n1017,n373,n1018);
nor (n1018,n1019,n1020);
and (n1019,n366,n344);
and (n1020,n348,n367);
nand (n1021,n1022,n1023);
or (n1022,n529,n544);
or (n1023,n530,n1024);
nor (n1024,n1025,n1026);
and (n1025,n378,n16);
and (n1026,n382,n17);
or (n1027,n1028,n1039);
and (n1028,n1029,n1038);
xor (n1029,n1030,n1037);
or (n1030,n1031,n1036);
and (n1031,n1032,n1035);
xor (n1032,n1033,n1034);
xor (n1033,n846,n859);
xor (n1034,n491,n508);
xor (n1035,n970,n977);
and (n1036,n1033,n1034);
xor (n1037,n949,n968);
xor (n1038,n487,n525);
and (n1039,n1030,n1037);
or (n1040,n1041,n1155);
and (n1041,n1042,n1142);
xor (n1042,n1043,n1141);
or (n1043,n1044,n1140);
and (n1044,n1045,n1096);
xor (n1045,n1046,n1095);
or (n1046,n1047,n1094);
and (n1047,n1048,n1072);
xor (n1048,n1049,n1050);
xor (n1049,n509,n515);
or (n1050,n1051,n1071);
and (n1051,n1052,n1065);
xor (n1052,n1053,n1059);
nand (n1053,n1054,n1058);
or (n1054,n603,n1055);
nor (n1055,n1056,n1057);
and (n1056,n617,n667);
and (n1057,n618,n671);
or (n1058,n631,n623);
nand (n1059,n1060,n1064);
or (n1060,n641,n1061);
nor (n1061,n1062,n1063);
and (n1062,n656,n319);
and (n1063,n652,n323);
or (n1064,n657,n643);
nand (n1065,n1066,n1070);
or (n1066,n678,n1067);
nor (n1067,n1068,n1069);
and (n1068,n433,n722);
and (n1069,n428,n726);
or (n1070,n690,n686);
and (n1071,n1053,n1059);
or (n1072,n1073,n1093);
and (n1073,n1074,n1087);
xor (n1074,n1075,n1081);
nand (n1075,n1076,n1080);
or (n1076,n1077,n406);
nor (n1077,n1078,n1079);
and (n1078,n472,n138);
and (n1079,n476,n139);
or (n1080,n703,n407);
nand (n1081,n1082,n1086);
or (n1082,n458,n1083);
nor (n1083,n1084,n1085);
and (n1084,n571,n261);
and (n1085,n575,n254);
or (n1086,n459,n762);
nand (n1087,n1088,n1092);
or (n1088,n422,n1089);
nor (n1089,n1090,n1091);
and (n1090,n440,n793);
and (n1091,n436,n797);
or (n1092,n423,n712);
and (n1093,n1075,n1081);
and (n1094,n1049,n1050);
xor (n1095,n591,n728);
or (n1096,n1097,n1139);
and (n1097,n1098,n1138);
xor (n1098,n1099,n1116);
or (n1099,n1100,n1115);
and (n1100,n1101,n1109);
xor (n1101,n1102,n1103);
nor (n1102,n373,n130);
nand (n1103,n1104,n1108);
or (n1104,n135,n1105);
nor (n1105,n1106,n1107);
and (n1106,n272,n149);
and (n1107,n276,n150);
or (n1108,n136,n517);
nand (n1109,n1110,n1114);
or (n1110,n251,n1111);
nor (n1111,n1112,n1113);
and (n1112,n443,n269);
and (n1113,n447,n265);
or (n1114,n597,n252);
and (n1115,n1102,n1103);
or (n1116,n1117,n1137);
and (n1117,n1118,n1131);
xor (n1118,n1119,n1125);
nand (n1119,n1120,n1124);
or (n1120,n771,n1121);
nor (n1121,n1122,n1123);
and (n1122,n607,n634);
and (n1123,n608,n638);
or (n1124,n790,n782);
nand (n1125,n1126,n1130);
or (n1126,n800,n1127);
nor (n1127,n1128,n1129);
and (n1128,n352,n293);
and (n1129,n356,n294);
or (n1130,n815,n811);
nand (n1131,n1132,n1136);
or (n1132,n290,n1133);
nor (n1133,n1134,n1135);
and (n1134,n386,n308);
and (n1135,n390,n304);
or (n1136,n291,n733);
and (n1137,n1119,n1125);
xor (n1138,n675,n710);
and (n1139,n1099,n1116);
and (n1140,n1046,n1095);
xor (n1141,n588,n842);
or (n1142,n1143,n1154);
and (n1143,n1144,n1153);
xor (n1144,n1145,n1146);
xor (n1145,n756,n840);
or (n1146,n1147,n1152);
and (n1147,n1148,n1151);
xor (n1148,n1149,n1150);
xor (n1149,n594,n639);
xor (n1150,n759,n798);
xor (n1151,n730,n746);
and (n1152,n1149,n1150);
xor (n1153,n1032,n1035);
and (n1154,n1145,n1146);
and (n1155,n1043,n1141);
or (n1156,n1157,n1278);
and (n1157,n1158,n1277);
xor (n1158,n1159,n1160);
xor (n1159,n1029,n1038);
or (n1160,n1161,n1276);
and (n1161,n1162,n1275);
xor (n1162,n1163,n1262);
or (n1163,n1164,n1261);
and (n1164,n1165,n1260);
xor (n1165,n1166,n1211);
or (n1166,n1167,n1210);
and (n1167,n1168,n1188);
xor (n1168,n1169,n1175);
nand (n1169,n1170,n1174);
or (n1170,n326,n1171);
nor (n1171,n1172,n1173);
and (n1172,n502,n337);
and (n1173,n506,n338);
or (n1174,n328,n742);
and (n1175,n1176,n1182);
nor (n1176,n1177,n337);
nor (n1177,n1178,n1181);
and (n1178,n1179,n308);
not (n1179,n1180);
and (n1180,n131,n331);
and (n1181,n330,n130);
nand (n1182,n1183,n1187);
or (n1183,n135,n1184);
nor (n1184,n1185,n1186);
and (n1185,n579,n149);
and (n1186,n583,n150);
or (n1187,n1105,n136);
or (n1188,n1189,n1209);
and (n1189,n1190,n1203);
xor (n1190,n1191,n1197);
nand (n1191,n1192,n1196);
or (n1192,n678,n1193);
nor (n1193,n1194,n1195);
and (n1194,n433,n714);
and (n1195,n428,n718);
or (n1196,n1067,n686);
nand (n1197,n1198,n1202);
or (n1198,n1199,n406);
nor (n1199,n1200,n1201);
and (n1200,n280,n138);
and (n1201,n284,n139);
or (n1202,n1077,n407);
nand (n1203,n1204,n1208);
or (n1204,n458,n1205);
nor (n1205,n1206,n1207);
and (n1206,n451,n261);
and (n1207,n455,n254);
or (n1208,n1083,n459);
and (n1209,n1191,n1197);
and (n1210,n1169,n1175);
or (n1211,n1212,n1259);
and (n1212,n1213,n1258);
xor (n1213,n1214,n1236);
or (n1214,n1215,n1235);
and (n1215,n1216,n1229);
xor (n1216,n1217,n1223);
nand (n1217,n1218,n1222);
or (n1218,n251,n1219);
nor (n1219,n1220,n1221);
and (n1220,n692,n269);
and (n1221,n696,n265);
or (n1222,n1111,n252);
nand (n1223,n1224,n1228);
or (n1224,n603,n1225);
nor (n1225,n1226,n1227);
and (n1226,n617,n659);
and (n1227,n618,n663);
or (n1228,n631,n1055);
nand (n1229,n1230,n1234);
or (n1230,n641,n1231);
nor (n1231,n1232,n1233);
and (n1232,n656,n311);
and (n1233,n652,n315);
or (n1234,n1061,n643);
and (n1235,n1217,n1223);
or (n1236,n1237,n1257);
and (n1237,n1238,n1251);
xor (n1238,n1239,n1245);
nand (n1239,n1240,n1244);
or (n1240,n422,n1241);
nor (n1241,n1242,n1243);
and (n1242,n440,n784);
and (n1243,n436,n788);
or (n1244,n423,n1089);
nand (n1245,n1246,n1250);
or (n1246,n771,n1247);
nor (n1247,n1248,n1249);
and (n1248,n607,n625);
and (n1249,n608,n629);
or (n1250,n790,n1121);
nand (n1251,n1252,n1256);
or (n1252,n800,n1253);
nor (n1253,n1254,n1255);
and (n1254,n293,n344);
and (n1255,n294,n348);
or (n1256,n815,n1127);
and (n1257,n1239,n1245);
xor (n1258,n1074,n1087);
and (n1259,n1214,n1236);
xor (n1260,n1048,n1072);
and (n1261,n1166,n1211);
or (n1262,n1263,n1274);
and (n1263,n1264,n1273);
xor (n1264,n1265,n1272);
or (n1265,n1266,n1271);
and (n1266,n1267,n1270);
xor (n1267,n1268,n1269);
xor (n1268,n1101,n1109);
xor (n1269,n1052,n1065);
xor (n1270,n1118,n1131);
and (n1271,n1268,n1269);
xor (n1272,n1148,n1151);
xor (n1273,n1098,n1138);
and (n1274,n1265,n1272);
xor (n1275,n1045,n1096);
and (n1276,n1163,n1262);
xor (n1277,n1042,n1142);
and (n1278,n1159,n1160);
nor (n1279,n5,n1156);
not (n1280,n1281);
nor (n1281,n1282,n2893);
and (n1282,n1283,n2886);
or (n1283,n1284,n2885);
and (n1284,n1285,n1528);
xor (n1285,n1286,n1521);
or (n1286,n1287,n1520);
and (n1287,n1288,n1505);
xor (n1288,n1289,n1290);
xor (n1289,n1264,n1273);
or (n1290,n1291,n1504);
and (n1291,n1292,n1445);
xor (n1292,n1293,n1395);
or (n1293,n1294,n1394);
and (n1294,n1295,n1312);
xor (n1295,n1296,n1297);
xor (n1296,n1216,n1229);
xor (n1297,n1298,n1311);
xor (n1298,n1299,n1305);
nand (n1299,n1300,n1304);
or (n1300,n290,n1301);
nor (n1301,n1302,n1303);
and (n1302,n378,n308);
and (n1303,n382,n304);
or (n1304,n291,n1133);
nand (n1305,n1306,n1310);
or (n1306,n326,n1307);
nor (n1307,n1308,n1309);
and (n1308,n338,n130);
and (n1309,n337,n131);
or (n1310,n328,n1171);
xor (n1311,n1176,n1182);
or (n1312,n1313,n1393);
and (n1313,n1314,n1362);
xor (n1314,n1315,n1331);
and (n1315,n1316,n1322);
nor (n1316,n1317,n308);
nor (n1317,n1318,n1321);
and (n1318,n1319,n293);
not (n1319,n1320);
and (n1320,n131,n297);
and (n1321,n301,n130);
nand (n1322,n1323,n1327);
or (n1323,n135,n1324);
nor (n1324,n1325,n1326);
and (n1325,n451,n149);
and (n1326,n455,n150);
or (n1327,n136,n1328);
nor (n1328,n1329,n1330);
and (n1329,n571,n149);
and (n1330,n575,n150);
or (n1331,n1332,n1361);
and (n1332,n1333,n1352);
xor (n1333,n1334,n1343);
nand (n1334,n1335,n1339);
or (n1335,n678,n1336);
nor (n1336,n1337,n1338);
and (n1337,n433,n784);
and (n1338,n428,n788);
or (n1339,n1340,n686);
nor (n1340,n1341,n1342);
and (n1341,n433,n793);
and (n1342,n428,n797);
nand (n1343,n1344,n1348);
or (n1344,n1345,n406);
nor (n1345,n1346,n1347);
and (n1346,n579,n138);
and (n1347,n583,n139);
or (n1348,n1349,n407);
nor (n1349,n1350,n1351);
and (n1350,n272,n138);
and (n1351,n276,n139);
nand (n1352,n1353,n1357);
or (n1353,n458,n1354);
nor (n1354,n1355,n1356);
and (n1355,n692,n261);
and (n1356,n696,n254);
or (n1357,n1358,n459);
nor (n1358,n1359,n1360);
and (n1359,n443,n261);
and (n1360,n447,n254);
and (n1361,n1334,n1343);
or (n1362,n1363,n1392);
and (n1363,n1364,n1383);
xor (n1364,n1365,n1374);
nand (n1365,n1366,n1370);
or (n1366,n251,n1367);
nor (n1367,n1368,n1369);
and (n1368,n714,n269);
and (n1369,n718,n265);
or (n1370,n252,n1371);
nor (n1371,n1372,n1373);
and (n1372,n722,n269);
and (n1373,n726,n265);
nand (n1374,n1375,n1379);
or (n1375,n603,n1376);
nor (n1376,n1377,n1378);
and (n1377,n617,n311);
and (n1378,n618,n315);
or (n1379,n1380,n631);
nor (n1380,n1381,n1382);
and (n1381,n617,n319);
and (n1382,n618,n323);
nand (n1383,n1384,n1388);
or (n1384,n641,n1385);
nor (n1385,n1386,n1387);
and (n1386,n656,n344);
and (n1387,n652,n348);
or (n1388,n1389,n643);
nor (n1389,n1390,n1391);
and (n1390,n656,n352);
and (n1391,n652,n356);
and (n1392,n1365,n1374);
and (n1393,n1315,n1331);
and (n1394,n1296,n1297);
xor (n1395,n1396,n1401);
xor (n1396,n1397,n1400);
or (n1397,n1398,n1399);
and (n1398,n1298,n1311);
and (n1399,n1299,n1305);
xor (n1400,n1168,n1188);
or (n1401,n1402,n1444);
and (n1402,n1403,n1431);
xor (n1403,n1404,n1420);
or (n1404,n1405,n1419);
and (n1405,n1406,n1413);
xor (n1406,n1407,n1410);
nand (n1407,n1408,n1409);
or (n1408,n1349,n406);
or (n1409,n1199,n407);
nand (n1410,n1411,n1412);
or (n1411,n458,n1358);
or (n1412,n1205,n459);
nand (n1413,n1414,n1418);
or (n1414,n422,n1415);
nor (n1415,n1416,n1417);
and (n1416,n440,n634);
and (n1417,n436,n638);
or (n1418,n423,n1241);
and (n1419,n1407,n1410);
or (n1420,n1421,n1430);
and (n1421,n1422,n1427);
xor (n1422,n1423,n1424);
nor (n1423,n328,n130);
nand (n1424,n1425,n1426);
or (n1425,n135,n1328);
or (n1426,n136,n1184);
nand (n1427,n1428,n1429);
or (n1428,n251,n1371);
or (n1429,n252,n1219);
and (n1430,n1423,n1424);
or (n1431,n1432,n1443);
and (n1432,n1433,n1440);
xor (n1433,n1434,n1437);
nand (n1434,n1435,n1436);
or (n1435,n603,n1380);
or (n1436,n631,n1225);
nand (n1437,n1438,n1439);
or (n1438,n641,n1389);
or (n1439,n1231,n643);
nand (n1440,n1441,n1442);
or (n1441,n678,n1340);
or (n1442,n1193,n686);
and (n1443,n1434,n1437);
and (n1444,n1404,n1420);
or (n1445,n1446,n1503);
and (n1446,n1447,n1483);
xor (n1447,n1448,n1482);
or (n1448,n1449,n1481);
and (n1449,n1450,n1480);
xor (n1450,n1451,n1479);
or (n1451,n1452,n1478);
and (n1452,n1453,n1469);
xor (n1453,n1454,n1460);
nand (n1454,n1455,n1459);
or (n1455,n422,n1456);
nor (n1456,n1457,n1458);
and (n1457,n440,n625);
and (n1458,n436,n629);
or (n1459,n423,n1415);
nand (n1460,n1461,n1465);
or (n1461,n771,n1462);
nor (n1462,n1463,n1464);
and (n1463,n607,n659);
and (n1464,n608,n663);
or (n1465,n790,n1466);
nor (n1466,n1467,n1468);
and (n1467,n607,n667);
and (n1468,n608,n671);
nand (n1469,n1470,n1474);
or (n1470,n800,n1471);
nor (n1471,n1472,n1473);
and (n1472,n378,n293);
and (n1473,n382,n294);
or (n1474,n815,n1475);
nor (n1475,n1476,n1477);
and (n1476,n386,n293);
and (n1477,n390,n294);
and (n1478,n1454,n1460);
xor (n1479,n1406,n1413);
xor (n1480,n1433,n1440);
and (n1481,n1451,n1479);
xor (n1482,n1403,n1431);
xor (n1483,n1484,n1487);
xor (n1484,n1485,n1486);
xor (n1485,n1238,n1251);
xor (n1486,n1190,n1203);
or (n1487,n1488,n1502);
and (n1488,n1489,n1496);
xor (n1489,n1490,n1493);
nand (n1490,n1491,n1492);
or (n1491,n771,n1466);
or (n1492,n790,n1247);
nand (n1493,n1494,n1495);
or (n1494,n800,n1475);
or (n1495,n815,n1253);
nand (n1496,n1497,n1501);
or (n1497,n290,n1498);
nor (n1498,n1499,n1500);
and (n1499,n502,n308);
and (n1500,n506,n304);
or (n1501,n291,n1301);
and (n1502,n1490,n1493);
and (n1503,n1448,n1482);
and (n1504,n1293,n1395);
xor (n1505,n1506,n1511);
xor (n1506,n1507,n1510);
or (n1507,n1508,n1509);
and (n1508,n1396,n1401);
and (n1509,n1397,n1400);
xor (n1510,n1165,n1260);
or (n1511,n1512,n1519);
and (n1512,n1513,n1518);
xor (n1513,n1514,n1517);
or (n1514,n1515,n1516);
and (n1515,n1484,n1487);
and (n1516,n1485,n1486);
xor (n1517,n1267,n1270);
xor (n1518,n1213,n1258);
and (n1519,n1514,n1517);
and (n1520,n1289,n1290);
xor (n1521,n1522,n1527);
xor (n1522,n1523,n1524);
xor (n1523,n1144,n1153);
or (n1524,n1525,n1526);
and (n1525,n1506,n1511);
and (n1526,n1507,n1510);
xor (n1527,n1162,n1275);
nand (n1528,n1529,n2879);
or (n1529,n1530,n2861,n2874);
nor (n1530,n1531,n2860);
and (n1531,n1532,n2839);
or (n1532,n1533,n2838);
and (n1533,n1534,n1888);
xor (n1534,n1535,n1861);
or (n1535,n1536,n1860);
and (n1536,n1537,n1775);
xor (n1537,n1538,n1662);
xor (n1538,n1539,n1632);
xor (n1539,n1540,n1571);
xor (n1540,n1541,n1549);
xor (n1541,n1542,n1548);
nand (n1542,n1543,n1547);
or (n1543,n290,n1544);
nor (n1544,n1545,n1546);
and (n1545,n304,n130);
and (n1546,n308,n131);
or (n1547,n291,n1498);
xor (n1548,n1316,n1322);
or (n1549,n1550,n1570);
and (n1550,n1551,n1564);
xor (n1551,n1552,n1558);
nand (n1552,n1553,n1557);
or (n1553,n678,n1554);
nor (n1554,n1555,n1556);
and (n1555,n433,n634);
and (n1556,n428,n638);
or (n1557,n1336,n686);
nand (n1558,n1559,n1563);
or (n1559,n458,n1560);
nor (n1560,n1561,n1562);
and (n1561,n722,n261);
and (n1562,n726,n254);
or (n1563,n459,n1354);
nand (n1564,n1565,n1569);
or (n1565,n422,n1566);
nor (n1566,n1567,n1568);
and (n1567,n440,n667);
and (n1568,n436,n671);
or (n1569,n423,n1456);
and (n1570,n1552,n1558);
or (n1571,n1572,n1631);
and (n1572,n1573,n1630);
xor (n1573,n1574,n1605);
or (n1574,n1575,n1604);
and (n1575,n1576,n1595);
xor (n1576,n1577,n1586);
nand (n1577,n1578,n1582);
or (n1578,n251,n1579);
nor (n1579,n1580,n1581);
and (n1580,n784,n269);
and (n1581,n788,n265);
or (n1582,n252,n1583);
nor (n1583,n1584,n1585);
and (n1584,n793,n269);
and (n1585,n797,n265);
nand (n1586,n1587,n1591);
or (n1587,n603,n1588);
nor (n1588,n1589,n1590);
and (n1589,n617,n344);
and (n1590,n348,n618);
or (n1591,n631,n1592);
nor (n1592,n1593,n1594);
and (n1593,n352,n617);
and (n1594,n356,n618);
nand (n1595,n1596,n1600);
or (n1596,n641,n1597);
nor (n1597,n1598,n1599);
and (n1598,n378,n656);
and (n1599,n382,n652);
or (n1600,n1601,n643);
nor (n1601,n1602,n1603);
and (n1602,n386,n656);
and (n1603,n390,n652);
and (n1604,n1577,n1586);
or (n1605,n1606,n1629);
and (n1606,n1607,n1623);
xor (n1607,n1608,n1617);
nand (n1608,n1609,n1613);
or (n1609,n135,n1610);
nor (n1610,n1611,n1612);
and (n1611,n149,n692);
and (n1612,n696,n150);
or (n1613,n1614,n136);
nor (n1614,n1615,n1616);
and (n1615,n443,n149);
and (n1616,n447,n150);
nand (n1617,n1618,n1622);
or (n1618,n678,n1619);
nor (n1619,n1620,n1621);
and (n1620,n433,n625);
and (n1621,n428,n629);
or (n1622,n1554,n686);
nand (n1623,n1624,n1628);
or (n1624,n458,n1625);
nor (n1625,n1626,n1627);
and (n1626,n714,n261);
and (n1627,n718,n254);
or (n1628,n459,n1560);
and (n1629,n1608,n1617);
xor (n1630,n1551,n1564);
and (n1631,n1574,n1605);
xor (n1632,n1633,n1661);
xor (n1633,n1634,n1648);
or (n1634,n1635,n1647);
and (n1635,n1636,n1644);
xor (n1636,n1637,n1638);
nor (n1637,n291,n130);
nand (n1638,n1639,n1643);
or (n1639,n1640,n406);
nor (n1640,n1641,n1642);
and (n1641,n571,n138);
and (n1642,n575,n139);
or (n1643,n1345,n407);
nand (n1644,n1645,n1646);
or (n1645,n251,n1583);
or (n1646,n252,n1367);
and (n1647,n1637,n1638);
or (n1648,n1649,n1660);
and (n1649,n1650,n1657);
xor (n1650,n1651,n1654);
nand (n1651,n1652,n1653);
or (n1652,n603,n1592);
or (n1653,n1376,n631);
nand (n1654,n1655,n1656);
or (n1655,n641,n1601);
or (n1656,n1385,n643);
nand (n1657,n1658,n1659);
or (n1658,n135,n1614);
or (n1659,n136,n1324);
and (n1660,n1651,n1654);
xor (n1661,n1333,n1352);
xor (n1662,n1663,n1725);
xor (n1663,n1664,n1698);
or (n1664,n1665,n1697);
and (n1665,n1666,n1669);
xor (n1666,n1667,n1668);
xor (n1667,n1636,n1644);
xor (n1668,n1650,n1657);
or (n1669,n1670,n1696);
and (n1670,n1671,n1687);
xor (n1671,n1672,n1678);
nand (n1672,n1673,n1677);
or (n1673,n422,n1674);
nor (n1674,n1675,n1676);
and (n1675,n440,n659);
and (n1676,n436,n663);
or (n1677,n423,n1566);
nand (n1678,n1679,n1683);
or (n1679,n771,n1680);
nor (n1680,n1681,n1682);
and (n1681,n607,n311);
and (n1682,n608,n315);
or (n1683,n1684,n790);
nor (n1684,n1685,n1686);
and (n1685,n607,n319);
and (n1686,n608,n323);
nand (n1687,n1688,n1692);
or (n1688,n800,n1689);
nor (n1689,n1690,n1691);
and (n1690,n294,n130);
and (n1691,n293,n131);
or (n1692,n815,n1693);
nor (n1693,n1694,n1695);
and (n1694,n502,n293);
and (n1695,n506,n294);
and (n1696,n1672,n1678);
and (n1697,n1667,n1668);
xor (n1698,n1699,n1702);
xor (n1699,n1700,n1701);
xor (n1700,n1364,n1383);
xor (n1701,n1453,n1469);
or (n1702,n1703,n1724);
and (n1703,n1704,n1711);
xor (n1704,n1705,n1708);
nand (n1705,n1706,n1707);
or (n1706,n771,n1684);
or (n1707,n790,n1462);
nand (n1708,n1709,n1710);
or (n1709,n800,n1693);
or (n1710,n815,n1471);
and (n1711,n1712,n1718);
nor (n1712,n1713,n293);
nor (n1713,n1714,n1717);
and (n1714,n1715,n656);
not (n1715,n1716);
and (n1716,n131,n803);
and (n1717,n807,n130);
nand (n1718,n1719,n1723);
or (n1719,n1720,n406);
nor (n1720,n1721,n1722);
and (n1721,n451,n138);
and (n1722,n455,n139);
or (n1723,n1640,n407);
and (n1724,n1705,n1708);
or (n1725,n1726,n1774);
and (n1726,n1727,n1773);
xor (n1727,n1728,n1729);
xor (n1728,n1704,n1711);
or (n1729,n1730,n1772);
and (n1730,n1731,n1750);
xor (n1731,n1732,n1733);
xor (n1732,n1712,n1718);
or (n1733,n1734,n1749);
and (n1734,n1735,n1743);
xor (n1735,n1736,n1737);
nor (n1736,n815,n130);
nand (n1737,n1738,n1742);
or (n1738,n1739,n406);
nor (n1739,n1740,n1741);
and (n1740,n443,n138);
and (n1741,n447,n139);
or (n1742,n1720,n407);
nand (n1743,n1744,n1745);
or (n1744,n1579,n252);
or (n1745,n251,n1746);
nor (n1746,n1747,n1748);
and (n1747,n634,n269);
and (n1748,n638,n265);
and (n1749,n1736,n1737);
or (n1750,n1751,n1771);
and (n1751,n1752,n1765);
xor (n1752,n1753,n1759);
nand (n1753,n1754,n1758);
or (n1754,n603,n1755);
nor (n1755,n1756,n1757);
and (n1756,n386,n617);
and (n1757,n390,n618);
or (n1758,n1588,n631);
nand (n1759,n1760,n1764);
or (n1760,n641,n1761);
nor (n1761,n1762,n1763);
and (n1762,n502,n656);
and (n1763,n506,n652);
or (n1764,n1597,n643);
nand (n1765,n1766,n1770);
or (n1766,n135,n1767);
nor (n1767,n1768,n1769);
and (n1768,n149,n722);
and (n1769,n726,n150);
or (n1770,n136,n1610);
and (n1771,n1753,n1759);
and (n1772,n1732,n1733);
xor (n1773,n1573,n1630);
and (n1774,n1728,n1729);
or (n1775,n1776,n1859);
and (n1776,n1777,n1807);
xor (n1777,n1778,n1806);
or (n1778,n1779,n1805);
and (n1779,n1780,n1804);
xor (n1780,n1781,n1803);
or (n1781,n1782,n1802);
and (n1782,n1783,n1796);
xor (n1783,n1784,n1790);
nand (n1784,n1785,n1789);
or (n1785,n678,n1786);
nor (n1786,n1787,n1788);
and (n1787,n433,n667);
and (n1788,n428,n671);
or (n1789,n1619,n686);
nand (n1790,n1791,n1795);
or (n1791,n458,n1792);
nor (n1792,n1793,n1794);
and (n1793,n793,n261);
and (n1794,n797,n254);
or (n1795,n459,n1625);
nand (n1796,n1797,n1801);
or (n1797,n422,n1798);
nor (n1798,n1799,n1800);
and (n1799,n440,n319);
and (n1800,n436,n323);
or (n1801,n423,n1674);
and (n1802,n1784,n1790);
xor (n1803,n1607,n1623);
xor (n1804,n1576,n1595);
and (n1805,n1781,n1803);
xor (n1806,n1666,n1669);
or (n1807,n1808,n1858);
and (n1808,n1809,n1857);
xor (n1809,n1810,n1811);
xor (n1810,n1671,n1687);
or (n1811,n1812,n1856);
and (n1812,n1813,n1833);
xor (n1813,n1814,n1820);
nand (n1814,n1815,n1819);
or (n1815,n771,n1816);
nor (n1816,n1817,n1818);
and (n1817,n607,n352);
and (n1818,n608,n356);
or (n1819,n1680,n790);
and (n1820,n1821,n1827);
nor (n1821,n1822,n656);
nor (n1822,n1823,n1826);
and (n1823,n617,n1824);
not (n1824,n1825);
and (n1825,n131,n646);
and (n1826,n645,n130);
nand (n1827,n1828,n1832);
or (n1828,n1829,n406);
nor (n1829,n1830,n1831);
and (n1830,n692,n138);
and (n1831,n696,n139);
or (n1832,n1739,n407);
or (n1833,n1834,n1855);
and (n1834,n1835,n1848);
xor (n1835,n1836,n1842);
nand (n1836,n1837,n1841);
or (n1837,n251,n1838);
nor (n1838,n1839,n1840);
and (n1839,n625,n269);
and (n1840,n629,n265);
or (n1841,n1746,n252);
nand (n1842,n1843,n1847);
or (n1843,n603,n1844);
nor (n1844,n1845,n1846);
and (n1845,n378,n617);
and (n1846,n382,n618);
or (n1847,n631,n1755);
nand (n1848,n1849,n1854);
or (n1849,n1850,n641);
not (n1850,n1851);
nand (n1851,n1852,n1853);
or (n1852,n656,n131);
or (n1853,n652,n130);
or (n1854,n1761,n643);
and (n1855,n1836,n1842);
and (n1856,n1814,n1820);
xor (n1857,n1731,n1750);
and (n1858,n1810,n1811);
and (n1859,n1778,n1806);
and (n1860,n1538,n1662);
xor (n1861,n1862,n1885);
xor (n1862,n1863,n1872);
xor (n1863,n1864,n1869);
xor (n1864,n1865,n1866);
xor (n1865,n1314,n1362);
or (n1866,n1867,n1868);
and (n1867,n1633,n1661);
and (n1868,n1634,n1648);
or (n1869,n1870,n1871);
and (n1870,n1699,n1702);
and (n1871,n1700,n1701);
xor (n1872,n1873,n1882);
xor (n1873,n1874,n1875);
xor (n1874,n1450,n1480);
xor (n1875,n1876,n1879);
xor (n1876,n1877,n1878);
xor (n1877,n1422,n1427);
xor (n1878,n1489,n1496);
or (n1879,n1880,n1881);
and (n1880,n1541,n1549);
and (n1881,n1542,n1548);
or (n1882,n1883,n1884);
and (n1883,n1539,n1632);
and (n1884,n1540,n1571);
or (n1885,n1886,n1887);
and (n1886,n1663,n1725);
and (n1887,n1664,n1698);
nand (n1888,n1889,n2832);
or (n1889,n1890,n2825);
nand (n1890,n1891,n2814);
not (n1891,n1892);
nor (n1892,n1893,n2803);
nor (n1893,n1894,n2752);
nand (n1894,n1895,n2626);
or (n1895,n1896,n2625);
and (n1896,n1897,n2215);
xor (n1897,n1898,n2129);
or (n1898,n1899,n2128);
and (n1899,n1900,n2077);
xor (n1900,n1901,n1984);
xor (n1901,n1902,n1953);
xor (n1902,n1903,n1924);
xor (n1903,n1904,n1915);
xor (n1904,n1905,n1906);
nor (n1905,n631,n130);
nand (n1906,n1907,n1911);
or (n1907,n1908,n406);
nor (n1908,n1909,n1910);
and (n1909,n138,n793);
and (n1910,n797,n139);
or (n1911,n1912,n407);
nor (n1912,n1913,n1914);
and (n1913,n714,n138);
and (n1914,n718,n139);
nand (n1915,n1916,n1920);
or (n1916,n135,n1917);
nor (n1917,n1918,n1919);
and (n1918,n149,n634);
and (n1919,n638,n150);
or (n1920,n136,n1921);
nor (n1921,n1922,n1923);
and (n1922,n784,n149);
and (n1923,n788,n150);
or (n1924,n1925,n1952);
and (n1925,n1926,n1942);
xor (n1926,n1927,n1933);
nand (n1927,n1928,n1932);
or (n1928,n135,n1929);
nor (n1929,n1930,n1931);
and (n1930,n149,n625);
and (n1931,n629,n150);
or (n1932,n136,n1917);
nand (n1933,n1934,n1938);
or (n1934,n251,n1935);
nor (n1935,n1936,n1937);
and (n1936,n311,n269);
and (n1937,n315,n265);
or (n1938,n252,n1939);
nor (n1939,n1940,n1941);
and (n1940,n319,n269);
and (n1941,n323,n265);
nand (n1942,n1943,n1948);
or (n1943,n1944,n678);
not (n1944,n1945);
nand (n1945,n1946,n1947);
or (n1946,n428,n348);
or (n1947,n433,n344);
or (n1948,n1949,n686);
nor (n1949,n1950,n1951);
and (n1950,n433,n352);
and (n1951,n428,n356);
and (n1952,n1927,n1933);
or (n1953,n1954,n1983);
and (n1954,n1955,n1974);
xor (n1955,n1956,n1965);
nand (n1956,n1957,n1961);
or (n1957,n458,n1958);
nor (n1958,n1959,n1960);
and (n1959,n659,n261);
and (n1960,n663,n254);
or (n1961,n1962,n459);
nor (n1962,n1963,n1964);
and (n1963,n667,n261);
and (n1964,n671,n254);
nand (n1965,n1966,n1970);
or (n1966,n422,n1967);
nor (n1967,n1968,n1969);
and (n1968,n378,n440);
and (n1969,n382,n436);
or (n1970,n1971,n423);
nor (n1971,n1972,n1973);
and (n1972,n386,n440);
and (n1973,n390,n436);
nand (n1974,n1975,n1979);
or (n1975,n790,n1976);
nor (n1976,n1977,n1978);
and (n1977,n502,n607);
and (n1978,n506,n608);
or (n1979,n771,n1980);
nor (n1980,n1981,n1982);
and (n1981,n608,n130);
and (n1982,n607,n131);
and (n1983,n1956,n1965);
xor (n1984,n1985,n2033);
xor (n1985,n1986,n2013);
xor (n1986,n1987,n2000);
xor (n1987,n1988,n1994);
nand (n1988,n1989,n1990);
or (n1989,n422,n1971);
or (n1990,n1991,n423);
nor (n1991,n1992,n1993);
and (n1992,n440,n344);
and (n1993,n436,n348);
nand (n1994,n1995,n1996);
or (n1995,n771,n1976);
or (n1996,n1997,n790);
nor (n1997,n1998,n1999);
and (n1998,n378,n607);
and (n1999,n382,n608);
and (n2000,n2001,n2007);
nand (n2001,n2002,n2006);
or (n2002,n2003,n406);
nor (n2003,n2004,n2005);
and (n2004,n138,n784);
and (n2005,n788,n139);
or (n2006,n1908,n407);
nor (n2007,n2008,n607);
nor (n2008,n2009,n2012);
and (n2009,n440,n2010);
not (n2010,n2011);
and (n2011,n131,n774);
and (n2012,n778,n130);
xor (n2013,n2014,n2027);
xor (n2014,n2015,n2021);
nand (n2015,n2016,n2017);
or (n2016,n251,n1939);
or (n2017,n2018,n252);
nor (n2018,n2019,n2020);
and (n2019,n659,n269);
and (n2020,n663,n265);
nand (n2021,n2022,n2023);
or (n2022,n678,n1949);
or (n2023,n2024,n686);
nor (n2024,n2025,n2026);
and (n2025,n433,n311);
and (n2026,n428,n315);
nand (n2027,n2028,n2032);
or (n2028,n459,n2029);
nor (n2029,n2030,n2031);
and (n2030,n625,n261);
and (n2031,n629,n254);
or (n2032,n458,n1962);
or (n2033,n2034,n2076);
and (n2034,n2035,n2054);
xor (n2035,n2036,n2037);
xor (n2036,n2001,n2007);
or (n2037,n2038,n2053);
and (n2038,n2039,n2047);
xor (n2039,n2040,n2041);
nor (n2040,n790,n130);
nand (n2041,n2042,n2046);
or (n2042,n2043,n406);
nor (n2043,n2044,n2045);
and (n2044,n138,n634);
and (n2045,n638,n139);
or (n2046,n2003,n407);
nand (n2047,n2048,n2049);
or (n2048,n136,n1929);
or (n2049,n135,n2050);
nor (n2050,n2051,n2052);
and (n2051,n667,n149);
and (n2052,n671,n150);
and (n2053,n2040,n2041);
or (n2054,n2055,n2075);
and (n2055,n2056,n2069);
xor (n2056,n2057,n2063);
nand (n2057,n2058,n2062);
or (n2058,n251,n2059);
nor (n2059,n2060,n2061);
and (n2060,n352,n269);
and (n2061,n356,n265);
or (n2062,n1935,n252);
nand (n2063,n2064,n2065);
or (n2064,n686,n1944);
or (n2065,n678,n2066);
nor (n2066,n2067,n2068);
and (n2067,n433,n386);
and (n2068,n428,n390);
nand (n2069,n2070,n2071);
or (n2070,n423,n1967);
or (n2071,n422,n2072);
nor (n2072,n2073,n2074);
and (n2073,n502,n440);
and (n2074,n506,n436);
and (n2075,n2057,n2063);
and (n2076,n2036,n2037);
or (n2077,n2078,n2127);
and (n2078,n2079,n2082);
xor (n2079,n2080,n2081);
xor (n2080,n1955,n1974);
xor (n2081,n1926,n1942);
or (n2082,n2083,n2126);
and (n2083,n2084,n2104);
xor (n2084,n2085,n2091);
nand (n2085,n2086,n2090);
or (n2086,n458,n2087);
nor (n2087,n2088,n2089);
and (n2088,n319,n261);
and (n2089,n323,n254);
or (n2090,n459,n1958);
and (n2091,n2092,n2098);
nand (n2092,n2093,n2097);
or (n2093,n2094,n406);
nor (n2094,n2095,n2096);
and (n2095,n625,n138);
and (n2096,n629,n139);
or (n2097,n2043,n407);
nor (n2098,n2099,n440);
nor (n2099,n2100,n2103);
and (n2100,n433,n2101);
not (n2101,n2102);
and (n2102,n131,n425);
and (n2103,n432,n130);
or (n2104,n2105,n2125);
and (n2105,n2106,n2119);
xor (n2106,n2107,n2113);
nand (n2107,n2108,n2112);
or (n2108,n135,n2109);
nor (n2109,n2110,n2111);
and (n2110,n659,n149);
and (n2111,n663,n150);
or (n2112,n136,n2050);
nand (n2113,n2114,n2118);
or (n2114,n251,n2115);
nor (n2115,n2116,n2117);
and (n2116,n344,n269);
and (n2117,n348,n265);
or (n2118,n2059,n252);
nand (n2119,n2120,n2124);
or (n2120,n678,n2121);
nor (n2121,n2122,n2123);
and (n2122,n378,n433);
and (n2123,n382,n428);
or (n2124,n2066,n686);
and (n2125,n2107,n2113);
and (n2126,n2085,n2091);
and (n2127,n2080,n2081);
and (n2128,n1901,n1984);
xor (n2129,n2130,n2163);
xor (n2130,n2131,n2160);
xor (n2131,n2132,n2139);
xor (n2132,n2133,n2136);
or (n2133,n2134,n2135);
and (n2134,n2014,n2027);
and (n2135,n2015,n2021);
or (n2136,n2137,n2138);
and (n2137,n1987,n2000);
and (n2138,n1988,n1994);
xor (n2139,n2140,n2153);
xor (n2140,n2141,n2147);
nand (n2141,n2142,n2143);
or (n2142,n678,n2024);
or (n2143,n2144,n686);
nor (n2144,n2145,n2146);
and (n2145,n433,n319);
and (n2146,n428,n323);
nand (n2147,n2148,n2149);
or (n2148,n458,n2029);
or (n2149,n459,n2150);
nor (n2150,n2151,n2152);
and (n2151,n634,n261);
and (n2152,n638,n254);
nand (n2153,n2154,n2159);
or (n2154,n423,n2155);
not (n2155,n2156);
nand (n2156,n2157,n2158);
or (n2157,n356,n436);
or (n2158,n440,n352);
or (n2159,n422,n1991);
or (n2160,n2161,n2162);
and (n2161,n1985,n2033);
and (n2162,n1986,n2013);
xor (n2163,n2164,n2191);
xor (n2164,n2165,n2188);
xor (n2165,n2166,n2182);
xor (n2166,n2167,n2173);
nand (n2167,n2168,n2169);
or (n2168,n135,n1921);
or (n2169,n136,n2170);
nor (n2170,n2171,n2172);
and (n2171,n149,n793);
and (n2172,n797,n150);
nand (n2173,n2174,n2178);
or (n2174,n603,n2175);
nor (n2175,n2176,n2177);
and (n2176,n618,n130);
and (n2177,n617,n131);
or (n2178,n2179,n631);
nor (n2179,n2180,n2181);
and (n2180,n502,n617);
and (n2181,n506,n618);
nand (n2182,n2183,n2187);
or (n2183,n2184,n252);
nor (n2184,n2185,n2186);
and (n2185,n667,n269);
and (n2186,n671,n265);
or (n2187,n251,n2018);
or (n2188,n2189,n2190);
and (n2189,n1902,n1953);
and (n2190,n1903,n1924);
xor (n2191,n2192,n2212);
xor (n2192,n2193,n2199);
nand (n2193,n2194,n2195);
or (n2194,n771,n1997);
or (n2195,n2196,n790);
nor (n2196,n2197,n2198);
and (n2197,n386,n607);
and (n2198,n390,n608);
xor (n2199,n2200,n2206);
nand (n2200,n2201,n2202);
or (n2201,n1912,n406);
or (n2202,n2203,n407);
nor (n2203,n2204,n2205);
and (n2204,n722,n138);
and (n2205,n726,n139);
nor (n2206,n2207,n617);
nor (n2207,n2208,n2211);
and (n2208,n607,n2209);
not (n2209,n2210);
and (n2210,n131,n611);
and (n2211,n622,n130);
or (n2212,n2213,n2214);
and (n2213,n1904,n1915);
and (n2214,n1905,n1906);
or (n2215,n2216,n2624);
and (n2216,n2217,n2248);
xor (n2217,n2218,n2247);
or (n2218,n2219,n2246);
and (n2219,n2220,n2245);
xor (n2220,n2221,n2244);
or (n2221,n2222,n2243);
and (n2222,n2223,n2226);
xor (n2223,n2224,n2225);
xor (n2224,n2039,n2047);
xor (n2225,n2056,n2069);
or (n2226,n2227,n2242);
and (n2227,n2228,n2241);
xor (n2228,n2229,n2235);
nand (n2229,n2230,n2234);
or (n2230,n422,n2231);
nor (n2231,n2232,n2233);
and (n2232,n436,n130);
and (n2233,n440,n131);
or (n2234,n2072,n423);
nand (n2235,n2236,n2240);
or (n2236,n458,n2237);
nor (n2237,n2238,n2239);
and (n2238,n311,n261);
and (n2239,n315,n254);
or (n2240,n2087,n459);
xor (n2241,n2092,n2098);
and (n2242,n2229,n2235);
and (n2243,n2224,n2225);
xor (n2244,n2035,n2054);
xor (n2245,n2079,n2082);
and (n2246,n2221,n2244);
xor (n2247,n1900,n2077);
nand (n2248,n2249,n2621,n2623);
or (n2249,n2250,n2616);
nand (n2250,n2251,n2605);
or (n2251,n2252,n2604);
and (n2252,n2253,n2374);
xor (n2253,n2254,n2359);
or (n2254,n2255,n2358);
and (n2255,n2256,n2324);
xor (n2256,n2257,n2279);
xor (n2257,n2258,n2273);
xor (n2258,n2259,n2266);
nand (n2259,n2260,n2265);
or (n2260,n251,n2261);
not (n2261,n2262);
nor (n2262,n2263,n2264);
and (n2263,n269,n390);
and (n2264,n386,n265);
or (n2265,n2115,n252);
nand (n2266,n2267,n2272);
or (n2267,n2268,n678);
not (n2268,n2269);
nand (n2269,n2270,n2271);
or (n2270,n506,n428);
or (n2271,n502,n433);
or (n2272,n2121,n686);
nand (n2273,n2274,n2278);
or (n2274,n458,n2275);
nor (n2275,n2276,n2277);
and (n2276,n352,n261);
and (n2277,n356,n254);
or (n2278,n459,n2237);
or (n2279,n2280,n2323);
and (n2280,n2281,n2303);
xor (n2281,n2282,n2288);
nand (n2282,n2283,n2287);
or (n2283,n458,n2284);
nor (n2284,n2285,n2286);
and (n2285,n344,n261);
and (n2286,n348,n254);
or (n2287,n2275,n459);
xor (n2288,n2289,n2295);
nor (n2289,n2290,n433);
nor (n2290,n2291,n2294);
and (n2291,n2292,n269);
not (n2292,n2293);
and (n2293,n131,n681);
and (n2294,n685,n130);
nand (n2295,n2296,n2299);
or (n2296,n406,n2297);
not (n2297,n2298);
xnor (n2298,n659,n138);
or (n2299,n2300,n407);
nor (n2300,n2301,n2302);
and (n2301,n138,n667);
and (n2302,n671,n139);
or (n2303,n2304,n2322);
and (n2304,n2305,n2313);
xor (n2305,n2306,n2307);
nor (n2306,n686,n130);
nand (n2307,n2308,n2309);
or (n2308,n407,n2297);
or (n2309,n2310,n406);
nor (n2310,n2311,n2312);
and (n2311,n138,n319);
and (n2312,n323,n139);
nand (n2313,n2314,n2318);
or (n2314,n251,n2315);
nor (n2315,n2316,n2317);
and (n2316,n502,n269);
and (n2317,n506,n265);
or (n2318,n2319,n252);
nor (n2319,n2320,n2321);
and (n2320,n378,n269);
and (n2321,n382,n265);
and (n2322,n2306,n2307);
and (n2323,n2282,n2288);
xor (n2324,n2325,n2339);
xor (n2325,n2326,n2327);
and (n2326,n2289,n2295);
xor (n2327,n2328,n2333);
xor (n2328,n2329,n2330);
nor (n2329,n423,n130);
nand (n2330,n2331,n2332);
or (n2331,n2300,n406);
or (n2332,n2094,n407);
nand (n2333,n2334,n2338);
or (n2334,n135,n2335);
nor (n2335,n2336,n2337);
and (n2336,n319,n149);
and (n2337,n323,n150);
or (n2338,n136,n2109);
or (n2339,n2340,n2357);
and (n2340,n2341,n2351);
xor (n2341,n2342,n2348);
nand (n2342,n2343,n2347);
or (n2343,n135,n2344);
nor (n2344,n2345,n2346);
and (n2345,n149,n311);
and (n2346,n315,n150);
or (n2347,n2335,n136);
nand (n2348,n2349,n2350);
or (n2349,n252,n2261);
or (n2350,n2319,n251);
nand (n2351,n2352,n2353);
or (n2352,n686,n2268);
or (n2353,n678,n2354);
nor (n2354,n2355,n2356);
and (n2355,n428,n130);
and (n2356,n433,n131);
and (n2357,n2342,n2348);
and (n2358,n2257,n2279);
xor (n2359,n2360,n2365);
xor (n2360,n2361,n2362);
xor (n2361,n2106,n2119);
or (n2362,n2363,n2364);
and (n2363,n2325,n2339);
and (n2364,n2326,n2327);
xor (n2365,n2366,n2373);
xor (n2366,n2367,n2370);
or (n2367,n2368,n2369);
and (n2368,n2328,n2333);
and (n2369,n2329,n2330);
or (n2370,n2371,n2372);
and (n2371,n2258,n2273);
and (n2372,n2259,n2266);
xor (n2373,n2228,n2241);
or (n2374,n2375,n2603);
and (n2375,n2376,n2413);
xor (n2376,n2377,n2412);
or (n2377,n2378,n2411);
and (n2378,n2379,n2410);
xor (n2379,n2380,n2409);
or (n2380,n2381,n2408);
and (n2381,n2382,n2395);
xor (n2382,n2383,n2389);
nand (n2383,n2384,n2388);
or (n2384,n135,n2385);
nor (n2385,n2386,n2387);
and (n2386,n352,n149);
and (n2387,n150,n356);
or (n2388,n2344,n136);
nand (n2389,n2390,n2394);
or (n2390,n458,n2391);
nor (n2391,n2392,n2393);
and (n2392,n386,n261);
and (n2393,n390,n254);
or (n2394,n2284,n459);
and (n2395,n2396,n2402);
nor (n2396,n2397,n269);
nor (n2397,n2398,n2401);
and (n2398,n2399,n261);
not (n2399,n2400);
and (n2400,n131,n257);
and (n2401,n262,n130);
nand (n2402,n2403,n2407);
or (n2403,n2404,n406);
nor (n2404,n2405,n2406);
and (n2405,n138,n311);
and (n2406,n315,n139);
or (n2407,n2310,n407);
and (n2408,n2383,n2389);
xor (n2409,n2341,n2351);
xor (n2410,n2281,n2303);
and (n2411,n2380,n2409);
xor (n2412,n2256,n2324);
nand (n2413,n2414,n2600,n2602);
or (n2414,n2415,n2473);
nand (n2415,n2416,n2468);
not (n2416,n2417);
nor (n2417,n2418,n2444);
xor (n2418,n2419,n2443);
xor (n2419,n2420,n2442);
or (n2420,n2421,n2441);
and (n2421,n2422,n2435);
xor (n2422,n2423,n2429);
nand (n2423,n2424,n2428);
or (n2424,n251,n2425);
nor (n2425,n2426,n2427);
and (n2426,n265,n130);
and (n2427,n269,n131);
or (n2428,n2315,n252);
nand (n2429,n2430,n2434);
or (n2430,n2431,n135);
nor (n2431,n2432,n2433);
and (n2432,n150,n348);
and (n2433,n149,n344);
or (n2434,n2385,n136);
nand (n2435,n2436,n2440);
or (n2436,n458,n2437);
nor (n2437,n2438,n2439);
and (n2438,n378,n261);
and (n2439,n382,n254);
or (n2440,n2391,n459);
and (n2441,n2423,n2429);
xor (n2442,n2305,n2313);
xor (n2443,n2382,n2395);
or (n2444,n2445,n2467);
and (n2445,n2446,n2466);
xor (n2446,n2447,n2448);
xor (n2447,n2396,n2402);
or (n2448,n2449,n2465);
and (n2449,n2450,n2459);
xor (n2450,n2451,n2452);
nor (n2451,n252,n130);
nand (n2452,n2453,n2458);
or (n2453,n2454,n406);
not (n2454,n2455);
nand (n2455,n2456,n2457);
or (n2456,n139,n356);
nand (n2457,n356,n139);
or (n2458,n2404,n407);
nand (n2459,n2460,n2464);
or (n2460,n135,n2461);
nor (n2461,n2462,n2463);
and (n2462,n149,n386);
and (n2463,n150,n390);
or (n2464,n2431,n136);
and (n2465,n2451,n2452);
xor (n2466,n2422,n2435);
and (n2467,n2447,n2448);
or (n2468,n2469,n2470);
xor (n2469,n2379,n2410);
or (n2470,n2471,n2472);
and (n2471,n2419,n2443);
and (n2472,n2420,n2442);
nor (n2473,n2474,n2599);
and (n2474,n2475,n2594);
or (n2475,n2476,n2593);
and (n2476,n2477,n2518);
xor (n2477,n2478,n2511);
or (n2478,n2479,n2510);
and (n2479,n2480,n2496);
xor (n2480,n2481,n2487);
nand (n2481,n2482,n2486);
or (n2482,n135,n2483);
nor (n2483,n2484,n2485);
and (n2484,n150,n382);
and (n2485,n149,n378);
or (n2486,n2461,n136);
or (n2487,n2488,n2492);
nor (n2488,n2489,n459);
nor (n2489,n2490,n2491);
and (n2490,n261,n502);
and (n2491,n254,n506);
nor (n2492,n458,n2493);
nor (n2493,n2494,n2495);
and (n2494,n254,n130);
and (n2495,n261,n131);
xor (n2496,n2497,n2503);
nor (n2497,n2498,n261);
nor (n2498,n2499,n2502);
and (n2499,n2500,n149);
not (n2500,n2501);
and (n2501,n131,n462);
and (n2502,n468,n130);
nand (n2503,n2504,n2509);
or (n2504,n406,n2505);
not (n2505,n2506);
nand (n2506,n2507,n2508);
or (n2507,n138,n344);
nand (n2508,n344,n138);
nand (n2509,n2455,n408);
and (n2510,n2481,n2487);
xor (n2511,n2512,n2517);
xor (n2512,n2513,n2516);
nand (n2513,n2514,n2515);
or (n2514,n458,n2489);
or (n2515,n2437,n459);
and (n2516,n2497,n2503);
xor (n2517,n2450,n2459);
or (n2518,n2519,n2592);
and (n2519,n2520,n2540);
xor (n2520,n2521,n2539);
or (n2521,n2522,n2538);
and (n2522,n2523,n2532);
xor (n2523,n2524,n2525);
and (n2524,n460,n131);
nand (n2525,n2526,n2531);
or (n2526,n406,n2527);
not (n2527,n2528);
nand (n2528,n2529,n2530);
or (n2529,n139,n390);
nand (n2530,n390,n139);
nand (n2531,n2506,n408);
nand (n2532,n2533,n2537);
or (n2533,n135,n2534);
nor (n2534,n2535,n2536);
and (n2535,n149,n502);
and (n2536,n150,n506);
or (n2537,n2483,n136);
and (n2538,n2524,n2525);
xor (n2539,n2480,n2496);
or (n2540,n2541,n2591);
and (n2541,n2542,n2559);
xor (n2542,n2543,n2558);
and (n2543,n2544,n2550);
and (n2544,n2545,n150);
nand (n2545,n2546,n2549);
nand (n2546,n2547,n138);
not (n2547,n2548);
and (n2548,n131,n142);
nand (n2549,n146,n130);
nand (n2550,n2551,n2552);
or (n2551,n407,n2527);
nand (n2552,n2553,n2557);
not (n2553,n2554);
nor (n2554,n2555,n2556);
and (n2555,n382,n139);
and (n2556,n378,n138);
not (n2557,n406);
xor (n2558,n2523,n2532);
or (n2559,n2560,n2590);
and (n2560,n2561,n2569);
xor (n2561,n2562,n2568);
nand (n2562,n2563,n2567);
or (n2563,n135,n2564);
nor (n2564,n2565,n2566);
and (n2565,n150,n130);
and (n2566,n149,n131);
or (n2567,n2534,n136);
xor (n2568,n2544,n2550);
or (n2569,n2570,n2589);
and (n2570,n2571,n2579);
xor (n2571,n2572,n2573);
nor (n2572,n136,n130);
nand (n2573,n2574,n2578);
or (n2574,n2575,n406);
or (n2575,n2576,n2577);
and (n2576,n138,n506);
and (n2577,n502,n139);
or (n2578,n2554,n407);
nor (n2579,n2580,n2587);
nor (n2580,n2581,n2583);
and (n2581,n2582,n408);
not (n2582,n2575);
and (n2583,n2584,n2557);
nand (n2584,n2585,n2586);
or (n2585,n138,n131);
or (n2586,n139,n130);
or (n2587,n138,n2588);
and (n2588,n131,n408);
and (n2589,n2572,n2573);
and (n2590,n2562,n2568);
and (n2591,n2543,n2558);
and (n2592,n2521,n2539);
and (n2593,n2478,n2511);
or (n2594,n2595,n2596);
xor (n2595,n2446,n2466);
or (n2596,n2597,n2598);
and (n2597,n2512,n2517);
and (n2598,n2513,n2516);
and (n2599,n2595,n2596);
nand (n2600,n2468,n2601);
and (n2601,n2418,n2444);
nand (n2602,n2469,n2470);
and (n2603,n2377,n2412);
and (n2604,n2254,n2359);
or (n2605,n2606,n2613);
xor (n2606,n2607,n2612);
xor (n2607,n2608,n2609);
xor (n2608,n2084,n2104);
or (n2609,n2610,n2611);
and (n2610,n2366,n2373);
and (n2611,n2367,n2370);
xor (n2612,n2223,n2226);
or (n2613,n2614,n2615);
and (n2614,n2360,n2365);
and (n2615,n2361,n2362);
nor (n2616,n2617,n2618);
xor (n2617,n2220,n2245);
or (n2618,n2619,n2620);
and (n2619,n2607,n2612);
and (n2620,n2608,n2609);
or (n2621,n2616,n2622);
nand (n2622,n2606,n2613);
nand (n2623,n2617,n2618);
and (n2624,n2218,n2247);
and (n2625,n1898,n2129);
nor (n2626,n2627,n2747);
nor (n2627,n2628,n2738);
xor (n2628,n2629,n2693);
xor (n2629,n2630,n2668);
xor (n2630,n2631,n2653);
xor (n2631,n2632,n2633);
xor (n2632,n1835,n1848);
xor (n2633,n2634,n2647);
xor (n2634,n2635,n2641);
nand (n2635,n2636,n2640);
or (n2636,n135,n2637);
nor (n2637,n2638,n2639);
and (n2638,n149,n714);
and (n2639,n718,n150);
or (n2640,n136,n1767);
nand (n2641,n2642,n2646);
or (n2642,n678,n2643);
nor (n2643,n2644,n2645);
and (n2644,n433,n659);
and (n2645,n428,n663);
or (n2646,n1786,n686);
nand (n2647,n2648,n2652);
or (n2648,n2649,n458);
nor (n2649,n2650,n2651);
and (n2650,n784,n261);
and (n2651,n788,n254);
or (n2652,n459,n1792);
xor (n2653,n2654,n2667);
xor (n2654,n2655,n2661);
nand (n2655,n2656,n2660);
or (n2656,n422,n2657);
nor (n2657,n2658,n2659);
and (n2658,n440,n311);
and (n2659,n436,n315);
or (n2660,n1798,n423);
nand (n2661,n2662,n2666);
or (n2662,n771,n2663);
nor (n2663,n2664,n2665);
and (n2664,n607,n344);
and (n2665,n348,n608);
or (n2666,n790,n1816);
xor (n2667,n1821,n1827);
or (n2668,n2669,n2692);
and (n2669,n2670,n2677);
xor (n2670,n2671,n2674);
or (n2671,n2672,n2673);
and (n2672,n2192,n2212);
and (n2673,n2193,n2199);
or (n2674,n2675,n2676);
and (n2675,n2132,n2139);
and (n2676,n2133,n2136);
xor (n2677,n2678,n2689);
xor (n2678,n2679,n2680);
and (n2679,n2200,n2206);
xor (n2680,n2681,n2686);
xor (n2681,n2682,n2683);
nor (n2682,n643,n130);
nand (n2683,n2684,n2685);
or (n2684,n2203,n406);
or (n2685,n1829,n407);
nand (n2686,n2687,n2688);
or (n2687,n135,n2170);
or (n2688,n136,n2637);
or (n2689,n2690,n2691);
and (n2690,n2166,n2182);
and (n2691,n2167,n2173);
and (n2692,n2671,n2674);
xor (n2693,n2694,n2729);
xor (n2694,n2695,n2698);
or (n2695,n2696,n2697);
and (n2696,n2678,n2689);
and (n2697,n2679,n2680);
xor (n2698,n2699,n2716);
xor (n2699,n2700,n2703);
or (n2700,n2701,n2702);
and (n2701,n2681,n2686);
and (n2702,n2682,n2683);
or (n2703,n2704,n2715);
and (n2704,n2705,n2712);
xor (n2705,n2706,n2709);
nand (n2706,n2707,n2708);
or (n2707,n458,n2150);
or (n2708,n459,n2649);
nand (n2709,n2710,n2711);
or (n2710,n2155,n422);
or (n2711,n2657,n423);
nand (n2712,n2713,n2714);
or (n2713,n771,n2196);
or (n2714,n2663,n790);
and (n2715,n2706,n2709);
or (n2716,n2717,n2728);
and (n2717,n2718,n2725);
xor (n2718,n2719,n2722);
nand (n2719,n2720,n2721);
or (n2720,n603,n2179);
or (n2721,n1844,n631);
nand (n2722,n2723,n2724);
or (n2723,n251,n2184);
or (n2724,n1838,n252);
nand (n2725,n2726,n2727);
or (n2726,n678,n2144);
or (n2727,n2643,n686);
and (n2728,n2719,n2722);
or (n2729,n2730,n2737);
and (n2730,n2731,n2736);
xor (n2731,n2732,n2735);
or (n2732,n2733,n2734);
and (n2733,n2140,n2153);
and (n2734,n2141,n2147);
xor (n2735,n2705,n2712);
xor (n2736,n2718,n2725);
and (n2737,n2732,n2735);
or (n2738,n2739,n2746);
and (n2739,n2740,n2745);
xor (n2740,n2741,n2742);
xor (n2741,n2731,n2736);
or (n2742,n2743,n2744);
and (n2743,n2164,n2191);
and (n2744,n2165,n2188);
xor (n2745,n2670,n2677);
and (n2746,n2741,n2742);
nor (n2747,n2748,n2749);
xor (n2748,n2740,n2745);
or (n2749,n2750,n2751);
and (n2750,n2130,n2163);
and (n2751,n2131,n2160);
or (n2752,n2753,n2798);
nor (n2753,n2754,n2789);
xor (n2754,n2755,n2774);
xor (n2755,n2756,n2757);
xor (n2756,n1809,n1857);
or (n2757,n2758,n2773);
and (n2758,n2759,n2766);
xor (n2759,n2760,n2763);
or (n2760,n2761,n2762);
and (n2761,n2699,n2716);
and (n2762,n2700,n2703);
or (n2763,n2764,n2765);
and (n2764,n2631,n2653);
and (n2765,n2632,n2633);
xor (n2766,n2767,n2772);
xor (n2767,n2768,n2771);
or (n2768,n2769,n2770);
and (n2769,n2634,n2647);
and (n2770,n2635,n2641);
xor (n2771,n1783,n1796);
xor (n2772,n1735,n1743);
and (n2773,n2760,n2763);
xor (n2774,n2775,n2780);
xor (n2775,n2776,n2779);
or (n2776,n2777,n2778);
and (n2777,n2767,n2772);
and (n2778,n2768,n2771);
xor (n2779,n1780,n1804);
or (n2780,n2781,n2788);
and (n2781,n2782,n2787);
xor (n2782,n2783,n2784);
xor (n2783,n1752,n1765);
or (n2784,n2785,n2786);
and (n2785,n2654,n2667);
and (n2786,n2655,n2661);
xor (n2787,n1813,n1833);
and (n2788,n2783,n2784);
or (n2789,n2790,n2797);
and (n2790,n2791,n2796);
xor (n2791,n2792,n2793);
xor (n2792,n2782,n2787);
or (n2793,n2794,n2795);
and (n2794,n2694,n2729);
and (n2795,n2695,n2698);
xor (n2796,n2759,n2766);
and (n2797,n2792,n2793);
nor (n2798,n2799,n2802);
or (n2799,n2800,n2801);
and (n2800,n2629,n2693);
and (n2801,n2630,n2668);
xor (n2802,n2791,n2796);
nand (n2803,n2804,n2813);
or (n2804,n2805,n2753);
nor (n2805,n2806,n2812);
and (n2806,n2807,n2811);
nand (n2807,n2808,n2810);
or (n2808,n2627,n2809);
nand (n2809,n2748,n2749);
nand (n2810,n2628,n2738);
not (n2811,n2798);
and (n2812,n2799,n2802);
nand (n2813,n2754,n2789);
or (n2814,n2815,n2822);
xor (n2815,n2816,n2821);
xor (n2816,n2817,n2818);
xor (n2817,n1727,n1773);
or (n2818,n2819,n2820);
and (n2819,n2775,n2780);
and (n2820,n2776,n2779);
xor (n2821,n1777,n1807);
or (n2822,n2823,n2824);
and (n2823,n2755,n2774);
and (n2824,n2756,n2757);
and (n2825,n2826,n2828);
not (n2826,n2827);
xor (n2827,n1537,n1775);
not (n2828,n2829);
or (n2829,n2830,n2831);
and (n2830,n2816,n2821);
and (n2831,n2817,n2818);
nor (n2832,n2833,n2837);
and (n2833,n2834,n2835);
not (n2834,n2825);
not (n2835,n2836);
nand (n2836,n2815,n2822);
nor (n2837,n2826,n2828);
and (n2838,n1535,n1861);
nand (n2839,n2840,n2844);
not (n2840,n2841);
or (n2841,n2842,n2843);
and (n2842,n1862,n1885);
and (n2843,n1863,n1872);
not (n2844,n2845);
xor (n2845,n2846,n2851);
xor (n2846,n2847,n2848);
xor (n2847,n1447,n1483);
or (n2848,n2849,n2850);
and (n2849,n1873,n1882);
and (n2850,n1874,n1875);
xor (n2851,n2852,n2857);
xor (n2852,n2853,n2854);
xor (n2853,n1295,n1312);
or (n2854,n2855,n2856);
and (n2855,n1876,n1879);
and (n2856,n1877,n1878);
or (n2857,n2858,n2859);
and (n2858,n1864,n1869);
and (n2859,n1865,n1866);
nor (n2860,n2844,n2840);
and (n2861,n2862,n2872);
not (n2862,n2863);
or (n2863,n2864,n2871);
and (n2864,n2865,n2868);
xor (n2865,n2866,n2867);
xor (n2866,n1513,n1518);
xor (n2867,n1292,n1445);
or (n2868,n2869,n2870);
and (n2869,n2852,n2857);
and (n2870,n2853,n2854);
and (n2871,n2866,n2867);
not (n2872,n2873);
xor (n2873,n1288,n1505);
nor (n2874,n2875,n2876);
xor (n2875,n2865,n2868);
or (n2876,n2877,n2878);
and (n2877,n2846,n2851);
and (n2878,n2847,n2848);
nor (n2879,n2880,n2884);
and (n2880,n2881,n2882);
not (n2881,n2861);
not (n2882,n2883);
nand (n2883,n2875,n2876);
nor (n2884,n2862,n2872);
and (n2885,n1286,n1521);
nand (n2886,n2887,n2889);
not (n2887,n2888);
xor (n2888,n1158,n1277);
not (n2889,n2890);
or (n2890,n2891,n2892);
and (n2891,n1522,n1527);
and (n2892,n1523,n1524);
nor (n2893,n2887,n2889);
or (n2894,n1281,n3);
xor (n2895,n2896,n5150);
xor (n2896,n2897,n5147);
xor (n2897,n2898,n5146);
xor (n2898,n2899,n5138);
xor (n2899,n2900,n5137);
xor (n2900,n2901,n5122);
xor (n2901,n2902,n5121);
xor (n2902,n2903,n5101);
xor (n2903,n2904,n5100);
xor (n2904,n2905,n5073);
xor (n2905,n2906,n5072);
xor (n2906,n2907,n5040);
xor (n2907,n2908,n5039);
xor (n2908,n2909,n5000);
xor (n2909,n2910,n4999);
xor (n2910,n2911,n4955);
xor (n2911,n2912,n4954);
xor (n2912,n2913,n4903);
xor (n2913,n2914,n4902);
xor (n2914,n2915,n4846);
xor (n2915,n2916,n4845);
xor (n2916,n2917,n4782);
xor (n2917,n2918,n4781);
xor (n2918,n2919,n4713);
xor (n2919,n2920,n4712);
xor (n2920,n2921,n4637);
xor (n2921,n2922,n4636);
xor (n2922,n2923,n4556);
xor (n2923,n2924,n4555);
xor (n2924,n2925,n4468);
xor (n2925,n2926,n4467);
xor (n2926,n2927,n4375);
xor (n2927,n2928,n4374);
xor (n2928,n2929,n4275);
xor (n2929,n2930,n4274);
xor (n2930,n2931,n4170);
xor (n2931,n2932,n4169);
xor (n2932,n2933,n4058);
xor (n2933,n2934,n4057);
xor (n2934,n2935,n3941);
xor (n2935,n2936,n3940);
xor (n2936,n2937,n3818);
xor (n2937,n2938,n3817);
xor (n2938,n2939,n3689);
xor (n2939,n2940,n3688);
xor (n2940,n2941,n3553);
xor (n2941,n2942,n3552);
xor (n2942,n2943,n3412);
xor (n2943,n2944,n3411);
xor (n2944,n2945,n3264);
xor (n2945,n2946,n3263);
xor (n2946,n2947,n3111);
xor (n2947,n2948,n3110);
xor (n2948,n2949,n2952);
xor (n2949,n2950,n2951);
and (n2950,n412,n408);
and (n2951,n398,n139);
or (n2952,n2953,n2956);
and (n2953,n2954,n2955);
and (n2954,n398,n408);
and (n2955,n241,n139);
and (n2956,n2957,n2958);
xor (n2957,n2954,n2955);
or (n2958,n2959,n2962);
and (n2959,n2960,n2961);
and (n2960,n241,n408);
and (n2961,n156,n139);
and (n2962,n2963,n2964);
xor (n2963,n2960,n2961);
or (n2964,n2965,n2968);
and (n2965,n2966,n2967);
and (n2966,n156,n408);
and (n2967,n480,n139);
and (n2968,n2969,n2970);
xor (n2969,n2966,n2967);
or (n2970,n2971,n2974);
and (n2971,n2972,n2973);
and (n2972,n480,n408);
and (n2973,n472,n139);
and (n2974,n2975,n2976);
xor (n2975,n2972,n2973);
or (n2976,n2977,n2980);
and (n2977,n2978,n2979);
and (n2978,n472,n408);
and (n2979,n280,n139);
and (n2980,n2981,n2982);
xor (n2981,n2978,n2979);
or (n2982,n2983,n2986);
and (n2983,n2984,n2985);
and (n2984,n280,n408);
and (n2985,n272,n139);
and (n2986,n2987,n2988);
xor (n2987,n2984,n2985);
or (n2988,n2989,n2992);
and (n2989,n2990,n2991);
and (n2990,n272,n408);
and (n2991,n579,n139);
and (n2992,n2993,n2994);
xor (n2993,n2990,n2991);
or (n2994,n2995,n2998);
and (n2995,n2996,n2997);
and (n2996,n579,n408);
and (n2997,n571,n139);
and (n2998,n2999,n3000);
xor (n2999,n2996,n2997);
or (n3000,n3001,n3004);
and (n3001,n3002,n3003);
and (n3002,n571,n408);
and (n3003,n451,n139);
and (n3004,n3005,n3006);
xor (n3005,n3002,n3003);
or (n3006,n3007,n3010);
and (n3007,n3008,n3009);
and (n3008,n451,n408);
and (n3009,n443,n139);
and (n3010,n3011,n3012);
xor (n3011,n3008,n3009);
or (n3012,n3013,n3016);
and (n3013,n3014,n3015);
and (n3014,n443,n408);
and (n3015,n692,n139);
and (n3016,n3017,n3018);
xor (n3017,n3014,n3015);
or (n3018,n3019,n3022);
and (n3019,n3020,n3021);
and (n3020,n692,n408);
and (n3021,n722,n139);
and (n3022,n3023,n3024);
xor (n3023,n3020,n3021);
or (n3024,n3025,n3028);
and (n3025,n3026,n3027);
and (n3026,n722,n408);
and (n3027,n714,n139);
and (n3028,n3029,n3030);
xor (n3029,n3026,n3027);
or (n3030,n3031,n3034);
and (n3031,n3032,n3033);
and (n3032,n714,n408);
and (n3033,n793,n139);
and (n3034,n3035,n3036);
xor (n3035,n3032,n3033);
or (n3036,n3037,n3040);
and (n3037,n3038,n3039);
and (n3038,n793,n408);
and (n3039,n784,n139);
and (n3040,n3041,n3042);
xor (n3041,n3038,n3039);
or (n3042,n3043,n3046);
and (n3043,n3044,n3045);
and (n3044,n784,n408);
and (n3045,n634,n139);
and (n3046,n3047,n3048);
xor (n3047,n3044,n3045);
or (n3048,n3049,n3052);
and (n3049,n3050,n3051);
and (n3050,n634,n408);
and (n3051,n625,n139);
and (n3052,n3053,n3054);
xor (n3053,n3050,n3051);
or (n3054,n3055,n3058);
and (n3055,n3056,n3057);
and (n3056,n625,n408);
and (n3057,n667,n139);
and (n3058,n3059,n3060);
xor (n3059,n3056,n3057);
or (n3060,n3061,n3064);
and (n3061,n3062,n3063);
and (n3062,n667,n408);
and (n3063,n659,n139);
and (n3064,n3065,n3066);
xor (n3065,n3062,n3063);
or (n3066,n3067,n3070);
and (n3067,n3068,n3069);
and (n3068,n659,n408);
and (n3069,n319,n139);
and (n3070,n3071,n3072);
xor (n3071,n3068,n3069);
or (n3072,n3073,n3076);
and (n3073,n3074,n3075);
and (n3074,n319,n408);
and (n3075,n311,n139);
and (n3076,n3077,n3078);
xor (n3077,n3074,n3075);
or (n3078,n3079,n3082);
and (n3079,n3080,n3081);
and (n3080,n311,n408);
and (n3081,n352,n139);
and (n3082,n3083,n3084);
xor (n3083,n3080,n3081);
or (n3084,n3085,n3088);
and (n3085,n3086,n3087);
and (n3086,n352,n408);
and (n3087,n344,n139);
and (n3088,n3089,n3090);
xor (n3089,n3086,n3087);
or (n3090,n3091,n3094);
and (n3091,n3092,n3093);
and (n3092,n344,n408);
and (n3093,n386,n139);
and (n3094,n3095,n3096);
xor (n3095,n3092,n3093);
or (n3096,n3097,n3100);
and (n3097,n3098,n3099);
and (n3098,n386,n408);
and (n3099,n378,n139);
and (n3100,n3101,n3102);
xor (n3101,n3098,n3099);
or (n3102,n3103,n3105);
and (n3103,n3104,n2577);
and (n3104,n378,n408);
and (n3105,n3106,n3107);
xor (n3106,n3104,n2577);
and (n3107,n3108,n3109);
and (n3108,n502,n408);
and (n3109,n131,n139);
and (n3110,n241,n142);
or (n3111,n3112,n3115);
and (n3112,n3113,n3114);
xor (n3113,n2957,n2958);
and (n3114,n156,n142);
and (n3115,n3116,n3117);
xor (n3116,n3113,n3114);
or (n3117,n3118,n3121);
and (n3118,n3119,n3120);
xor (n3119,n2963,n2964);
and (n3120,n480,n142);
and (n3121,n3122,n3123);
xor (n3122,n3119,n3120);
or (n3123,n3124,n3127);
and (n3124,n3125,n3126);
xor (n3125,n2969,n2970);
and (n3126,n472,n142);
and (n3127,n3128,n3129);
xor (n3128,n3125,n3126);
or (n3129,n3130,n3133);
and (n3130,n3131,n3132);
xor (n3131,n2975,n2976);
and (n3132,n280,n142);
and (n3133,n3134,n3135);
xor (n3134,n3131,n3132);
or (n3135,n3136,n3139);
and (n3136,n3137,n3138);
xor (n3137,n2981,n2982);
and (n3138,n272,n142);
and (n3139,n3140,n3141);
xor (n3140,n3137,n3138);
or (n3141,n3142,n3145);
and (n3142,n3143,n3144);
xor (n3143,n2987,n2988);
and (n3144,n579,n142);
and (n3145,n3146,n3147);
xor (n3146,n3143,n3144);
or (n3147,n3148,n3151);
and (n3148,n3149,n3150);
xor (n3149,n2993,n2994);
and (n3150,n571,n142);
and (n3151,n3152,n3153);
xor (n3152,n3149,n3150);
or (n3153,n3154,n3157);
and (n3154,n3155,n3156);
xor (n3155,n2999,n3000);
and (n3156,n451,n142);
and (n3157,n3158,n3159);
xor (n3158,n3155,n3156);
or (n3159,n3160,n3163);
and (n3160,n3161,n3162);
xor (n3161,n3005,n3006);
and (n3162,n443,n142);
and (n3163,n3164,n3165);
xor (n3164,n3161,n3162);
or (n3165,n3166,n3169);
and (n3166,n3167,n3168);
xor (n3167,n3011,n3012);
and (n3168,n692,n142);
and (n3169,n3170,n3171);
xor (n3170,n3167,n3168);
or (n3171,n3172,n3175);
and (n3172,n3173,n3174);
xor (n3173,n3017,n3018);
and (n3174,n722,n142);
and (n3175,n3176,n3177);
xor (n3176,n3173,n3174);
or (n3177,n3178,n3181);
and (n3178,n3179,n3180);
xor (n3179,n3023,n3024);
and (n3180,n714,n142);
and (n3181,n3182,n3183);
xor (n3182,n3179,n3180);
or (n3183,n3184,n3187);
and (n3184,n3185,n3186);
xor (n3185,n3029,n3030);
and (n3186,n793,n142);
and (n3187,n3188,n3189);
xor (n3188,n3185,n3186);
or (n3189,n3190,n3193);
and (n3190,n3191,n3192);
xor (n3191,n3035,n3036);
and (n3192,n784,n142);
and (n3193,n3194,n3195);
xor (n3194,n3191,n3192);
or (n3195,n3196,n3199);
and (n3196,n3197,n3198);
xor (n3197,n3041,n3042);
and (n3198,n634,n142);
and (n3199,n3200,n3201);
xor (n3200,n3197,n3198);
or (n3201,n3202,n3205);
and (n3202,n3203,n3204);
xor (n3203,n3047,n3048);
and (n3204,n625,n142);
and (n3205,n3206,n3207);
xor (n3206,n3203,n3204);
or (n3207,n3208,n3211);
and (n3208,n3209,n3210);
xor (n3209,n3053,n3054);
and (n3210,n667,n142);
and (n3211,n3212,n3213);
xor (n3212,n3209,n3210);
or (n3213,n3214,n3217);
and (n3214,n3215,n3216);
xor (n3215,n3059,n3060);
and (n3216,n659,n142);
and (n3217,n3218,n3219);
xor (n3218,n3215,n3216);
or (n3219,n3220,n3223);
and (n3220,n3221,n3222);
xor (n3221,n3065,n3066);
and (n3222,n319,n142);
and (n3223,n3224,n3225);
xor (n3224,n3221,n3222);
or (n3225,n3226,n3229);
and (n3226,n3227,n3228);
xor (n3227,n3071,n3072);
and (n3228,n311,n142);
and (n3229,n3230,n3231);
xor (n3230,n3227,n3228);
or (n3231,n3232,n3235);
and (n3232,n3233,n3234);
xor (n3233,n3077,n3078);
and (n3234,n352,n142);
and (n3235,n3236,n3237);
xor (n3236,n3233,n3234);
or (n3237,n3238,n3241);
and (n3238,n3239,n3240);
xor (n3239,n3083,n3084);
and (n3240,n344,n142);
and (n3241,n3242,n3243);
xor (n3242,n3239,n3240);
or (n3243,n3244,n3247);
and (n3244,n3245,n3246);
xor (n3245,n3089,n3090);
and (n3246,n386,n142);
and (n3247,n3248,n3249);
xor (n3248,n3245,n3246);
or (n3249,n3250,n3253);
and (n3250,n3251,n3252);
xor (n3251,n3095,n3096);
and (n3252,n378,n142);
and (n3253,n3254,n3255);
xor (n3254,n3251,n3252);
or (n3255,n3256,n3259);
and (n3256,n3257,n3258);
xor (n3257,n3101,n3102);
and (n3258,n502,n142);
and (n3259,n3260,n3261);
xor (n3260,n3257,n3258);
and (n3261,n3262,n2548);
xor (n3262,n3106,n3107);
and (n3263,n156,n150);
or (n3264,n3265,n3268);
and (n3265,n3266,n3267);
xor (n3266,n3116,n3117);
and (n3267,n480,n150);
and (n3268,n3269,n3270);
xor (n3269,n3266,n3267);
or (n3270,n3271,n3274);
and (n3271,n3272,n3273);
xor (n3272,n3122,n3123);
and (n3273,n472,n150);
and (n3274,n3275,n3276);
xor (n3275,n3272,n3273);
or (n3276,n3277,n3280);
and (n3277,n3278,n3279);
xor (n3278,n3128,n3129);
and (n3279,n280,n150);
and (n3280,n3281,n3282);
xor (n3281,n3278,n3279);
or (n3282,n3283,n3286);
and (n3283,n3284,n3285);
xor (n3284,n3134,n3135);
and (n3285,n272,n150);
and (n3286,n3287,n3288);
xor (n3287,n3284,n3285);
or (n3288,n3289,n3292);
and (n3289,n3290,n3291);
xor (n3290,n3140,n3141);
and (n3291,n579,n150);
and (n3292,n3293,n3294);
xor (n3293,n3290,n3291);
or (n3294,n3295,n3298);
and (n3295,n3296,n3297);
xor (n3296,n3146,n3147);
and (n3297,n571,n150);
and (n3298,n3299,n3300);
xor (n3299,n3296,n3297);
or (n3300,n3301,n3304);
and (n3301,n3302,n3303);
xor (n3302,n3152,n3153);
and (n3303,n451,n150);
and (n3304,n3305,n3306);
xor (n3305,n3302,n3303);
or (n3306,n3307,n3310);
and (n3307,n3308,n3309);
xor (n3308,n3158,n3159);
and (n3309,n443,n150);
and (n3310,n3311,n3312);
xor (n3311,n3308,n3309);
or (n3312,n3313,n3316);
and (n3313,n3314,n3315);
xor (n3314,n3164,n3165);
and (n3315,n692,n150);
and (n3316,n3317,n3318);
xor (n3317,n3314,n3315);
or (n3318,n3319,n3322);
and (n3319,n3320,n3321);
xor (n3320,n3170,n3171);
and (n3321,n722,n150);
and (n3322,n3323,n3324);
xor (n3323,n3320,n3321);
or (n3324,n3325,n3328);
and (n3325,n3326,n3327);
xor (n3326,n3176,n3177);
and (n3327,n714,n150);
and (n3328,n3329,n3330);
xor (n3329,n3326,n3327);
or (n3330,n3331,n3334);
and (n3331,n3332,n3333);
xor (n3332,n3182,n3183);
and (n3333,n793,n150);
and (n3334,n3335,n3336);
xor (n3335,n3332,n3333);
or (n3336,n3337,n3340);
and (n3337,n3338,n3339);
xor (n3338,n3188,n3189);
and (n3339,n784,n150);
and (n3340,n3341,n3342);
xor (n3341,n3338,n3339);
or (n3342,n3343,n3346);
and (n3343,n3344,n3345);
xor (n3344,n3194,n3195);
and (n3345,n634,n150);
and (n3346,n3347,n3348);
xor (n3347,n3344,n3345);
or (n3348,n3349,n3352);
and (n3349,n3350,n3351);
xor (n3350,n3200,n3201);
and (n3351,n625,n150);
and (n3352,n3353,n3354);
xor (n3353,n3350,n3351);
or (n3354,n3355,n3358);
and (n3355,n3356,n3357);
xor (n3356,n3206,n3207);
and (n3357,n667,n150);
and (n3358,n3359,n3360);
xor (n3359,n3356,n3357);
or (n3360,n3361,n3364);
and (n3361,n3362,n3363);
xor (n3362,n3212,n3213);
and (n3363,n659,n150);
and (n3364,n3365,n3366);
xor (n3365,n3362,n3363);
or (n3366,n3367,n3370);
and (n3367,n3368,n3369);
xor (n3368,n3218,n3219);
and (n3369,n319,n150);
and (n3370,n3371,n3372);
xor (n3371,n3368,n3369);
or (n3372,n3373,n3376);
and (n3373,n3374,n3375);
xor (n3374,n3224,n3225);
and (n3375,n311,n150);
and (n3376,n3377,n3378);
xor (n3377,n3374,n3375);
or (n3378,n3379,n3382);
and (n3379,n3380,n3381);
xor (n3380,n3230,n3231);
and (n3381,n352,n150);
and (n3382,n3383,n3384);
xor (n3383,n3380,n3381);
or (n3384,n3385,n3388);
and (n3385,n3386,n3387);
xor (n3386,n3236,n3237);
and (n3387,n344,n150);
and (n3388,n3389,n3390);
xor (n3389,n3386,n3387);
or (n3390,n3391,n3394);
and (n3391,n3392,n3393);
xor (n3392,n3242,n3243);
and (n3393,n386,n150);
and (n3394,n3395,n3396);
xor (n3395,n3392,n3393);
or (n3396,n3397,n3400);
and (n3397,n3398,n3399);
xor (n3398,n3248,n3249);
and (n3399,n378,n150);
and (n3400,n3401,n3402);
xor (n3401,n3398,n3399);
or (n3402,n3403,n3406);
and (n3403,n3404,n3405);
xor (n3404,n3254,n3255);
and (n3405,n502,n150);
and (n3406,n3407,n3408);
xor (n3407,n3404,n3405);
and (n3408,n3409,n3410);
xor (n3409,n3260,n3261);
and (n3410,n131,n150);
and (n3411,n480,n462);
or (n3412,n3413,n3416);
and (n3413,n3414,n3415);
xor (n3414,n3269,n3270);
and (n3415,n472,n462);
and (n3416,n3417,n3418);
xor (n3417,n3414,n3415);
or (n3418,n3419,n3422);
and (n3419,n3420,n3421);
xor (n3420,n3275,n3276);
and (n3421,n280,n462);
and (n3422,n3423,n3424);
xor (n3423,n3420,n3421);
or (n3424,n3425,n3428);
and (n3425,n3426,n3427);
xor (n3426,n3281,n3282);
and (n3427,n272,n462);
and (n3428,n3429,n3430);
xor (n3429,n3426,n3427);
or (n3430,n3431,n3434);
and (n3431,n3432,n3433);
xor (n3432,n3287,n3288);
and (n3433,n579,n462);
and (n3434,n3435,n3436);
xor (n3435,n3432,n3433);
or (n3436,n3437,n3440);
and (n3437,n3438,n3439);
xor (n3438,n3293,n3294);
and (n3439,n571,n462);
and (n3440,n3441,n3442);
xor (n3441,n3438,n3439);
or (n3442,n3443,n3446);
and (n3443,n3444,n3445);
xor (n3444,n3299,n3300);
and (n3445,n451,n462);
and (n3446,n3447,n3448);
xor (n3447,n3444,n3445);
or (n3448,n3449,n3452);
and (n3449,n3450,n3451);
xor (n3450,n3305,n3306);
and (n3451,n443,n462);
and (n3452,n3453,n3454);
xor (n3453,n3450,n3451);
or (n3454,n3455,n3458);
and (n3455,n3456,n3457);
xor (n3456,n3311,n3312);
and (n3457,n692,n462);
and (n3458,n3459,n3460);
xor (n3459,n3456,n3457);
or (n3460,n3461,n3464);
and (n3461,n3462,n3463);
xor (n3462,n3317,n3318);
and (n3463,n722,n462);
and (n3464,n3465,n3466);
xor (n3465,n3462,n3463);
or (n3466,n3467,n3470);
and (n3467,n3468,n3469);
xor (n3468,n3323,n3324);
and (n3469,n714,n462);
and (n3470,n3471,n3472);
xor (n3471,n3468,n3469);
or (n3472,n3473,n3476);
and (n3473,n3474,n3475);
xor (n3474,n3329,n3330);
and (n3475,n793,n462);
and (n3476,n3477,n3478);
xor (n3477,n3474,n3475);
or (n3478,n3479,n3482);
and (n3479,n3480,n3481);
xor (n3480,n3335,n3336);
and (n3481,n784,n462);
and (n3482,n3483,n3484);
xor (n3483,n3480,n3481);
or (n3484,n3485,n3488);
and (n3485,n3486,n3487);
xor (n3486,n3341,n3342);
and (n3487,n634,n462);
and (n3488,n3489,n3490);
xor (n3489,n3486,n3487);
or (n3490,n3491,n3494);
and (n3491,n3492,n3493);
xor (n3492,n3347,n3348);
and (n3493,n625,n462);
and (n3494,n3495,n3496);
xor (n3495,n3492,n3493);
or (n3496,n3497,n3500);
and (n3497,n3498,n3499);
xor (n3498,n3353,n3354);
and (n3499,n667,n462);
and (n3500,n3501,n3502);
xor (n3501,n3498,n3499);
or (n3502,n3503,n3506);
and (n3503,n3504,n3505);
xor (n3504,n3359,n3360);
and (n3505,n659,n462);
and (n3506,n3507,n3508);
xor (n3507,n3504,n3505);
or (n3508,n3509,n3512);
and (n3509,n3510,n3511);
xor (n3510,n3365,n3366);
and (n3511,n319,n462);
and (n3512,n3513,n3514);
xor (n3513,n3510,n3511);
or (n3514,n3515,n3518);
and (n3515,n3516,n3517);
xor (n3516,n3371,n3372);
and (n3517,n311,n462);
and (n3518,n3519,n3520);
xor (n3519,n3516,n3517);
or (n3520,n3521,n3524);
and (n3521,n3522,n3523);
xor (n3522,n3377,n3378);
and (n3523,n352,n462);
and (n3524,n3525,n3526);
xor (n3525,n3522,n3523);
or (n3526,n3527,n3530);
and (n3527,n3528,n3529);
xor (n3528,n3383,n3384);
and (n3529,n344,n462);
and (n3530,n3531,n3532);
xor (n3531,n3528,n3529);
or (n3532,n3533,n3536);
and (n3533,n3534,n3535);
xor (n3534,n3389,n3390);
and (n3535,n386,n462);
and (n3536,n3537,n3538);
xor (n3537,n3534,n3535);
or (n3538,n3539,n3542);
and (n3539,n3540,n3541);
xor (n3540,n3395,n3396);
and (n3541,n378,n462);
and (n3542,n3543,n3544);
xor (n3543,n3540,n3541);
or (n3544,n3545,n3548);
and (n3545,n3546,n3547);
xor (n3546,n3401,n3402);
and (n3547,n502,n462);
and (n3548,n3549,n3550);
xor (n3549,n3546,n3547);
and (n3550,n3551,n2501);
xor (n3551,n3407,n3408);
and (n3552,n472,n254);
or (n3553,n3554,n3557);
and (n3554,n3555,n3556);
xor (n3555,n3417,n3418);
and (n3556,n280,n254);
and (n3557,n3558,n3559);
xor (n3558,n3555,n3556);
or (n3559,n3560,n3563);
and (n3560,n3561,n3562);
xor (n3561,n3423,n3424);
and (n3562,n272,n254);
and (n3563,n3564,n3565);
xor (n3564,n3561,n3562);
or (n3565,n3566,n3569);
and (n3566,n3567,n3568);
xor (n3567,n3429,n3430);
and (n3568,n579,n254);
and (n3569,n3570,n3571);
xor (n3570,n3567,n3568);
or (n3571,n3572,n3575);
and (n3572,n3573,n3574);
xor (n3573,n3435,n3436);
and (n3574,n571,n254);
and (n3575,n3576,n3577);
xor (n3576,n3573,n3574);
or (n3577,n3578,n3581);
and (n3578,n3579,n3580);
xor (n3579,n3441,n3442);
and (n3580,n451,n254);
and (n3581,n3582,n3583);
xor (n3582,n3579,n3580);
or (n3583,n3584,n3587);
and (n3584,n3585,n3586);
xor (n3585,n3447,n3448);
and (n3586,n443,n254);
and (n3587,n3588,n3589);
xor (n3588,n3585,n3586);
or (n3589,n3590,n3593);
and (n3590,n3591,n3592);
xor (n3591,n3453,n3454);
and (n3592,n692,n254);
and (n3593,n3594,n3595);
xor (n3594,n3591,n3592);
or (n3595,n3596,n3599);
and (n3596,n3597,n3598);
xor (n3597,n3459,n3460);
and (n3598,n722,n254);
and (n3599,n3600,n3601);
xor (n3600,n3597,n3598);
or (n3601,n3602,n3605);
and (n3602,n3603,n3604);
xor (n3603,n3465,n3466);
and (n3604,n714,n254);
and (n3605,n3606,n3607);
xor (n3606,n3603,n3604);
or (n3607,n3608,n3611);
and (n3608,n3609,n3610);
xor (n3609,n3471,n3472);
and (n3610,n793,n254);
and (n3611,n3612,n3613);
xor (n3612,n3609,n3610);
or (n3613,n3614,n3617);
and (n3614,n3615,n3616);
xor (n3615,n3477,n3478);
and (n3616,n784,n254);
and (n3617,n3618,n3619);
xor (n3618,n3615,n3616);
or (n3619,n3620,n3623);
and (n3620,n3621,n3622);
xor (n3621,n3483,n3484);
and (n3622,n634,n254);
and (n3623,n3624,n3625);
xor (n3624,n3621,n3622);
or (n3625,n3626,n3629);
and (n3626,n3627,n3628);
xor (n3627,n3489,n3490);
and (n3628,n625,n254);
and (n3629,n3630,n3631);
xor (n3630,n3627,n3628);
or (n3631,n3632,n3635);
and (n3632,n3633,n3634);
xor (n3633,n3495,n3496);
and (n3634,n667,n254);
and (n3635,n3636,n3637);
xor (n3636,n3633,n3634);
or (n3637,n3638,n3641);
and (n3638,n3639,n3640);
xor (n3639,n3501,n3502);
and (n3640,n659,n254);
and (n3641,n3642,n3643);
xor (n3642,n3639,n3640);
or (n3643,n3644,n3647);
and (n3644,n3645,n3646);
xor (n3645,n3507,n3508);
and (n3646,n319,n254);
and (n3647,n3648,n3649);
xor (n3648,n3645,n3646);
or (n3649,n3650,n3653);
and (n3650,n3651,n3652);
xor (n3651,n3513,n3514);
and (n3652,n311,n254);
and (n3653,n3654,n3655);
xor (n3654,n3651,n3652);
or (n3655,n3656,n3659);
and (n3656,n3657,n3658);
xor (n3657,n3519,n3520);
and (n3658,n352,n254);
and (n3659,n3660,n3661);
xor (n3660,n3657,n3658);
or (n3661,n3662,n3665);
and (n3662,n3663,n3664);
xor (n3663,n3525,n3526);
and (n3664,n344,n254);
and (n3665,n3666,n3667);
xor (n3666,n3663,n3664);
or (n3667,n3668,n3671);
and (n3668,n3669,n3670);
xor (n3669,n3531,n3532);
and (n3670,n386,n254);
and (n3671,n3672,n3673);
xor (n3672,n3669,n3670);
or (n3673,n3674,n3677);
and (n3674,n3675,n3676);
xor (n3675,n3537,n3538);
and (n3676,n378,n254);
and (n3677,n3678,n3679);
xor (n3678,n3675,n3676);
or (n3679,n3680,n3683);
and (n3680,n3681,n3682);
xor (n3681,n3543,n3544);
and (n3682,n502,n254);
and (n3683,n3684,n3685);
xor (n3684,n3681,n3682);
and (n3685,n3686,n3687);
xor (n3686,n3549,n3550);
and (n3687,n131,n254);
and (n3688,n280,n257);
or (n3689,n3690,n3693);
and (n3690,n3691,n3692);
xor (n3691,n3558,n3559);
and (n3692,n272,n257);
and (n3693,n3694,n3695);
xor (n3694,n3691,n3692);
or (n3695,n3696,n3699);
and (n3696,n3697,n3698);
xor (n3697,n3564,n3565);
and (n3698,n579,n257);
and (n3699,n3700,n3701);
xor (n3700,n3697,n3698);
or (n3701,n3702,n3705);
and (n3702,n3703,n3704);
xor (n3703,n3570,n3571);
and (n3704,n571,n257);
and (n3705,n3706,n3707);
xor (n3706,n3703,n3704);
or (n3707,n3708,n3711);
and (n3708,n3709,n3710);
xor (n3709,n3576,n3577);
and (n3710,n451,n257);
and (n3711,n3712,n3713);
xor (n3712,n3709,n3710);
or (n3713,n3714,n3717);
and (n3714,n3715,n3716);
xor (n3715,n3582,n3583);
and (n3716,n443,n257);
and (n3717,n3718,n3719);
xor (n3718,n3715,n3716);
or (n3719,n3720,n3723);
and (n3720,n3721,n3722);
xor (n3721,n3588,n3589);
and (n3722,n692,n257);
and (n3723,n3724,n3725);
xor (n3724,n3721,n3722);
or (n3725,n3726,n3729);
and (n3726,n3727,n3728);
xor (n3727,n3594,n3595);
and (n3728,n722,n257);
and (n3729,n3730,n3731);
xor (n3730,n3727,n3728);
or (n3731,n3732,n3735);
and (n3732,n3733,n3734);
xor (n3733,n3600,n3601);
and (n3734,n714,n257);
and (n3735,n3736,n3737);
xor (n3736,n3733,n3734);
or (n3737,n3738,n3741);
and (n3738,n3739,n3740);
xor (n3739,n3606,n3607);
and (n3740,n793,n257);
and (n3741,n3742,n3743);
xor (n3742,n3739,n3740);
or (n3743,n3744,n3747);
and (n3744,n3745,n3746);
xor (n3745,n3612,n3613);
and (n3746,n784,n257);
and (n3747,n3748,n3749);
xor (n3748,n3745,n3746);
or (n3749,n3750,n3753);
and (n3750,n3751,n3752);
xor (n3751,n3618,n3619);
and (n3752,n634,n257);
and (n3753,n3754,n3755);
xor (n3754,n3751,n3752);
or (n3755,n3756,n3759);
and (n3756,n3757,n3758);
xor (n3757,n3624,n3625);
and (n3758,n625,n257);
and (n3759,n3760,n3761);
xor (n3760,n3757,n3758);
or (n3761,n3762,n3765);
and (n3762,n3763,n3764);
xor (n3763,n3630,n3631);
and (n3764,n667,n257);
and (n3765,n3766,n3767);
xor (n3766,n3763,n3764);
or (n3767,n3768,n3771);
and (n3768,n3769,n3770);
xor (n3769,n3636,n3637);
and (n3770,n659,n257);
and (n3771,n3772,n3773);
xor (n3772,n3769,n3770);
or (n3773,n3774,n3777);
and (n3774,n3775,n3776);
xor (n3775,n3642,n3643);
and (n3776,n319,n257);
and (n3777,n3778,n3779);
xor (n3778,n3775,n3776);
or (n3779,n3780,n3783);
and (n3780,n3781,n3782);
xor (n3781,n3648,n3649);
and (n3782,n311,n257);
and (n3783,n3784,n3785);
xor (n3784,n3781,n3782);
or (n3785,n3786,n3789);
and (n3786,n3787,n3788);
xor (n3787,n3654,n3655);
and (n3788,n352,n257);
and (n3789,n3790,n3791);
xor (n3790,n3787,n3788);
or (n3791,n3792,n3795);
and (n3792,n3793,n3794);
xor (n3793,n3660,n3661);
and (n3794,n344,n257);
and (n3795,n3796,n3797);
xor (n3796,n3793,n3794);
or (n3797,n3798,n3801);
and (n3798,n3799,n3800);
xor (n3799,n3666,n3667);
and (n3800,n386,n257);
and (n3801,n3802,n3803);
xor (n3802,n3799,n3800);
or (n3803,n3804,n3807);
and (n3804,n3805,n3806);
xor (n3805,n3672,n3673);
and (n3806,n378,n257);
and (n3807,n3808,n3809);
xor (n3808,n3805,n3806);
or (n3809,n3810,n3813);
and (n3810,n3811,n3812);
xor (n3811,n3678,n3679);
and (n3812,n502,n257);
and (n3813,n3814,n3815);
xor (n3814,n3811,n3812);
and (n3815,n3816,n2400);
xor (n3816,n3684,n3685);
and (n3817,n272,n265);
or (n3818,n3819,n3822);
and (n3819,n3820,n3821);
xor (n3820,n3694,n3695);
and (n3821,n579,n265);
and (n3822,n3823,n3824);
xor (n3823,n3820,n3821);
or (n3824,n3825,n3828);
and (n3825,n3826,n3827);
xor (n3826,n3700,n3701);
and (n3827,n571,n265);
and (n3828,n3829,n3830);
xor (n3829,n3826,n3827);
or (n3830,n3831,n3834);
and (n3831,n3832,n3833);
xor (n3832,n3706,n3707);
and (n3833,n451,n265);
and (n3834,n3835,n3836);
xor (n3835,n3832,n3833);
or (n3836,n3837,n3840);
and (n3837,n3838,n3839);
xor (n3838,n3712,n3713);
and (n3839,n443,n265);
and (n3840,n3841,n3842);
xor (n3841,n3838,n3839);
or (n3842,n3843,n3846);
and (n3843,n3844,n3845);
xor (n3844,n3718,n3719);
and (n3845,n692,n265);
and (n3846,n3847,n3848);
xor (n3847,n3844,n3845);
or (n3848,n3849,n3852);
and (n3849,n3850,n3851);
xor (n3850,n3724,n3725);
and (n3851,n722,n265);
and (n3852,n3853,n3854);
xor (n3853,n3850,n3851);
or (n3854,n3855,n3858);
and (n3855,n3856,n3857);
xor (n3856,n3730,n3731);
and (n3857,n714,n265);
and (n3858,n3859,n3860);
xor (n3859,n3856,n3857);
or (n3860,n3861,n3864);
and (n3861,n3862,n3863);
xor (n3862,n3736,n3737);
and (n3863,n793,n265);
and (n3864,n3865,n3866);
xor (n3865,n3862,n3863);
or (n3866,n3867,n3870);
and (n3867,n3868,n3869);
xor (n3868,n3742,n3743);
and (n3869,n784,n265);
and (n3870,n3871,n3872);
xor (n3871,n3868,n3869);
or (n3872,n3873,n3876);
and (n3873,n3874,n3875);
xor (n3874,n3748,n3749);
and (n3875,n634,n265);
and (n3876,n3877,n3878);
xor (n3877,n3874,n3875);
or (n3878,n3879,n3882);
and (n3879,n3880,n3881);
xor (n3880,n3754,n3755);
and (n3881,n625,n265);
and (n3882,n3883,n3884);
xor (n3883,n3880,n3881);
or (n3884,n3885,n3888);
and (n3885,n3886,n3887);
xor (n3886,n3760,n3761);
and (n3887,n667,n265);
and (n3888,n3889,n3890);
xor (n3889,n3886,n3887);
or (n3890,n3891,n3894);
and (n3891,n3892,n3893);
xor (n3892,n3766,n3767);
and (n3893,n659,n265);
and (n3894,n3895,n3896);
xor (n3895,n3892,n3893);
or (n3896,n3897,n3900);
and (n3897,n3898,n3899);
xor (n3898,n3772,n3773);
and (n3899,n319,n265);
and (n3900,n3901,n3902);
xor (n3901,n3898,n3899);
or (n3902,n3903,n3906);
and (n3903,n3904,n3905);
xor (n3904,n3778,n3779);
and (n3905,n311,n265);
and (n3906,n3907,n3908);
xor (n3907,n3904,n3905);
or (n3908,n3909,n3912);
and (n3909,n3910,n3911);
xor (n3910,n3784,n3785);
and (n3911,n352,n265);
and (n3912,n3913,n3914);
xor (n3913,n3910,n3911);
or (n3914,n3915,n3918);
and (n3915,n3916,n3917);
xor (n3916,n3790,n3791);
and (n3917,n344,n265);
and (n3918,n3919,n3920);
xor (n3919,n3916,n3917);
or (n3920,n3921,n3923);
and (n3921,n3922,n2264);
xor (n3922,n3796,n3797);
and (n3923,n3924,n3925);
xor (n3924,n3922,n2264);
or (n3925,n3926,n3929);
and (n3926,n3927,n3928);
xor (n3927,n3802,n3803);
and (n3928,n378,n265);
and (n3929,n3930,n3931);
xor (n3930,n3927,n3928);
or (n3931,n3932,n3935);
and (n3932,n3933,n3934);
xor (n3933,n3808,n3809);
and (n3934,n502,n265);
and (n3935,n3936,n3937);
xor (n3936,n3933,n3934);
and (n3937,n3938,n3939);
xor (n3938,n3814,n3815);
and (n3939,n131,n265);
and (n3940,n579,n681);
or (n3941,n3942,n3945);
and (n3942,n3943,n3944);
xor (n3943,n3823,n3824);
and (n3944,n571,n681);
and (n3945,n3946,n3947);
xor (n3946,n3943,n3944);
or (n3947,n3948,n3951);
and (n3948,n3949,n3950);
xor (n3949,n3829,n3830);
and (n3950,n451,n681);
and (n3951,n3952,n3953);
xor (n3952,n3949,n3950);
or (n3953,n3954,n3957);
and (n3954,n3955,n3956);
xor (n3955,n3835,n3836);
and (n3956,n443,n681);
and (n3957,n3958,n3959);
xor (n3958,n3955,n3956);
or (n3959,n3960,n3963);
and (n3960,n3961,n3962);
xor (n3961,n3841,n3842);
and (n3962,n692,n681);
and (n3963,n3964,n3965);
xor (n3964,n3961,n3962);
or (n3965,n3966,n3969);
and (n3966,n3967,n3968);
xor (n3967,n3847,n3848);
and (n3968,n722,n681);
and (n3969,n3970,n3971);
xor (n3970,n3967,n3968);
or (n3971,n3972,n3975);
and (n3972,n3973,n3974);
xor (n3973,n3853,n3854);
and (n3974,n714,n681);
and (n3975,n3976,n3977);
xor (n3976,n3973,n3974);
or (n3977,n3978,n3981);
and (n3978,n3979,n3980);
xor (n3979,n3859,n3860);
and (n3980,n793,n681);
and (n3981,n3982,n3983);
xor (n3982,n3979,n3980);
or (n3983,n3984,n3987);
and (n3984,n3985,n3986);
xor (n3985,n3865,n3866);
and (n3986,n784,n681);
and (n3987,n3988,n3989);
xor (n3988,n3985,n3986);
or (n3989,n3990,n3993);
and (n3990,n3991,n3992);
xor (n3991,n3871,n3872);
and (n3992,n634,n681);
and (n3993,n3994,n3995);
xor (n3994,n3991,n3992);
or (n3995,n3996,n3999);
and (n3996,n3997,n3998);
xor (n3997,n3877,n3878);
and (n3998,n625,n681);
and (n3999,n4000,n4001);
xor (n4000,n3997,n3998);
or (n4001,n4002,n4005);
and (n4002,n4003,n4004);
xor (n4003,n3883,n3884);
and (n4004,n667,n681);
and (n4005,n4006,n4007);
xor (n4006,n4003,n4004);
or (n4007,n4008,n4011);
and (n4008,n4009,n4010);
xor (n4009,n3889,n3890);
and (n4010,n659,n681);
and (n4011,n4012,n4013);
xor (n4012,n4009,n4010);
or (n4013,n4014,n4017);
and (n4014,n4015,n4016);
xor (n4015,n3895,n3896);
and (n4016,n319,n681);
and (n4017,n4018,n4019);
xor (n4018,n4015,n4016);
or (n4019,n4020,n4023);
and (n4020,n4021,n4022);
xor (n4021,n3901,n3902);
and (n4022,n311,n681);
and (n4023,n4024,n4025);
xor (n4024,n4021,n4022);
or (n4025,n4026,n4029);
and (n4026,n4027,n4028);
xor (n4027,n3907,n3908);
and (n4028,n352,n681);
and (n4029,n4030,n4031);
xor (n4030,n4027,n4028);
or (n4031,n4032,n4035);
and (n4032,n4033,n4034);
xor (n4033,n3913,n3914);
and (n4034,n344,n681);
and (n4035,n4036,n4037);
xor (n4036,n4033,n4034);
or (n4037,n4038,n4041);
and (n4038,n4039,n4040);
xor (n4039,n3919,n3920);
and (n4040,n386,n681);
and (n4041,n4042,n4043);
xor (n4042,n4039,n4040);
or (n4043,n4044,n4047);
and (n4044,n4045,n4046);
xor (n4045,n3924,n3925);
and (n4046,n378,n681);
and (n4047,n4048,n4049);
xor (n4048,n4045,n4046);
or (n4049,n4050,n4053);
and (n4050,n4051,n4052);
xor (n4051,n3930,n3931);
and (n4052,n502,n681);
and (n4053,n4054,n4055);
xor (n4054,n4051,n4052);
and (n4055,n4056,n2293);
xor (n4056,n3936,n3937);
and (n4057,n571,n428);
or (n4058,n4059,n4062);
and (n4059,n4060,n4061);
xor (n4060,n3946,n3947);
and (n4061,n451,n428);
and (n4062,n4063,n4064);
xor (n4063,n4060,n4061);
or (n4064,n4065,n4068);
and (n4065,n4066,n4067);
xor (n4066,n3952,n3953);
and (n4067,n443,n428);
and (n4068,n4069,n4070);
xor (n4069,n4066,n4067);
or (n4070,n4071,n4074);
and (n4071,n4072,n4073);
xor (n4072,n3958,n3959);
and (n4073,n692,n428);
and (n4074,n4075,n4076);
xor (n4075,n4072,n4073);
or (n4076,n4077,n4080);
and (n4077,n4078,n4079);
xor (n4078,n3964,n3965);
and (n4079,n722,n428);
and (n4080,n4081,n4082);
xor (n4081,n4078,n4079);
or (n4082,n4083,n4086);
and (n4083,n4084,n4085);
xor (n4084,n3970,n3971);
and (n4085,n714,n428);
and (n4086,n4087,n4088);
xor (n4087,n4084,n4085);
or (n4088,n4089,n4092);
and (n4089,n4090,n4091);
xor (n4090,n3976,n3977);
and (n4091,n793,n428);
and (n4092,n4093,n4094);
xor (n4093,n4090,n4091);
or (n4094,n4095,n4098);
and (n4095,n4096,n4097);
xor (n4096,n3982,n3983);
and (n4097,n784,n428);
and (n4098,n4099,n4100);
xor (n4099,n4096,n4097);
or (n4100,n4101,n4104);
and (n4101,n4102,n4103);
xor (n4102,n3988,n3989);
and (n4103,n634,n428);
and (n4104,n4105,n4106);
xor (n4105,n4102,n4103);
or (n4106,n4107,n4110);
and (n4107,n4108,n4109);
xor (n4108,n3994,n3995);
and (n4109,n625,n428);
and (n4110,n4111,n4112);
xor (n4111,n4108,n4109);
or (n4112,n4113,n4116);
and (n4113,n4114,n4115);
xor (n4114,n4000,n4001);
and (n4115,n667,n428);
and (n4116,n4117,n4118);
xor (n4117,n4114,n4115);
or (n4118,n4119,n4122);
and (n4119,n4120,n4121);
xor (n4120,n4006,n4007);
and (n4121,n659,n428);
and (n4122,n4123,n4124);
xor (n4123,n4120,n4121);
or (n4124,n4125,n4128);
and (n4125,n4126,n4127);
xor (n4126,n4012,n4013);
and (n4127,n319,n428);
and (n4128,n4129,n4130);
xor (n4129,n4126,n4127);
or (n4130,n4131,n4134);
and (n4131,n4132,n4133);
xor (n4132,n4018,n4019);
and (n4133,n311,n428);
and (n4134,n4135,n4136);
xor (n4135,n4132,n4133);
or (n4136,n4137,n4140);
and (n4137,n4138,n4139);
xor (n4138,n4024,n4025);
and (n4139,n352,n428);
and (n4140,n4141,n4142);
xor (n4141,n4138,n4139);
or (n4142,n4143,n4146);
and (n4143,n4144,n4145);
xor (n4144,n4030,n4031);
and (n4145,n344,n428);
and (n4146,n4147,n4148);
xor (n4147,n4144,n4145);
or (n4148,n4149,n4152);
and (n4149,n4150,n4151);
xor (n4150,n4036,n4037);
and (n4151,n386,n428);
and (n4152,n4153,n4154);
xor (n4153,n4150,n4151);
or (n4154,n4155,n4158);
and (n4155,n4156,n4157);
xor (n4156,n4042,n4043);
and (n4157,n378,n428);
and (n4158,n4159,n4160);
xor (n4159,n4156,n4157);
or (n4160,n4161,n4164);
and (n4161,n4162,n4163);
xor (n4162,n4048,n4049);
and (n4163,n502,n428);
and (n4164,n4165,n4166);
xor (n4165,n4162,n4163);
and (n4166,n4167,n4168);
xor (n4167,n4054,n4055);
and (n4168,n131,n428);
and (n4169,n451,n425);
or (n4170,n4171,n4174);
and (n4171,n4172,n4173);
xor (n4172,n4063,n4064);
and (n4173,n443,n425);
and (n4174,n4175,n4176);
xor (n4175,n4172,n4173);
or (n4176,n4177,n4180);
and (n4177,n4178,n4179);
xor (n4178,n4069,n4070);
and (n4179,n692,n425);
and (n4180,n4181,n4182);
xor (n4181,n4178,n4179);
or (n4182,n4183,n4186);
and (n4183,n4184,n4185);
xor (n4184,n4075,n4076);
and (n4185,n722,n425);
and (n4186,n4187,n4188);
xor (n4187,n4184,n4185);
or (n4188,n4189,n4192);
and (n4189,n4190,n4191);
xor (n4190,n4081,n4082);
and (n4191,n714,n425);
and (n4192,n4193,n4194);
xor (n4193,n4190,n4191);
or (n4194,n4195,n4198);
and (n4195,n4196,n4197);
xor (n4196,n4087,n4088);
and (n4197,n793,n425);
and (n4198,n4199,n4200);
xor (n4199,n4196,n4197);
or (n4200,n4201,n4204);
and (n4201,n4202,n4203);
xor (n4202,n4093,n4094);
and (n4203,n784,n425);
and (n4204,n4205,n4206);
xor (n4205,n4202,n4203);
or (n4206,n4207,n4210);
and (n4207,n4208,n4209);
xor (n4208,n4099,n4100);
and (n4209,n634,n425);
and (n4210,n4211,n4212);
xor (n4211,n4208,n4209);
or (n4212,n4213,n4216);
and (n4213,n4214,n4215);
xor (n4214,n4105,n4106);
and (n4215,n625,n425);
and (n4216,n4217,n4218);
xor (n4217,n4214,n4215);
or (n4218,n4219,n4222);
and (n4219,n4220,n4221);
xor (n4220,n4111,n4112);
and (n4221,n667,n425);
and (n4222,n4223,n4224);
xor (n4223,n4220,n4221);
or (n4224,n4225,n4228);
and (n4225,n4226,n4227);
xor (n4226,n4117,n4118);
and (n4227,n659,n425);
and (n4228,n4229,n4230);
xor (n4229,n4226,n4227);
or (n4230,n4231,n4234);
and (n4231,n4232,n4233);
xor (n4232,n4123,n4124);
and (n4233,n319,n425);
and (n4234,n4235,n4236);
xor (n4235,n4232,n4233);
or (n4236,n4237,n4240);
and (n4237,n4238,n4239);
xor (n4238,n4129,n4130);
and (n4239,n311,n425);
and (n4240,n4241,n4242);
xor (n4241,n4238,n4239);
or (n4242,n4243,n4246);
and (n4243,n4244,n4245);
xor (n4244,n4135,n4136);
and (n4245,n352,n425);
and (n4246,n4247,n4248);
xor (n4247,n4244,n4245);
or (n4248,n4249,n4252);
and (n4249,n4250,n4251);
xor (n4250,n4141,n4142);
and (n4251,n344,n425);
and (n4252,n4253,n4254);
xor (n4253,n4250,n4251);
or (n4254,n4255,n4258);
and (n4255,n4256,n4257);
xor (n4256,n4147,n4148);
and (n4257,n386,n425);
and (n4258,n4259,n4260);
xor (n4259,n4256,n4257);
or (n4260,n4261,n4264);
and (n4261,n4262,n4263);
xor (n4262,n4153,n4154);
and (n4263,n378,n425);
and (n4264,n4265,n4266);
xor (n4265,n4262,n4263);
or (n4266,n4267,n4270);
and (n4267,n4268,n4269);
xor (n4268,n4159,n4160);
and (n4269,n502,n425);
and (n4270,n4271,n4272);
xor (n4271,n4268,n4269);
and (n4272,n4273,n2102);
xor (n4273,n4165,n4166);
and (n4274,n443,n436);
or (n4275,n4276,n4279);
and (n4276,n4277,n4278);
xor (n4277,n4175,n4176);
and (n4278,n692,n436);
and (n4279,n4280,n4281);
xor (n4280,n4277,n4278);
or (n4281,n4282,n4285);
and (n4282,n4283,n4284);
xor (n4283,n4181,n4182);
and (n4284,n722,n436);
and (n4285,n4286,n4287);
xor (n4286,n4283,n4284);
or (n4287,n4288,n4291);
and (n4288,n4289,n4290);
xor (n4289,n4187,n4188);
and (n4290,n714,n436);
and (n4291,n4292,n4293);
xor (n4292,n4289,n4290);
or (n4293,n4294,n4297);
and (n4294,n4295,n4296);
xor (n4295,n4193,n4194);
and (n4296,n793,n436);
and (n4297,n4298,n4299);
xor (n4298,n4295,n4296);
or (n4299,n4300,n4303);
and (n4300,n4301,n4302);
xor (n4301,n4199,n4200);
and (n4302,n784,n436);
and (n4303,n4304,n4305);
xor (n4304,n4301,n4302);
or (n4305,n4306,n4309);
and (n4306,n4307,n4308);
xor (n4307,n4205,n4206);
and (n4308,n634,n436);
and (n4309,n4310,n4311);
xor (n4310,n4307,n4308);
or (n4311,n4312,n4315);
and (n4312,n4313,n4314);
xor (n4313,n4211,n4212);
and (n4314,n625,n436);
and (n4315,n4316,n4317);
xor (n4316,n4313,n4314);
or (n4317,n4318,n4321);
and (n4318,n4319,n4320);
xor (n4319,n4217,n4218);
and (n4320,n667,n436);
and (n4321,n4322,n4323);
xor (n4322,n4319,n4320);
or (n4323,n4324,n4327);
and (n4324,n4325,n4326);
xor (n4325,n4223,n4224);
and (n4326,n659,n436);
and (n4327,n4328,n4329);
xor (n4328,n4325,n4326);
or (n4329,n4330,n4333);
and (n4330,n4331,n4332);
xor (n4331,n4229,n4230);
and (n4332,n319,n436);
and (n4333,n4334,n4335);
xor (n4334,n4331,n4332);
or (n4335,n4336,n4339);
and (n4336,n4337,n4338);
xor (n4337,n4235,n4236);
and (n4338,n311,n436);
and (n4339,n4340,n4341);
xor (n4340,n4337,n4338);
or (n4341,n4342,n4345);
and (n4342,n4343,n4344);
xor (n4343,n4241,n4242);
and (n4344,n352,n436);
and (n4345,n4346,n4347);
xor (n4346,n4343,n4344);
or (n4347,n4348,n4351);
and (n4348,n4349,n4350);
xor (n4349,n4247,n4248);
and (n4350,n344,n436);
and (n4351,n4352,n4353);
xor (n4352,n4349,n4350);
or (n4353,n4354,n4357);
and (n4354,n4355,n4356);
xor (n4355,n4253,n4254);
and (n4356,n386,n436);
and (n4357,n4358,n4359);
xor (n4358,n4355,n4356);
or (n4359,n4360,n4363);
and (n4360,n4361,n4362);
xor (n4361,n4259,n4260);
and (n4362,n378,n436);
and (n4363,n4364,n4365);
xor (n4364,n4361,n4362);
or (n4365,n4366,n4369);
and (n4366,n4367,n4368);
xor (n4367,n4265,n4266);
and (n4368,n502,n436);
and (n4369,n4370,n4371);
xor (n4370,n4367,n4368);
and (n4371,n4372,n4373);
xor (n4372,n4271,n4272);
and (n4373,n131,n436);
and (n4374,n692,n774);
or (n4375,n4376,n4379);
and (n4376,n4377,n4378);
xor (n4377,n4280,n4281);
and (n4378,n722,n774);
and (n4379,n4380,n4381);
xor (n4380,n4377,n4378);
or (n4381,n4382,n4385);
and (n4382,n4383,n4384);
xor (n4383,n4286,n4287);
and (n4384,n714,n774);
and (n4385,n4386,n4387);
xor (n4386,n4383,n4384);
or (n4387,n4388,n4391);
and (n4388,n4389,n4390);
xor (n4389,n4292,n4293);
and (n4390,n793,n774);
and (n4391,n4392,n4393);
xor (n4392,n4389,n4390);
or (n4393,n4394,n4397);
and (n4394,n4395,n4396);
xor (n4395,n4298,n4299);
and (n4396,n784,n774);
and (n4397,n4398,n4399);
xor (n4398,n4395,n4396);
or (n4399,n4400,n4403);
and (n4400,n4401,n4402);
xor (n4401,n4304,n4305);
and (n4402,n634,n774);
and (n4403,n4404,n4405);
xor (n4404,n4401,n4402);
or (n4405,n4406,n4409);
and (n4406,n4407,n4408);
xor (n4407,n4310,n4311);
and (n4408,n625,n774);
and (n4409,n4410,n4411);
xor (n4410,n4407,n4408);
or (n4411,n4412,n4415);
and (n4412,n4413,n4414);
xor (n4413,n4316,n4317);
and (n4414,n667,n774);
and (n4415,n4416,n4417);
xor (n4416,n4413,n4414);
or (n4417,n4418,n4421);
and (n4418,n4419,n4420);
xor (n4419,n4322,n4323);
and (n4420,n659,n774);
and (n4421,n4422,n4423);
xor (n4422,n4419,n4420);
or (n4423,n4424,n4427);
and (n4424,n4425,n4426);
xor (n4425,n4328,n4329);
and (n4426,n319,n774);
and (n4427,n4428,n4429);
xor (n4428,n4425,n4426);
or (n4429,n4430,n4433);
and (n4430,n4431,n4432);
xor (n4431,n4334,n4335);
and (n4432,n311,n774);
and (n4433,n4434,n4435);
xor (n4434,n4431,n4432);
or (n4435,n4436,n4439);
and (n4436,n4437,n4438);
xor (n4437,n4340,n4341);
and (n4438,n352,n774);
and (n4439,n4440,n4441);
xor (n4440,n4437,n4438);
or (n4441,n4442,n4445);
and (n4442,n4443,n4444);
xor (n4443,n4346,n4347);
and (n4444,n344,n774);
and (n4445,n4446,n4447);
xor (n4446,n4443,n4444);
or (n4447,n4448,n4451);
and (n4448,n4449,n4450);
xor (n4449,n4352,n4353);
and (n4450,n386,n774);
and (n4451,n4452,n4453);
xor (n4452,n4449,n4450);
or (n4453,n4454,n4457);
and (n4454,n4455,n4456);
xor (n4455,n4358,n4359);
and (n4456,n378,n774);
and (n4457,n4458,n4459);
xor (n4458,n4455,n4456);
or (n4459,n4460,n4463);
and (n4460,n4461,n4462);
xor (n4461,n4364,n4365);
and (n4462,n502,n774);
and (n4463,n4464,n4465);
xor (n4464,n4461,n4462);
and (n4465,n4466,n2011);
xor (n4466,n4370,n4371);
and (n4467,n722,n608);
or (n4468,n4469,n4472);
and (n4469,n4470,n4471);
xor (n4470,n4380,n4381);
and (n4471,n714,n608);
and (n4472,n4473,n4474);
xor (n4473,n4470,n4471);
or (n4474,n4475,n4478);
and (n4475,n4476,n4477);
xor (n4476,n4386,n4387);
and (n4477,n793,n608);
and (n4478,n4479,n4480);
xor (n4479,n4476,n4477);
or (n4480,n4481,n4484);
and (n4481,n4482,n4483);
xor (n4482,n4392,n4393);
and (n4483,n784,n608);
and (n4484,n4485,n4486);
xor (n4485,n4482,n4483);
or (n4486,n4487,n4490);
and (n4487,n4488,n4489);
xor (n4488,n4398,n4399);
and (n4489,n634,n608);
and (n4490,n4491,n4492);
xor (n4491,n4488,n4489);
or (n4492,n4493,n4496);
and (n4493,n4494,n4495);
xor (n4494,n4404,n4405);
and (n4495,n625,n608);
and (n4496,n4497,n4498);
xor (n4497,n4494,n4495);
or (n4498,n4499,n4502);
and (n4499,n4500,n4501);
xor (n4500,n4410,n4411);
and (n4501,n667,n608);
and (n4502,n4503,n4504);
xor (n4503,n4500,n4501);
or (n4504,n4505,n4508);
and (n4505,n4506,n4507);
xor (n4506,n4416,n4417);
and (n4507,n659,n608);
and (n4508,n4509,n4510);
xor (n4509,n4506,n4507);
or (n4510,n4511,n4514);
and (n4511,n4512,n4513);
xor (n4512,n4422,n4423);
and (n4513,n319,n608);
and (n4514,n4515,n4516);
xor (n4515,n4512,n4513);
or (n4516,n4517,n4520);
and (n4517,n4518,n4519);
xor (n4518,n4428,n4429);
and (n4519,n311,n608);
and (n4520,n4521,n4522);
xor (n4521,n4518,n4519);
or (n4522,n4523,n4526);
and (n4523,n4524,n4525);
xor (n4524,n4434,n4435);
and (n4525,n352,n608);
and (n4526,n4527,n4528);
xor (n4527,n4524,n4525);
or (n4528,n4529,n4532);
and (n4529,n4530,n4531);
xor (n4530,n4440,n4441);
and (n4531,n344,n608);
and (n4532,n4533,n4534);
xor (n4533,n4530,n4531);
or (n4534,n4535,n4538);
and (n4535,n4536,n4537);
xor (n4536,n4446,n4447);
and (n4537,n386,n608);
and (n4538,n4539,n4540);
xor (n4539,n4536,n4537);
or (n4540,n4541,n4544);
and (n4541,n4542,n4543);
xor (n4542,n4452,n4453);
and (n4543,n378,n608);
and (n4544,n4545,n4546);
xor (n4545,n4542,n4543);
or (n4546,n4547,n4550);
and (n4547,n4548,n4549);
xor (n4548,n4458,n4459);
and (n4549,n502,n608);
and (n4550,n4551,n4552);
xor (n4551,n4548,n4549);
and (n4552,n4553,n4554);
xor (n4553,n4464,n4465);
and (n4554,n131,n608);
and (n4555,n714,n611);
or (n4556,n4557,n4560);
and (n4557,n4558,n4559);
xor (n4558,n4473,n4474);
and (n4559,n793,n611);
and (n4560,n4561,n4562);
xor (n4561,n4558,n4559);
or (n4562,n4563,n4566);
and (n4563,n4564,n4565);
xor (n4564,n4479,n4480);
and (n4565,n784,n611);
and (n4566,n4567,n4568);
xor (n4567,n4564,n4565);
or (n4568,n4569,n4572);
and (n4569,n4570,n4571);
xor (n4570,n4485,n4486);
and (n4571,n634,n611);
and (n4572,n4573,n4574);
xor (n4573,n4570,n4571);
or (n4574,n4575,n4578);
and (n4575,n4576,n4577);
xor (n4576,n4491,n4492);
and (n4577,n625,n611);
and (n4578,n4579,n4580);
xor (n4579,n4576,n4577);
or (n4580,n4581,n4584);
and (n4581,n4582,n4583);
xor (n4582,n4497,n4498);
and (n4583,n667,n611);
and (n4584,n4585,n4586);
xor (n4585,n4582,n4583);
or (n4586,n4587,n4590);
and (n4587,n4588,n4589);
xor (n4588,n4503,n4504);
and (n4589,n659,n611);
and (n4590,n4591,n4592);
xor (n4591,n4588,n4589);
or (n4592,n4593,n4596);
and (n4593,n4594,n4595);
xor (n4594,n4509,n4510);
and (n4595,n319,n611);
and (n4596,n4597,n4598);
xor (n4597,n4594,n4595);
or (n4598,n4599,n4602);
and (n4599,n4600,n4601);
xor (n4600,n4515,n4516);
and (n4601,n311,n611);
and (n4602,n4603,n4604);
xor (n4603,n4600,n4601);
or (n4604,n4605,n4608);
and (n4605,n4606,n4607);
xor (n4606,n4521,n4522);
and (n4607,n352,n611);
and (n4608,n4609,n4610);
xor (n4609,n4606,n4607);
or (n4610,n4611,n4614);
and (n4611,n4612,n4613);
xor (n4612,n4527,n4528);
and (n4613,n344,n611);
and (n4614,n4615,n4616);
xor (n4615,n4612,n4613);
or (n4616,n4617,n4620);
and (n4617,n4618,n4619);
xor (n4618,n4533,n4534);
and (n4619,n386,n611);
and (n4620,n4621,n4622);
xor (n4621,n4618,n4619);
or (n4622,n4623,n4626);
and (n4623,n4624,n4625);
xor (n4624,n4539,n4540);
and (n4625,n378,n611);
and (n4626,n4627,n4628);
xor (n4627,n4624,n4625);
or (n4628,n4629,n4632);
and (n4629,n4630,n4631);
xor (n4630,n4545,n4546);
and (n4631,n502,n611);
and (n4632,n4633,n4634);
xor (n4633,n4630,n4631);
and (n4634,n4635,n2210);
xor (n4635,n4551,n4552);
and (n4636,n793,n618);
or (n4637,n4638,n4641);
and (n4638,n4639,n4640);
xor (n4639,n4561,n4562);
and (n4640,n784,n618);
and (n4641,n4642,n4643);
xor (n4642,n4639,n4640);
or (n4643,n4644,n4647);
and (n4644,n4645,n4646);
xor (n4645,n4567,n4568);
and (n4646,n634,n618);
and (n4647,n4648,n4649);
xor (n4648,n4645,n4646);
or (n4649,n4650,n4653);
and (n4650,n4651,n4652);
xor (n4651,n4573,n4574);
and (n4652,n625,n618);
and (n4653,n4654,n4655);
xor (n4654,n4651,n4652);
or (n4655,n4656,n4659);
and (n4656,n4657,n4658);
xor (n4657,n4579,n4580);
and (n4658,n667,n618);
and (n4659,n4660,n4661);
xor (n4660,n4657,n4658);
or (n4661,n4662,n4665);
and (n4662,n4663,n4664);
xor (n4663,n4585,n4586);
and (n4664,n659,n618);
and (n4665,n4666,n4667);
xor (n4666,n4663,n4664);
or (n4667,n4668,n4671);
and (n4668,n4669,n4670);
xor (n4669,n4591,n4592);
and (n4670,n319,n618);
and (n4671,n4672,n4673);
xor (n4672,n4669,n4670);
or (n4673,n4674,n4677);
and (n4674,n4675,n4676);
xor (n4675,n4597,n4598);
and (n4676,n311,n618);
and (n4677,n4678,n4679);
xor (n4678,n4675,n4676);
or (n4679,n4680,n4683);
and (n4680,n4681,n4682);
xor (n4681,n4603,n4604);
and (n4682,n352,n618);
and (n4683,n4684,n4685);
xor (n4684,n4681,n4682);
or (n4685,n4686,n4689);
and (n4686,n4687,n4688);
xor (n4687,n4609,n4610);
and (n4688,n344,n618);
and (n4689,n4690,n4691);
xor (n4690,n4687,n4688);
or (n4691,n4692,n4695);
and (n4692,n4693,n4694);
xor (n4693,n4615,n4616);
and (n4694,n386,n618);
and (n4695,n4696,n4697);
xor (n4696,n4693,n4694);
or (n4697,n4698,n4701);
and (n4698,n4699,n4700);
xor (n4699,n4621,n4622);
and (n4700,n378,n618);
and (n4701,n4702,n4703);
xor (n4702,n4699,n4700);
or (n4703,n4704,n4707);
and (n4704,n4705,n4706);
xor (n4705,n4627,n4628);
and (n4706,n502,n618);
and (n4707,n4708,n4709);
xor (n4708,n4705,n4706);
and (n4709,n4710,n4711);
xor (n4710,n4633,n4634);
and (n4711,n131,n618);
and (n4712,n784,n646);
or (n4713,n4714,n4717);
and (n4714,n4715,n4716);
xor (n4715,n4642,n4643);
and (n4716,n634,n646);
and (n4717,n4718,n4719);
xor (n4718,n4715,n4716);
or (n4719,n4720,n4723);
and (n4720,n4721,n4722);
xor (n4721,n4648,n4649);
and (n4722,n625,n646);
and (n4723,n4724,n4725);
xor (n4724,n4721,n4722);
or (n4725,n4726,n4729);
and (n4726,n4727,n4728);
xor (n4727,n4654,n4655);
and (n4728,n667,n646);
and (n4729,n4730,n4731);
xor (n4730,n4727,n4728);
or (n4731,n4732,n4735);
and (n4732,n4733,n4734);
xor (n4733,n4660,n4661);
and (n4734,n659,n646);
and (n4735,n4736,n4737);
xor (n4736,n4733,n4734);
or (n4737,n4738,n4741);
and (n4738,n4739,n4740);
xor (n4739,n4666,n4667);
and (n4740,n319,n646);
and (n4741,n4742,n4743);
xor (n4742,n4739,n4740);
or (n4743,n4744,n4747);
and (n4744,n4745,n4746);
xor (n4745,n4672,n4673);
and (n4746,n311,n646);
and (n4747,n4748,n4749);
xor (n4748,n4745,n4746);
or (n4749,n4750,n4753);
and (n4750,n4751,n4752);
xor (n4751,n4678,n4679);
and (n4752,n352,n646);
and (n4753,n4754,n4755);
xor (n4754,n4751,n4752);
or (n4755,n4756,n4759);
and (n4756,n4757,n4758);
xor (n4757,n4684,n4685);
and (n4758,n344,n646);
and (n4759,n4760,n4761);
xor (n4760,n4757,n4758);
or (n4761,n4762,n4765);
and (n4762,n4763,n4764);
xor (n4763,n4690,n4691);
and (n4764,n386,n646);
and (n4765,n4766,n4767);
xor (n4766,n4763,n4764);
or (n4767,n4768,n4771);
and (n4768,n4769,n4770);
xor (n4769,n4696,n4697);
and (n4770,n378,n646);
and (n4771,n4772,n4773);
xor (n4772,n4769,n4770);
or (n4773,n4774,n4777);
and (n4774,n4775,n4776);
xor (n4775,n4702,n4703);
and (n4776,n502,n646);
and (n4777,n4778,n4779);
xor (n4778,n4775,n4776);
and (n4779,n4780,n1825);
xor (n4780,n4708,n4709);
and (n4781,n634,n652);
or (n4782,n4783,n4786);
and (n4783,n4784,n4785);
xor (n4784,n4718,n4719);
and (n4785,n625,n652);
and (n4786,n4787,n4788);
xor (n4787,n4784,n4785);
or (n4788,n4789,n4792);
and (n4789,n4790,n4791);
xor (n4790,n4724,n4725);
and (n4791,n667,n652);
and (n4792,n4793,n4794);
xor (n4793,n4790,n4791);
or (n4794,n4795,n4798);
and (n4795,n4796,n4797);
xor (n4796,n4730,n4731);
and (n4797,n659,n652);
and (n4798,n4799,n4800);
xor (n4799,n4796,n4797);
or (n4800,n4801,n4804);
and (n4801,n4802,n4803);
xor (n4802,n4736,n4737);
and (n4803,n319,n652);
and (n4804,n4805,n4806);
xor (n4805,n4802,n4803);
or (n4806,n4807,n4810);
and (n4807,n4808,n4809);
xor (n4808,n4742,n4743);
and (n4809,n311,n652);
and (n4810,n4811,n4812);
xor (n4811,n4808,n4809);
or (n4812,n4813,n4816);
and (n4813,n4814,n4815);
xor (n4814,n4748,n4749);
and (n4815,n352,n652);
and (n4816,n4817,n4818);
xor (n4817,n4814,n4815);
or (n4818,n4819,n4822);
and (n4819,n4820,n4821);
xor (n4820,n4754,n4755);
and (n4821,n344,n652);
and (n4822,n4823,n4824);
xor (n4823,n4820,n4821);
or (n4824,n4825,n4828);
and (n4825,n4826,n4827);
xor (n4826,n4760,n4761);
and (n4827,n386,n652);
and (n4828,n4829,n4830);
xor (n4829,n4826,n4827);
or (n4830,n4831,n4834);
and (n4831,n4832,n4833);
xor (n4832,n4766,n4767);
and (n4833,n378,n652);
and (n4834,n4835,n4836);
xor (n4835,n4832,n4833);
or (n4836,n4837,n4840);
and (n4837,n4838,n4839);
xor (n4838,n4772,n4773);
and (n4839,n502,n652);
and (n4840,n4841,n4842);
xor (n4841,n4838,n4839);
and (n4842,n4843,n4844);
xor (n4843,n4778,n4779);
and (n4844,n131,n652);
and (n4845,n625,n803);
or (n4846,n4847,n4850);
and (n4847,n4848,n4849);
xor (n4848,n4787,n4788);
and (n4849,n667,n803);
and (n4850,n4851,n4852);
xor (n4851,n4848,n4849);
or (n4852,n4853,n4856);
and (n4853,n4854,n4855);
xor (n4854,n4793,n4794);
and (n4855,n659,n803);
and (n4856,n4857,n4858);
xor (n4857,n4854,n4855);
or (n4858,n4859,n4862);
and (n4859,n4860,n4861);
xor (n4860,n4799,n4800);
and (n4861,n319,n803);
and (n4862,n4863,n4864);
xor (n4863,n4860,n4861);
or (n4864,n4865,n4868);
and (n4865,n4866,n4867);
xor (n4866,n4805,n4806);
and (n4867,n311,n803);
and (n4868,n4869,n4870);
xor (n4869,n4866,n4867);
or (n4870,n4871,n4874);
and (n4871,n4872,n4873);
xor (n4872,n4811,n4812);
and (n4873,n352,n803);
and (n4874,n4875,n4876);
xor (n4875,n4872,n4873);
or (n4876,n4877,n4880);
and (n4877,n4878,n4879);
xor (n4878,n4817,n4818);
and (n4879,n344,n803);
and (n4880,n4881,n4882);
xor (n4881,n4878,n4879);
or (n4882,n4883,n4886);
and (n4883,n4884,n4885);
xor (n4884,n4823,n4824);
and (n4885,n386,n803);
and (n4886,n4887,n4888);
xor (n4887,n4884,n4885);
or (n4888,n4889,n4892);
and (n4889,n4890,n4891);
xor (n4890,n4829,n4830);
and (n4891,n378,n803);
and (n4892,n4893,n4894);
xor (n4893,n4890,n4891);
or (n4894,n4895,n4898);
and (n4895,n4896,n4897);
xor (n4896,n4835,n4836);
and (n4897,n502,n803);
and (n4898,n4899,n4900);
xor (n4899,n4896,n4897);
and (n4900,n4901,n1716);
xor (n4901,n4841,n4842);
and (n4902,n667,n294);
or (n4903,n4904,n4907);
and (n4904,n4905,n4906);
xor (n4905,n4851,n4852);
and (n4906,n659,n294);
and (n4907,n4908,n4909);
xor (n4908,n4905,n4906);
or (n4909,n4910,n4913);
and (n4910,n4911,n4912);
xor (n4911,n4857,n4858);
and (n4912,n319,n294);
and (n4913,n4914,n4915);
xor (n4914,n4911,n4912);
or (n4915,n4916,n4919);
and (n4916,n4917,n4918);
xor (n4917,n4863,n4864);
and (n4918,n311,n294);
and (n4919,n4920,n4921);
xor (n4920,n4917,n4918);
or (n4921,n4922,n4925);
and (n4922,n4923,n4924);
xor (n4923,n4869,n4870);
and (n4924,n352,n294);
and (n4925,n4926,n4927);
xor (n4926,n4923,n4924);
or (n4927,n4928,n4931);
and (n4928,n4929,n4930);
xor (n4929,n4875,n4876);
and (n4930,n344,n294);
and (n4931,n4932,n4933);
xor (n4932,n4929,n4930);
or (n4933,n4934,n4937);
and (n4934,n4935,n4936);
xor (n4935,n4881,n4882);
and (n4936,n386,n294);
and (n4937,n4938,n4939);
xor (n4938,n4935,n4936);
or (n4939,n4940,n4943);
and (n4940,n4941,n4942);
xor (n4941,n4887,n4888);
and (n4942,n378,n294);
and (n4943,n4944,n4945);
xor (n4944,n4941,n4942);
or (n4945,n4946,n4949);
and (n4946,n4947,n4948);
xor (n4947,n4893,n4894);
and (n4948,n502,n294);
and (n4949,n4950,n4951);
xor (n4950,n4947,n4948);
and (n4951,n4952,n4953);
xor (n4952,n4899,n4900);
and (n4953,n131,n294);
and (n4954,n659,n297);
or (n4955,n4956,n4959);
and (n4956,n4957,n4958);
xor (n4957,n4908,n4909);
and (n4958,n319,n297);
and (n4959,n4960,n4961);
xor (n4960,n4957,n4958);
or (n4961,n4962,n4965);
and (n4962,n4963,n4964);
xor (n4963,n4914,n4915);
and (n4964,n311,n297);
and (n4965,n4966,n4967);
xor (n4966,n4963,n4964);
or (n4967,n4968,n4971);
and (n4968,n4969,n4970);
xor (n4969,n4920,n4921);
and (n4970,n352,n297);
and (n4971,n4972,n4973);
xor (n4972,n4969,n4970);
or (n4973,n4974,n4977);
and (n4974,n4975,n4976);
xor (n4975,n4926,n4927);
and (n4976,n344,n297);
and (n4977,n4978,n4979);
xor (n4978,n4975,n4976);
or (n4979,n4980,n4983);
and (n4980,n4981,n4982);
xor (n4981,n4932,n4933);
and (n4982,n386,n297);
and (n4983,n4984,n4985);
xor (n4984,n4981,n4982);
or (n4985,n4986,n4989);
and (n4986,n4987,n4988);
xor (n4987,n4938,n4939);
and (n4988,n378,n297);
and (n4989,n4990,n4991);
xor (n4990,n4987,n4988);
or (n4991,n4992,n4995);
and (n4992,n4993,n4994);
xor (n4993,n4944,n4945);
and (n4994,n502,n297);
and (n4995,n4996,n4997);
xor (n4996,n4993,n4994);
and (n4997,n4998,n1320);
xor (n4998,n4950,n4951);
and (n4999,n319,n304);
or (n5000,n5001,n5004);
and (n5001,n5002,n5003);
xor (n5002,n4960,n4961);
and (n5003,n311,n304);
and (n5004,n5005,n5006);
xor (n5005,n5002,n5003);
or (n5006,n5007,n5010);
and (n5007,n5008,n5009);
xor (n5008,n4966,n4967);
and (n5009,n352,n304);
and (n5010,n5011,n5012);
xor (n5011,n5008,n5009);
or (n5012,n5013,n5016);
and (n5013,n5014,n5015);
xor (n5014,n4972,n4973);
and (n5015,n344,n304);
and (n5016,n5017,n5018);
xor (n5017,n5014,n5015);
or (n5018,n5019,n5022);
and (n5019,n5020,n5021);
xor (n5020,n4978,n4979);
and (n5021,n386,n304);
and (n5022,n5023,n5024);
xor (n5023,n5020,n5021);
or (n5024,n5025,n5028);
and (n5025,n5026,n5027);
xor (n5026,n4984,n4985);
and (n5027,n378,n304);
and (n5028,n5029,n5030);
xor (n5029,n5026,n5027);
or (n5030,n5031,n5034);
and (n5031,n5032,n5033);
xor (n5032,n4990,n4991);
and (n5033,n502,n304);
and (n5034,n5035,n5036);
xor (n5035,n5032,n5033);
and (n5036,n5037,n5038);
xor (n5037,n4996,n4997);
and (n5038,n131,n304);
and (n5039,n311,n331);
or (n5040,n5041,n5044);
and (n5041,n5042,n5043);
xor (n5042,n5005,n5006);
and (n5043,n352,n331);
and (n5044,n5045,n5046);
xor (n5045,n5042,n5043);
or (n5046,n5047,n5050);
and (n5047,n5048,n5049);
xor (n5048,n5011,n5012);
and (n5049,n344,n331);
and (n5050,n5051,n5052);
xor (n5051,n5048,n5049);
or (n5052,n5053,n5056);
and (n5053,n5054,n5055);
xor (n5054,n5017,n5018);
and (n5055,n386,n331);
and (n5056,n5057,n5058);
xor (n5057,n5054,n5055);
or (n5058,n5059,n5062);
and (n5059,n5060,n5061);
xor (n5060,n5023,n5024);
and (n5061,n378,n331);
and (n5062,n5063,n5064);
xor (n5063,n5060,n5061);
or (n5064,n5065,n5068);
and (n5065,n5066,n5067);
xor (n5066,n5029,n5030);
and (n5067,n502,n331);
and (n5068,n5069,n5070);
xor (n5069,n5066,n5067);
and (n5070,n5071,n1180);
xor (n5071,n5035,n5036);
and (n5072,n352,n338);
or (n5073,n5074,n5077);
and (n5074,n5075,n5076);
xor (n5075,n5045,n5046);
and (n5076,n344,n338);
and (n5077,n5078,n5079);
xor (n5078,n5075,n5076);
or (n5079,n5080,n5083);
and (n5080,n5081,n5082);
xor (n5081,n5051,n5052);
and (n5082,n386,n338);
and (n5083,n5084,n5085);
xor (n5084,n5081,n5082);
or (n5085,n5086,n5089);
and (n5086,n5087,n5088);
xor (n5087,n5057,n5058);
and (n5088,n378,n338);
and (n5089,n5090,n5091);
xor (n5090,n5087,n5088);
or (n5091,n5092,n5095);
and (n5092,n5093,n5094);
xor (n5093,n5063,n5064);
and (n5094,n502,n338);
and (n5095,n5096,n5097);
xor (n5096,n5093,n5094);
and (n5097,n5098,n5099);
xor (n5098,n5069,n5070);
and (n5099,n131,n338);
and (n5100,n344,n363);
or (n5101,n5102,n5105);
and (n5102,n5103,n5104);
xor (n5103,n5078,n5079);
and (n5104,n386,n363);
and (n5105,n5106,n5107);
xor (n5106,n5103,n5104);
or (n5107,n5108,n5111);
and (n5108,n5109,n5110);
xor (n5109,n5084,n5085);
and (n5110,n378,n363);
and (n5111,n5112,n5113);
xor (n5112,n5109,n5110);
or (n5113,n5114,n5117);
and (n5114,n5115,n5116);
xor (n5115,n5090,n5091);
and (n5116,n502,n363);
and (n5117,n5118,n5119);
xor (n5118,n5115,n5116);
and (n5119,n5120,n513);
xor (n5120,n5096,n5097);
and (n5121,n386,n367);
or (n5122,n5123,n5126);
and (n5123,n5124,n5125);
xor (n5124,n5106,n5107);
and (n5125,n378,n367);
and (n5126,n5127,n5128);
xor (n5127,n5124,n5125);
or (n5128,n5129,n5132);
and (n5129,n5130,n5131);
xor (n5130,n5112,n5113);
and (n5131,n502,n367);
and (n5132,n5133,n5134);
xor (n5133,n5130,n5131);
and (n5134,n5135,n5136);
xor (n5135,n5118,n5119);
and (n5136,n131,n367);
and (n5137,n378,n532);
or (n5138,n5139,n5142);
and (n5139,n5140,n5141);
xor (n5140,n5127,n5128);
and (n5141,n502,n532);
and (n5142,n5143,n5144);
xor (n5143,n5140,n5141);
and (n5144,n5145,n552);
xor (n5145,n5133,n5134);
and (n5146,n502,n17);
and (n5147,n5148,n5149);
xor (n5148,n5143,n5144);
and (n5149,n131,n17);
and (n5150,n131,n122);
endmodule
