module top (out,n24,n27,n28,n29,n37,n38,n44,n45,n50
        ,n58,n60,n61,n70,n71,n81,n96,n97,n100,n106
        ,n128,n129,n136,n246,n247,n255,n295,n302,n306,n370
        ,n376,n382,n388,n393,n431,n451,n457,n464,n470,n619
        ,n631,n646,n657,n699,n727);
output out;
input n24;
input n27;
input n28;
input n29;
input n37;
input n38;
input n44;
input n45;
input n50;
input n58;
input n60;
input n61;
input n70;
input n71;
input n81;
input n96;
input n97;
input n100;
input n106;
input n128;
input n129;
input n136;
input n246;
input n247;
input n255;
input n295;
input n302;
input n306;
input n370;
input n376;
input n382;
input n388;
input n393;
input n431;
input n451;
input n457;
input n464;
input n470;
input n619;
input n631;
input n646;
input n657;
input n699;
input n727;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n25;
wire n26;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n46;
wire n47;
wire n48;
wire n49;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n59;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n98;
wire n99;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n303;
wire n304;
wire n305;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n367;
wire n368;
wire n369;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n389;
wire n390;
wire n391;
wire n392;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
xor (out,n0,n740);
nand (n0,n1,n728,n739);
or (n1,n2,n658);
nand (n2,n3,n402,n632);
not (n3,n4);
not (n4,n5);
or (n5,n6,n296,n401);
not (n6,n7);
nand (n7,n8,n295);
and (n8,n9,n294);
nand (n9,n10,n293);
or (n10,n11,n233);
not (n11,n12);
or (n12,n13,n232);
and (n13,n14,n148);
xor (n14,n15,n111);
or (n15,n16,n110);
and (n16,n17,n84);
xor (n17,n18,n53);
nand (n18,n19,n47);
or (n19,n20,n31);
not (n20,n21);
nor (n21,n22,n30);
and (n22,n23,n25);
not (n23,n24);
not (n25,n26);
wire s0n26,s1n26,notn26;
or (n26,s0n26,s1n26);
not(notn26,n29);
and (s0n26,notn26,n27);
and (s1n26,n29,n28);
and (n30,n24,n26);
not (n31,n32);
and (n32,n33,n40);
nand (n33,n34,n39);
or (n34,n35,n26);
not (n35,n36);
wire s0n36,s1n36,notn36;
or (n36,s0n36,s1n36);
not(notn36,n29);
and (s0n36,notn36,n37);
and (s1n36,n29,n38);
nand (n39,n26,n35);
not (n40,n41);
nand (n41,n42,n46);
or (n42,n35,n43);
wire s0n43,s1n43,notn43;
or (n43,s0n43,s1n43);
not(notn43,n29);
and (s0n43,notn43,n44);
and (s1n43,n29,n45);
nand (n46,n43,n35);
nand (n47,n41,n48);
nor (n48,n49,n51);
and (n49,n50,n26);
and (n51,n25,n52);
not (n52,n50);
nand (n53,n54,n73);
or (n54,n55,n65);
not (n55,n56);
nor (n56,n57,n62);
and (n57,n58,n59);
wire s0n59,s1n59,notn59;
or (n59,s0n59,s1n59);
not(notn59,n29);
and (s0n59,notn59,n60);
and (s1n59,n29,n61);
and (n62,n63,n64);
not (n63,n58);
not (n64,n59);
not (n65,n66);
nand (n66,n67,n72);
or (n67,n68,n26);
not (n68,n69);
wire s0n69,s1n69,notn69;
or (n69,s0n69,s1n69);
not(notn69,n29);
and (s0n69,notn69,n70);
and (s1n69,n29,n71);
nand (n72,n26,n68);
nand (n73,n74,n79);
not (n74,n75);
nand (n75,n65,n76);
nand (n76,n77,n78);
or (n77,n68,n59);
nand (n78,n59,n68);
nand (n79,n80,n82);
or (n80,n64,n81);
or (n82,n59,n83);
not (n83,n81);
xor (n84,n85,n90);
and (n85,n86,n59);
nand (n86,n87,n89);
or (n87,n26,n88);
and (n88,n81,n69);
or (n89,n69,n81);
nand (n90,n91,n103);
or (n91,n92,n98);
not (n92,n93);
nor (n93,n94,n95);
not (n94,n43);
wire s0n95,s1n95,notn95;
or (n95,s0n95,s1n95);
not(notn95,n29);
and (s0n95,notn95,n96);
and (s1n95,n29,n97);
nor (n98,n99,n101);
and (n99,n94,n100);
and (n101,n43,n102);
not (n102,n100);
or (n103,n104,n109);
nor (n104,n105,n107);
and (n105,n106,n94);
and (n107,n108,n43);
not (n108,n106);
not (n109,n95);
and (n110,n18,n53);
xor (n111,n112,n120);
xor (n112,n113,n119);
nand (n113,n114,n115);
or (n114,n55,n75);
or (n115,n65,n116);
nor (n116,n117,n118);
and (n117,n64,n24);
and (n118,n59,n23);
and (n119,n85,n90);
xor (n120,n121,n141);
xor (n121,n122,n131);
and (n122,n123,n81);
not (n123,n124);
nor (n124,n125,n130);
and (n125,n126,n59);
not (n126,n127);
wire s0n127,s1n127,notn127;
or (n127,s0n127,s1n127);
not(notn127,n29);
and (s0n127,notn127,n128);
and (s1n127,n29,n129);
and (n130,n127,n64);
nand (n131,n132,n139);
or (n132,n109,n133);
not (n133,n134);
nor (n134,n135,n137);
and (n135,n136,n43);
and (n137,n138,n94);
not (n138,n136);
nand (n139,n140,n93);
not (n140,n104);
nand (n141,n142,n144);
or (n142,n143,n31);
not (n143,n48);
nand (n144,n41,n145);
nand (n145,n146,n147);
or (n146,n26,n102);
or (n147,n25,n100);
or (n148,n149,n231);
and (n149,n150,n171);
xor (n150,n151,n170);
or (n151,n152,n169);
and (n152,n153,n162);
xor (n153,n154,n155);
and (n154,n66,n81);
nand (n155,n156,n161);
or (n156,n157,n31);
not (n157,n158);
nor (n158,n159,n160);
and (n159,n58,n26);
and (n160,n63,n25);
nand (n161,n21,n41);
nand (n162,n163,n168);
or (n163,n92,n164);
not (n164,n165);
nor (n165,n166,n167);
and (n166,n52,n94);
and (n167,n50,n43);
or (n168,n98,n109);
and (n169,n154,n155);
xor (n170,n17,n84);
or (n171,n172,n230);
and (n172,n173,n229);
xor (n173,n174,n188);
nor (n174,n175,n183);
not (n175,n176);
nand (n176,n177,n182);
or (n177,n178,n92);
not (n178,n179);
nand (n179,n180,n181);
or (n180,n23,n43);
nand (n181,n43,n23);
nand (n182,n165,n95);
nand (n183,n184,n26);
nand (n184,n185,n187);
or (n185,n43,n186);
and (n186,n81,n36);
or (n187,n36,n81);
nand (n188,n189,n227);
or (n189,n190,n213);
not (n190,n191);
nand (n191,n192,n212);
or (n192,n193,n202);
nor (n193,n194,n201);
nand (n194,n195,n200);
or (n195,n196,n92);
not (n196,n197);
nand (n197,n198,n199);
or (n198,n63,n43);
nand (n199,n43,n63);
nand (n200,n179,n95);
nor (n201,n40,n83);
nand (n202,n203,n210);
nand (n203,n204,n209);
or (n204,n205,n92);
not (n205,n206);
nand (n206,n207,n208);
or (n207,n94,n81);
or (n208,n43,n83);
nand (n209,n197,n95);
nor (n210,n211,n94);
and (n211,n81,n95);
nand (n212,n194,n201);
not (n213,n214);
nand (n214,n215,n223);
not (n215,n216);
nand (n216,n217,n222);
or (n217,n218,n31);
not (n218,n219);
nand (n219,n220,n221);
or (n220,n25,n81);
or (n221,n26,n83);
nand (n222,n41,n158);
nor (n223,n224,n226);
and (n224,n175,n225);
not (n225,n183);
and (n226,n176,n183);
nand (n227,n228,n216);
not (n228,n223);
xor (n229,n153,n162);
and (n230,n174,n188);
and (n231,n151,n170);
and (n232,n15,n111);
not (n233,n234);
nand (n234,n235,n292);
or (n235,n236,n289);
xor (n236,n237,n260);
xor (n237,n238,n257);
xor (n238,n239,n248);
nor (n239,n240,n244);
nor (n240,n241,n243);
and (n241,n64,n242);
nand (n242,n127,n81);
and (n243,n126,n83);
not (n244,n245);
wire s0n245,s1n245,notn245;
or (n245,s0n245,s1n245);
not(notn245,n29);
and (s0n245,notn245,n246);
and (s1n245,n29,n247);
nand (n248,n249,n250);
or (n249,n133,n92);
nand (n250,n251,n95);
not (n251,n252);
nor (n252,n253,n256);
and (n253,n254,n43);
not (n254,n255);
and (n256,n255,n94);
or (n257,n258,n259);
and (n258,n121,n141);
and (n259,n122,n131);
xor (n260,n261,n283);
xor (n261,n262,n276);
nand (n262,n263,n272);
or (n263,n264,n268);
not (n264,n265);
nand (n265,n266,n267);
or (n266,n244,n81);
or (n267,n245,n83);
nand (n268,n124,n269);
nand (n269,n270,n271);
or (n270,n126,n245);
nand (n271,n245,n126);
or (n272,n124,n273);
nor (n273,n274,n275);
and (n274,n58,n244);
and (n275,n63,n245);
nand (n276,n277,n279);
or (n277,n278,n31);
not (n278,n145);
nand (n279,n41,n280);
nor (n280,n281,n282);
and (n281,n106,n26);
and (n282,n108,n25);
nand (n283,n284,n285);
or (n284,n75,n116);
or (n285,n65,n286);
nor (n286,n287,n288);
and (n287,n64,n50);
and (n288,n59,n52);
or (n289,n290,n291);
and (n290,n112,n120);
and (n291,n113,n119);
nand (n292,n236,n289);
or (n293,n234,n12);
not (n294,n29);
and (n296,n8,n297);
or (n297,n298,n303,n400);
not (n298,n299);
nand (n299,n300,n302);
and (n300,n301,n294);
xor (n301,n14,n148);
and (n303,n300,n304);
or (n304,n305,n367,n399);
and (n305,n306,n307);
wire s0n307,s1n307,notn307;
or (n307,s0n307,s1n307);
not(notn307,n29);
and (s0n307,notn307,n308);
and (s1n307,n29,1'b0);
xor (n308,n309,n365);
xor (n309,n310,n363);
xor (n310,n311,n362);
xor (n311,n312,n354);
xor (n312,n313,n30);
xor (n313,n314,n340);
xor (n314,n315,n339);
xor (n315,n316,n319);
xor (n316,n317,n318);
and (n317,n106,n95);
and (n318,n100,n43);
or (n319,n320,n322);
and (n320,n321,n167);
and (n321,n100,n95);
and (n322,n323,n324);
xor (n323,n321,n167);
or (n324,n325,n328);
and (n325,n326,n327);
and (n326,n50,n95);
and (n327,n24,n43);
and (n328,n329,n330);
xor (n329,n326,n327);
or (n330,n331,n334);
and (n331,n332,n333);
and (n332,n24,n95);
and (n333,n58,n43);
and (n334,n335,n336);
xor (n335,n332,n333);
and (n336,n337,n338);
and (n337,n58,n95);
and (n338,n81,n43);
and (n339,n50,n36);
or (n340,n341,n344);
and (n341,n342,n343);
xor (n342,n323,n324);
and (n343,n24,n36);
and (n344,n345,n346);
xor (n345,n342,n343);
or (n346,n347,n350);
and (n347,n348,n349);
xor (n348,n329,n330);
and (n349,n58,n36);
and (n350,n351,n352);
xor (n351,n348,n349);
and (n352,n353,n186);
xor (n353,n335,n336);
or (n354,n355,n357);
and (n355,n356,n159);
xor (n356,n345,n346);
and (n357,n358,n359);
xor (n358,n356,n159);
and (n359,n360,n361);
xor (n360,n351,n352);
and (n361,n81,n26);
and (n362,n58,n69);
and (n363,n364,n88);
xor (n364,n358,n359);
and (n365,n81,n59);
and (n367,n307,n368);
or (n368,n369,n373,n398);
and (n369,n370,n371);
wire s0n371,s1n371,notn371;
or (n371,s0n371,s1n371);
not(notn371,n29);
and (s0n371,notn371,n372);
and (s1n371,n29,1'b0);
xor (n372,n364,n88);
and (n373,n371,n374);
or (n374,n375,n379,n397);
and (n375,n376,n377);
wire s0n377,s1n377,notn377;
or (n377,s0n377,s1n377);
not(notn377,n29);
and (s0n377,notn377,n378);
and (s1n377,n29,1'b0);
xor (n378,n360,n361);
and (n379,n377,n380);
or (n380,n381,n385,n396);
and (n381,n382,n383);
wire s0n383,s1n383,notn383;
or (n383,s0n383,s1n383);
not(notn383,n29);
and (s0n383,notn383,n384);
and (s1n383,n29,1'b0);
xor (n384,n353,n186);
and (n385,n383,n386);
or (n386,n387,n391,n395);
and (n387,n388,n389);
wire s0n389,s1n389,notn389;
or (n389,s0n389,s1n389);
not(notn389,n29);
and (s0n389,notn389,n390);
and (s1n389,n29,1'b0);
xor (n390,n337,n338);
and (n391,n389,n392);
and (n392,n393,n394);
wire s0n394,s1n394,notn394;
or (n394,s0n394,s1n394);
not(notn394,n29);
and (s0n394,notn394,n211);
and (s1n394,n29,1'b0);
and (n395,n388,n392);
and (n396,n382,n386);
and (n397,n376,n380);
and (n398,n370,n374);
and (n399,n306,n368);
and (n400,n302,n304);
and (n401,n295,n297);
nor (n402,n403,n620);
nor (n403,n404,n619);
nand (n404,n405,n407);
or (n405,n294,n406);
not (n406,n378);
nand (n407,n408,n294);
xnor (n408,n409,n565);
nand (n409,n410,n564);
nand (n410,n411,n529);
not (n411,n412);
xor (n412,n413,n507);
xor (n413,n414,n444);
xor (n414,n415,n435);
xor (n415,n416,n426);
nand (n416,n417,n422);
or (n417,n418,n268);
not (n418,n419);
nor (n419,n420,n421);
and (n420,n100,n245);
and (n421,n102,n244);
nand (n422,n123,n423);
nor (n423,n424,n425);
and (n424,n106,n245);
and (n425,n108,n244);
nor (n426,n427,n432);
nand (n427,n245,n428);
not (n428,n429);
wire s0n429,s1n429,notn429;
or (n429,s0n429,s1n429);
not(notn429,n29);
and (s0n429,notn429,1'b0);
and (s1n429,n29,n430);
and (n430,n431,n247);
nor (n432,n433,n434);
and (n433,n429,n52);
and (n434,n428,n50);
nand (n435,n436,n440);
or (n436,n75,n437);
nor (n437,n438,n439);
and (n438,n64,n136);
and (n439,n59,n138);
or (n440,n65,n441);
nor (n441,n442,n443);
and (n442,n64,n255);
and (n443,n59,n254);
xor (n444,n445,n486);
xor (n445,n446,n473);
xor (n446,n447,n460);
nand (n447,n448,n454);
or (n448,n92,n449);
nor (n449,n450,n452);
and (n450,n94,n451);
and (n452,n43,n453);
not (n453,n451);
or (n454,n455,n109);
nor (n455,n456,n458);
and (n456,n94,n457);
and (n458,n43,n459);
not (n459,n457);
nand (n460,n461,n467);
or (n461,n31,n462);
nor (n462,n463,n465);
and (n463,n25,n464);
and (n465,n26,n466);
not (n466,n464);
or (n467,n40,n468);
nor (n468,n469,n471);
and (n469,n25,n470);
and (n471,n26,n472);
not (n472,n470);
and (n473,n474,n480);
nand (n474,n475,n479);
or (n475,n92,n476);
nor (n476,n477,n478);
and (n477,n94,n470);
and (n478,n43,n472);
or (n479,n449,n109);
nand (n480,n481,n485);
or (n481,n31,n482);
nor (n482,n483,n484);
and (n483,n25,n255);
and (n484,n26,n254);
or (n485,n462,n40);
or (n486,n487,n506);
and (n487,n488,n500);
xor (n488,n489,n496);
nand (n489,n490,n495);
or (n490,n491,n268);
not (n491,n492);
nor (n492,n493,n494);
and (n493,n50,n245);
and (n494,n52,n244);
nand (n495,n123,n419);
nor (n496,n427,n497);
nor (n497,n498,n499);
and (n498,n429,n23);
and (n499,n428,n24);
nand (n500,n501,n505);
or (n501,n75,n502);
nor (n502,n503,n504);
and (n503,n64,n106);
and (n504,n59,n108);
or (n505,n65,n437);
and (n506,n489,n496);
and (n507,n508,n509);
xor (n508,n474,n480);
or (n509,n510,n528);
and (n510,n511,n522);
xor (n511,n512,n518);
nand (n512,n513,n517);
or (n513,n514,n268);
nor (n514,n515,n516);
and (n515,n24,n244);
and (n516,n23,n245);
nand (n517,n492,n123);
nor (n518,n427,n519);
nor (n519,n520,n521);
and (n520,n429,n63);
and (n521,n428,n58);
nand (n522,n523,n527);
or (n523,n92,n524);
nor (n524,n525,n526);
and (n525,n94,n464);
and (n526,n43,n466);
or (n527,n476,n109);
and (n528,n512,n518);
not (n529,n530);
or (n530,n531,n563);
and (n531,n532,n535);
xor (n532,n533,n534);
xor (n533,n488,n500);
xor (n534,n508,n509);
or (n535,n536,n562);
and (n536,n537,n550);
xor (n537,n538,n544);
nand (n538,n539,n543);
or (n539,n75,n540);
nor (n540,n541,n542);
and (n541,n64,n100);
and (n542,n59,n102);
or (n543,n65,n502);
nand (n544,n545,n549);
or (n545,n31,n546);
nor (n546,n547,n548);
and (n547,n25,n136);
and (n548,n26,n138);
or (n549,n482,n40);
or (n550,n551,n561);
and (n551,n552,n558);
xor (n552,n553,n555);
and (n553,n554,n81);
not (n554,n427);
nand (n555,n556,n557);
or (n556,n92,n252);
or (n557,n524,n109);
nand (n558,n559,n560);
or (n559,n268,n273);
or (n560,n124,n514);
and (n561,n553,n555);
and (n562,n538,n544);
and (n563,n533,n534);
nand (n564,n412,n530);
nand (n565,n566,n618);
or (n566,n567,n587);
nor (n567,n568,n569);
xor (n568,n532,n535);
or (n569,n570,n586);
and (n570,n571,n585);
xor (n571,n572,n573);
xor (n572,n511,n522);
or (n573,n574,n584);
and (n574,n575,n583);
xor (n575,n576,n580);
nand (n576,n577,n579);
or (n577,n31,n578);
not (n578,n280);
or (n579,n40,n546);
nand (n580,n581,n582);
or (n581,n75,n286);
or (n582,n65,n540);
and (n583,n239,n248);
and (n584,n576,n580);
xor (n585,n537,n550);
and (n586,n572,n573);
not (n587,n588);
nand (n588,n589,n613);
not (n589,n590);
nor (n590,n591,n594);
nor (n591,n592,n593);
and (n592,n12,n235);
not (n593,n292);
nand (n594,n595,n607);
not (n595,n596);
nor (n596,n597,n604);
xor (n597,n598,n603);
xor (n598,n599,n602);
or (n599,n600,n601);
and (n600,n261,n283);
and (n601,n262,n276);
xor (n602,n552,n558);
xor (n603,n575,n583);
or (n604,n605,n606);
and (n605,n237,n260);
and (n606,n238,n257);
not (n607,n608);
nor (n608,n609,n612);
or (n609,n610,n611);
and (n610,n598,n603);
and (n611,n599,n602);
xor (n612,n571,n585);
nor (n613,n614,n617);
and (n614,n607,n615);
not (n615,n616);
nand (n616,n597,n604);
and (n617,n609,n612);
nand (n618,n568,n569);
nor (n620,n621,n631);
nand (n621,n622,n624);
or (n622,n294,n623);
not (n623,n384);
nand (n624,n625,n294);
nand (n625,n626,n630);
or (n626,n627,n587);
not (n627,n628);
nand (n628,n629,n618);
not (n629,n567);
or (n630,n588,n628);
nor (n632,n633,n647);
nor (n633,n634,n646);
nand (n634,n635,n637);
or (n635,n294,n636);
not (n636,n390);
nand (n637,n638,n294);
nand (n638,n639,n645);
or (n639,n640,n642);
not (n640,n641);
or (n641,n617,n608);
not (n642,n643);
nand (n643,n644,n616);
or (n644,n591,n596);
or (n645,n643,n641);
nor (n647,n648,n657);
or (n648,n649,n650);
and (n649,n29,n211);
and (n650,n294,n651);
nand (n651,n652,n656);
or (n652,n653,n654);
not (n653,n591);
not (n654,n655);
nor (n655,n615,n596);
or (n656,n655,n591);
nor (n658,n659,n727);
nand (n659,n660,n662);
or (n660,n294,n661);
not (n661,n372);
nand (n662,n663,n294);
nand (n663,n664,n726);
or (n664,n665,n720);
not (n665,n666);
nand (n666,n667,n719);
nand (n667,n668,n715);
not (n668,n669);
xor (n669,n670,n712);
xor (n670,n671,n691);
xor (n671,n672,n685);
xor (n672,n673,n681);
nand (n673,n674,n676);
or (n674,n675,n268);
not (n675,n423);
nand (n676,n677,n123);
not (n677,n678);
nor (n678,n679,n680);
and (n679,n244,n136);
and (n680,n245,n138);
nor (n681,n427,n682);
nor (n682,n683,n684);
and (n683,n429,n102);
and (n684,n428,n100);
nand (n685,n686,n687);
or (n686,n75,n441);
or (n687,n65,n688);
nor (n688,n689,n690);
and (n689,n64,n464);
and (n690,n59,n466);
xor (n691,n692,n709);
xor (n692,n693,n708);
xor (n693,n694,n702);
nand (n694,n695,n696);
or (n695,n92,n455);
or (n696,n697,n109);
nor (n697,n698,n700);
and (n698,n94,n699);
and (n700,n43,n701);
not (n701,n699);
nand (n702,n703,n704);
or (n703,n31,n468);
or (n704,n705,n40);
nor (n705,n706,n707);
and (n706,n25,n451);
and (n707,n26,n453);
and (n708,n447,n460);
or (n709,n710,n711);
and (n710,n415,n435);
and (n711,n416,n426);
or (n712,n713,n714);
and (n713,n445,n486);
and (n714,n446,n473);
not (n715,n716);
or (n716,n717,n718);
and (n717,n413,n507);
and (n718,n414,n444);
nand (n719,n669,n716);
not (n720,n721);
nand (n721,n722,n725,n564);
nand (n722,n723,n410);
nand (n723,n724,n618);
or (n724,n613,n567);
nand (n725,n410,n590,n629);
or (n726,n721,n666);
or (n728,n658,n729);
nor (n729,n730,n735);
and (n730,n402,n731);
nand (n731,n732,n734);
or (n732,n633,n733);
nand (n733,n648,n657);
nand (n734,n634,n646);
nand (n735,n736,n738);
or (n736,n403,n737);
nand (n737,n621,n631);
nand (n738,n404,n619);
nand (n739,n659,n727);
or (n740,n741,n1063,n1088);
and (n741,n727,n742);
wire s0n742,s1n742,notn742;
or (n742,s0n742,s1n742);
not(notn742,n29);
and (s0n742,notn742,n743);
and (s1n742,n29,n372);
xor (n743,n744,n1041);
xor (n744,n745,n1061);
xor (n745,n746,n1036);
xor (n746,n747,n1054);
xor (n747,n748,n1030);
xor (n748,n749,n1042);
xor (n749,n750,n1024);
xor (n750,n751,n1021);
xor (n751,n752,n1020);
xor (n752,n753,n995);
xor (n753,n754,n424);
xor (n754,n755,n962);
xor (n755,n756,n961);
xor (n756,n757,n925);
xor (n757,n758,n924);
xor (n758,n759,n885);
xor (n759,n760,n884);
xor (n760,n761,n847);
xor (n761,n762,n846);
xor (n762,n763,n807);
xor (n763,n764,n806);
xor (n764,n765,n768);
xor (n765,n766,n767);
and (n766,n699,n95);
and (n767,n457,n43);
or (n768,n769,n772);
and (n769,n770,n771);
and (n770,n457,n95);
and (n771,n451,n43);
and (n772,n773,n774);
xor (n773,n770,n771);
or (n774,n775,n778);
and (n775,n776,n777);
and (n776,n451,n95);
and (n777,n470,n43);
and (n778,n779,n780);
xor (n779,n776,n777);
or (n780,n781,n784);
and (n781,n782,n783);
and (n782,n470,n95);
and (n783,n464,n43);
and (n784,n785,n786);
xor (n785,n782,n783);
or (n786,n787,n790);
and (n787,n788,n789);
and (n788,n464,n95);
and (n789,n255,n43);
and (n790,n791,n792);
xor (n791,n788,n789);
or (n792,n793,n795);
and (n793,n794,n135);
and (n794,n255,n95);
and (n795,n796,n797);
xor (n796,n794,n135);
or (n797,n798,n801);
and (n798,n799,n800);
and (n799,n136,n95);
and (n800,n106,n43);
and (n801,n802,n803);
xor (n802,n799,n800);
or (n803,n804,n805);
and (n804,n317,n318);
and (n805,n316,n319);
and (n806,n451,n36);
or (n807,n808,n811);
and (n808,n809,n810);
xor (n809,n773,n774);
and (n810,n470,n36);
and (n811,n812,n813);
xor (n812,n809,n810);
or (n813,n814,n817);
and (n814,n815,n816);
xor (n815,n779,n780);
and (n816,n464,n36);
and (n817,n818,n819);
xor (n818,n815,n816);
or (n819,n820,n823);
and (n820,n821,n822);
xor (n821,n785,n786);
and (n822,n255,n36);
and (n823,n824,n825);
xor (n824,n821,n822);
or (n825,n826,n829);
and (n826,n827,n828);
xor (n827,n791,n792);
and (n828,n136,n36);
and (n829,n830,n831);
xor (n830,n827,n828);
or (n831,n832,n835);
and (n832,n833,n834);
xor (n833,n796,n797);
and (n834,n106,n36);
and (n835,n836,n837);
xor (n836,n833,n834);
or (n837,n838,n841);
and (n838,n839,n840);
xor (n839,n802,n803);
and (n840,n100,n36);
and (n841,n842,n843);
xor (n842,n839,n840);
or (n843,n844,n845);
and (n844,n315,n339);
and (n845,n314,n340);
and (n846,n470,n26);
or (n847,n848,n851);
and (n848,n849,n850);
xor (n849,n812,n813);
and (n850,n464,n26);
and (n851,n852,n853);
xor (n852,n849,n850);
or (n853,n854,n857);
and (n854,n855,n856);
xor (n855,n818,n819);
and (n856,n255,n26);
and (n857,n858,n859);
xor (n858,n855,n856);
or (n859,n860,n863);
and (n860,n861,n862);
xor (n861,n824,n825);
and (n862,n136,n26);
and (n863,n864,n865);
xor (n864,n861,n862);
or (n865,n866,n868);
and (n866,n867,n281);
xor (n867,n830,n831);
and (n868,n869,n870);
xor (n869,n867,n281);
or (n870,n871,n874);
and (n871,n872,n873);
xor (n872,n836,n837);
and (n873,n100,n26);
and (n874,n875,n876);
xor (n875,n872,n873);
or (n876,n877,n879);
and (n877,n878,n49);
xor (n878,n842,n843);
and (n879,n880,n881);
xor (n880,n878,n49);
or (n881,n882,n883);
and (n882,n313,n30);
and (n883,n312,n354);
and (n884,n464,n69);
or (n885,n886,n889);
and (n886,n887,n888);
xor (n887,n852,n853);
and (n888,n255,n69);
and (n889,n890,n891);
xor (n890,n887,n888);
or (n891,n892,n895);
and (n892,n893,n894);
xor (n893,n858,n859);
and (n894,n136,n69);
and (n895,n896,n897);
xor (n896,n893,n894);
or (n897,n898,n901);
and (n898,n899,n900);
xor (n899,n864,n865);
and (n900,n106,n69);
and (n901,n902,n903);
xor (n902,n899,n900);
or (n903,n904,n907);
and (n904,n905,n906);
xor (n905,n869,n870);
and (n906,n100,n69);
and (n907,n908,n909);
xor (n908,n905,n906);
or (n909,n910,n913);
and (n910,n911,n912);
xor (n911,n875,n876);
and (n912,n50,n69);
and (n913,n914,n915);
xor (n914,n911,n912);
or (n915,n916,n919);
and (n916,n917,n918);
xor (n917,n880,n881);
and (n918,n24,n69);
and (n919,n920,n921);
xor (n920,n917,n918);
or (n921,n922,n923);
and (n922,n311,n362);
and (n923,n310,n363);
and (n924,n255,n59);
or (n925,n926,n929);
and (n926,n927,n928);
xor (n927,n890,n891);
and (n928,n136,n59);
and (n929,n930,n931);
xor (n930,n927,n928);
or (n931,n932,n935);
and (n932,n933,n934);
xor (n933,n896,n897);
and (n934,n106,n59);
and (n935,n936,n937);
xor (n936,n933,n934);
or (n937,n938,n941);
and (n938,n939,n940);
xor (n939,n902,n903);
and (n940,n100,n59);
and (n941,n942,n943);
xor (n942,n939,n940);
or (n943,n944,n947);
and (n944,n945,n946);
xor (n945,n908,n909);
and (n946,n50,n59);
and (n947,n948,n949);
xor (n948,n945,n946);
or (n949,n950,n953);
and (n950,n951,n952);
xor (n951,n914,n915);
and (n952,n24,n59);
and (n953,n954,n955);
xor (n954,n951,n952);
or (n955,n956,n958);
and (n956,n957,n57);
xor (n957,n920,n921);
and (n958,n959,n960);
xor (n959,n957,n57);
and (n960,n309,n365);
and (n961,n136,n127);
or (n962,n963,n966);
and (n963,n964,n965);
xor (n964,n930,n931);
and (n965,n106,n127);
and (n966,n967,n968);
xor (n967,n964,n965);
or (n968,n969,n972);
and (n969,n970,n971);
xor (n970,n936,n937);
and (n971,n100,n127);
and (n972,n973,n974);
xor (n973,n970,n971);
or (n974,n975,n978);
and (n975,n976,n977);
xor (n976,n942,n943);
and (n977,n50,n127);
and (n978,n979,n980);
xor (n979,n976,n977);
or (n980,n981,n984);
and (n981,n982,n983);
xor (n982,n948,n949);
and (n983,n24,n127);
and (n984,n985,n986);
xor (n985,n982,n983);
or (n986,n987,n990);
and (n987,n988,n989);
xor (n988,n954,n955);
and (n989,n58,n127);
and (n990,n991,n992);
xor (n991,n988,n989);
and (n992,n993,n994);
xor (n993,n959,n960);
not (n994,n242);
or (n995,n996,n998);
and (n996,n997,n420);
xor (n997,n967,n968);
and (n998,n999,n1000);
xor (n999,n997,n420);
or (n1000,n1001,n1003);
and (n1001,n1002,n493);
xor (n1002,n973,n974);
and (n1003,n1004,n1005);
xor (n1004,n1002,n493);
or (n1005,n1006,n1009);
and (n1006,n1007,n1008);
xor (n1007,n979,n980);
and (n1008,n24,n245);
and (n1009,n1010,n1011);
xor (n1010,n1007,n1008);
or (n1011,n1012,n1015);
and (n1012,n1013,n1014);
xor (n1013,n985,n986);
and (n1014,n58,n245);
and (n1015,n1016,n1017);
xor (n1016,n1013,n1014);
and (n1017,n1018,n1019);
xor (n1018,n991,n992);
and (n1019,n81,n245);
and (n1020,n100,n429);
or (n1021,n1022,n1025);
and (n1022,n1023,n1024);
xor (n1023,n999,n1000);
and (n1024,n50,n429);
and (n1025,n1026,n1027);
xor (n1026,n1023,n1024);
or (n1027,n1028,n1031);
and (n1028,n1029,n1030);
xor (n1029,n1004,n1005);
and (n1030,n24,n429);
and (n1031,n1032,n1033);
xor (n1032,n1029,n1030);
or (n1033,n1034,n1037);
and (n1034,n1035,n1036);
xor (n1035,n1010,n1011);
and (n1036,n58,n429);
and (n1037,n1038,n1039);
xor (n1038,n1035,n1036);
and (n1039,n1040,n1041);
xor (n1040,n1016,n1017);
and (n1041,n81,n429);
or (n1042,n1043,n1045);
and (n1043,n1044,n1030);
xor (n1044,n1026,n1027);
and (n1045,n1046,n1047);
xor (n1046,n1044,n1030);
or (n1047,n1048,n1050);
and (n1048,n1049,n1036);
xor (n1049,n1032,n1033);
and (n1050,n1051,n1052);
xor (n1051,n1049,n1036);
and (n1052,n1053,n1041);
xor (n1053,n1038,n1039);
or (n1054,n1055,n1057);
and (n1055,n1056,n1036);
xor (n1056,n1046,n1047);
and (n1057,n1058,n1059);
xor (n1058,n1056,n1036);
and (n1059,n1060,n1041);
xor (n1060,n1051,n1052);
and (n1061,n1062,n1041);
xor (n1062,n1058,n1059);
and (n1063,n742,n1064);
or (n1064,n1065,n1068,n1087);
and (n1065,n619,n1066);
wire s0n1066,s1n1066,notn1066;
or (n1066,s0n1066,s1n1066);
not(notn1066,n29);
and (s0n1066,notn1066,n1067);
and (s1n1066,n29,n378);
xor (n1067,n1062,n1041);
and (n1068,n1066,n1069);
or (n1069,n1070,n1073,n1086);
and (n1070,n631,n1071);
wire s0n1071,s1n1071,notn1071;
or (n1071,s0n1071,s1n1071);
not(notn1071,n29);
and (s0n1071,notn1071,n1072);
and (s1n1071,n29,n384);
xor (n1072,n1060,n1041);
and (n1073,n1071,n1074);
or (n1074,n1075,n1078,n1085);
and (n1075,n646,n1076);
wire s0n1076,s1n1076,notn1076;
or (n1076,s0n1076,s1n1076);
not(notn1076,n29);
and (s0n1076,notn1076,n1077);
and (s1n1076,n29,n390);
xor (n1077,n1053,n1041);
and (n1078,n1076,n1079);
or (n1079,n1080,n1083,n1084);
and (n1080,n657,n1081);
wire s0n1081,s1n1081,notn1081;
or (n1081,s0n1081,s1n1081);
not(notn1081,n29);
and (s0n1081,notn1081,n1082);
and (s1n1081,n29,n211);
xor (n1082,n1040,n1041);
and (n1083,n1081,n5);
and (n1084,n657,n5);
and (n1085,n646,n1079);
and (n1086,n631,n1074);
and (n1087,n619,n1069);
and (n1088,n727,n1064);
endmodule
