module top (out,n27,n28,n33,n42,n43,n48,n53,n59,n68
        ,n69,n75,n79,n85,n99,n100,n107,n114,n116,n122
        ,n128,n134,n143,n144,n151,n156,n162,n175,n180,n186
        ,n193,n203,n204,n215,n222,n237,n259,n266,n279,n286
        ,n291,n297,n313,n319,n328,n335,n341,n348,n358,n371
        ,n378,n383,n389,n396,n397,n404,n407,n416,n417,n434
        ,n441,n442,n453,n459,n466,n477,n483,n489,n928,n935
        ,n956,n1125,n1131,n1142,n1146,n1163,n1169,n1175,n1177,n1192
        ,n1197,n1210,n1215,n1227,n1244,n1250,n1289,n1305,n1317,n1323
        ,n1344,n1357,n1377,n1463,n1470,n1475,n1595,n1639,n5179,n5180
        ,n5183);
output out;
input n27;
input n28;
input n33;
input n42;
input n43;
input n48;
input n53;
input n59;
input n68;
input n69;
input n75;
input n79;
input n85;
input n99;
input n100;
input n107;
input n114;
input n116;
input n122;
input n128;
input n134;
input n143;
input n144;
input n151;
input n156;
input n162;
input n175;
input n180;
input n186;
input n193;
input n203;
input n204;
input n215;
input n222;
input n237;
input n259;
input n266;
input n279;
input n286;
input n291;
input n297;
input n313;
input n319;
input n328;
input n335;
input n341;
input n348;
input n358;
input n371;
input n378;
input n383;
input n389;
input n396;
input n397;
input n404;
input n407;
input n416;
input n417;
input n434;
input n441;
input n442;
input n453;
input n459;
input n466;
input n477;
input n483;
input n489;
input n928;
input n935;
input n956;
input n1125;
input n1131;
input n1142;
input n1146;
input n1163;
input n1169;
input n1175;
input n1177;
input n1192;
input n1197;
input n1210;
input n1215;
input n1227;
input n1244;
input n1250;
input n1289;
input n1305;
input n1317;
input n1323;
input n1344;
input n1357;
input n1377;
input n1463;
input n1470;
input n1475;
input n1595;
input n1639;
input n5179;
input n5180;
input n5183;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n24;
wire n25;
wire n26;
wire n29;
wire n30;
wire n31;
wire n32;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n44;
wire n45;
wire n46;
wire n47;
wire n49;
wire n50;
wire n51;
wire n52;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n76;
wire n77;
wire n78;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n115;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n152;
wire n153;
wire n154;
wire n155;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n176;
wire n177;
wire n178;
wire n179;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n287;
wire n288;
wire n289;
wire n290;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n379;
wire n380;
wire n381;
wire n382;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n405;
wire n406;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1143;
wire n1144;
wire n1145;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1176;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2988;
wire n2989;
wire n2990;
wire n2991;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2996;
wire n2997;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3003;
wire n3004;
wire n3005;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3010;
wire n3011;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3038;
wire n3039;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
wire n3056;
wire n3057;
wire n3058;
wire n3059;
wire n3060;
wire n3061;
wire n3062;
wire n3063;
wire n3064;
wire n3065;
wire n3066;
wire n3067;
wire n3068;
wire n3069;
wire n3070;
wire n3071;
wire n3072;
wire n3073;
wire n3074;
wire n3075;
wire n3076;
wire n3077;
wire n3078;
wire n3079;
wire n3080;
wire n3081;
wire n3082;
wire n3083;
wire n3084;
wire n3085;
wire n3086;
wire n3087;
wire n3088;
wire n3089;
wire n3090;
wire n3091;
wire n3092;
wire n3093;
wire n3094;
wire n3095;
wire n3096;
wire n3097;
wire n3098;
wire n3099;
wire n3100;
wire n3101;
wire n3102;
wire n3103;
wire n3104;
wire n3105;
wire n3106;
wire n3107;
wire n3108;
wire n3109;
wire n3110;
wire n3111;
wire n3112;
wire n3113;
wire n3114;
wire n3115;
wire n3116;
wire n3117;
wire n3118;
wire n3119;
wire n3120;
wire n3121;
wire n3122;
wire n3123;
wire n3124;
wire n3125;
wire n3126;
wire n3127;
wire n3128;
wire n3129;
wire n3130;
wire n3131;
wire n3132;
wire n3133;
wire n3134;
wire n3135;
wire n3136;
wire n3137;
wire n3138;
wire n3139;
wire n3140;
wire n3141;
wire n3142;
wire n3143;
wire n3144;
wire n3145;
wire n3146;
wire n3147;
wire n3148;
wire n3149;
wire n3150;
wire n3151;
wire n3152;
wire n3153;
wire n3154;
wire n3155;
wire n3156;
wire n3157;
wire n3158;
wire n3159;
wire n3160;
wire n3161;
wire n3162;
wire n3163;
wire n3164;
wire n3165;
wire n3166;
wire n3167;
wire n3168;
wire n3169;
wire n3170;
wire n3171;
wire n3172;
wire n3173;
wire n3174;
wire n3175;
wire n3176;
wire n3177;
wire n3178;
wire n3179;
wire n3180;
wire n3181;
wire n3182;
wire n3183;
wire n3184;
wire n3185;
wire n3186;
wire n3187;
wire n3188;
wire n3189;
wire n3190;
wire n3191;
wire n3192;
wire n3193;
wire n3194;
wire n3195;
wire n3196;
wire n3197;
wire n3198;
wire n3199;
wire n3200;
wire n3201;
wire n3202;
wire n3203;
wire n3204;
wire n3205;
wire n3206;
wire n3207;
wire n3208;
wire n3209;
wire n3210;
wire n3211;
wire n3212;
wire n3213;
wire n3214;
wire n3215;
wire n3216;
wire n3217;
wire n3218;
wire n3219;
wire n3220;
wire n3221;
wire n3222;
wire n3223;
wire n3224;
wire n3225;
wire n3226;
wire n3227;
wire n3228;
wire n3229;
wire n3230;
wire n3231;
wire n3232;
wire n3233;
wire n3234;
wire n3235;
wire n3236;
wire n3237;
wire n3238;
wire n3239;
wire n3240;
wire n3241;
wire n3242;
wire n3243;
wire n3244;
wire n3245;
wire n3246;
wire n3247;
wire n3248;
wire n3249;
wire n3250;
wire n3251;
wire n3252;
wire n3253;
wire n3254;
wire n3255;
wire n3256;
wire n3257;
wire n3258;
wire n3259;
wire n3260;
wire n3261;
wire n3262;
wire n3263;
wire n3264;
wire n3265;
wire n3266;
wire n3267;
wire n3268;
wire n3269;
wire n3270;
wire n3271;
wire n3272;
wire n3273;
wire n3274;
wire n3275;
wire n3276;
wire n3277;
wire n3278;
wire n3279;
wire n3280;
wire n3281;
wire n3282;
wire n3283;
wire n3284;
wire n3285;
wire n3286;
wire n3287;
wire n3288;
wire n3289;
wire n3290;
wire n3291;
wire n3292;
wire n3293;
wire n3294;
wire n3295;
wire n3296;
wire n3297;
wire n3298;
wire n3299;
wire n3300;
wire n3301;
wire n3302;
wire n3303;
wire n3304;
wire n3305;
wire n3306;
wire n3307;
wire n3308;
wire n3309;
wire n3310;
wire n3311;
wire n3312;
wire n3313;
wire n3314;
wire n3315;
wire n3316;
wire n3317;
wire n3318;
wire n3319;
wire n3320;
wire n3321;
wire n3322;
wire n3323;
wire n3324;
wire n3325;
wire n3326;
wire n3327;
wire n3328;
wire n3329;
wire n3330;
wire n3331;
wire n3332;
wire n3333;
wire n3334;
wire n3335;
wire n3336;
wire n3337;
wire n3338;
wire n3339;
wire n3340;
wire n3341;
wire n3342;
wire n3343;
wire n3344;
wire n3345;
wire n3346;
wire n3347;
wire n3348;
wire n3349;
wire n3350;
wire n3351;
wire n3352;
wire n3353;
wire n3354;
wire n3355;
wire n3356;
wire n3357;
wire n3358;
wire n3359;
wire n3360;
wire n3361;
wire n3362;
wire n3363;
wire n3364;
wire n3365;
wire n3366;
wire n3367;
wire n3368;
wire n3369;
wire n3370;
wire n3371;
wire n3372;
wire n3373;
wire n3374;
wire n3375;
wire n3376;
wire n3377;
wire n3378;
wire n3379;
wire n3380;
wire n3381;
wire n3382;
wire n3383;
wire n3384;
wire n3385;
wire n3386;
wire n3387;
wire n3388;
wire n3389;
wire n3390;
wire n3391;
wire n3392;
wire n3393;
wire n3394;
wire n3395;
wire n3396;
wire n3397;
wire n3398;
wire n3399;
wire n3400;
wire n3401;
wire n3402;
wire n3403;
wire n3404;
wire n3405;
wire n3406;
wire n3407;
wire n3408;
wire n3409;
wire n3410;
wire n3411;
wire n3412;
wire n3413;
wire n3414;
wire n3415;
wire n3416;
wire n3417;
wire n3418;
wire n3419;
wire n3420;
wire n3421;
wire n3422;
wire n3423;
wire n3424;
wire n3425;
wire n3426;
wire n3427;
wire n3428;
wire n3429;
wire n3430;
wire n3431;
wire n3432;
wire n3433;
wire n3434;
wire n3435;
wire n3436;
wire n3437;
wire n3438;
wire n3439;
wire n3440;
wire n3441;
wire n3442;
wire n3443;
wire n3444;
wire n3445;
wire n3446;
wire n3447;
wire n3448;
wire n3449;
wire n3450;
wire n3451;
wire n3452;
wire n3453;
wire n3454;
wire n3455;
wire n3456;
wire n3457;
wire n3458;
wire n3459;
wire n3460;
wire n3461;
wire n3462;
wire n3463;
wire n3464;
wire n3465;
wire n3466;
wire n3467;
wire n3468;
wire n3469;
wire n3470;
wire n3471;
wire n3472;
wire n3473;
wire n3474;
wire n3475;
wire n3476;
wire n3477;
wire n3478;
wire n3479;
wire n3480;
wire n3481;
wire n3482;
wire n3483;
wire n3484;
wire n3485;
wire n3486;
wire n3487;
wire n3488;
wire n3489;
wire n3490;
wire n3491;
wire n3492;
wire n3493;
wire n3494;
wire n3495;
wire n3496;
wire n3497;
wire n3498;
wire n3499;
wire n3500;
wire n3501;
wire n3502;
wire n3503;
wire n3504;
wire n3505;
wire n3506;
wire n3507;
wire n3508;
wire n3509;
wire n3510;
wire n3511;
wire n3512;
wire n3513;
wire n3514;
wire n3515;
wire n3516;
wire n3517;
wire n3518;
wire n3519;
wire n3520;
wire n3521;
wire n3522;
wire n3523;
wire n3524;
wire n3525;
wire n3526;
wire n3527;
wire n3528;
wire n3529;
wire n3530;
wire n3531;
wire n3532;
wire n3533;
wire n3534;
wire n3535;
wire n3536;
wire n3537;
wire n3538;
wire n3539;
wire n3540;
wire n3541;
wire n3542;
wire n3543;
wire n3544;
wire n3545;
wire n3546;
wire n3547;
wire n3548;
wire n3549;
wire n3550;
wire n3551;
wire n3552;
wire n3553;
wire n3554;
wire n3555;
wire n3556;
wire n3557;
wire n3558;
wire n3559;
wire n3560;
wire n3561;
wire n3562;
wire n3563;
wire n3564;
wire n3565;
wire n3566;
wire n3567;
wire n3568;
wire n3569;
wire n3570;
wire n3571;
wire n3572;
wire n3573;
wire n3574;
wire n3575;
wire n3576;
wire n3577;
wire n3578;
wire n3579;
wire n3580;
wire n3581;
wire n3582;
wire n3583;
wire n3584;
wire n3585;
wire n3586;
wire n3587;
wire n3588;
wire n3589;
wire n3590;
wire n3591;
wire n3592;
wire n3593;
wire n3594;
wire n3595;
wire n3596;
wire n3597;
wire n3598;
wire n3599;
wire n3600;
wire n3601;
wire n3602;
wire n3603;
wire n3604;
wire n3605;
wire n3606;
wire n3607;
wire n3608;
wire n3609;
wire n3610;
wire n3611;
wire n3612;
wire n3613;
wire n3614;
wire n3615;
wire n3616;
wire n3617;
wire n3618;
wire n3619;
wire n3620;
wire n3621;
wire n3622;
wire n3623;
wire n3624;
wire n3625;
wire n3626;
wire n3627;
wire n3628;
wire n3629;
wire n3630;
wire n3631;
wire n3632;
wire n3633;
wire n3634;
wire n3635;
wire n3636;
wire n3637;
wire n3638;
wire n3639;
wire n3640;
wire n3641;
wire n3642;
wire n3643;
wire n3644;
wire n3645;
wire n3646;
wire n3647;
wire n3648;
wire n3649;
wire n3650;
wire n3651;
wire n3652;
wire n3653;
wire n3654;
wire n3655;
wire n3656;
wire n3657;
wire n3658;
wire n3659;
wire n3660;
wire n3661;
wire n3662;
wire n3663;
wire n3664;
wire n3665;
wire n3666;
wire n3667;
wire n3668;
wire n3669;
wire n3670;
wire n3671;
wire n3672;
wire n3673;
wire n3674;
wire n3675;
wire n3676;
wire n3677;
wire n3678;
wire n3679;
wire n3680;
wire n3681;
wire n3682;
wire n3683;
wire n3684;
wire n3685;
wire n3686;
wire n3687;
wire n3688;
wire n3689;
wire n3690;
wire n3691;
wire n3692;
wire n3693;
wire n3694;
wire n3695;
wire n3696;
wire n3697;
wire n3698;
wire n3699;
wire n3700;
wire n3701;
wire n3702;
wire n3703;
wire n3704;
wire n3705;
wire n3706;
wire n3707;
wire n3708;
wire n3709;
wire n3710;
wire n3711;
wire n3712;
wire n3713;
wire n3714;
wire n3715;
wire n3716;
wire n3717;
wire n3718;
wire n3719;
wire n3720;
wire n3721;
wire n3722;
wire n3723;
wire n3724;
wire n3725;
wire n3726;
wire n3727;
wire n3728;
wire n3729;
wire n3730;
wire n3731;
wire n3732;
wire n3733;
wire n3734;
wire n3735;
wire n3736;
wire n3737;
wire n3738;
wire n3739;
wire n3740;
wire n3741;
wire n3742;
wire n3743;
wire n3744;
wire n3745;
wire n3746;
wire n3747;
wire n3748;
wire n3749;
wire n3750;
wire n3751;
wire n3752;
wire n3753;
wire n3754;
wire n3755;
wire n3756;
wire n3757;
wire n3758;
wire n3759;
wire n3760;
wire n3761;
wire n3762;
wire n3763;
wire n3764;
wire n3765;
wire n3766;
wire n3767;
wire n3768;
wire n3769;
wire n3770;
wire n3771;
wire n3772;
wire n3773;
wire n3774;
wire n3775;
wire n3776;
wire n3777;
wire n3778;
wire n3779;
wire n3780;
wire n3781;
wire n3782;
wire n3783;
wire n3784;
wire n3785;
wire n3786;
wire n3787;
wire n3788;
wire n3789;
wire n3790;
wire n3791;
wire n3792;
wire n3793;
wire n3794;
wire n3795;
wire n3796;
wire n3797;
wire n3798;
wire n3799;
wire n3800;
wire n3801;
wire n3802;
wire n3803;
wire n3804;
wire n3805;
wire n3806;
wire n3807;
wire n3808;
wire n3809;
wire n3810;
wire n3811;
wire n3812;
wire n3813;
wire n3814;
wire n3815;
wire n3816;
wire n3817;
wire n3818;
wire n3819;
wire n3820;
wire n3821;
wire n3822;
wire n3823;
wire n3824;
wire n3825;
wire n3826;
wire n3827;
wire n3828;
wire n3829;
wire n3830;
wire n3831;
wire n3832;
wire n3833;
wire n3834;
wire n3835;
wire n3836;
wire n3837;
wire n3838;
wire n3839;
wire n3840;
wire n3841;
wire n3842;
wire n3843;
wire n3844;
wire n3845;
wire n3846;
wire n3847;
wire n3848;
wire n3849;
wire n3850;
wire n3851;
wire n3852;
wire n3853;
wire n3854;
wire n3855;
wire n3856;
wire n3857;
wire n3858;
wire n3859;
wire n3860;
wire n3861;
wire n3862;
wire n3863;
wire n3864;
wire n3865;
wire n3866;
wire n3867;
wire n3868;
wire n3869;
wire n3870;
wire n3871;
wire n3872;
wire n3873;
wire n3874;
wire n3875;
wire n3876;
wire n3877;
wire n3878;
wire n3879;
wire n3880;
wire n3881;
wire n3882;
wire n3883;
wire n3884;
wire n3885;
wire n3886;
wire n3887;
wire n3888;
wire n3889;
wire n3890;
wire n3891;
wire n3892;
wire n3893;
wire n3894;
wire n3895;
wire n3896;
wire n3897;
wire n3898;
wire n3899;
wire n3900;
wire n3901;
wire n3902;
wire n3903;
wire n3904;
wire n3905;
wire n3906;
wire n3907;
wire n3908;
wire n3909;
wire n3910;
wire n3911;
wire n3912;
wire n3913;
wire n3914;
wire n3915;
wire n3916;
wire n3917;
wire n3918;
wire n3919;
wire n3920;
wire n3921;
wire n3922;
wire n3923;
wire n3924;
wire n3925;
wire n3926;
wire n3927;
wire n3928;
wire n3929;
wire n3930;
wire n3931;
wire n3932;
wire n3933;
wire n3934;
wire n3935;
wire n3936;
wire n3937;
wire n3938;
wire n3939;
wire n3940;
wire n3941;
wire n3942;
wire n3943;
wire n3944;
wire n3945;
wire n3946;
wire n3947;
wire n3948;
wire n3949;
wire n3950;
wire n3951;
wire n3952;
wire n3953;
wire n3954;
wire n3955;
wire n3956;
wire n3957;
wire n3958;
wire n3959;
wire n3960;
wire n3961;
wire n3962;
wire n3963;
wire n3964;
wire n3965;
wire n3966;
wire n3967;
wire n3968;
wire n3969;
wire n3970;
wire n3971;
wire n3972;
wire n3973;
wire n3974;
wire n3975;
wire n3976;
wire n3977;
wire n3978;
wire n3979;
wire n3980;
wire n3981;
wire n3982;
wire n3983;
wire n3984;
wire n3985;
wire n3986;
wire n3987;
wire n3988;
wire n3989;
wire n3990;
wire n3991;
wire n3992;
wire n3993;
wire n3994;
wire n3995;
wire n3996;
wire n3997;
wire n3998;
wire n3999;
wire n4000;
wire n4001;
wire n4002;
wire n4003;
wire n4004;
wire n4005;
wire n4006;
wire n4007;
wire n4008;
wire n4009;
wire n4010;
wire n4011;
wire n4012;
wire n4013;
wire n4014;
wire n4015;
wire n4016;
wire n4017;
wire n4018;
wire n4019;
wire n4020;
wire n4021;
wire n4022;
wire n4023;
wire n4024;
wire n4025;
wire n4026;
wire n4027;
wire n4028;
wire n4029;
wire n4030;
wire n4031;
wire n4032;
wire n4033;
wire n4034;
wire n4035;
wire n4036;
wire n4037;
wire n4038;
wire n4039;
wire n4040;
wire n4041;
wire n4042;
wire n4043;
wire n4044;
wire n4045;
wire n4046;
wire n4047;
wire n4048;
wire n4049;
wire n4050;
wire n4051;
wire n4052;
wire n4053;
wire n4054;
wire n4055;
wire n4056;
wire n4057;
wire n4058;
wire n4059;
wire n4060;
wire n4061;
wire n4062;
wire n4063;
wire n4064;
wire n4065;
wire n4066;
wire n4067;
wire n4068;
wire n4069;
wire n4070;
wire n4071;
wire n4072;
wire n4073;
wire n4074;
wire n4075;
wire n4076;
wire n4077;
wire n4078;
wire n4079;
wire n4080;
wire n4081;
wire n4082;
wire n4083;
wire n4084;
wire n4085;
wire n4086;
wire n4087;
wire n4088;
wire n4089;
wire n4090;
wire n4091;
wire n4092;
wire n4093;
wire n4094;
wire n4095;
wire n4096;
wire n4097;
wire n4098;
wire n4099;
wire n4100;
wire n4101;
wire n4102;
wire n4103;
wire n4104;
wire n4105;
wire n4106;
wire n4107;
wire n4108;
wire n4109;
wire n4110;
wire n4111;
wire n4112;
wire n4113;
wire n4114;
wire n4115;
wire n4116;
wire n4117;
wire n4118;
wire n4119;
wire n4120;
wire n4121;
wire n4122;
wire n4123;
wire n4124;
wire n4125;
wire n4126;
wire n4127;
wire n4128;
wire n4129;
wire n4130;
wire n4131;
wire n4132;
wire n4133;
wire n4134;
wire n4135;
wire n4136;
wire n4137;
wire n4138;
wire n4139;
wire n4140;
wire n4141;
wire n4142;
wire n4143;
wire n4144;
wire n4145;
wire n4146;
wire n4147;
wire n4148;
wire n4149;
wire n4150;
wire n4151;
wire n4152;
wire n4153;
wire n4154;
wire n4155;
wire n4156;
wire n4157;
wire n4158;
wire n4159;
wire n4160;
wire n4161;
wire n4162;
wire n4163;
wire n4164;
wire n4165;
wire n4166;
wire n4167;
wire n4168;
wire n4169;
wire n4170;
wire n4171;
wire n4172;
wire n4173;
wire n4174;
wire n4175;
wire n4176;
wire n4177;
wire n4178;
wire n4179;
wire n4180;
wire n4181;
wire n4182;
wire n4183;
wire n4184;
wire n4185;
wire n4186;
wire n4187;
wire n4188;
wire n4189;
wire n4190;
wire n4191;
wire n4192;
wire n4193;
wire n4194;
wire n4195;
wire n4196;
wire n4197;
wire n4198;
wire n4199;
wire n4200;
wire n4201;
wire n4202;
wire n4203;
wire n4204;
wire n4205;
wire n4206;
wire n4207;
wire n4208;
wire n4209;
wire n4210;
wire n4211;
wire n4212;
wire n4213;
wire n4214;
wire n4215;
wire n4216;
wire n4217;
wire n4218;
wire n4219;
wire n4220;
wire n4221;
wire n4222;
wire n4223;
wire n4224;
wire n4225;
wire n4226;
wire n4227;
wire n4228;
wire n4229;
wire n4230;
wire n4231;
wire n4232;
wire n4233;
wire n4234;
wire n4235;
wire n4236;
wire n4237;
wire n4238;
wire n4239;
wire n4240;
wire n4241;
wire n4242;
wire n4243;
wire n4244;
wire n4245;
wire n4246;
wire n4247;
wire n4248;
wire n4249;
wire n4250;
wire n4251;
wire n4252;
wire n4253;
wire n4254;
wire n4255;
wire n4256;
wire n4257;
wire n4258;
wire n4259;
wire n4260;
wire n4261;
wire n4262;
wire n4263;
wire n4264;
wire n4265;
wire n4266;
wire n4267;
wire n4268;
wire n4269;
wire n4270;
wire n4271;
wire n4272;
wire n4273;
wire n4274;
wire n4275;
wire n4276;
wire n4277;
wire n4278;
wire n4279;
wire n4280;
wire n4281;
wire n4282;
wire n4283;
wire n4284;
wire n4285;
wire n4286;
wire n4287;
wire n4288;
wire n4289;
wire n4290;
wire n4291;
wire n4292;
wire n4293;
wire n4294;
wire n4295;
wire n4296;
wire n4297;
wire n4298;
wire n4299;
wire n4300;
wire n4301;
wire n4302;
wire n4303;
wire n4304;
wire n4305;
wire n4306;
wire n4307;
wire n4308;
wire n4309;
wire n4310;
wire n4311;
wire n4312;
wire n4313;
wire n4314;
wire n4315;
wire n4316;
wire n4317;
wire n4318;
wire n4319;
wire n4320;
wire n4321;
wire n4322;
wire n4323;
wire n4324;
wire n4325;
wire n4326;
wire n4327;
wire n4328;
wire n4329;
wire n4330;
wire n4331;
wire n4332;
wire n4333;
wire n4334;
wire n4335;
wire n4336;
wire n4337;
wire n4338;
wire n4339;
wire n4340;
wire n4341;
wire n4342;
wire n4343;
wire n4344;
wire n4345;
wire n4346;
wire n4347;
wire n4348;
wire n4349;
wire n4350;
wire n4351;
wire n4352;
wire n4353;
wire n4354;
wire n4355;
wire n4356;
wire n4357;
wire n4358;
wire n4359;
wire n4360;
wire n4361;
wire n4362;
wire n4363;
wire n4364;
wire n4365;
wire n4366;
wire n4367;
wire n4368;
wire n4369;
wire n4370;
wire n4371;
wire n4372;
wire n4373;
wire n4374;
wire n4375;
wire n4376;
wire n4377;
wire n4378;
wire n4379;
wire n4380;
wire n4381;
wire n4382;
wire n4383;
wire n4384;
wire n4385;
wire n4386;
wire n4387;
wire n4388;
wire n4389;
wire n4390;
wire n4391;
wire n4392;
wire n4393;
wire n4394;
wire n4395;
wire n4396;
wire n4397;
wire n4398;
wire n4399;
wire n4400;
wire n4401;
wire n4402;
wire n4403;
wire n4404;
wire n4405;
wire n4406;
wire n4407;
wire n4408;
wire n4409;
wire n4410;
wire n4411;
wire n4412;
wire n4413;
wire n4414;
wire n4415;
wire n4416;
wire n4417;
wire n4418;
wire n4419;
wire n4420;
wire n4421;
wire n4422;
wire n4423;
wire n4424;
wire n4425;
wire n4426;
wire n4427;
wire n4428;
wire n4429;
wire n4430;
wire n4431;
wire n4432;
wire n4433;
wire n4434;
wire n4435;
wire n4436;
wire n4437;
wire n4438;
wire n4439;
wire n4440;
wire n4441;
wire n4442;
wire n4443;
wire n4444;
wire n4445;
wire n4446;
wire n4447;
wire n4448;
wire n4449;
wire n4450;
wire n4451;
wire n4452;
wire n4453;
wire n4454;
wire n4455;
wire n4456;
wire n4457;
wire n4458;
wire n4459;
wire n4460;
wire n4461;
wire n4462;
wire n4463;
wire n4464;
wire n4465;
wire n4466;
wire n4467;
wire n4468;
wire n4469;
wire n4470;
wire n4471;
wire n4472;
wire n4473;
wire n4474;
wire n4475;
wire n4476;
wire n4477;
wire n4478;
wire n4479;
wire n4480;
wire n4481;
wire n4482;
wire n4483;
wire n4484;
wire n4485;
wire n4486;
wire n4487;
wire n4488;
wire n4489;
wire n4490;
wire n4491;
wire n4492;
wire n4493;
wire n4494;
wire n4495;
wire n4496;
wire n4497;
wire n4498;
wire n4499;
wire n4500;
wire n4501;
wire n4502;
wire n4503;
wire n4504;
wire n4505;
wire n4506;
wire n4507;
wire n4508;
wire n4509;
wire n4510;
wire n4511;
wire n4512;
wire n4513;
wire n4514;
wire n4515;
wire n4516;
wire n4517;
wire n4518;
wire n4519;
wire n4520;
wire n4521;
wire n4522;
wire n4523;
wire n4524;
wire n4525;
wire n4526;
wire n4527;
wire n4528;
wire n4529;
wire n4530;
wire n4531;
wire n4532;
wire n4533;
wire n4534;
wire n4535;
wire n4536;
wire n4537;
wire n4538;
wire n4539;
wire n4540;
wire n4541;
wire n4542;
wire n4543;
wire n4544;
wire n4545;
wire n4546;
wire n4547;
wire n4548;
wire n4549;
wire n4550;
wire n4551;
wire n4552;
wire n4553;
wire n4554;
wire n4555;
wire n4556;
wire n4557;
wire n4558;
wire n4559;
wire n4560;
wire n4561;
wire n4562;
wire n4563;
wire n4564;
wire n4565;
wire n4566;
wire n4567;
wire n4568;
wire n4569;
wire n4570;
wire n4571;
wire n4572;
wire n4573;
wire n4574;
wire n4575;
wire n4576;
wire n4577;
wire n4578;
wire n4579;
wire n4580;
wire n4581;
wire n4582;
wire n4583;
wire n4584;
wire n4585;
wire n4586;
wire n4587;
wire n4588;
wire n4589;
wire n4590;
wire n4591;
wire n4592;
wire n4593;
wire n4594;
wire n4595;
wire n4596;
wire n4597;
wire n4598;
wire n4599;
wire n4600;
wire n4601;
wire n4602;
wire n4603;
wire n4604;
wire n4605;
wire n4606;
wire n4607;
wire n4608;
wire n4609;
wire n4610;
wire n4611;
wire n4612;
wire n4613;
wire n4614;
wire n4615;
wire n4616;
wire n4617;
wire n4618;
wire n4619;
wire n4620;
wire n4621;
wire n4622;
wire n4623;
wire n4624;
wire n4625;
wire n4626;
wire n4627;
wire n4628;
wire n4629;
wire n4630;
wire n4631;
wire n4632;
wire n4633;
wire n4634;
wire n4635;
wire n4636;
wire n4637;
wire n4638;
wire n4639;
wire n4640;
wire n4641;
wire n4642;
wire n4643;
wire n4644;
wire n4645;
wire n4646;
wire n4647;
wire n4648;
wire n4649;
wire n4650;
wire n4651;
wire n4652;
wire n4653;
wire n4654;
wire n4655;
wire n4656;
wire n4657;
wire n4658;
wire n4659;
wire n4660;
wire n4661;
wire n4662;
wire n4663;
wire n4664;
wire n4665;
wire n4666;
wire n4667;
wire n4668;
wire n4669;
wire n4670;
wire n4671;
wire n4672;
wire n4673;
wire n4674;
wire n4675;
wire n4676;
wire n4677;
wire n4678;
wire n4679;
wire n4680;
wire n4681;
wire n4682;
wire n4683;
wire n4684;
wire n4685;
wire n4686;
wire n4687;
wire n4688;
wire n4689;
wire n4690;
wire n4691;
wire n4692;
wire n4693;
wire n4694;
wire n4695;
wire n4696;
wire n4697;
wire n4698;
wire n4699;
wire n4700;
wire n4701;
wire n4702;
wire n4703;
wire n4704;
wire n4705;
wire n4706;
wire n4707;
wire n4708;
wire n4709;
wire n4710;
wire n4711;
wire n4712;
wire n4713;
wire n4714;
wire n4715;
wire n4716;
wire n4717;
wire n4718;
wire n4719;
wire n4720;
wire n4721;
wire n4722;
wire n4723;
wire n4724;
wire n4725;
wire n4726;
wire n4727;
wire n4728;
wire n4729;
wire n4730;
wire n4731;
wire n4732;
wire n4733;
wire n4734;
wire n4735;
wire n4736;
wire n4737;
wire n4738;
wire n4739;
wire n4740;
wire n4741;
wire n4742;
wire n4743;
wire n4744;
wire n4745;
wire n4746;
wire n4747;
wire n4748;
wire n4749;
wire n4750;
wire n4751;
wire n4752;
wire n4753;
wire n4754;
wire n4755;
wire n4756;
wire n4757;
wire n4758;
wire n4759;
wire n4760;
wire n4761;
wire n4762;
wire n4763;
wire n4764;
wire n4765;
wire n4766;
wire n4767;
wire n4768;
wire n4769;
wire n4770;
wire n4771;
wire n4772;
wire n4773;
wire n4774;
wire n4775;
wire n4776;
wire n4777;
wire n4778;
wire n4779;
wire n4780;
wire n4781;
wire n4782;
wire n4783;
wire n4784;
wire n4785;
wire n4786;
wire n4787;
wire n4788;
wire n4789;
wire n4790;
wire n4791;
wire n4792;
wire n4793;
wire n4794;
wire n4795;
wire n4796;
wire n4797;
wire n4798;
wire n4799;
wire n4800;
wire n4801;
wire n4802;
wire n4803;
wire n4804;
wire n4805;
wire n4806;
wire n4807;
wire n4808;
wire n4809;
wire n4810;
wire n4811;
wire n4812;
wire n4813;
wire n4814;
wire n4815;
wire n4816;
wire n4817;
wire n4818;
wire n4819;
wire n4820;
wire n4821;
wire n4822;
wire n4823;
wire n4824;
wire n4825;
wire n4826;
wire n4827;
wire n4828;
wire n4829;
wire n4830;
wire n4831;
wire n4832;
wire n4833;
wire n4834;
wire n4835;
wire n4836;
wire n4837;
wire n4838;
wire n4839;
wire n4840;
wire n4841;
wire n4842;
wire n4843;
wire n4844;
wire n4845;
wire n4846;
wire n4847;
wire n4848;
wire n4849;
wire n4850;
wire n4851;
wire n4852;
wire n4853;
wire n4854;
wire n4855;
wire n4856;
wire n4857;
wire n4858;
wire n4859;
wire n4860;
wire n4861;
wire n4862;
wire n4863;
wire n4864;
wire n4865;
wire n4866;
wire n4867;
wire n4868;
wire n4869;
wire n4870;
wire n4871;
wire n4872;
wire n4873;
wire n4874;
wire n4875;
wire n4876;
wire n4877;
wire n4878;
wire n4879;
wire n4880;
wire n4881;
wire n4882;
wire n4883;
wire n4884;
wire n4885;
wire n4886;
wire n4887;
wire n4888;
wire n4889;
wire n4890;
wire n4891;
wire n4892;
wire n4893;
wire n4894;
wire n4895;
wire n4896;
wire n4897;
wire n4898;
wire n4899;
wire n4900;
wire n4901;
wire n4902;
wire n4903;
wire n4904;
wire n4905;
wire n4906;
wire n4907;
wire n4908;
wire n4909;
wire n4910;
wire n4911;
wire n4912;
wire n4913;
wire n4914;
wire n4915;
wire n4916;
wire n4917;
wire n4918;
wire n4919;
wire n4920;
wire n4921;
wire n4922;
wire n4923;
wire n4924;
wire n4925;
wire n4926;
wire n4927;
wire n4928;
wire n4929;
wire n4930;
wire n4931;
wire n4932;
wire n4933;
wire n4934;
wire n4935;
wire n4936;
wire n4937;
wire n4938;
wire n4939;
wire n4940;
wire n4941;
wire n4942;
wire n4943;
wire n4944;
wire n4945;
wire n4946;
wire n4947;
wire n4948;
wire n4949;
wire n4950;
wire n4951;
wire n4952;
wire n4953;
wire n4954;
wire n4955;
wire n4956;
wire n4957;
wire n4958;
wire n4959;
wire n4960;
wire n4961;
wire n4962;
wire n4963;
wire n4964;
wire n4965;
wire n4966;
wire n4967;
wire n4968;
wire n4969;
wire n4970;
wire n4971;
wire n4972;
wire n4973;
wire n4974;
wire n4975;
wire n4976;
wire n4977;
wire n4978;
wire n4979;
wire n4980;
wire n4981;
wire n4982;
wire n4983;
wire n4984;
wire n4985;
wire n4986;
wire n4987;
wire n4988;
wire n4989;
wire n4990;
wire n4991;
wire n4992;
wire n4993;
wire n4994;
wire n4995;
wire n4996;
wire n4997;
wire n4998;
wire n4999;
wire n5000;
wire n5001;
wire n5002;
wire n5003;
wire n5004;
wire n5005;
wire n5006;
wire n5007;
wire n5008;
wire n5009;
wire n5010;
wire n5011;
wire n5012;
wire n5013;
wire n5014;
wire n5015;
wire n5016;
wire n5017;
wire n5018;
wire n5019;
wire n5020;
wire n5021;
wire n5022;
wire n5023;
wire n5024;
wire n5025;
wire n5026;
wire n5027;
wire n5028;
wire n5029;
wire n5030;
wire n5031;
wire n5032;
wire n5033;
wire n5034;
wire n5035;
wire n5036;
wire n5037;
wire n5038;
wire n5039;
wire n5040;
wire n5041;
wire n5042;
wire n5043;
wire n5044;
wire n5045;
wire n5046;
wire n5047;
wire n5048;
wire n5049;
wire n5050;
wire n5051;
wire n5052;
wire n5053;
wire n5054;
wire n5055;
wire n5056;
wire n5057;
wire n5058;
wire n5059;
wire n5060;
wire n5061;
wire n5062;
wire n5063;
wire n5064;
wire n5065;
wire n5066;
wire n5067;
wire n5068;
wire n5069;
wire n5070;
wire n5071;
wire n5072;
wire n5073;
wire n5074;
wire n5075;
wire n5076;
wire n5077;
wire n5078;
wire n5079;
wire n5080;
wire n5081;
wire n5082;
wire n5083;
wire n5084;
wire n5085;
wire n5086;
wire n5087;
wire n5088;
wire n5089;
wire n5090;
wire n5091;
wire n5092;
wire n5093;
wire n5094;
wire n5095;
wire n5096;
wire n5097;
wire n5098;
wire n5099;
wire n5100;
wire n5101;
wire n5102;
wire n5103;
wire n5104;
wire n5105;
wire n5106;
wire n5107;
wire n5108;
wire n5109;
wire n5110;
wire n5111;
wire n5112;
wire n5113;
wire n5114;
wire n5115;
wire n5116;
wire n5117;
wire n5118;
wire n5119;
wire n5120;
wire n5121;
wire n5122;
wire n5123;
wire n5124;
wire n5125;
wire n5126;
wire n5127;
wire n5128;
wire n5129;
wire n5130;
wire n5131;
wire n5132;
wire n5133;
wire n5134;
wire n5135;
wire n5136;
wire n5137;
wire n5138;
wire n5139;
wire n5140;
wire n5141;
wire n5142;
wire n5143;
wire n5144;
wire n5145;
wire n5146;
wire n5147;
wire n5148;
wire n5149;
wire n5150;
wire n5151;
wire n5152;
wire n5153;
wire n5154;
wire n5155;
wire n5156;
wire n5157;
wire n5158;
wire n5159;
wire n5160;
wire n5161;
wire n5162;
wire n5163;
wire n5164;
wire n5165;
wire n5166;
wire n5167;
wire n5168;
wire n5169;
wire n5170;
wire n5171;
wire n5172;
wire n5173;
wire n5174;
wire n5175;
wire n5176;
wire n5177;
wire n5178;
wire n5181;
wire n5182;
wire n5184;
wire n5185;
wire n5186;
wire n5187;
wire n5188;
wire n5189;
wire n5190;
wire n5191;
wire n5192;
wire n5193;
wire n5194;
wire n5195;
wire n5196;
wire n5197;
wire n5198;
wire n5199;
wire n5200;
wire n5201;
wire n5202;
wire n5203;
wire n5204;
wire n5205;
wire n5206;
wire n5207;
wire n5208;
wire n5209;
wire n5210;
wire n5211;
wire n5212;
wire n5213;
wire n5214;
wire n5215;
wire n5216;
wire n5217;
wire n5218;
wire n5219;
wire n5220;
wire n5221;
wire n5222;
wire n5223;
wire n5224;
wire n5225;
wire n5226;
wire n5227;
wire n5228;
wire n5229;
wire n5230;
wire n5231;
wire n5232;
wire n5233;
wire n5234;
wire n5235;
wire n5236;
wire n5237;
wire n5238;
wire n5239;
wire n5240;
wire n5241;
wire n5242;
wire n5243;
wire n5244;
wire n5245;
wire n5246;
wire n5247;
wire n5248;
wire n5249;
wire n5250;
wire n5251;
wire n5252;
wire n5253;
wire n5254;
wire n5255;
wire n5256;
wire n5257;
wire n5258;
wire n5259;
wire n5260;
wire n5261;
wire n5262;
wire n5263;
wire n5264;
wire n5265;
wire n5266;
wire n5267;
wire n5268;
wire n5269;
wire n5270;
wire n5271;
wire n5272;
wire n5273;
wire n5274;
wire n5275;
wire n5276;
wire n5277;
wire n5278;
wire n5279;
wire n5280;
wire n5281;
wire n5282;
wire n5283;
wire n5284;
wire n5285;
wire n5286;
wire n5287;
wire n5288;
wire n5289;
wire n5290;
wire n5291;
wire n5292;
wire n5293;
wire n5294;
wire n5295;
wire n5296;
wire n5297;
wire n5298;
wire n5299;
wire n5300;
wire n5301;
wire n5302;
wire n5303;
wire n5304;
wire n5305;
wire n5306;
wire n5307;
wire n5308;
wire n5309;
wire n5310;
wire n5311;
wire n5312;
wire n5313;
wire n5314;
wire n5315;
wire n5316;
wire n5317;
wire n5318;
wire n5319;
wire n5320;
wire n5321;
wire n5322;
wire n5323;
wire n5324;
wire n5325;
wire n5326;
wire n5327;
wire n5328;
wire n5329;
wire n5330;
wire n5331;
wire n5332;
wire n5333;
wire n5334;
wire n5335;
wire n5336;
wire n5337;
wire n5338;
wire n5339;
wire n5340;
wire n5341;
wire n5342;
wire n5343;
wire n5344;
wire n5345;
wire n5346;
wire n5347;
wire n5348;
wire n5349;
wire n5350;
wire n5351;
wire n5352;
wire n5353;
wire n5354;
wire n5355;
wire n5356;
wire n5357;
wire n5358;
wire n5359;
wire n5360;
wire n5361;
wire n5362;
wire n5363;
wire n5364;
wire n5365;
wire n5366;
wire n5367;
wire n5368;
wire n5369;
wire n5370;
wire n5371;
wire n5372;
wire n5373;
wire n5374;
wire n5375;
wire n5376;
wire n5377;
wire n5378;
wire n5379;
wire n5380;
wire n5381;
wire n5382;
wire n5383;
wire n5384;
wire n5385;
wire n5386;
wire n5387;
wire n5388;
wire n5389;
wire n5390;
wire n5391;
wire n5392;
wire n5393;
wire n5394;
wire n5395;
wire n5396;
wire n5397;
wire n5398;
wire n5399;
wire n5400;
wire n5401;
wire n5402;
wire n5403;
wire n5404;
wire n5405;
wire n5406;
wire n5407;
wire n5408;
wire n5409;
wire n5410;
wire n5411;
wire n5412;
wire n5413;
wire n5414;
wire n5415;
wire n5416;
wire n5417;
wire n5418;
wire n5419;
wire n5420;
wire n5421;
wire n5422;
wire n5423;
wire n5424;
wire n5425;
wire n5426;
wire n5427;
wire n5428;
wire n5429;
wire n5430;
wire n5431;
wire n5432;
wire n5433;
wire n5434;
wire n5435;
wire n5436;
wire n5437;
wire n5438;
wire n5439;
wire n5440;
wire n5441;
wire n5442;
wire n5443;
wire n5444;
wire n5445;
wire n5446;
wire n5447;
wire n5448;
wire n5449;
wire n5450;
wire n5451;
wire n5452;
wire n5453;
wire n5454;
wire n5455;
wire n5456;
wire n5457;
wire n5458;
wire n5459;
wire n5460;
wire n5461;
wire n5462;
wire n5463;
wire n5464;
wire n5465;
wire n5466;
wire n5467;
wire n5468;
wire n5469;
wire n5470;
wire n5471;
wire n5472;
wire n5473;
wire n5474;
wire n5475;
wire n5476;
wire n5477;
wire n5478;
wire n5479;
wire n5480;
wire n5481;
wire n5482;
wire n5483;
wire n5484;
wire n5485;
wire n5486;
wire n5487;
wire n5488;
wire n5489;
wire n5490;
wire n5491;
wire n5492;
wire n5493;
wire n5494;
wire n5495;
wire n5496;
wire n5497;
wire n5498;
wire n5499;
wire n5500;
wire n5501;
wire n5502;
wire n5503;
wire n5504;
wire n5505;
wire n5506;
wire n5507;
wire n5508;
wire n5509;
wire n5510;
wire n5511;
wire n5512;
wire n5513;
wire n5514;
wire n5515;
wire n5516;
wire n5517;
wire n5518;
wire n5519;
wire n5520;
wire n5521;
wire n5522;
wire n5523;
wire n5524;
wire n5525;
wire n5526;
wire n5527;
wire n5528;
wire n5529;
wire n5530;
wire n5531;
wire n5532;
wire n5533;
wire n5534;
wire n5535;
wire n5536;
wire n5537;
wire n5538;
wire n5539;
wire n5540;
wire n5541;
wire n5542;
wire n5543;
wire n5544;
wire n5545;
wire n5546;
wire n5547;
wire n5548;
wire n5549;
wire n5550;
wire n5551;
wire n5552;
wire n5553;
wire n5554;
wire n5555;
wire n5556;
wire n5557;
wire n5558;
wire n5559;
wire n5560;
wire n5561;
wire n5562;
wire n5563;
wire n5564;
wire n5565;
wire n5566;
wire n5567;
wire n5568;
wire n5569;
wire n5570;
wire n5571;
wire n5572;
wire n5573;
wire n5574;
wire n5575;
wire n5576;
wire n5577;
wire n5578;
wire n5579;
wire n5580;
wire n5581;
wire n5582;
wire n5583;
wire n5584;
wire n5585;
wire n5586;
wire n5587;
wire n5588;
wire n5589;
wire n5590;
wire n5591;
wire n5592;
wire n5593;
wire n5594;
wire n5595;
wire n5596;
wire n5597;
wire n5598;
wire n5599;
wire n5600;
wire n5601;
wire n5602;
wire n5603;
wire n5604;
wire n5605;
wire n5606;
wire n5607;
wire n5608;
wire n5609;
wire n5610;
wire n5611;
wire n5612;
wire n5613;
wire n5614;
wire n5615;
wire n5616;
wire n5617;
wire n5618;
wire n5619;
wire n5620;
wire n5621;
wire n5622;
wire n5623;
wire n5624;
wire n5625;
wire n5626;
wire n5627;
wire n5628;
wire n5629;
wire n5630;
wire n5631;
wire n5632;
wire n5633;
wire n5634;
wire n5635;
wire n5636;
wire n5637;
wire n5638;
wire n5639;
wire n5640;
wire n5641;
wire n5642;
wire n5643;
wire n5644;
wire n5645;
wire n5646;
wire n5647;
wire n5648;
wire n5649;
wire n5650;
wire n5651;
wire n5652;
wire n5653;
wire n5654;
wire n5655;
wire n5656;
wire n5657;
wire n5658;
wire n5659;
wire n5660;
wire n5661;
wire n5662;
wire n5663;
wire n5664;
wire n5665;
wire n5666;
wire n5667;
wire n5668;
wire n5669;
wire n5670;
wire n5671;
wire n5672;
wire n5673;
wire n5674;
wire n5675;
wire n5676;
wire n5677;
wire n5678;
wire n5679;
wire n5680;
wire n5681;
wire n5682;
wire n5683;
wire n5684;
wire n5685;
wire n5686;
wire n5687;
wire n5688;
wire n5689;
wire n5690;
wire n5691;
wire n5692;
wire n5693;
wire n5694;
wire n5695;
wire n5696;
wire n5697;
wire n5698;
wire n5699;
wire n5700;
wire n5701;
wire n5702;
wire n5703;
wire n5704;
wire n5705;
wire n5706;
wire n5707;
wire n5708;
wire n5709;
wire n5710;
wire n5711;
wire n5712;
wire n5713;
wire n5714;
wire n5715;
wire n5716;
wire n5717;
wire n5718;
wire n5719;
wire n5720;
wire n5721;
wire n5722;
wire n5723;
wire n5724;
wire n5725;
wire n5726;
wire n5727;
wire n5728;
wire n5729;
wire n5730;
wire n5731;
wire n5732;
wire n5733;
wire n5734;
wire n5735;
wire n5736;
wire n5737;
wire n5738;
wire n5739;
wire n5740;
wire n5741;
wire n5742;
wire n5743;
wire n5744;
wire n5745;
wire n5746;
wire n5747;
wire n5748;
wire n5749;
wire n5750;
wire n5751;
wire n5752;
wire n5753;
wire n5754;
wire n5755;
wire n5756;
wire n5757;
wire n5758;
wire n5759;
wire n5760;
wire n5761;
wire n5762;
wire n5763;
wire n5764;
wire n5765;
wire n5766;
wire n5767;
wire n5768;
wire n5769;
wire n5770;
wire n5771;
wire n5772;
wire n5773;
wire n5774;
wire n5775;
wire n5776;
wire n5777;
wire n5778;
wire n5779;
wire n5780;
wire n5781;
wire n5782;
wire n5783;
wire n5784;
wire n5785;
wire n5786;
wire n5787;
wire n5788;
wire n5789;
wire n5790;
wire n5791;
wire n5792;
wire n5793;
wire n5794;
wire n5795;
wire n5796;
wire n5797;
wire n5798;
wire n5799;
wire n5800;
wire n5801;
wire n5802;
wire n5803;
wire n5804;
wire n5805;
wire n5806;
wire n5807;
wire n5808;
wire n5809;
wire n5810;
wire n5811;
wire n5812;
wire n5813;
wire n5814;
wire n5815;
wire n5816;
wire n5817;
wire n5818;
wire n5819;
wire n5820;
wire n5821;
wire n5822;
wire n5823;
wire n5824;
wire n5825;
wire n5826;
wire n5827;
wire n5828;
wire n5829;
wire n5830;
wire n5831;
wire n5832;
wire n5833;
wire n5834;
wire n5835;
wire n5836;
wire n5837;
wire n5838;
wire n5839;
wire n5840;
wire n5841;
wire n5842;
wire n5843;
wire n5844;
wire n5845;
wire n5846;
wire n5847;
wire n5848;
wire n5849;
wire n5850;
wire n5851;
wire n5852;
wire n5853;
wire n5854;
wire n5855;
wire n5856;
wire n5857;
wire n5858;
wire n5859;
wire n5860;
wire n5861;
wire n5862;
wire n5863;
wire n5864;
wire n5865;
wire n5866;
wire n5867;
wire n5868;
wire n5869;
wire n5870;
wire n5871;
wire n5872;
wire n5873;
wire n5874;
wire n5875;
wire n5876;
wire n5877;
wire n5878;
wire n5879;
wire n5880;
wire n5881;
wire n5882;
wire n5883;
wire n5884;
wire n5885;
wire n5886;
wire n5887;
wire n5888;
wire n5889;
wire n5890;
wire n5891;
wire n5892;
wire n5893;
wire n5894;
wire n5895;
wire n5896;
wire n5897;
wire n5898;
wire n5899;
wire n5900;
wire n5901;
wire n5902;
wire n5903;
wire n5904;
wire n5905;
wire n5906;
wire n5907;
wire n5908;
wire n5909;
wire n5910;
wire n5911;
wire n5912;
wire n5913;
wire n5914;
wire n5915;
wire n5916;
wire n5917;
wire n5918;
wire n5919;
wire n5920;
wire n5921;
wire n5922;
wire n5923;
wire n5924;
wire n5925;
wire n5926;
wire n5927;
wire n5928;
wire n5929;
wire n5930;
wire n5931;
wire n5932;
wire n5933;
wire n5934;
wire n5935;
wire n5936;
wire n5937;
wire n5938;
wire n5939;
wire n5940;
wire n5941;
wire n5942;
wire n5943;
wire n5944;
wire n5945;
wire n5946;
wire n5947;
wire n5948;
wire n5949;
wire n5950;
wire n5951;
wire n5952;
wire n5953;
wire n5954;
wire n5955;
wire n5956;
wire n5957;
wire n5958;
wire n5959;
wire n5960;
wire n5961;
wire n5962;
wire n5963;
wire n5964;
wire n5965;
wire n5966;
wire n5967;
wire n5968;
wire n5969;
wire n5970;
wire n5971;
wire n5972;
wire n5973;
wire n5974;
wire n5975;
wire n5976;
wire n5977;
wire n5978;
wire n5979;
wire n5980;
wire n5981;
wire n5982;
wire n5983;
wire n5984;
wire n5985;
wire n5986;
wire n5987;
wire n5988;
wire n5989;
wire n5990;
wire n5991;
wire n5992;
wire n5993;
wire n5994;
wire n5995;
wire n5996;
wire n5997;
wire n5998;
wire n5999;
wire n6000;
wire n6001;
wire n6002;
wire n6003;
wire n6004;
wire n6005;
wire n6006;
wire n6007;
wire n6008;
wire n6009;
wire n6010;
wire n6011;
wire n6012;
wire n6013;
wire n6014;
wire n6015;
wire n6016;
wire n6017;
wire n6018;
wire n6019;
wire n6020;
wire n6021;
wire n6022;
wire n6023;
wire n6024;
wire n6025;
wire n6026;
wire n6027;
wire n6028;
wire n6029;
wire n6030;
wire n6031;
wire n6032;
wire n6033;
wire n6034;
wire n6035;
wire n6036;
wire n6037;
wire n6038;
wire n6039;
wire n6040;
wire n6041;
wire n6042;
wire n6043;
wire n6044;
wire n6045;
wire n6046;
wire n6047;
wire n6048;
wire n6049;
wire n6050;
wire n6051;
wire n6052;
wire n6053;
wire n6054;
wire n6055;
wire n6056;
wire n6057;
wire n6058;
wire n6059;
wire n6060;
wire n6061;
wire n6062;
wire n6063;
wire n6064;
wire n6065;
wire n6066;
wire n6067;
wire n6068;
wire n6069;
wire n6070;
wire n6071;
wire n6072;
wire n6073;
wire n6074;
wire n6075;
wire n6076;
wire n6077;
wire n6078;
wire n6079;
wire n6080;
wire n6081;
wire n6082;
wire n6083;
wire n6084;
wire n6085;
wire n6086;
wire n6087;
wire n6088;
wire n6089;
wire n6090;
wire n6091;
wire n6092;
wire n6093;
wire n6094;
wire n6095;
wire n6096;
wire n6097;
wire n6098;
wire n6099;
wire n6100;
wire n6101;
wire n6102;
wire n6103;
wire n6104;
wire n6105;
wire n6106;
wire n6107;
wire n6108;
wire n6109;
wire n6110;
wire n6111;
wire n6112;
wire n6113;
wire n6114;
wire n6115;
wire n6116;
wire n6117;
wire n6118;
wire n6119;
wire n6120;
wire n6121;
wire n6122;
wire n6123;
wire n6124;
wire n6125;
wire n6126;
wire n6127;
wire n6128;
wire n6129;
wire n6130;
wire n6131;
wire n6132;
wire n6133;
wire n6134;
wire n6135;
wire n6136;
wire n6137;
wire n6138;
wire n6139;
wire n6140;
wire n6141;
wire n6142;
wire n6143;
wire n6144;
wire n6145;
wire n6146;
wire n6147;
wire n6148;
wire n6149;
wire n6150;
wire n6151;
wire n6152;
wire n6153;
wire n6154;
wire n6155;
wire n6156;
wire n6157;
wire n6158;
wire n6159;
wire n6160;
wire n6161;
wire n6162;
wire n6163;
wire n6164;
wire n6165;
wire n6166;
wire n6167;
wire n6168;
wire n6169;
wire n6170;
wire n6171;
wire n6172;
wire n6173;
wire n6174;
wire n6175;
wire n6176;
wire n6177;
wire n6178;
wire n6179;
wire n6180;
wire n6181;
wire n6182;
wire n6183;
wire n6184;
wire n6185;
wire n6186;
wire n6187;
wire n6188;
wire n6189;
wire n6190;
wire n6191;
wire n6192;
wire n6193;
wire n6194;
wire n6195;
wire n6196;
wire n6197;
wire n6198;
wire n6199;
wire n6200;
wire n6201;
wire n6202;
wire n6203;
wire n6204;
wire n6205;
wire n6206;
wire n6207;
wire n6208;
wire n6209;
wire n6210;
wire n6211;
wire n6212;
wire n6213;
wire n6214;
wire n6215;
wire n6216;
wire n6217;
wire n6218;
wire n6219;
wire n6220;
wire n6221;
wire n6222;
wire n6223;
wire n6224;
wire n6225;
wire n6226;
wire n6227;
wire n6228;
wire n6229;
wire n6230;
wire n6231;
wire n6232;
wire n6233;
wire n6234;
wire n6235;
wire n6236;
wire n6237;
wire n6238;
wire n6239;
wire n6240;
wire n6241;
wire n6242;
wire n6243;
wire n6244;
wire n6245;
wire n6246;
wire n6247;
wire n6248;
wire n6249;
wire n6250;
wire n6251;
wire n6252;
wire n6253;
wire n6254;
wire n6255;
wire n6256;
wire n6257;
wire n6258;
wire n6259;
wire n6260;
wire n6261;
wire n6262;
wire n6263;
wire n6264;
wire n6265;
wire n6266;
wire n6267;
wire n6268;
wire n6269;
wire n6270;
wire n6271;
wire n6272;
wire n6273;
wire n6274;
wire n6275;
wire n6276;
wire n6277;
wire n6278;
wire n6279;
wire n6280;
wire n6281;
wire n6282;
wire n6283;
wire n6284;
wire n6285;
wire n6286;
wire n6287;
wire n6288;
wire n6289;
wire n6290;
wire n6291;
wire n6292;
wire n6293;
wire n6294;
wire n6295;
wire n6296;
wire n6297;
wire n6298;
wire n6299;
wire n6300;
wire n6301;
wire n6302;
wire n6303;
wire n6304;
wire n6305;
wire n6306;
wire n6307;
wire n6308;
wire n6309;
wire n6310;
wire n6311;
wire n6312;
wire n6313;
wire n6314;
wire n6315;
wire n6316;
wire n6317;
wire n6318;
wire n6319;
wire n6320;
wire n6321;
wire n6322;
wire n6323;
wire n6324;
wire n6325;
wire n6326;
wire n6327;
wire n6328;
wire n6329;
wire n6330;
wire n6331;
wire n6332;
wire n6333;
wire n6334;
wire n6335;
wire n6336;
wire n6337;
wire n6338;
wire n6339;
wire n6340;
wire n6341;
wire n6342;
wire n6343;
wire n6344;
wire n6345;
wire n6346;
wire n6347;
wire n6348;
wire n6349;
wire n6350;
wire n6351;
wire n6352;
wire n6353;
wire n6354;
wire n6355;
wire n6356;
wire n6357;
wire n6358;
wire n6359;
wire n6360;
wire n6361;
wire n6362;
wire n6363;
wire n6364;
wire n6365;
wire n6366;
wire n6367;
wire n6368;
wire n6369;
wire n6370;
wire n6371;
wire n6372;
wire n6373;
wire n6374;
wire n6375;
wire n6376;
wire n6377;
wire n6378;
wire n6379;
wire n6380;
wire n6381;
wire n6382;
wire n6383;
wire n6384;
wire n6385;
wire n6386;
wire n6387;
wire n6388;
wire n6389;
wire n6390;
wire n6391;
wire n6392;
wire n6393;
wire n6394;
wire n6395;
wire n6396;
wire n6397;
wire n6398;
wire n6399;
wire n6400;
wire n6401;
wire n6402;
wire n6403;
wire n6404;
wire n6405;
wire n6406;
wire n6407;
wire n6408;
wire n6409;
wire n6410;
wire n6411;
wire n6412;
wire n6413;
wire n6414;
wire n6415;
wire n6416;
wire n6417;
wire n6418;
wire n6419;
wire n6420;
wire n6421;
wire n6422;
wire n6423;
wire n6424;
wire n6425;
wire n6426;
wire n6427;
wire n6428;
wire n6429;
wire n6430;
wire n6431;
wire n6432;
wire n6433;
wire n6434;
wire n6435;
wire n6436;
wire n6437;
wire n6438;
wire n6439;
wire n6440;
wire n6441;
wire n6442;
wire n6443;
wire n6444;
wire n6445;
wire n6446;
wire n6447;
wire n6448;
wire n6449;
wire n6450;
wire n6451;
wire n6452;
wire n6453;
wire n6454;
wire n6455;
wire n6456;
wire n6457;
wire n6458;
wire n6459;
wire n6460;
wire n6461;
wire n6462;
wire n6463;
wire n6464;
wire n6465;
wire n6466;
wire n6467;
wire n6468;
wire n6469;
wire n6470;
wire n6471;
wire n6472;
wire n6473;
wire n6474;
wire n6475;
wire n6476;
wire n6477;
wire n6478;
wire n6479;
wire n6480;
wire n6481;
wire n6482;
wire n6483;
wire n6484;
wire n6485;
wire n6486;
wire n6487;
wire n6488;
wire n6489;
wire n6490;
wire n6491;
wire n6492;
wire n6493;
wire n6494;
wire n6495;
wire n6496;
wire n6497;
wire n6498;
wire n6499;
wire n6500;
wire n6501;
wire n6502;
wire n6503;
wire n6504;
wire n6505;
wire n6506;
wire n6507;
wire n6508;
wire n6509;
wire n6510;
wire n6511;
wire n6512;
wire n6513;
wire n6514;
wire n6515;
wire n6516;
wire n6517;
wire n6518;
wire n6519;
wire n6520;
wire n6521;
wire n6522;
wire n6523;
wire n6524;
wire n6525;
wire n6526;
wire n6527;
wire n6528;
wire n6529;
wire n6530;
wire n6531;
wire n6532;
wire n6533;
wire n6534;
wire n6535;
wire n6536;
wire n6537;
wire n6538;
wire n6539;
wire n6540;
wire n6541;
wire n6542;
wire n6543;
wire n6544;
wire n6545;
wire n6546;
wire n6547;
wire n6548;
wire n6549;
wire n6550;
wire n6551;
wire n6552;
wire n6553;
wire n6554;
wire n6555;
wire n6556;
wire n6557;
wire n6558;
wire n6559;
wire n6560;
wire n6561;
wire n6562;
wire n6563;
wire n6564;
wire n6565;
wire n6566;
wire n6567;
wire n6568;
wire n6569;
wire n6570;
wire n6571;
wire n6572;
wire n6573;
wire n6574;
wire n6575;
wire n6576;
wire n6577;
wire n6578;
wire n6579;
wire n6580;
wire n6581;
wire n6582;
wire n6583;
wire n6584;
wire n6585;
wire n6586;
wire n6587;
wire n6588;
wire n6589;
wire n6590;
wire n6591;
wire n6592;
wire n6593;
wire n6594;
wire n6595;
wire n6596;
wire n6597;
wire n6598;
wire n6599;
wire n6600;
wire n6601;
wire n6602;
wire n6603;
wire n6604;
wire n6605;
wire n6606;
wire n6607;
wire n6608;
wire n6609;
wire n6610;
wire n6611;
wire n6612;
wire n6613;
wire n6614;
wire n6615;
wire n6616;
wire n6617;
wire n6618;
wire n6619;
wire n6620;
wire n6621;
wire n6622;
wire n6623;
wire n6624;
wire n6625;
wire n6626;
wire n6627;
wire n6628;
wire n6629;
wire n6630;
wire n6631;
wire n6632;
wire n6633;
wire n6634;
wire n6635;
wire n6636;
wire n6637;
wire n6638;
wire n6639;
wire n6640;
wire n6641;
wire n6642;
wire n6643;
wire n6644;
wire n6645;
wire n6646;
wire n6647;
wire n6648;
wire n6649;
wire n6650;
wire n6651;
wire n6652;
wire n6653;
wire n6654;
wire n6655;
wire n6656;
wire n6657;
wire n6658;
wire n6659;
wire n6660;
wire n6661;
wire n6662;
wire n6663;
wire n6664;
wire n6665;
wire n6666;
wire n6667;
wire n6668;
wire n6669;
wire n6670;
wire n6671;
wire n6672;
wire n6673;
wire n6674;
wire n6675;
wire n6676;
wire n6677;
wire n6678;
wire n6679;
wire n6680;
wire n6681;
wire n6682;
wire n6683;
wire n6684;
wire n6685;
wire n6686;
wire n6687;
wire n6688;
wire n6689;
wire n6690;
wire n6691;
wire n6692;
wire n6693;
wire n6694;
wire n6695;
wire n6696;
wire n6697;
wire n6698;
wire n6699;
wire n6700;
wire n6701;
wire n6702;
wire n6703;
wire n6704;
wire n6705;
wire n6706;
wire n6707;
wire n6708;
wire n6709;
wire n6710;
wire n6711;
wire n6712;
wire n6713;
wire n6714;
wire n6715;
wire n6716;
wire n6717;
wire n6718;
wire n6719;
wire n6720;
wire n6721;
wire n6722;
wire n6723;
wire n6724;
wire n6725;
wire n6726;
wire n6727;
wire n6728;
wire n6729;
wire n6730;
wire n6731;
wire n6732;
wire n6733;
wire n6734;
wire n6735;
wire n6736;
wire n6737;
wire n6738;
wire n6739;
wire n6740;
wire n6741;
wire n6742;
wire n6743;
wire n6744;
wire n6745;
wire n6746;
wire n6747;
wire n6748;
wire n6749;
wire n6750;
wire n6751;
wire n6752;
wire n6753;
wire n6754;
wire n6755;
wire n6756;
wire n6757;
wire n6758;
wire n6759;
wire n6760;
wire n6761;
wire n6762;
wire n6763;
wire n6764;
wire n6765;
wire n6766;
wire n6767;
wire n6768;
wire n6769;
wire n6770;
wire n6771;
wire n6772;
wire n6773;
wire n6774;
wire n6775;
wire n6776;
wire n6777;
wire n6778;
wire n6779;
wire n6780;
wire n6781;
wire n6782;
wire n6783;
wire n6784;
wire n6785;
wire n6786;
wire n6787;
wire n6788;
wire n6789;
wire n6790;
wire n6791;
wire n6792;
wire n6793;
wire n6794;
wire n6795;
wire n6796;
wire n6797;
wire n6798;
wire n6799;
wire n6800;
wire n6801;
wire n6802;
wire n6803;
wire n6804;
wire n6805;
wire n6806;
wire n6807;
wire n6808;
wire n6809;
wire n6810;
wire n6811;
wire n6812;
wire n6813;
wire n6814;
wire n6815;
wire n6816;
wire n6817;
wire n6818;
wire n6819;
wire n6820;
wire n6821;
wire n6822;
wire n6823;
wire n6824;
wire n6825;
wire n6826;
wire n6827;
wire n6828;
wire n6829;
wire n6830;
wire n6831;
wire n6832;
wire n6833;
wire n6834;
wire n6835;
wire n6836;
wire n6837;
wire n6838;
wire n6839;
wire n6840;
wire n6841;
wire n6842;
wire n6843;
wire n6844;
wire n6845;
wire n6846;
wire n6847;
wire n6848;
wire n6849;
wire n6850;
wire n6851;
wire n6852;
wire n6853;
wire n6854;
wire n6855;
wire n6856;
wire n6857;
wire n6858;
wire n6859;
wire n6860;
wire n6861;
wire n6862;
wire n6863;
wire n6864;
wire n6865;
wire n6866;
wire n6867;
wire n6868;
wire n6869;
wire n6870;
wire n6871;
wire n6872;
wire n6873;
wire n6874;
wire n6875;
wire n6876;
wire n6877;
wire n6878;
wire n6879;
wire n6880;
wire n6881;
wire n6882;
wire n6883;
wire n6884;
wire n6885;
wire n6886;
wire n6887;
wire n6888;
wire n6889;
wire n6890;
wire n6891;
wire n6892;
wire n6893;
wire n6894;
wire n6895;
wire n6896;
wire n6897;
wire n6898;
wire n6899;
wire n6900;
wire n6901;
wire n6902;
wire n6903;
wire n6904;
wire n6905;
wire n6906;
wire n6907;
wire n6908;
wire n6909;
wire n6910;
wire n6911;
wire n6912;
wire n6913;
wire n6914;
wire n6915;
wire n6916;
wire n6917;
wire n6918;
wire n6919;
wire n6920;
wire n6921;
wire n6922;
wire n6923;
wire n6924;
wire n6925;
wire n6926;
wire n6927;
wire n6928;
wire n6929;
wire n6930;
wire n6931;
wire n6932;
wire n6933;
wire n6934;
wire n6935;
wire n6936;
wire n6937;
wire n6938;
wire n6939;
wire n6940;
wire n6941;
wire n6942;
wire n6943;
wire n6944;
wire n6945;
wire n6946;
wire n6947;
wire n6948;
wire n6949;
wire n6950;
wire n6951;
wire n6952;
wire n6953;
wire n6954;
wire n6955;
wire n6956;
wire n6957;
wire n6958;
wire n6959;
wire n6960;
wire n6961;
wire n6962;
wire n6963;
wire n6964;
wire n6965;
wire n6966;
wire n6967;
wire n6968;
wire n6969;
wire n6970;
wire n6971;
wire n6972;
wire n6973;
wire n6974;
wire n6975;
wire n6976;
wire n6977;
wire n6978;
wire n6979;
wire n6980;
wire n6981;
wire n6982;
wire n6983;
wire n6984;
wire n6985;
wire n6986;
wire n6987;
wire n6988;
wire n6989;
wire n6990;
wire n6991;
wire n6992;
wire n6993;
wire n6994;
wire n6995;
wire n6996;
wire n6997;
wire n6998;
wire n6999;
wire n7000;
wire n7001;
wire n7002;
wire n7003;
wire n7004;
wire n7005;
wire n7006;
wire n7007;
wire n7008;
wire n7009;
wire n7010;
wire n7011;
wire n7012;
wire n7013;
wire n7014;
wire n7015;
wire n7016;
wire n7017;
wire n7018;
wire n7019;
wire n7020;
wire n7021;
wire n7022;
wire n7023;
wire n7024;
wire n7025;
wire n7026;
wire n7027;
wire n7028;
wire n7029;
wire n7030;
wire n7031;
wire n7032;
wire n7033;
wire n7034;
wire n7035;
wire n7036;
wire n7037;
wire n7038;
wire n7039;
wire n7040;
wire n7041;
wire n7042;
wire n7043;
wire n7044;
wire n7045;
wire n7046;
wire n7047;
wire n7048;
wire n7049;
wire n7050;
wire n7051;
wire n7052;
wire n7053;
wire n7054;
wire n7055;
wire n7056;
wire n7057;
wire n7058;
wire n7059;
wire n7060;
wire n7061;
wire n7062;
wire n7063;
wire n7064;
wire n7065;
wire n7066;
wire n7067;
wire n7068;
wire n7069;
wire n7070;
wire n7071;
wire n7072;
wire n7073;
wire n7074;
wire n7075;
wire n7076;
wire n7077;
wire n7078;
wire n7079;
wire n7080;
wire n7081;
wire n7082;
wire n7083;
wire n7084;
wire n7085;
wire n7086;
wire n7087;
wire n7088;
wire n7089;
wire n7090;
wire n7091;
wire n7092;
wire n7093;
wire n7094;
wire n7095;
wire n7096;
wire n7097;
wire n7098;
wire n7099;
wire n7100;
wire n7101;
wire n7102;
wire n7103;
wire n7104;
wire n7105;
wire n7106;
wire n7107;
wire n7108;
wire n7109;
wire n7110;
wire n7111;
wire n7112;
wire n7113;
wire n7114;
wire n7115;
wire n7116;
wire n7117;
wire n7118;
wire n7119;
wire n7120;
wire n7121;
wire n7122;
wire n7123;
wire n7124;
wire n7125;
wire n7126;
wire n7127;
wire n7128;
wire n7129;
wire n7130;
wire n7131;
wire n7132;
wire n7133;
wire n7134;
wire n7135;
wire n7136;
wire n7137;
wire n7138;
wire n7139;
wire n7140;
wire n7141;
wire n7142;
wire n7143;
wire n7144;
wire n7145;
wire n7146;
wire n7147;
wire n7148;
wire n7149;
wire n7150;
wire n7151;
wire n7152;
wire n7153;
wire n7154;
wire n7155;
wire n7156;
wire n7157;
wire n7158;
wire n7159;
wire n7160;
wire n7161;
wire n7162;
wire n7163;
wire n7164;
wire n7165;
wire n7166;
wire n7167;
wire n7168;
wire n7169;
wire n7170;
wire n7171;
wire n7172;
wire n7173;
wire n7174;
wire n7175;
wire n7176;
wire n7177;
wire n7178;
wire n7179;
wire n7180;
wire n7181;
wire n7182;
wire n7183;
wire n7184;
wire n7185;
wire n7186;
wire n7187;
wire n7188;
wire n7189;
wire n7190;
wire n7191;
wire n7192;
wire n7193;
wire n7194;
wire n7195;
wire n7196;
wire n7197;
wire n7198;
wire n7199;
wire n7200;
wire n7201;
wire n7202;
wire n7203;
wire n7204;
wire n7205;
wire n7206;
wire n7207;
wire n7208;
wire n7209;
wire n7210;
wire n7211;
wire n7212;
wire n7213;
wire n7214;
wire n7215;
wire n7216;
wire n7217;
wire n7218;
wire n7219;
wire n7220;
wire n7221;
wire n7222;
wire n7223;
wire n7224;
wire n7225;
wire n7226;
wire n7227;
wire n7228;
wire n7229;
wire n7230;
wire n7231;
wire n7232;
wire n7233;
wire n7234;
wire n7235;
wire n7236;
wire n7237;
wire n7238;
wire n7239;
wire n7240;
wire n7241;
wire n7242;
wire n7243;
wire n7244;
wire n7245;
wire n7246;
wire n7247;
wire n7248;
wire n7249;
wire n7250;
wire n7251;
wire n7252;
wire n7253;
wire n7254;
wire n7255;
wire n7256;
wire n7257;
wire n7258;
wire n7259;
wire n7260;
wire n7261;
wire n7262;
wire n7263;
wire n7264;
wire n7265;
wire n7266;
wire n7267;
wire n7268;
wire n7269;
wire n7270;
wire n7271;
wire n7272;
wire n7273;
wire n7274;
wire n7275;
wire n7276;
wire n7277;
wire n7278;
wire n7279;
wire n7280;
wire n7281;
wire n7282;
wire n7283;
wire n7284;
wire n7285;
wire n7286;
wire n7287;
wire n7288;
wire n7289;
wire n7290;
wire n7291;
wire n7292;
wire n7293;
wire n7294;
wire n7295;
wire n7296;
wire n7297;
wire n7298;
wire n7299;
wire n7300;
wire n7301;
wire n7302;
wire n7303;
wire n7304;
wire n7305;
wire n7306;
wire n7307;
wire n7308;
wire n7309;
wire n7310;
wire n7311;
wire n7312;
wire n7313;
wire n7314;
wire n7315;
wire n7316;
wire n7317;
wire n7318;
wire n7319;
wire n7320;
wire n7321;
wire n7322;
wire n7323;
wire n7324;
wire n7325;
wire n7326;
wire n7327;
wire n7328;
wire n7329;
wire n7330;
wire n7331;
wire n7332;
wire n7333;
wire n7334;
wire n7335;
wire n7336;
wire n7337;
wire n7338;
wire n7339;
wire n7340;
wire n7341;
wire n7342;
wire n7343;
wire n7344;
wire n7345;
wire n7346;
wire n7347;
wire n7348;
wire n7349;
wire n7350;
wire n7351;
wire n7352;
wire n7353;
wire n7354;
wire n7355;
wire n7356;
wire n7357;
wire n7358;
wire n7359;
wire n7360;
wire n7361;
wire n7362;
wire n7363;
wire n7364;
wire n7365;
wire n7366;
wire n7367;
wire n7368;
wire n7369;
wire n7370;
wire n7371;
wire n7372;
wire n7373;
wire n7374;
wire n7375;
wire n7376;
wire n7377;
wire n7378;
wire n7379;
wire n7380;
wire n7381;
wire n7382;
wire n7383;
wire n7384;
wire n7385;
wire n7386;
wire n7387;
wire n7388;
wire n7389;
wire n7390;
wire n7391;
wire n7392;
wire n7393;
wire n7394;
wire n7395;
wire n7396;
wire n7397;
wire n7398;
wire n7399;
wire n7400;
wire n7401;
wire n7402;
wire n7403;
wire n7404;
wire n7405;
wire n7406;
wire n7407;
wire n7408;
wire n7409;
wire n7410;
wire n7411;
wire n7412;
wire n7413;
wire n7414;
wire n7415;
wire n7416;
wire n7417;
wire n7418;
wire n7419;
wire n7420;
wire n7421;
wire n7422;
wire n7423;
wire n7424;
wire n7425;
wire n7426;
wire n7427;
wire n7428;
wire n7429;
wire n7430;
wire n7431;
wire n7432;
wire n7433;
wire n7434;
wire n7435;
wire n7436;
wire n7437;
wire n7438;
wire n7439;
wire n7440;
wire n7441;
wire n7442;
wire n7443;
wire n7444;
wire n7445;
wire n7446;
wire n7447;
wire n7448;
wire n7449;
wire n7450;
wire n7451;
wire n7452;
wire n7453;
wire n7454;
wire n7455;
wire n7456;
wire n7457;
wire n7458;
wire n7459;
wire n7460;
wire n7461;
wire n7462;
wire n7463;
wire n7464;
wire n7465;
wire n7466;
wire n7467;
wire n7468;
wire n7469;
wire n7470;
wire n7471;
wire n7472;
wire n7473;
wire n7474;
wire n7475;
wire n7476;
wire n7477;
wire n7478;
wire n7479;
wire n7480;
wire n7481;
wire n7482;
wire n7483;
wire n7484;
wire n7485;
wire n7486;
wire n7487;
wire n7488;
wire n7489;
wire n7490;
wire n7491;
wire n7492;
wire n7493;
wire n7494;
wire n7495;
wire n7496;
wire n7497;
wire n7498;
wire n7499;
wire n7500;
wire n7501;
wire n7502;
wire n7503;
wire n7504;
wire n7505;
wire n7506;
wire n7507;
wire n7508;
wire n7509;
wire n7510;
wire n7511;
wire n7512;
wire n7513;
wire n7514;
wire n7515;
wire n7516;
wire n7517;
wire n7518;
wire n7519;
wire n7520;
wire n7521;
wire n7522;
wire n7523;
wire n7524;
wire n7525;
wire n7526;
wire n7527;
wire n7528;
wire n7529;
wire n7530;
wire n7531;
wire n7532;
wire n7533;
wire n7534;
wire n7535;
wire n7536;
wire n7537;
wire n7538;
wire n7539;
wire n7540;
wire n7541;
wire n7542;
wire n7543;
wire n7544;
wire n7545;
wire n7546;
wire n7547;
wire n7548;
wire n7549;
wire n7550;
wire n7551;
wire n7552;
wire n7553;
wire n7554;
wire n7555;
wire n7556;
wire n7557;
wire n7558;
wire n7559;
wire n7560;
wire n7561;
wire n7562;
wire n7563;
wire n7564;
wire n7565;
wire n7566;
wire n7567;
wire n7568;
wire n7569;
wire n7570;
wire n7571;
wire n7572;
wire n7573;
wire n7574;
wire n7575;
wire n7576;
wire n7577;
wire n7578;
wire n7579;
wire n7580;
wire n7581;
wire n7582;
wire n7583;
wire n7584;
wire n7585;
wire n7586;
wire n7587;
wire n7588;
wire n7589;
wire n7590;
wire n7591;
wire n7592;
wire n7593;
wire n7594;
wire n7595;
wire n7596;
wire n7597;
wire n7598;
wire n7599;
wire n7600;
wire n7601;
wire n7602;
wire n7603;
wire n7604;
wire n7605;
wire n7606;
wire n7607;
wire n7608;
wire n7609;
wire n7610;
wire n7611;
wire n7612;
wire n7613;
wire n7614;
wire n7615;
wire n7616;
wire n7617;
wire n7618;
wire n7619;
wire n7620;
wire n7621;
wire n7622;
wire n7623;
wire n7624;
wire n7625;
wire n7626;
wire n7627;
wire n7628;
wire n7629;
wire n7630;
wire n7631;
wire n7632;
wire n7633;
wire n7634;
wire n7635;
wire n7636;
wire n7637;
wire n7638;
wire n7639;
wire n7640;
wire n7641;
wire n7642;
wire n7643;
wire n7644;
wire n7645;
wire n7646;
wire n7647;
wire n7648;
wire n7649;
wire n7650;
wire n7651;
wire n7652;
wire n7653;
wire n7654;
wire n7655;
wire n7656;
wire n7657;
wire n7658;
wire n7659;
wire n7660;
wire n7661;
wire n7662;
wire n7663;
wire n7664;
wire n7665;
wire n7666;
wire n7667;
wire n7668;
wire n7669;
wire n7670;
wire n7671;
wire n7672;
wire n7673;
wire n7674;
wire n7675;
wire n7676;
wire n7677;
wire n7678;
wire n7679;
wire n7680;
wire n7681;
wire n7682;
wire n7683;
wire n7684;
wire n7685;
wire n7686;
wire n7687;
wire n7688;
wire n7689;
wire n7690;
wire n7691;
wire n7692;
wire n7693;
wire n7694;
wire n7695;
wire n7696;
wire n7697;
wire n7698;
wire n7699;
wire n7700;
wire n7701;
wire n7702;
wire n7703;
wire n7704;
wire n7705;
wire n7706;
wire n7707;
wire n7708;
wire n7709;
wire n7710;
wire n7711;
wire n7712;
wire n7713;
wire n7714;
wire n7715;
wire n7716;
wire n7717;
wire n7718;
wire n7719;
wire n7720;
wire n7721;
wire n7722;
wire n7723;
wire n7724;
wire n7725;
wire n7726;
wire n7727;
wire n7728;
wire n7729;
wire n7730;
wire n7731;
wire n7732;
wire n7733;
wire n7734;
wire n7735;
wire n7736;
wire n7737;
wire n7738;
wire n7739;
wire n7740;
wire n7741;
wire n7742;
wire n7743;
wire n7744;
wire n7745;
wire n7746;
wire n7747;
wire n7748;
wire n7749;
wire n7750;
wire n7751;
wire n7752;
wire n7753;
wire n7754;
wire n7755;
wire n7756;
wire n7757;
wire n7758;
wire n7759;
wire n7760;
wire n7761;
wire n7762;
wire n7763;
wire n7764;
wire n7765;
wire n7766;
wire n7767;
wire n7768;
wire n7769;
wire n7770;
wire n7771;
wire n7772;
wire n7773;
wire n7774;
wire n7775;
wire n7776;
wire n7777;
wire n7778;
wire n7779;
wire n7780;
wire n7781;
wire n7782;
wire n7783;
wire n7784;
wire n7785;
wire n7786;
wire n7787;
wire n7788;
wire n7789;
wire n7790;
wire n7791;
wire n7792;
wire n7793;
wire n7794;
wire n7795;
wire n7796;
wire n7797;
wire n7798;
wire n7799;
wire n7800;
wire n7801;
wire n7802;
wire n7803;
wire n7804;
wire n7805;
wire n7806;
wire n7807;
wire n7808;
wire n7809;
wire n7810;
wire n7811;
wire n7812;
wire n7813;
wire n7814;
wire n7815;
wire n7816;
wire n7817;
wire n7818;
wire n7819;
wire n7820;
wire n7821;
wire n7822;
wire n7823;
wire n7824;
wire n7825;
wire n7826;
wire n7827;
wire n7828;
wire n7829;
wire n7830;
wire n7831;
wire n7832;
wire n7833;
wire n7834;
wire n7835;
wire n7836;
wire n7837;
wire n7838;
wire n7839;
wire n7840;
wire n7841;
wire n7842;
wire n7843;
wire n7844;
wire n7845;
wire n7846;
wire n7847;
wire n7848;
wire n7849;
wire n7850;
wire n7851;
wire n7852;
wire n7853;
wire n7854;
wire n7855;
wire n7856;
wire n7857;
wire n7858;
wire n7859;
wire n7860;
wire n7861;
wire n7862;
wire n7863;
wire n7864;
wire n7865;
wire n7866;
wire n7867;
wire n7868;
wire n7869;
wire n7870;
wire n7871;
wire n7872;
wire n7873;
wire n7874;
wire n7875;
wire n7876;
wire n7877;
wire n7878;
wire n7879;
wire n7880;
wire n7881;
wire n7882;
wire n7883;
wire n7884;
wire n7885;
wire n7886;
wire n7887;
wire n7888;
wire n7889;
wire n7890;
wire n7891;
wire n7892;
wire n7893;
wire n7894;
wire n7895;
wire n7896;
wire n7897;
wire n7898;
wire n7899;
wire n7900;
wire n7901;
wire n7902;
wire n7903;
wire n7904;
wire n7905;
wire n7906;
wire n7907;
wire n7908;
wire n7909;
wire n7910;
wire n7911;
wire n7912;
wire n7913;
wire n7914;
wire n7915;
wire n7916;
wire n7917;
wire n7918;
wire n7919;
wire n7920;
wire n7921;
wire n7922;
wire n7923;
wire n7924;
wire n7925;
wire n7926;
wire n7927;
wire n7928;
wire n7929;
wire n7930;
wire n7931;
wire n7932;
wire n7933;
wire n7934;
wire n7935;
wire n7936;
wire n7937;
wire n7938;
wire n7939;
wire n7940;
wire n7941;
wire n7942;
wire n7943;
wire n7944;
wire n7945;
wire n7946;
wire n7947;
wire n7948;
wire n7949;
wire n7950;
wire n7951;
wire n7952;
wire n7953;
wire n7954;
wire n7955;
wire n7956;
wire n7957;
wire n7958;
wire n7959;
wire n7960;
wire n7961;
wire n7962;
wire n7963;
wire n7964;
wire n7965;
wire n7966;
wire n7967;
wire n7968;
wire n7969;
wire n7970;
wire n7971;
wire n7972;
wire n7973;
wire n7974;
wire n7975;
wire n7976;
wire n7977;
wire n7978;
wire n7979;
wire n7980;
wire n7981;
wire n7982;
wire n7983;
wire n7984;
wire n7985;
wire n7986;
wire n7987;
wire n7988;
wire n7989;
wire n7990;
wire n7991;
wire n7992;
wire n7993;
wire n7994;
wire n7995;
wire n7996;
wire n7997;
wire n7998;
wire n7999;
wire n8000;
wire n8001;
wire n8002;
wire n8003;
wire n8004;
wire n8005;
wire n8006;
wire n8007;
wire n8008;
wire n8009;
wire n8010;
wire n8011;
wire n8012;
wire n8013;
wire n8014;
wire n8015;
wire n8016;
wire n8017;
wire n8018;
wire n8019;
wire n8020;
wire n8021;
wire n8022;
wire n8023;
wire n8024;
wire n8025;
wire n8026;
wire n8027;
wire n8028;
wire n8029;
wire n8030;
wire n8031;
wire n8032;
wire n8033;
wire n8034;
wire n8035;
wire n8036;
wire n8037;
wire n8038;
wire n8039;
wire n8040;
wire n8041;
wire n8042;
wire n8043;
wire n8044;
wire n8045;
wire n8046;
wire n8047;
wire n8048;
wire n8049;
wire n8050;
wire n8051;
wire n8052;
wire n8053;
wire n8054;
wire n8055;
wire n8056;
wire n8057;
wire n8058;
wire n8059;
wire n8060;
wire n8061;
wire n8062;
wire n8063;
wire n8064;
wire n8065;
wire n8066;
wire n8067;
wire n8068;
wire n8069;
wire n8070;
wire n8071;
wire n8072;
wire n8073;
wire n8074;
wire n8075;
wire n8076;
wire n8077;
wire n8078;
wire n8079;
wire n8080;
wire n8081;
wire n8082;
wire n8083;
wire n8084;
wire n8085;
wire n8086;
wire n8087;
wire n8088;
wire n8089;
wire n8090;
wire n8091;
wire n8092;
wire n8093;
wire n8094;
wire n8095;
wire n8096;
wire n8097;
wire n8098;
wire n8099;
wire n8100;
wire n8101;
wire n8102;
wire n8103;
wire n8104;
wire n8105;
wire n8106;
wire n8107;
wire n8108;
wire n8109;
wire n8110;
wire n8111;
wire n8112;
wire n8113;
wire n8114;
wire n8115;
wire n8116;
wire n8117;
wire n8118;
wire n8119;
wire n8120;
wire n8121;
wire n8122;
wire n8123;
wire n8124;
wire n8125;
wire n8126;
wire n8127;
wire n8128;
wire n8129;
wire n8130;
wire n8131;
wire n8132;
wire n8133;
wire n8134;
wire n8135;
wire n8136;
wire n8137;
wire n8138;
wire n8139;
wire n8140;
wire n8141;
wire n8142;
wire n8143;
wire n8144;
wire n8145;
wire n8146;
wire n8147;
wire n8148;
wire n8149;
wire n8150;
wire n8151;
wire n8152;
wire n8153;
wire n8154;
wire n8155;
wire n8156;
wire n8157;
wire n8158;
wire n8159;
wire n8160;
wire n8161;
wire n8162;
wire n8163;
wire n8164;
wire n8165;
wire n8166;
wire n8167;
wire n8168;
wire n8169;
wire n8170;
wire n8171;
wire n8172;
wire n8173;
wire n8174;
wire n8175;
wire n8176;
wire n8177;
wire n8178;
wire n8179;
wire n8180;
wire n8181;
wire n8182;
wire n8183;
wire n8184;
wire n8185;
wire n8186;
wire n8187;
wire n8188;
wire n8189;
wire n8190;
wire n8191;
wire n8192;
wire n8193;
wire n8194;
wire n8195;
wire n8196;
wire n8197;
wire n8198;
wire n8199;
wire n8200;
wire n8201;
wire n8202;
wire n8203;
wire n8204;
wire n8205;
wire n8206;
wire n8207;
wire n8208;
wire n8209;
wire n8210;
wire n8211;
wire n8212;
wire n8213;
wire n8214;
wire n8215;
wire n8216;
wire n8217;
wire n8218;
wire n8219;
wire n8220;
wire n8221;
wire n8222;
wire n8223;
wire n8224;
wire n8225;
wire n8226;
wire n8227;
wire n8228;
wire n8229;
wire n8230;
wire n8231;
wire n8232;
wire n8233;
wire n8234;
wire n8235;
wire n8236;
wire n8237;
wire n8238;
wire n8239;
wire n8240;
wire n8241;
wire n8242;
wire n8243;
wire n8244;
wire n8245;
wire n8246;
wire n8247;
wire n8248;
wire n8249;
wire n8250;
wire n8251;
wire n8252;
wire n8253;
wire n8254;
wire n8255;
wire n8256;
wire n8257;
wire n8258;
wire n8259;
wire n8260;
wire n8261;
wire n8262;
wire n8263;
wire n8264;
wire n8265;
wire n8266;
wire n8267;
wire n8268;
wire n8269;
wire n8270;
wire n8271;
wire n8272;
wire n8273;
wire n8274;
wire n8275;
wire n8276;
wire n8277;
wire n8278;
wire n8279;
wire n8280;
wire n8281;
wire n8282;
wire n8283;
wire n8284;
wire n8285;
wire n8286;
wire n8287;
wire n8288;
wire n8289;
wire n8290;
wire n8291;
wire n8292;
wire n8293;
wire n8294;
wire n8295;
wire n8296;
wire n8297;
wire n8298;
wire n8299;
wire n8300;
wire n8301;
wire n8302;
wire n8303;
wire n8304;
wire n8305;
wire n8306;
wire n8307;
wire n8308;
wire n8309;
wire n8310;
wire n8311;
wire n8312;
wire n8313;
wire n8314;
wire n8315;
wire n8316;
wire n8317;
wire n8318;
wire n8319;
wire n8320;
wire n8321;
wire n8322;
wire n8323;
wire n8324;
wire n8325;
wire n8326;
wire n8327;
wire n8328;
wire n8329;
wire n8330;
wire n8331;
wire n8332;
wire n8333;
wire n8334;
wire n8335;
wire n8336;
wire n8337;
wire n8338;
wire n8339;
wire n8340;
wire n8341;
wire n8342;
wire n8343;
wire n8344;
wire n8345;
wire n8346;
wire n8347;
wire n8348;
wire n8349;
wire n8350;
wire n8351;
wire n8352;
wire n8353;
wire n8354;
wire n8355;
wire n8356;
wire n8357;
wire n8358;
wire n8359;
wire n8360;
wire n8361;
wire n8362;
wire n8363;
wire n8364;
wire n8365;
wire n8366;
wire n8367;
wire n8368;
wire n8369;
wire n8370;
wire n8371;
wire n8372;
wire n8373;
wire n8374;
wire n8375;
wire n8376;
wire n8377;
wire n8378;
wire n8379;
wire n8380;
wire n8381;
wire n8382;
wire n8383;
wire n8384;
wire n8385;
wire n8386;
wire n8387;
wire n8388;
wire n8389;
wire n8390;
wire n8391;
wire n8392;
wire n8393;
wire n8394;
wire n8395;
wire n8396;
wire n8397;
wire n8398;
wire n8399;
wire n8400;
wire n8401;
wire n8402;
wire n8403;
wire n8404;
wire n8405;
wire n8406;
wire n8407;
wire n8408;
wire n8409;
wire n8410;
wire n8411;
wire n8412;
wire n8413;
wire n8414;
wire n8415;
wire n8416;
wire n8417;
wire n8418;
wire n8419;
wire n8420;
wire n8421;
wire n8422;
wire n8423;
wire n8424;
wire n8425;
wire n8426;
wire n8427;
wire n8428;
wire n8429;
wire n8430;
wire n8431;
wire n8432;
wire n8433;
wire n8434;
wire n8435;
wire n8436;
wire n8437;
wire n8438;
wire n8439;
wire n8440;
wire n8441;
wire n8442;
wire n8443;
wire n8444;
wire n8445;
wire n8446;
wire n8447;
wire n8448;
wire n8449;
wire n8450;
wire n8451;
wire n8452;
wire n8453;
wire n8454;
wire n8455;
wire n8456;
wire n8457;
wire n8458;
wire n8459;
wire n8460;
wire n8461;
wire n8462;
wire n8463;
wire n8464;
wire n8465;
wire n8466;
wire n8467;
wire n8468;
wire n8469;
wire n8470;
wire n8471;
wire n8472;
wire n8473;
wire n8474;
wire n8475;
wire n8476;
wire n8477;
wire n8478;
wire n8479;
wire n8480;
wire n8481;
wire n8482;
wire n8483;
wire n8484;
wire n8485;
wire n8486;
wire n8487;
wire n8488;
wire n8489;
wire n8490;
wire n8491;
wire n8492;
wire n8493;
wire n8494;
wire n8495;
wire n8496;
wire n8497;
wire n8498;
wire n8499;
wire n8500;
wire n8501;
wire n8502;
wire n8503;
wire n8504;
wire n8505;
wire n8506;
wire n8507;
wire n8508;
wire n8509;
wire n8510;
wire n8511;
wire n8512;
wire n8513;
wire n8514;
wire n8515;
wire n8516;
wire n8517;
wire n8518;
wire n8519;
wire n8520;
wire n8521;
wire n8522;
wire n8523;
wire n8524;
wire n8525;
wire n8526;
wire n8527;
wire n8528;
wire n8529;
wire n8530;
wire n8531;
wire n8532;
wire n8533;
wire n8534;
wire n8535;
wire n8536;
wire n8537;
wire n8538;
wire n8539;
wire n8540;
wire n8541;
wire n8542;
wire n8543;
wire n8544;
wire n8545;
wire n8546;
wire n8547;
wire n8548;
wire n8549;
wire n8550;
wire n8551;
wire n8552;
wire n8553;
wire n8554;
wire n8555;
wire n8556;
wire n8557;
wire n8558;
wire n8559;
wire n8560;
wire n8561;
wire n8562;
wire n8563;
wire n8564;
wire n8565;
wire n8566;
wire n8567;
wire n8568;
wire n8569;
wire n8570;
wire n8571;
wire n8572;
wire n8573;
wire n8574;
wire n8575;
wire n8576;
wire n8577;
wire n8578;
wire n8579;
wire n8580;
wire n8581;
wire n8582;
wire n8583;
wire n8584;
wire n8585;
wire n8586;
wire n8587;
wire n8588;
wire n8589;
wire n8590;
wire n8591;
wire n8592;
wire n8593;
wire n8594;
wire n8595;
wire n8596;
wire n8597;
wire n8598;
wire n8599;
wire n8600;
wire n8601;
wire n8602;
wire n8603;
wire n8604;
wire n8605;
wire n8606;
wire n8607;
wire n8608;
wire n8609;
wire n8610;
wire n8611;
wire n8612;
wire n8613;
wire n8614;
wire n8615;
wire n8616;
wire n8617;
wire n8618;
wire n8619;
wire n8620;
wire n8621;
wire n8622;
wire n8623;
wire n8624;
wire n8625;
wire n8626;
wire n8627;
wire n8628;
wire n8629;
wire n8630;
wire n8631;
wire n8632;
wire n8633;
wire n8634;
wire n8635;
wire n8636;
wire n8637;
wire n8638;
wire n8639;
wire n8640;
wire n8641;
wire n8642;
wire n8643;
wire n8644;
wire n8645;
wire n8646;
wire n8647;
wire n8648;
wire n8649;
wire n8650;
wire n8651;
wire n8652;
wire n8653;
wire n8654;
wire n8655;
wire n8656;
wire n8657;
wire n8658;
wire n8659;
wire n8660;
wire n8661;
wire n8662;
wire n8663;
wire n8664;
wire n8665;
wire n8666;
wire n8667;
wire n8668;
wire n8669;
wire n8670;
wire n8671;
wire n8672;
wire n8673;
wire n8674;
wire n8675;
wire n8676;
wire n8677;
wire n8678;
wire n8679;
wire n8680;
wire n8681;
wire n8682;
wire n8683;
wire n8684;
wire n8685;
wire n8686;
wire n8687;
wire n8688;
wire n8689;
wire n8690;
wire n8691;
wire n8692;
wire n8693;
wire n8694;
wire n8695;
wire n8696;
wire n8697;
wire n8698;
wire n8699;
wire n8700;
wire n8701;
wire n8702;
wire n8703;
wire n8704;
wire n8705;
wire n8706;
wire n8707;
wire n8708;
wire n8709;
wire n8710;
wire n8711;
wire n8712;
wire n8713;
wire n8714;
wire n8715;
wire n8716;
wire n8717;
wire n8718;
wire n8719;
wire n8720;
wire n8721;
wire n8722;
wire n8723;
wire n8724;
wire n8725;
wire n8726;
wire n8727;
wire n8728;
wire n8729;
wire n8730;
wire n8731;
wire n8732;
wire n8733;
wire n8734;
wire n8735;
wire n8736;
wire n8737;
wire n8738;
wire n8739;
wire n8740;
wire n8741;
wire n8742;
wire n8743;
wire n8744;
wire n8745;
wire n8746;
wire n8747;
wire n8748;
wire n8749;
wire n8750;
wire n8751;
wire n8752;
wire n8753;
wire n8754;
wire n8755;
wire n8756;
wire n8757;
wire n8758;
wire n8759;
wire n8760;
wire n8761;
wire n8762;
wire n8763;
wire n8764;
wire n8765;
wire n8766;
wire n8767;
wire n8768;
wire n8769;
wire n8770;
wire n8771;
wire n8772;
wire n8773;
wire n8774;
wire n8775;
wire n8776;
wire n8777;
wire n8778;
wire n8779;
wire n8780;
wire n8781;
wire n8782;
wire n8783;
wire n8784;
wire n8785;
wire n8786;
wire n8787;
wire n8788;
wire n8789;
wire n8790;
wire n8791;
wire n8792;
wire n8793;
wire n8794;
wire n8795;
wire n8796;
wire n8797;
wire n8798;
wire n8799;
wire n8800;
wire n8801;
wire n8802;
wire n8803;
wire n8804;
wire n8805;
wire n8806;
wire n8807;
wire n8808;
wire n8809;
wire n8810;
wire n8811;
wire n8812;
wire n8813;
wire n8814;
wire n8815;
wire n8816;
wire n8817;
wire n8818;
wire n8819;
wire n8820;
wire n8821;
wire n8822;
wire n8823;
wire n8824;
wire n8825;
wire n8826;
wire n8827;
wire n8828;
wire n8829;
wire n8830;
wire n8831;
wire n8832;
wire n8833;
wire n8834;
wire n8835;
wire n8836;
wire n8837;
wire n8838;
wire n8839;
wire n8840;
wire n8841;
wire n8842;
wire n8843;
wire n8844;
wire n8845;
wire n8846;
wire n8847;
wire n8848;
wire n8849;
wire n8850;
wire n8851;
wire n8852;
wire n8853;
wire n8854;
wire n8855;
wire n8856;
wire n8857;
wire n8858;
wire n8859;
wire n8860;
wire n8861;
wire n8862;
wire n8863;
wire n8864;
wire n8865;
wire n8866;
wire n8867;
wire n8868;
wire n8869;
wire n8870;
wire n8871;
wire n8872;
wire n8873;
wire n8874;
wire n8875;
wire n8876;
wire n8877;
wire n8878;
wire n8879;
wire n8880;
wire n8881;
wire n8882;
wire n8883;
wire n8884;
wire n8885;
wire n8886;
wire n8887;
wire n8888;
wire n8889;
wire n8890;
wire n8891;
wire n8892;
wire n8893;
wire n8894;
wire n8895;
wire n8896;
wire n8897;
wire n8898;
wire n8899;
wire n8900;
wire n8901;
wire n8902;
wire n8903;
wire n8904;
wire n8905;
wire n8906;
wire n8907;
wire n8908;
wire n8909;
wire n8910;
wire n8911;
wire n8912;
wire n8913;
wire n8914;
wire n8915;
wire n8916;
wire n8917;
wire n8918;
wire n8919;
wire n8920;
wire n8921;
wire n8922;
wire n8923;
wire n8924;
wire n8925;
wire n8926;
wire n8927;
wire n8928;
wire n8929;
wire n8930;
wire n8931;
wire n8932;
wire n8933;
wire n8934;
wire n8935;
wire n8936;
wire n8937;
wire n8938;
wire n8939;
wire n8940;
wire n8941;
wire n8942;
wire n8943;
wire n8944;
wire n8945;
wire n8946;
wire n8947;
wire n8948;
wire n8949;
wire n8950;
wire n8951;
wire n8952;
wire n8953;
wire n8954;
wire n8955;
wire n8956;
wire n8957;
wire n8958;
wire n8959;
wire n8960;
wire n8961;
wire n8962;
wire n8963;
wire n8964;
wire n8965;
wire n8966;
wire n8967;
wire n8968;
wire n8969;
wire n8970;
wire n8971;
wire n8972;
wire n8973;
wire n8974;
wire n8975;
wire n8976;
wire n8977;
wire n8978;
wire n8979;
wire n8980;
wire n8981;
wire n8982;
wire n8983;
wire n8984;
wire n8985;
wire n8986;
wire n8987;
wire n8988;
wire n8989;
wire n8990;
wire n8991;
wire n8992;
wire n8993;
wire n8994;
wire n8995;
wire n8996;
wire n8997;
wire n8998;
wire n8999;
wire n9000;
wire n9001;
wire n9002;
wire n9003;
wire n9004;
wire n9005;
wire n9006;
wire n9007;
wire n9008;
wire n9009;
wire n9010;
wire n9011;
wire n9012;
wire n9013;
wire n9014;
wire n9015;
wire n9016;
wire n9017;
wire n9018;
wire n9019;
wire n9020;
wire n9021;
wire n9022;
wire n9023;
wire n9024;
wire n9025;
wire n9026;
wire n9027;
wire n9028;
wire n9029;
wire n9030;
wire n9031;
wire n9032;
wire n9033;
wire n9034;
wire n9035;
wire n9036;
wire n9037;
wire n9038;
wire n9039;
wire n9040;
wire n9041;
wire n9042;
wire n9043;
wire n9044;
wire n9045;
wire n9046;
wire n9047;
wire n9048;
wire n9049;
wire n9050;
wire n9051;
wire n9052;
wire n9053;
wire n9054;
wire n9055;
wire n9056;
wire n9057;
wire n9058;
wire n9059;
wire n9060;
wire n9061;
wire n9062;
wire n9063;
wire n9064;
wire n9065;
wire n9066;
wire n9067;
wire n9068;
wire n9069;
wire n9070;
wire n9071;
wire n9072;
wire n9073;
wire n9074;
wire n9075;
wire n9076;
wire n9077;
wire n9078;
wire n9079;
wire n9080;
wire n9081;
wire n9082;
wire n9083;
wire n9084;
wire n9085;
wire n9086;
wire n9087;
wire n9088;
wire n9089;
wire n9090;
wire n9091;
wire n9092;
wire n9093;
wire n9094;
wire n9095;
wire n9096;
wire n9097;
wire n9098;
wire n9099;
wire n9100;
wire n9101;
wire n9102;
wire n9103;
wire n9104;
wire n9105;
wire n9106;
wire n9107;
wire n9108;
wire n9109;
wire n9110;
wire n9111;
wire n9112;
wire n9113;
wire n9114;
wire n9115;
wire n9116;
wire n9117;
wire n9118;
wire n9119;
wire n9120;
wire n9121;
wire n9122;
wire n9123;
wire n9124;
wire n9125;
wire n9126;
wire n9127;
wire n9128;
wire n9129;
wire n9130;
wire n9131;
wire n9132;
wire n9133;
wire n9134;
wire n9135;
wire n9136;
wire n9137;
wire n9138;
wire n9139;
wire n9140;
wire n9141;
wire n9142;
wire n9143;
wire n9144;
wire n9145;
wire n9146;
wire n9147;
wire n9148;
wire n9149;
wire n9150;
wire n9151;
wire n9152;
wire n9153;
wire n9154;
wire n9155;
wire n9156;
wire n9157;
wire n9158;
wire n9159;
wire n9160;
wire n9161;
wire n9162;
wire n9163;
wire n9164;
wire n9165;
wire n9166;
wire n9167;
wire n9168;
wire n9169;
wire n9170;
wire n9171;
wire n9172;
wire n9173;
wire n9174;
wire n9175;
wire n9176;
wire n9177;
wire n9178;
wire n9179;
wire n9180;
wire n9181;
wire n9182;
wire n9183;
wire n9184;
wire n9185;
wire n9186;
wire n9187;
wire n9188;
wire n9189;
wire n9190;
wire n9191;
wire n9192;
wire n9193;
wire n9194;
wire n9195;
wire n9196;
wire n9197;
wire n9198;
wire n9199;
wire n9200;
wire n9201;
wire n9202;
wire n9203;
wire n9204;
wire n9205;
wire n9206;
wire n9207;
wire n9208;
wire n9209;
wire n9210;
wire n9211;
wire n9212;
wire n9213;
wire n9214;
wire n9215;
wire n9216;
wire n9217;
wire n9218;
wire n9219;
wire n9220;
wire n9221;
wire n9222;
wire n9223;
wire n9224;
wire n9225;
wire n9226;
wire n9227;
wire n9228;
wire n9229;
wire n9230;
wire n9231;
wire n9232;
wire n9233;
wire n9234;
wire n9235;
wire n9236;
wire n9237;
wire n9238;
wire n9239;
wire n9240;
wire n9241;
wire n9242;
wire n9243;
wire n9244;
wire n9245;
wire n9246;
wire n9247;
wire n9248;
wire n9249;
wire n9250;
wire n9251;
wire n9252;
wire n9253;
wire n9254;
wire n9255;
wire n9256;
wire n9257;
wire n9258;
wire n9259;
wire n9260;
wire n9261;
wire n9262;
wire n9263;
wire n9264;
wire n9265;
wire n9266;
wire n9267;
wire n9268;
wire n9269;
wire n9270;
wire n9271;
wire n9272;
wire n9273;
wire n9274;
wire n9275;
wire n9276;
wire n9277;
wire n9278;
wire n9279;
wire n9280;
wire n9281;
wire n9282;
wire n9283;
wire n9284;
wire n9285;
wire n9286;
wire n9287;
wire n9288;
wire n9289;
wire n9290;
wire n9291;
wire n9292;
wire n9293;
wire n9294;
wire n9295;
wire n9296;
wire n9297;
wire n9298;
wire n9299;
wire n9300;
wire n9301;
wire n9302;
wire n9303;
wire n9304;
wire n9305;
wire n9306;
wire n9307;
wire n9308;
wire n9309;
wire n9310;
wire n9311;
wire n9312;
wire n9313;
wire n9314;
wire n9315;
wire n9316;
wire n9317;
wire n9318;
wire n9319;
wire n9320;
wire n9321;
wire n9322;
wire n9323;
wire n9324;
wire n9325;
wire n9326;
wire n9327;
wire n9328;
wire n9329;
wire n9330;
wire n9331;
wire n9332;
wire n9333;
wire n9334;
wire n9335;
wire n9336;
wire n9337;
wire n9338;
wire n9339;
wire n9340;
wire n9341;
wire n9342;
wire n9343;
wire n9344;
wire n9345;
wire n9346;
wire n9347;
wire n9348;
wire n9349;
wire n9350;
wire n9351;
wire n9352;
wire n9353;
wire n9354;
wire n9355;
wire n9356;
wire n9357;
wire n9358;
wire n9359;
wire n9360;
wire n9361;
wire n9362;
wire n9363;
wire n9364;
wire n9365;
wire n9366;
wire n9367;
wire n9368;
wire n9369;
wire n9370;
wire n9371;
wire n9372;
wire n9373;
wire n9374;
wire n9375;
wire n9376;
wire n9377;
wire n9378;
wire n9379;
wire n9380;
wire n9381;
wire n9382;
wire n9383;
wire n9384;
wire n9385;
wire n9386;
wire n9387;
wire n9388;
wire n9389;
wire n9390;
wire n9391;
wire n9392;
wire n9393;
wire n9394;
wire n9395;
wire n9396;
wire n9397;
wire n9398;
wire n9399;
wire n9400;
wire n9401;
wire n9402;
wire n9403;
wire n9404;
wire n9405;
wire n9406;
wire n9407;
wire n9408;
wire n9409;
wire n9410;
wire n9411;
wire n9412;
wire n9413;
wire n9414;
wire n9415;
wire n9416;
wire n9417;
wire n9418;
wire n9419;
wire n9420;
wire n9421;
wire n9422;
wire n9423;
wire n9424;
wire n9425;
wire n9426;
wire n9427;
wire n9428;
wire n9429;
wire n9430;
wire n9431;
wire n9432;
wire n9433;
wire n9434;
wire n9435;
wire n9436;
wire n9437;
wire n9438;
wire n9439;
wire n9440;
wire n9441;
wire n9442;
wire n9443;
wire n9444;
wire n9445;
wire n9446;
wire n9447;
wire n9448;
wire n9449;
wire n9450;
wire n9451;
wire n9452;
wire n9453;
wire n9454;
wire n9455;
wire n9456;
wire n9457;
wire n9458;
wire n9459;
wire n9460;
wire n9461;
wire n9462;
wire n9463;
wire n9464;
wire n9465;
wire n9466;
wire n9467;
wire n9468;
wire n9469;
wire n9470;
wire n9471;
wire n9472;
wire n9473;
wire n9474;
wire n9475;
wire n9476;
wire n9477;
wire n9478;
wire n9479;
wire n9480;
wire n9481;
wire n9482;
wire n9483;
wire n9484;
wire n9485;
wire n9486;
wire n9487;
wire n9488;
wire n9489;
wire n9490;
wire n9491;
wire n9492;
wire n9493;
wire n9494;
wire n9495;
wire n9496;
wire n9497;
wire n9498;
wire n9499;
wire n9500;
wire n9501;
wire n9502;
wire n9503;
wire n9504;
wire n9505;
wire n9506;
wire n9507;
wire n9508;
wire n9509;
wire n9510;
wire n9511;
wire n9512;
wire n9513;
wire n9514;
wire n9515;
wire n9516;
wire n9517;
wire n9518;
wire n9519;
wire n9520;
wire n9521;
wire n9522;
wire n9523;
wire n9524;
wire n9525;
wire n9526;
wire n9527;
wire n9528;
wire n9529;
wire n9530;
wire n9531;
wire n9532;
wire n9533;
wire n9534;
wire n9535;
wire n9536;
wire n9537;
wire n9538;
wire n9539;
wire n9540;
wire n9541;
wire n9542;
wire n9543;
wire n9544;
wire n9545;
wire n9546;
wire n9547;
wire n9548;
wire n9549;
wire n9550;
wire n9551;
wire n9552;
wire n9553;
wire n9554;
wire n9555;
wire n9556;
wire n9557;
wire n9558;
wire n9559;
wire n9560;
wire n9561;
wire n9562;
wire n9563;
wire n9564;
wire n9565;
wire n9566;
wire n9567;
wire n9568;
wire n9569;
wire n9570;
wire n9571;
wire n9572;
wire n9573;
wire n9574;
wire n9575;
wire n9576;
wire n9577;
wire n9578;
wire n9579;
wire n9580;
wire n9581;
wire n9582;
wire n9583;
wire n9584;
wire n9585;
wire n9586;
wire n9587;
wire n9588;
wire n9589;
wire n9590;
wire n9591;
wire n9592;
wire n9593;
wire n9594;
wire n9595;
wire n9596;
wire n9597;
wire n9598;
wire n9599;
wire n9600;
wire n9601;
wire n9602;
wire n9603;
wire n9604;
wire n9605;
wire n9606;
wire n9607;
wire n9608;
wire n9609;
wire n9610;
wire n9611;
wire n9612;
wire n9613;
wire n9614;
wire n9615;
wire n9616;
wire n9617;
wire n9618;
wire n9619;
wire n9620;
wire n9621;
wire n9622;
wire n9623;
wire n9624;
wire n9625;
wire n9626;
wire n9627;
wire n9628;
wire n9629;
wire n9630;
wire n9631;
wire n9632;
wire n9633;
wire n9634;
wire n9635;
wire n9636;
wire n9637;
wire n9638;
wire n9639;
wire n9640;
wire n9641;
wire n9642;
wire n9643;
wire n9644;
wire n9645;
wire n9646;
wire n9647;
wire n9648;
wire n9649;
wire n9650;
wire n9651;
wire n9652;
wire n9653;
wire n9654;
wire n9655;
wire n9656;
wire n9657;
wire n9658;
wire n9659;
wire n9660;
wire n9661;
wire n9662;
wire n9663;
wire n9664;
wire n9665;
wire n9666;
wire n9667;
wire n9668;
wire n9669;
wire n9670;
wire n9671;
wire n9672;
wire n9673;
wire n9674;
wire n9675;
wire n9676;
wire n9677;
wire n9678;
wire n9679;
wire n9680;
wire n9681;
wire n9682;
wire n9683;
wire n9684;
wire n9685;
wire n9686;
wire n9687;
wire n9688;
wire n9689;
wire n9690;
wire n9691;
wire n9692;
wire n9693;
wire n9694;
wire n9695;
wire n9696;
wire n9697;
wire n9698;
wire n9699;
wire n9700;
wire n9701;
wire n9702;
wire n9703;
wire n9704;
wire n9705;
wire n9706;
wire n9707;
wire n9708;
wire n9709;
wire n9710;
wire n9711;
wire n9712;
wire n9713;
wire n9714;
wire n9715;
wire n9716;
wire n9717;
wire n9718;
wire n9719;
wire n9720;
wire n9721;
wire n9722;
wire n9723;
wire n9724;
wire n9725;
wire n9726;
wire n9727;
wire n9728;
wire n9729;
wire n9730;
wire n9731;
wire n9732;
wire n9733;
wire n9734;
wire n9735;
wire n9736;
wire n9737;
wire n9738;
wire n9739;
wire n9740;
wire n9741;
wire n9742;
wire n9743;
wire n9744;
wire n9745;
wire n9746;
wire n9747;
wire n9748;
wire n9749;
wire n9750;
wire n9751;
wire n9752;
wire n9753;
wire n9754;
wire n9755;
wire n9756;
wire n9757;
wire n9758;
wire n9759;
wire n9760;
wire n9761;
wire n9762;
wire n9763;
wire n9764;
wire n9765;
wire n9766;
wire n9767;
wire n9768;
wire n9769;
wire n9770;
wire n9771;
wire n9772;
wire n9773;
wire n9774;
wire n9775;
wire n9776;
wire n9777;
wire n9778;
wire n9779;
wire n9780;
wire n9781;
wire n9782;
wire n9783;
wire n9784;
wire n9785;
wire n9786;
wire n9787;
wire n9788;
wire n9789;
wire n9790;
wire n9791;
wire n9792;
wire n9793;
wire n9794;
wire n9795;
wire n9796;
wire n9797;
wire n9798;
wire n9799;
wire n9800;
wire n9801;
wire n9802;
wire n9803;
wire n9804;
wire n9805;
wire n9806;
wire n9807;
wire n9808;
wire n9809;
wire n9810;
wire n9811;
wire n9812;
wire n9813;
wire n9814;
wire n9815;
wire n9816;
wire n9817;
wire n9818;
wire n9819;
wire n9820;
wire n9821;
wire n9822;
wire n9823;
wire n9824;
wire n9825;
wire n9826;
wire n9827;
wire n9828;
wire n9829;
wire n9830;
wire n9831;
wire n9832;
wire n9833;
wire n9834;
wire n9835;
wire n9836;
wire n9837;
wire n9838;
wire n9839;
wire n9840;
wire n9841;
wire n9842;
wire n9843;
wire n9844;
wire n9845;
wire n9846;
wire n9847;
wire n9848;
wire n9849;
wire n9850;
wire n9851;
wire n9852;
wire n9853;
wire n9854;
wire n9855;
wire n9856;
wire n9857;
wire n9858;
wire n9859;
wire n9860;
wire n9861;
wire n9862;
wire n9863;
wire n9864;
wire n9865;
wire n9866;
wire n9867;
wire n9868;
wire n9869;
wire n9870;
wire n9871;
wire n9872;
wire n9873;
wire n9874;
wire n9875;
wire n9876;
wire n9877;
wire n9878;
wire n9879;
wire n9880;
wire n9881;
wire n9882;
wire n9883;
wire n9884;
wire n9885;
wire n9886;
wire n9887;
wire n9888;
wire n9889;
wire n9890;
wire n9891;
wire n9892;
wire n9893;
wire n9894;
wire n9895;
wire n9896;
wire n9897;
wire n9898;
wire n9899;
wire n9900;
wire n9901;
wire n9902;
wire n9903;
wire n9904;
wire n9905;
wire n9906;
wire n9907;
wire n9908;
wire n9909;
wire n9910;
wire n9911;
wire n9912;
wire n9913;
wire n9914;
wire n9915;
wire n9916;
wire n9917;
wire n9918;
wire n9919;
wire n9920;
wire n9921;
wire n9922;
wire n9923;
wire n9924;
wire n9925;
wire n9926;
wire n9927;
wire n9928;
wire n9929;
wire n9930;
wire n9931;
wire n9932;
wire n9933;
wire n9934;
wire n9935;
wire n9936;
wire n9937;
wire n9938;
wire n9939;
wire n9940;
wire n9941;
wire n9942;
wire n9943;
wire n9944;
wire n9945;
wire n9946;
wire n9947;
wire n9948;
wire n9949;
wire n9950;
wire n9951;
wire n9952;
wire n9953;
wire n9954;
wire n9955;
wire n9956;
wire n9957;
wire n9958;
wire n9959;
wire n9960;
wire n9961;
wire n9962;
wire n9963;
wire n9964;
wire n9965;
wire n9966;
wire n9967;
wire n9968;
wire n9969;
wire n9970;
wire n9971;
wire n9972;
wire n9973;
wire n9974;
wire n9975;
wire n9976;
wire n9977;
wire n9978;
wire n9979;
wire n9980;
wire n9981;
wire n9982;
wire n9983;
wire n9984;
wire n9985;
wire n9986;
wire n9987;
wire n9988;
wire n9989;
wire n9990;
wire n9991;
wire n9992;
wire n9993;
wire n9994;
wire n9995;
wire n9996;
wire n9997;
wire n9998;
wire n9999;
wire n10000;
wire n10001;
wire n10002;
wire n10003;
wire n10004;
wire n10005;
wire n10006;
wire n10007;
wire n10008;
wire n10009;
wire n10010;
wire n10011;
wire n10012;
wire n10013;
wire n10014;
wire n10015;
wire n10016;
wire n10017;
wire n10018;
wire n10019;
wire n10020;
wire n10021;
wire n10022;
wire n10023;
wire n10024;
wire n10025;
wire n10026;
wire n10027;
wire n10028;
wire n10029;
wire n10030;
wire n10031;
wire n10032;
wire n10033;
wire n10034;
wire n10035;
wire n10036;
wire n10037;
wire n10038;
wire n10039;
wire n10040;
wire n10041;
wire n10042;
wire n10043;
wire n10044;
wire n10045;
wire n10046;
wire n10047;
wire n10048;
wire n10049;
wire n10050;
wire n10051;
wire n10052;
wire n10053;
wire n10054;
wire n10055;
wire n10056;
wire n10057;
wire n10058;
wire n10059;
wire n10060;
wire n10061;
wire n10062;
wire n10063;
wire n10064;
wire n10065;
wire n10066;
wire n10067;
wire n10068;
wire n10069;
wire n10070;
wire n10071;
wire n10072;
wire n10073;
wire n10074;
wire n10075;
wire n10076;
wire n10077;
wire n10078;
wire n10079;
wire n10080;
wire n10081;
wire n10082;
wire n10083;
wire n10084;
wire n10085;
wire n10086;
wire n10087;
wire n10088;
wire n10089;
wire n10090;
wire n10091;
wire n10092;
wire n10093;
wire n10094;
wire n10095;
wire n10096;
wire n10097;
wire n10098;
wire n10099;
wire n10100;
wire n10101;
wire n10102;
wire n10103;
wire n10104;
wire n10105;
wire n10106;
wire n10107;
wire n10108;
wire n10109;
wire n10110;
wire n10111;
wire n10112;
wire n10113;
wire n10114;
wire n10115;
wire n10116;
wire n10117;
wire n10118;
wire n10119;
wire n10120;
wire n10121;
wire n10122;
wire n10123;
wire n10124;
wire n10125;
wire n10126;
wire n10127;
wire n10128;
wire n10129;
wire n10130;
wire n10131;
wire n10132;
wire n10133;
wire n10134;
wire n10135;
wire n10136;
wire n10137;
wire n10138;
wire n10139;
wire n10140;
wire n10141;
wire n10142;
wire n10143;
wire n10144;
wire n10145;
wire n10146;
wire n10147;
wire n10148;
wire n10149;
wire n10150;
wire n10151;
wire n10152;
wire n10153;
wire n10154;
wire n10155;
wire n10156;
wire n10157;
wire n10158;
wire n10159;
wire n10160;
wire n10161;
wire n10162;
wire n10163;
wire n10164;
wire n10165;
wire n10166;
wire n10167;
wire n10168;
wire n10169;
wire n10170;
wire n10171;
wire n10172;
wire n10173;
wire n10174;
wire n10175;
wire n10176;
wire n10177;
wire n10178;
wire n10179;
wire n10180;
wire n10181;
wire n10182;
wire n10183;
wire n10184;
wire n10185;
wire n10186;
wire n10187;
wire n10188;
wire n10189;
wire n10190;
wire n10191;
wire n10192;
wire n10193;
wire n10194;
wire n10195;
wire n10196;
wire n10197;
wire n10198;
wire n10199;
wire n10200;
wire n10201;
wire n10202;
wire n10203;
wire n10204;
wire n10205;
wire n10206;
wire n10207;
wire n10208;
wire n10209;
wire n10210;
wire n10211;
wire n10212;
wire n10213;
wire n10214;
wire n10215;
wire n10216;
wire n10217;
wire n10218;
wire n10219;
wire n10220;
wire n10221;
wire n10222;
wire n10223;
wire n10224;
wire n10225;
wire n10226;
wire n10227;
wire n10228;
wire n10229;
wire n10230;
wire n10231;
wire n10232;
wire n10233;
wire n10234;
wire n10235;
wire n10236;
wire n10237;
wire n10238;
wire n10239;
wire n10240;
wire n10241;
wire n10242;
wire n10243;
wire n10244;
wire n10245;
wire n10246;
wire n10247;
wire n10248;
wire n10249;
wire n10250;
wire n10251;
wire n10252;
wire n10253;
wire n10254;
wire n10255;
wire n10256;
wire n10257;
wire n10258;
wire n10259;
wire n10260;
wire n10261;
wire n10262;
wire n10263;
wire n10264;
wire n10265;
wire n10266;
wire n10267;
wire n10268;
wire n10269;
wire n10270;
wire n10271;
wire n10272;
wire n10273;
wire n10274;
wire n10275;
wire n10276;
wire n10277;
wire n10278;
wire n10279;
wire n10280;
wire n10281;
wire n10282;
wire n10283;
wire n10284;
wire n10285;
wire n10286;
wire n10287;
wire n10288;
wire n10289;
wire n10290;
wire n10291;
wire n10292;
wire n10293;
wire n10294;
wire n10295;
wire n10296;
wire n10297;
wire n10298;
wire n10299;
wire n10300;
wire n10301;
wire n10302;
wire n10303;
wire n10304;
wire n10305;
wire n10306;
wire n10307;
wire n10308;
wire n10309;
wire n10310;
wire n10311;
wire n10312;
wire n10313;
wire n10314;
wire n10315;
wire n10316;
wire n10317;
wire n10318;
wire n10319;
wire n10320;
wire n10321;
wire n10322;
wire n10323;
wire n10324;
wire n10325;
wire n10326;
wire n10327;
wire n10328;
wire n10329;
wire n10330;
wire n10331;
wire n10332;
wire n10333;
wire n10334;
wire n10335;
wire n10336;
wire n10337;
wire n10338;
wire n10339;
wire n10340;
wire n10341;
wire n10342;
wire n10343;
wire n10344;
wire n10345;
wire n10346;
wire n10347;
wire n10348;
wire n10349;
wire n10350;
wire n10351;
wire n10352;
wire n10353;
wire n10354;
wire n10355;
wire n10356;
wire n10357;
wire n10358;
wire n10359;
wire n10360;
wire n10361;
wire n10362;
wire n10363;
wire n10364;
wire n10365;
wire n10366;
wire n10367;
wire n10368;
wire n10369;
wire n10370;
wire n10371;
wire n10372;
wire n10373;
wire n10374;
wire n10375;
wire n10376;
wire n10377;
wire n10378;
wire n10379;
wire n10380;
wire n10381;
wire n10382;
wire n10383;
wire n10384;
wire n10385;
wire n10386;
wire n10387;
wire n10388;
wire n10389;
wire n10390;
wire n10391;
wire n10392;
wire n10393;
wire n10394;
wire n10395;
wire n10396;
wire n10397;
wire n10398;
wire n10399;
wire n10400;
wire n10401;
wire n10402;
wire n10403;
wire n10404;
wire n10405;
wire n10406;
wire n10407;
wire n10408;
wire n10409;
wire n10410;
wire n10411;
wire n10412;
wire n10413;
wire n10414;
wire n10415;
xor (out,n0,n5184);
nand (n0,n1,n5181);
or (n1,n2,n5176);
not (n2,n3);
nand (n3,n4,n5175);
or (n4,n5,n1087);
nand (n5,n6,n1086);
not (n6,n7);
nor (n7,n8,n992);
or (n8,n9,n991);
and (n9,n10,n897);
xor (n10,n11,n757);
or (n11,n12,n756);
and (n12,n13,n630);
xor (n13,n14,n495);
or (n14,n15,n494);
and (n15,n16,n301);
xor (n16,n17,n88);
xor (n17,n18,n62);
xor (n18,n19,n35);
not (n19,n20);
nor (n20,n21,n32);
and (n21,n22,n23);
nand (n22,n23,n30);
not (n23,n24);
nand (n24,n25,n29);
or (n25,n26,n28);
not (n26,n27);
nand (n29,n26,n28);
nand (n30,n31,n34);
or (n31,n27,n32);
not (n32,n33);
nand (n34,n32,n27);
nand (n35,n36,n55);
or (n36,n37,n50);
not (n37,n38);
nor (n38,n39,n46);
nor (n39,n40,n44);
and (n40,n41,n43);
not (n41,n42);
and (n44,n45,n42);
not (n45,n43);
nand (n46,n47,n49);
or (n47,n45,n48);
nand (n49,n45,n48);
nor (n50,n51,n54);
and (n51,n42,n52);
not (n52,n53);
and (n54,n41,n53);
or (n55,n56,n57);
not (n56,n46);
nor (n57,n58,n60);
and (n58,n41,n59);
and (n60,n61,n42);
not (n61,n59);
nand (n62,n63,n82);
or (n63,n64,n77);
nand (n64,n65,n72);
nor (n65,n66,n70);
and (n66,n67,n69);
not (n67,n68);
and (n70,n68,n71);
not (n71,n69);
nand (n72,n73,n76);
or (n73,n69,n74);
not (n74,n75);
nand (n76,n74,n69);
nor (n77,n78,n80);
and (n78,n74,n79);
and (n80,n75,n81);
not (n81,n79);
or (n82,n65,n83);
nor (n83,n84,n86);
and (n84,n74,n85);
and (n86,n75,n87);
not (n87,n85);
or (n88,n89,n300);
and (n89,n90,n225);
xor (n90,n91,n166);
or (n91,n92,n165);
and (n92,n93,n136);
xor (n93,n94,n109);
nand (n94,n95,n107);
or (n95,n96,n102);
nand (n96,n97,n101);
or (n97,n98,n100);
not (n98,n99);
nand (n101,n98,n100);
not (n102,n103);
nand (n103,n104,n105);
not (n104,n96);
nand (n105,n106,n108);
or (n106,n98,n107);
nand (n108,n98,n107);
nand (n109,n110,n130);
or (n110,n111,n118);
not (n111,n112);
nand (n112,n113,n117);
or (n113,n114,n115);
not (n115,n116);
nand (n117,n114,n115);
not (n118,n119);
nor (n119,n120,n125);
nor (n120,n121,n123);
and (n121,n115,n122);
and (n123,n124,n116);
not (n124,n122);
nand (n125,n126,n129);
or (n126,n127,n122);
not (n127,n128);
nand (n129,n127,n122);
nand (n130,n131,n125);
nor (n131,n132,n135);
and (n132,n115,n133);
not (n133,n134);
and (n135,n116,n134);
nand (n136,n137,n159);
or (n137,n138,n154);
not (n138,n139);
nor (n139,n140,n148);
not (n140,n141);
nor (n141,n142,n145);
and (n142,n143,n144);
and (n145,n146,n147);
not (n146,n143);
not (n147,n144);
not (n148,n149);
or (n149,n150,n152);
and (n150,n143,n151);
and (n152,n146,n153);
not (n153,n151);
nor (n154,n155,n157);
and (n155,n147,n156);
and (n157,n144,n158);
not (n158,n156);
or (n159,n160,n149);
nor (n160,n161,n163);
and (n161,n162,n147);
and (n163,n164,n144);
not (n164,n162);
and (n165,n94,n109);
or (n166,n167,n224);
and (n167,n168,n211);
xor (n168,n169,n196);
nand (n169,n170,n188);
or (n170,n171,n182);
nand (n171,n172,n178);
nor (n172,n173,n176);
and (n173,n107,n174);
not (n174,n175);
and (n176,n177,n175);
not (n177,n107);
nand (n178,n179,n181);
or (n179,n174,n180);
nand (n181,n180,n174);
not (n182,n183);
nand (n183,n184,n187);
or (n184,n180,n185);
not (n185,n186);
nand (n187,n180,n185);
nand (n188,n189,n190);
not (n189,n172);
nand (n190,n191,n194);
or (n191,n192,n180);
not (n192,n193);
or (n194,n195,n193);
not (n195,n180);
not (n196,n197);
nor (n197,n198,n209);
and (n198,n199,n200);
nand (n199,n200,n207);
nor (n200,n201,n205);
and (n201,n202,n204);
not (n202,n203);
and (n205,n203,n206);
not (n206,n204);
nand (n207,n208,n210);
or (n208,n204,n209);
not (n209,n28);
nand (n210,n209,n204);
nand (n211,n212,n218);
or (n212,n37,n213);
nor (n213,n214,n216);
and (n214,n215,n41);
and (n216,n42,n217);
not (n217,n215);
or (n218,n219,n56);
nor (n219,n220,n223);
and (n220,n42,n221);
not (n221,n222);
and (n223,n41,n222);
and (n224,n169,n196);
or (n225,n226,n299);
and (n226,n227,n273);
xor (n227,n228,n248);
nand (n228,n229,n243);
or (n229,n230,n234);
not (n230,n231);
nor (n231,n232,n233);
and (n232,n67,n81);
and (n233,n68,n79);
nand (n234,n235,n240);
nor (n235,n236,n238);
and (n236,n32,n237);
and (n238,n33,n239);
not (n239,n237);
nand (n240,n241,n242);
or (n241,n239,n68);
nand (n242,n68,n239);
nand (n243,n244,n247);
nor (n244,n245,n246);
and (n245,n67,n87);
and (n246,n68,n85);
not (n247,n235);
nand (n248,n249,n268);
or (n249,n250,n255);
not (n250,n251);
nor (n251,n252,n254);
and (n252,n253,n52);
not (n253,n48);
and (n254,n48,n53);
nand (n255,n256,n263);
or (n256,n257,n260);
not (n257,n258);
nand (n258,n253,n259);
not (n260,n261);
nand (n261,n48,n262);
not (n262,n259);
nor (n263,n264,n267);
and (n264,n265,n259);
not (n265,n266);
and (n267,n266,n262);
nand (n268,n269,n272);
nor (n269,n270,n271);
and (n270,n253,n61);
and (n271,n48,n59);
not (n272,n263);
nand (n273,n274,n293);
or (n274,n275,n281);
not (n275,n276);
nor (n276,n277,n280);
and (n277,n265,n278);
not (n278,n279);
and (n280,n266,n279);
not (n281,n282);
nor (n282,n283,n288);
nor (n283,n284,n287);
and (n284,n266,n285);
not (n285,n286);
and (n287,n265,n286);
nand (n288,n289,n292);
or (n289,n290,n286);
not (n290,n291);
nand (n292,n290,n286);
nand (n293,n288,n294);
nor (n294,n295,n298);
and (n295,n296,n265);
not (n296,n297);
and (n298,n297,n266);
and (n299,n228,n248);
and (n300,n91,n166);
or (n301,n302,n493);
and (n302,n303,n426);
xor (n303,n304,n363);
or (n304,n305,n362);
and (n305,n306,n354);
xor (n306,n307,n330);
nand (n307,n308,n324);
or (n308,n309,n315);
not (n309,n310);
nor (n310,n311,n314);
and (n311,n290,n312);
not (n312,n313);
and (n314,n291,n313);
nand (n315,n316,n321);
not (n316,n317);
nand (n317,n318,n320);
or (n318,n195,n319);
nand (n320,n195,n319);
nand (n321,n322,n323);
or (n322,n319,n290);
nand (n323,n290,n319);
nand (n324,n325,n317);
nor (n325,n326,n329);
and (n326,n290,n327);
not (n327,n328);
and (n329,n291,n328);
nand (n330,n331,n343);
or (n331,n332,n337);
not (n332,n333);
nand (n333,n334,n336);
or (n334,n74,n335);
nand (n336,n74,n335);
not (n337,n338);
nand (n338,n339,n342);
or (n339,n340,n128);
not (n340,n341);
or (n342,n127,n341);
nand (n343,n344,n350);
not (n344,n345);
nor (n345,n346,n349);
and (n346,n128,n347);
not (n347,n348);
and (n349,n127,n348);
and (n350,n332,n351);
nand (n351,n352,n353);
or (n352,n335,n127);
nand (n353,n127,n335);
nand (n354,n355,n361);
or (n355,n22,n356);
nor (n356,n357,n359);
and (n357,n32,n358);
and (n359,n33,n360);
not (n360,n358);
or (n361,n23,n32);
and (n362,n307,n330);
or (n363,n364,n425);
and (n364,n365,n411);
xor (n365,n366,n391);
nand (n366,n367,n385);
or (n367,n368,n373);
nor (n368,n369,n372);
and (n369,n370,n151);
not (n370,n371);
and (n372,n153,n371);
not (n373,n374);
nor (n374,n375,n380);
nor (n375,n376,n379);
and (n376,n151,n377);
not (n377,n378);
nor (n379,n151,n377);
nand (n380,n381,n384);
or (n381,n382,n378);
not (n382,n383);
nand (n384,n382,n378);
nand (n385,n386,n380);
nor (n386,n387,n390);
and (n387,n153,n388);
not (n388,n389);
and (n390,n151,n389);
nand (n391,n392,n410);
or (n392,n393,n400);
nor (n393,n394,n398);
and (n394,n395,n397);
not (n395,n396);
and (n398,n399,n396);
not (n399,n397);
not (n400,n401);
nor (n401,n402,n405);
xnor (n402,n395,n403);
not (n403,n404);
nor (n405,n406,n408);
and (n406,n407,n404);
and (n408,n409,n403);
not (n409,n407);
nand (n410,n405,n396);
nand (n411,n412,n407);
or (n412,n413,n419);
nand (n413,n414,n418);
or (n414,n415,n417);
not (n415,n416);
nand (n418,n415,n417);
not (n419,n420);
nand (n420,n421,n424);
nand (n421,n422,n423);
or (n422,n417,n409);
nand (n423,n409,n417);
not (n424,n413);
and (n425,n366,n391);
or (n426,n427,n492);
and (n427,n428,n479);
xor (n428,n429,n455);
nand (n429,n430,n448);
or (n430,n431,n436);
not (n431,n432);
nand (n432,n433,n435);
or (n433,n434,n382);
nand (n435,n434,n382);
not (n436,n437);
and (n437,n438,n445);
nor (n438,n439,n443);
and (n439,n440,n442);
not (n440,n441);
and (n443,n441,n444);
not (n444,n442);
nand (n445,n446,n447);
or (n446,n442,n382);
nand (n447,n382,n442);
nand (n448,n449,n450);
not (n449,n438);
nor (n450,n451,n454);
and (n451,n452,n382);
not (n452,n453);
and (n454,n453,n383);
nand (n455,n456,n468);
or (n456,n457,n462);
nor (n457,n458,n460);
and (n458,n395,n459);
and (n460,n396,n461);
not (n461,n459);
not (n462,n463);
nor (n463,n464,n467);
and (n464,n465,n440);
not (n465,n466);
and (n467,n466,n441);
nand (n468,n469,n474);
not (n469,n470);
nand (n470,n457,n471);
nand (n471,n472,n473);
or (n472,n459,n440);
nand (n473,n440,n459);
nor (n474,n475,n478);
and (n475,n476,n440);
not (n476,n477);
and (n478,n477,n441);
nand (n479,n480,n486);
or (n480,n64,n481);
nor (n481,n482,n484);
and (n482,n483,n74);
and (n484,n485,n75);
not (n485,n483);
or (n486,n487,n65);
nor (n487,n488,n490);
and (n488,n489,n74);
and (n490,n491,n75);
not (n491,n489);
and (n492,n429,n455);
and (n493,n304,n363);
and (n494,n17,n88);
or (n495,n496,n629);
and (n496,n497,n622);
xor (n497,n498,n555);
xor (n498,n499,n545);
xor (n499,n500,n524);
or (n500,n501,n523);
and (n501,n502,n514);
xor (n502,n503,n507);
nand (n503,n504,n506);
or (n504,n505,n171);
not (n505,n190);
nand (n506,n189,n180);
nand (n507,n508,n510);
or (n508,n509,n118);
not (n509,n131);
nand (n510,n511,n125);
nor (n511,n512,n513);
and (n512,n115,n347);
and (n513,n116,n348);
nand (n514,n515,n517);
or (n515,n373,n516);
not (n516,n386);
or (n517,n518,n522);
nor (n518,n519,n520);
and (n519,n434,n153);
and (n520,n521,n151);
not (n521,n434);
not (n522,n380);
and (n523,n503,n507);
or (n524,n525,n544);
and (n525,n526,n537);
xor (n526,n527,n530);
nor (n527,n528,n395);
and (n528,n400,n529);
not (n529,n405);
nand (n530,n531,n533);
or (n531,n337,n532);
not (n532,n350);
nand (n533,n534,n333);
nor (n534,n535,n536);
and (n535,n127,n485);
and (n536,n128,n483);
nand (n537,n538,n540);
or (n538,n436,n539);
not (n539,n450);
or (n540,n438,n541);
nor (n541,n542,n543);
and (n542,n382,n477);
and (n543,n383,n476);
and (n544,n527,n530);
or (n545,n546,n554);
and (n546,n547,n551);
xor (n547,n20,n548);
nand (n548,n549,n550);
or (n549,n37,n219);
or (n550,n50,n56);
nand (n551,n552,n553);
or (n552,n64,n487);
or (n553,n77,n65);
and (n554,n20,n548);
xor (n555,n556,n606);
xor (n556,n557,n582);
or (n557,n558,n581);
and (n558,n559,n574);
xor (n559,n560,n567);
nand (n560,n561,n562);
or (n561,n462,n470);
nand (n562,n563,n566);
nor (n563,n564,n565);
and (n564,n399,n440);
and (n565,n397,n441);
not (n566,n457);
nand (n567,n568,n570);
or (n568,n569,n281);
not (n569,n294);
nand (n570,n288,n571);
nand (n571,n572,n573);
or (n572,n266,n312);
or (n573,n265,n313);
nand (n574,n575,n577);
or (n575,n315,n576);
not (n576,n325);
or (n577,n578,n316);
nor (n578,n579,n580);
and (n579,n290,n186);
and (n580,n291,n185);
and (n581,n560,n567);
or (n582,n583,n605);
and (n583,n584,n599);
xor (n584,n585,n592);
nand (n585,n586,n588);
or (n586,n587,n234);
not (n587,n244);
nand (n588,n589,n247);
nor (n589,n590,n591);
and (n590,n360,n67);
and (n591,n358,n68);
nand (n592,n593,n595);
or (n593,n594,n255);
not (n594,n269);
nand (n595,n596,n272);
nor (n596,n597,n598);
and (n597,n253,n278);
and (n598,n48,n279);
nand (n599,n600,n601);
or (n600,n138,n160);
or (n601,n602,n149);
nor (n602,n603,n604);
and (n603,n371,n147);
and (n604,n370,n144);
and (n605,n585,n592);
xor (n606,n607,n616);
xor (n607,n608,n609);
not (n608,n527);
nand (n609,n610,n612);
or (n610,n532,n611);
not (n611,n534);
or (n612,n613,n332);
nor (n613,n614,n615);
and (n614,n489,n127);
and (n615,n491,n128);
nand (n616,n617,n618);
or (n617,n436,n541);
or (n618,n438,n619);
nor (n619,n620,n621);
and (n620,n382,n466);
and (n621,n383,n465);
or (n622,n623,n628);
and (n623,n624,n627);
xor (n624,n625,n626);
xor (n625,n526,n537);
xor (n626,n502,n514);
xor (n627,n559,n574);
and (n628,n625,n626);
and (n629,n498,n555);
xor (n630,n631,n699);
xor (n631,n632,n696);
or (n632,n633,n695);
and (n633,n634,n676);
xor (n634,n635,n657);
xor (n635,n636,n648);
xor (n636,n637,n641);
nand (n637,n638,n640);
or (n638,n639,n470);
not (n639,n563);
nand (n640,n566,n441);
nand (n641,n642,n644);
or (n642,n643,n281);
not (n643,n571);
nand (n644,n645,n288);
nor (n645,n646,n647);
and (n646,n328,n266);
and (n647,n327,n265);
nand (n648,n649,n654);
or (n649,n316,n650);
not (n650,n651);
nor (n651,n652,n653);
and (n652,n290,n192);
and (n653,n291,n193);
nand (n654,n655,n656);
not (n655,n578);
not (n656,n315);
xor (n657,n658,n670);
xor (n658,n659,n662);
nand (n659,n660,n180);
or (n660,n189,n661);
not (n661,n171);
nand (n662,n663,n669);
or (n663,n664,n665);
not (n664,n125);
not (n665,n666);
nand (n666,n667,n668);
or (n667,n340,n116);
or (n668,n341,n115);
nand (n669,n119,n511);
nand (n670,n671,n672);
or (n671,n373,n518);
or (n672,n673,n522);
nor (n673,n674,n675);
and (n674,n153,n453);
and (n675,n151,n452);
xor (n676,n677,n689);
xor (n677,n678,n682);
nand (n678,n679,n681);
or (n679,n234,n680);
not (n680,n589);
or (n681,n235,n67);
nand (n682,n683,n685);
or (n683,n255,n684);
not (n684,n596);
or (n685,n686,n263);
nor (n686,n687,n688);
and (n687,n253,n297);
and (n688,n48,n296);
nand (n689,n690,n691);
or (n690,n138,n602);
or (n691,n692,n149);
nor (n692,n693,n694);
and (n693,n389,n147);
and (n694,n388,n144);
and (n695,n635,n657);
or (n696,n697,n698);
and (n697,n556,n606);
and (n698,n557,n582);
xor (n699,n700,n740);
xor (n700,n701,n718);
xor (n701,n702,n712);
xor (n702,n703,n706);
nand (n703,n704,n705);
or (n704,n650,n315);
nand (n705,n317,n291);
nand (n706,n707,n708);
or (n707,n665,n118);
or (n708,n709,n664);
nor (n709,n710,n711);
and (n710,n483,n115);
and (n711,n485,n116);
nand (n712,n713,n714);
or (n713,n436,n619);
or (n714,n715,n438);
nor (n715,n716,n717);
and (n716,n382,n397);
and (n717,n383,n399);
xor (n718,n719,n734);
xor (n719,n720,n726);
nand (n720,n721,n722);
or (n721,n138,n692);
or (n722,n723,n149);
nor (n723,n724,n725);
and (n724,n434,n147);
and (n725,n521,n144);
nand (n726,n727,n729);
or (n727,n281,n728);
not (n728,n645);
or (n729,n730,n731);
not (n730,n288);
nor (n731,n732,n733);
and (n732,n265,n186);
and (n733,n266,n185);
nand (n734,n735,n736);
or (n735,n64,n83);
or (n736,n737,n65);
nor (n737,n738,n739);
and (n738,n74,n358);
and (n739,n75,n360);
xor (n740,n741,n754);
xor (n741,n742,n748);
nand (n742,n743,n744);
or (n743,n255,n686);
or (n744,n745,n263);
nor (n745,n746,n747);
and (n746,n253,n313);
and (n747,n48,n312);
nand (n748,n749,n750);
or (n749,n613,n532);
nand (n750,n333,n751);
nor (n751,n752,n753);
and (n752,n79,n128);
and (n753,n81,n127);
nor (n754,n755,n440);
and (n755,n470,n457);
and (n756,n14,n495);
xor (n757,n758,n804);
xor (n758,n759,n801);
xor (n759,n760,n790);
xor (n760,n761,n787);
xor (n761,n762,n784);
xor (n762,n763,n766);
or (n763,n764,n765);
and (n764,n719,n734);
and (n765,n720,n726);
or (n766,n767,n783);
and (n767,n768,n777);
xor (n768,n769,n771);
nor (n769,n770,n67);
and (n770,n234,n235);
nand (n771,n772,n773);
or (n772,n373,n673);
or (n773,n774,n522);
nor (n774,n775,n776);
and (n775,n153,n477);
and (n776,n151,n476);
nand (n777,n778,n779);
or (n778,n37,n57);
or (n779,n56,n780);
nor (n780,n781,n782);
and (n781,n41,n279);
and (n782,n278,n42);
and (n783,n769,n771);
or (n784,n785,n786);
and (n785,n741,n754);
and (n786,n742,n748);
or (n787,n788,n789);
and (n788,n700,n740);
and (n789,n701,n718);
or (n790,n791,n800);
and (n791,n792,n799);
xor (n792,n793,n796);
or (n793,n794,n795);
and (n794,n677,n689);
and (n795,n678,n682);
or (n796,n797,n798);
and (n797,n636,n648);
and (n798,n637,n641);
xor (n799,n768,n777);
and (n800,n793,n796);
or (n801,n802,n803);
and (n802,n631,n699);
and (n803,n632,n696);
xor (n804,n805,n888);
xor (n805,n806,n844);
xor (n806,n807,n828);
xor (n807,n808,n811);
or (n808,n809,n810);
and (n809,n702,n712);
and (n810,n703,n706);
xor (n811,n812,n825);
xor (n812,n813,n819);
nand (n813,n814,n815);
or (n814,n138,n723);
or (n815,n816,n149);
nor (n816,n817,n818);
and (n817,n147,n453);
and (n818,n452,n144);
nand (n819,n820,n821);
or (n820,n281,n731);
or (n821,n730,n822);
nor (n822,n823,n824);
and (n823,n265,n193);
and (n824,n266,n192);
nand (n825,n826,n827);
or (n826,n64,n737);
or (n827,n65,n74);
xor (n828,n829,n837);
xor (n829,n830,n831);
not (n830,n769);
nand (n831,n832,n833);
or (n832,n373,n774);
or (n833,n522,n834);
nor (n834,n835,n836);
and (n835,n153,n466);
and (n836,n151,n465);
nand (n837,n838,n843);
or (n838,n839,n56);
not (n839,n840);
nand (n840,n841,n842);
or (n841,n296,n42);
or (n842,n41,n297);
or (n843,n37,n780);
xor (n844,n845,n875);
xor (n845,n846,n859);
xor (n846,n847,n856);
xor (n847,n848,n850);
nand (n848,n849,n291);
or (n849,n317,n656);
nand (n850,n851,n852);
or (n851,n118,n709);
or (n852,n853,n664);
nor (n853,n854,n855);
and (n854,n115,n489);
and (n855,n491,n116);
nand (n856,n857,n858);
or (n857,n436,n715);
or (n858,n438,n382);
xor (n859,n860,n874);
xor (n860,n861,n867);
nand (n861,n862,n863);
or (n862,n255,n745);
or (n863,n864,n263);
nor (n864,n865,n866);
and (n865,n253,n328);
and (n866,n48,n327);
nand (n867,n868,n870);
or (n868,n532,n869);
not (n869,n751);
or (n870,n871,n332);
nor (n871,n872,n873);
and (n872,n127,n85);
and (n873,n128,n87);
not (n874,n754);
or (n875,n876,n887);
and (n876,n877,n884);
xor (n877,n878,n881);
or (n878,n879,n880);
and (n879,n658,n670);
and (n880,n659,n662);
or (n881,n882,n883);
and (n882,n607,n616);
and (n883,n608,n609);
or (n884,n885,n886);
and (n885,n18,n62);
and (n886,n19,n35);
and (n887,n878,n881);
or (n888,n889,n896);
and (n889,n890,n895);
xor (n890,n891,n894);
or (n891,n892,n893);
and (n892,n499,n545);
and (n893,n500,n524);
xor (n894,n877,n884);
xor (n895,n792,n799);
and (n896,n891,n894);
or (n897,n898,n990);
and (n898,n899,n989);
xor (n899,n900,n901);
xor (n900,n890,n895);
or (n901,n902,n988);
and (n902,n903,n987);
xor (n903,n904,n905);
xor (n904,n634,n676);
or (n905,n906,n986);
and (n906,n907,n910);
xor (n907,n908,n909);
xor (n908,n547,n551);
xor (n909,n584,n599);
or (n910,n911,n985);
and (n911,n912,n960);
xor (n912,n913,n940);
or (n913,n914,n939);
and (n914,n915,n931);
xor (n915,n916,n922);
nand (n916,n917,n921);
nand (n917,n104,n918,n105);
nand (n918,n919,n920);
or (n919,n193,n177);
nand (n920,n193,n177);
nand (n921,n96,n107);
nand (n922,n923,n930);
or (n923,n924,n118);
not (n924,n925);
nor (n925,n926,n929);
and (n926,n115,n927);
not (n927,n928);
and (n929,n116,n928);
nand (n930,n112,n125);
nand (n931,n932,n938);
or (n932,n138,n933);
nor (n933,n934,n936);
and (n934,n935,n147);
and (n936,n937,n144);
not (n937,n935);
or (n938,n154,n149);
and (n939,n916,n922);
or (n940,n941,n959);
and (n941,n942,n950);
xor (n942,n943,n197);
nand (n943,n944,n949);
or (n944,n945,n171);
not (n945,n946);
nor (n946,n947,n948);
and (n947,n195,n327);
and (n948,n180,n328);
nand (n949,n183,n189);
nand (n950,n951,n958);
or (n951,n37,n952);
not (n952,n953);
nor (n953,n954,n957);
and (n954,n41,n955);
not (n955,n956);
and (n957,n42,n956);
or (n958,n213,n56);
and (n959,n943,n197);
or (n960,n961,n984);
and (n961,n962,n977);
xor (n962,n963,n970);
nand (n963,n964,n969);
or (n964,n965,n234);
not (n965,n966);
nor (n966,n967,n968);
and (n967,n67,n491);
and (n968,n68,n489);
nand (n969,n231,n247);
nand (n970,n971,n976);
or (n971,n972,n255);
not (n972,n973);
nor (n973,n974,n975);
and (n974,n253,n221);
and (n975,n48,n222);
nand (n976,n272,n251);
nand (n977,n978,n983);
or (n978,n281,n979);
not (n979,n980);
nor (n980,n981,n982);
and (n981,n61,n265);
and (n982,n59,n266);
or (n983,n275,n730);
and (n984,n963,n970);
and (n985,n913,n940);
and (n986,n908,n909);
xor (n987,n16,n301);
and (n988,n904,n905);
xor (n989,n13,n630);
and (n990,n900,n901);
and (n991,n11,n757);
xor (n992,n993,n1083);
xor (n993,n994,n997);
or (n994,n995,n996);
and (n995,n805,n888);
and (n996,n806,n844);
xor (n997,n998,n1037);
xor (n998,n999,n1034);
xor (n999,n1000,n1023);
xor (n1000,n1001,n1020);
xor (n1001,n1002,n1014);
xor (n1002,n1003,n1008);
not (n1003,n1004);
nand (n1004,n1005,n75);
or (n1005,n1006,n1007);
not (n1006,n65);
not (n1007,n64);
nand (n1008,n1009,n1010);
or (n1009,n138,n816);
or (n1010,n1011,n149);
nor (n1011,n1012,n1013);
and (n1012,n147,n477);
and (n1013,n144,n476);
nand (n1014,n1015,n1019);
or (n1015,n1016,n332);
nor (n1016,n1017,n1018);
and (n1017,n127,n358);
and (n1018,n128,n360);
or (n1019,n532,n871);
or (n1020,n1021,n1022);
and (n1021,n762,n784);
and (n1022,n763,n766);
xor (n1023,n1024,n1031);
xor (n1024,n1025,n1028);
or (n1025,n1026,n1027);
and (n1026,n847,n856);
and (n1027,n848,n850);
or (n1028,n1029,n1030);
and (n1029,n860,n874);
and (n1030,n861,n867);
or (n1031,n1032,n1033);
and (n1032,n829,n837);
and (n1033,n830,n831);
or (n1034,n1035,n1036);
and (n1035,n760,n790);
and (n1036,n761,n787);
xor (n1037,n1038,n1080);
xor (n1038,n1039,n1042);
or (n1039,n1040,n1041);
and (n1040,n807,n828);
and (n1041,n808,n811);
xor (n1042,n1043,n1064);
xor (n1043,n1044,n1047);
or (n1044,n1045,n1046);
and (n1045,n812,n825);
and (n1046,n813,n819);
xor (n1047,n1048,n1058);
xor (n1048,n1049,n1052);
nand (n1049,n1050,n1051);
or (n1050,n281,n822);
or (n1051,n730,n265);
nand (n1052,n1053,n1054);
or (n1053,n118,n853);
or (n1054,n1055,n664);
nor (n1055,n1056,n1057);
and (n1056,n115,n79);
and (n1057,n81,n116);
nand (n1058,n1059,n1060);
or (n1059,n839,n37);
or (n1060,n1061,n56);
nor (n1061,n1062,n1063);
and (n1062,n41,n313);
and (n1063,n42,n312);
xor (n1064,n1065,n1074);
xor (n1065,n1066,n1072);
nand (n1066,n1067,n1068);
or (n1067,n373,n834);
or (n1068,n522,n1069);
nor (n1069,n1070,n1071);
and (n1070,n153,n397);
and (n1071,n151,n399);
nor (n1072,n1073,n382);
and (n1073,n436,n438);
nand (n1074,n1075,n1076);
or (n1075,n255,n864);
or (n1076,n1077,n263);
nor (n1077,n1078,n1079);
and (n1078,n253,n186);
and (n1079,n48,n185);
or (n1080,n1081,n1082);
and (n1081,n845,n875);
and (n1082,n846,n859);
or (n1083,n1084,n1085);
and (n1084,n758,n804);
and (n1085,n759,n801);
nand (n1086,n8,n992);
nand (n1087,n1088,n5133,n5168);
nand (n1088,n1089,n5085);
not (n1089,n1090);
nand (n1090,n1091,n4145,n4945,n4964);
not (n1091,n1092);
nand (n1092,n1093,n3611);
nand (n1093,n1094,n3598,n3604);
nand (n1094,n1095,n2697);
nor (n1095,n1096,n2676);
nor (n1096,n1097,n2480);
xor (n1097,n1098,n2297);
xor (n1098,n1099,n2127);
xor (n1099,n1100,n1805);
xor (n1100,n1101,n1617);
or (n1101,n1102,n1616);
and (n1102,n1103,n1363);
xor (n1103,n1104,n1252);
xor (n1104,n1105,n1203);
xor (n1105,n1106,n1155);
xor (n1106,n1107,n1133);
xor (n1107,n1108,n1119);
nand (n1108,n1109,n1114);
or (n1109,n1110,n199);
not (n1110,n1111);
nand (n1111,n1112,n1113);
or (n1112,n347,n28);
nand (n1113,n28,n347);
nand (n1114,n1115,n1118);
nand (n1115,n1116,n1117);
or (n1116,n341,n209);
nand (n1117,n209,n341);
not (n1118,n200);
nand (n1119,n1120,n1127);
or (n1120,n1121,n281);
not (n1121,n1122);
nor (n1122,n1123,n1126);
and (n1123,n1124,n265);
not (n1124,n1125);
and (n1126,n1125,n266);
nand (n1127,n288,n1128);
nand (n1128,n1129,n1132);
or (n1129,n266,n1130);
not (n1130,n1131);
nand (n1132,n266,n1130);
nand (n1133,n1134,n1150);
or (n1134,n1135,n1138);
nor (n1135,n1136,n1137);
and (n1136,n415,n434);
and (n1137,n416,n521);
not (n1138,n1139);
and (n1139,n1140,n1144);
nand (n1140,n1141,n1143);
or (n1141,n1142,n415);
nand (n1143,n415,n1142);
nor (n1144,n1145,n1148);
and (n1145,n1146,n1147);
not (n1147,n1142);
and (n1148,n1149,n1142);
not (n1149,n1146);
nand (n1150,n1151,n1154);
nor (n1151,n1152,n1153);
and (n1152,n453,n416);
and (n1153,n452,n415);
not (n1154,n1144);
xor (n1155,n1156,n1187);
xor (n1156,n1157,n1171);
nand (n1157,n1158,n1165);
or (n1158,n1159,n64);
not (n1159,n1160);
nor (n1160,n1161,n1164);
and (n1161,n74,n1162);
not (n1162,n1163);
and (n1164,n1163,n75);
nand (n1165,n1166,n1006);
nand (n1166,n1167,n1170);
or (n1167,n75,n1168);
not (n1168,n1169);
nand (n1170,n75,n1168);
nand (n1171,n1172,n1183);
or (n1172,n1173,n1178);
not (n1173,n1174);
and (n1174,n1175,n1176);
not (n1176,n1177);
not (n1178,n1179);
nor (n1179,n1180,n1182);
and (n1180,n1181,n81);
not (n1181,n1175);
and (n1182,n79,n1175);
nand (n1183,n1184,n1177);
nor (n1184,n1185,n1186);
and (n1185,n1181,n87);
and (n1186,n85,n1175);
nand (n1187,n1188,n1198);
or (n1188,n1189,n1194);
nor (n1189,n1190,n1193);
and (n1190,n313,n1191);
not (n1191,n1192);
and (n1193,n1192,n312);
not (n1194,n1195);
and (n1195,n1192,n1196);
not (n1196,n1197);
or (n1198,n1199,n1196);
not (n1199,n1200);
nor (n1200,n1201,n1202);
and (n1201,n1191,n327);
and (n1202,n328,n1192);
xor (n1203,n1204,n1239);
xor (n1204,n1205,n1217);
nand (n1205,n1206,n1212);
or (n1206,n1207,n436);
not (n1207,n1208);
nand (n1208,n1209,n1211);
or (n1209,n1210,n382);
nand (n1211,n382,n1210);
nand (n1212,n449,n1213);
nand (n1213,n1214,n1216);
or (n1214,n1215,n382);
nand (n1216,n1215,n382);
nand (n1217,n1218,n1234);
or (n1218,n1219,n1223);
not (n1219,n1220);
nand (n1220,n1221,n1222);
or (n1221,n483,n202);
nand (n1222,n202,n483);
nand (n1223,n1224,n1231);
or (n1224,n1225,n1228);
not (n1225,n1226);
nand (n1226,n202,n1227);
not (n1228,n1229);
nand (n1229,n203,n1230);
not (n1230,n1227);
nor (n1231,n1232,n1233);
and (n1232,n1181,n1227);
and (n1233,n1175,n1230);
nand (n1234,n1235,n1238);
nand (n1235,n1236,n1237);
or (n1236,n203,n491);
nand (n1237,n203,n491);
not (n1238,n1231);
nand (n1239,n1240,n1246);
or (n1240,n255,n1241);
not (n1241,n1242);
nand (n1242,n1243,n1245);
or (n1243,n1244,n253);
nand (n1245,n253,n1244);
or (n1246,n1247,n263);
nor (n1247,n1248,n1251);
and (n1248,n1249,n48);
not (n1249,n1250);
and (n1251,n1250,n253);
xor (n1252,n1253,n1326);
xor (n1253,n1254,n1284);
xor (n1254,n1255,n1274);
xor (n1255,n1256,n1266);
nand (n1256,n1257,n1262);
or (n1257,n1258,n171);
not (n1258,n1259);
nor (n1259,n1260,n1261);
and (n1260,n195,n217);
and (n1261,n215,n180);
nand (n1262,n1263,n189);
nand (n1263,n1264,n1265);
or (n1264,n222,n195);
nand (n1265,n222,n195);
nand (n1266,n1267,n1272);
or (n1267,n1268,n420);
not (n1268,n1269);
nor (n1269,n1270,n1271);
and (n1270,n370,n409);
and (n1271,n371,n407);
nand (n1272,n1273,n413);
xnor (n1273,n409,n389);
nand (n1274,n1275,n1279);
or (n1275,n103,n1276);
nor (n1276,n1277,n1278);
and (n1277,n107,n52);
and (n1278,n177,n53);
or (n1279,n104,n1280);
not (n1280,n1281);
nor (n1281,n1282,n1283);
and (n1282,n177,n61);
and (n1283,n59,n107);
xor (n1284,n1285,n1311);
xor (n1285,n1286,n1299);
nand (n1286,n1287,n1294);
or (n1287,n1288,n1290);
not (n1288,n1289);
not (n1290,n1291);
nor (n1291,n1292,n1293);
and (n1292,n1149,n465);
and (n1293,n466,n1146);
nand (n1294,n1295,n1298);
nor (n1295,n1296,n1297);
and (n1296,n1149,n476);
and (n1297,n477,n1146);
nor (n1298,n1149,n1289);
nand (n1299,n1300,n1307);
or (n1300,n1301,n315);
not (n1301,n1302);
nor (n1302,n1303,n1306);
and (n1303,n290,n1304);
not (n1304,n1305);
and (n1306,n1305,n291);
nand (n1307,n317,n1308);
nand (n1308,n1309,n1310);
or (n1309,n291,n955);
nand (n1310,n291,n955);
nand (n1311,n1312,n1319);
or (n1312,n1313,n522);
not (n1313,n1314);
nand (n1314,n1315,n1318);
or (n1315,n151,n1316);
not (n1316,n1317);
nand (n1318,n1316,n151);
nand (n1319,n1320,n374);
not (n1320,n1321);
nor (n1321,n1322,n1324);
and (n1322,n1323,n153);
and (n1324,n1325,n151);
not (n1325,n1323);
xor (n1326,n1327,n1351);
xor (n1327,n1328,n1339);
nand (n1328,n1329,n1334);
or (n1329,n400,n1330);
not (n1330,n1331);
nand (n1331,n1332,n1333);
or (n1332,n156,n395);
nand (n1333,n395,n156);
or (n1334,n1335,n529);
not (n1335,n1336);
nand (n1336,n1337,n1338);
or (n1337,n162,n395);
nand (n1338,n162,n395);
nand (n1339,n1340,n1346);
or (n1340,n470,n1341);
not (n1341,n1342);
nand (n1342,n1343,n1345);
or (n1343,n1344,n440);
nand (n1345,n1344,n440);
or (n1346,n457,n1347);
not (n1347,n1348);
nor (n1348,n1349,n1350);
and (n1349,n440,n937);
and (n1350,n935,n441);
nand (n1351,n1352,n1359);
or (n1352,n234,n1353);
not (n1353,n1354);
nor (n1354,n1355,n1358);
and (n1355,n1356,n67);
not (n1356,n1357);
and (n1358,n1357,n68);
or (n1359,n1360,n235);
nor (n1360,n1361,n1362);
and (n1361,n67,n928);
and (n1362,n68,n927);
or (n1363,n1364,n1615);
and (n1364,n1365,n1543);
xor (n1365,n1366,n1480);
or (n1366,n1367,n1479);
and (n1367,n1368,n1440);
xor (n1368,n1369,n1406);
or (n1369,n1370,n1405);
and (n1370,n1371,n1394);
xor (n1371,n1372,n1384);
nand (n1372,n1373,n1380);
or (n1373,n1374,n281);
not (n1374,n1375);
nand (n1375,n1376,n1378);
or (n1376,n1377,n265);
or (n1378,n266,n1379);
not (n1379,n1377);
nand (n1380,n1381,n288);
nand (n1381,n1382,n1383);
or (n1382,n1244,n265);
nand (n1383,n1244,n265);
nand (n1384,n1385,n1390);
or (n1385,n420,n1386);
not (n1386,n1387);
nor (n1387,n1388,n1389);
and (n1388,n409,n937);
and (n1389,n935,n407);
nand (n1390,n1391,n413);
nand (n1391,n1392,n1393);
or (n1392,n156,n409);
nand (n1393,n156,n409);
nand (n1394,n1395,n1401);
or (n1395,n457,n1396);
not (n1396,n1397);
nand (n1397,n1398,n1400);
or (n1398,n1399,n441);
not (n1399,n1210);
or (n1400,n440,n1210);
or (n1401,n470,n1402);
nor (n1402,n1403,n1404);
and (n1403,n440,n1317);
and (n1404,n441,n1316);
and (n1405,n1372,n1384);
or (n1406,n1407,n1439);
and (n1407,n1408,n1429);
xor (n1408,n1409,n1419);
nand (n1409,n1410,n1415);
or (n1410,n1144,n1411);
not (n1411,n1412);
nand (n1412,n1413,n1414);
or (n1413,n415,n371);
nand (n1414,n371,n415);
or (n1415,n1138,n1416);
nor (n1416,n1417,n1418);
and (n1417,n415,n162);
and (n1418,n416,n164);
nand (n1419,n1420,n1425);
or (n1420,n1421,n1424);
nor (n1421,n1422,n1423);
and (n1422,n1149,n389);
and (n1423,n1146,n388);
not (n1424,n1298);
or (n1425,n1426,n1288);
nor (n1426,n1427,n1428);
and (n1427,n1149,n434);
and (n1428,n1146,n521);
nand (n1429,n1430,n1435);
or (n1430,n22,n1431);
not (n1431,n1432);
nor (n1432,n1433,n1434);
and (n1433,n32,n1168);
and (n1434,n1169,n33);
or (n1435,n1436,n23);
nor (n1436,n1437,n1438);
and (n1437,n1357,n32);
and (n1438,n33,n1356);
and (n1439,n1409,n1419);
or (n1440,n1441,n1478);
and (n1441,n1442,n1465);
xor (n1442,n1443,n1453);
nand (n1443,n1444,n1449);
or (n1444,n1445,n1194);
not (n1445,n1446);
nand (n1446,n1447,n1448);
or (n1447,n1191,n59);
nand (n1448,n59,n1191);
or (n1449,n1450,n1196);
nor (n1450,n1451,n1452);
and (n1451,n1191,n279);
and (n1452,n1192,n278);
nand (n1453,n1454,n1459);
or (n1454,n438,n1455);
not (n1455,n1456);
nand (n1456,n1457,n1458);
or (n1457,n383,n1325);
or (n1458,n382,n1323);
or (n1459,n436,n1460);
nor (n1460,n1461,n1464);
and (n1461,n383,n1462);
not (n1462,n1463);
and (n1464,n382,n1463);
nand (n1465,n1466,n1472);
or (n1466,n64,n1467);
nor (n1467,n1468,n1471);
and (n1468,n1469,n75);
not (n1469,n1470);
and (n1471,n1470,n74);
or (n1472,n1473,n65);
nor (n1473,n1474,n1476);
and (n1474,n74,n1475);
and (n1476,n75,n1477);
not (n1477,n1475);
and (n1478,n1443,n1453);
and (n1479,n1369,n1406);
or (n1480,n1481,n1542);
and (n1481,n1482,n1508);
xor (n1482,n1483,n1503);
or (n1483,n1484,n1502);
and (n1484,n1485,n1497);
xor (n1485,n1486,n1491);
nor (n1486,n1487,n265);
nor (n1487,n1488,n1490);
nor (n1488,n1489,n291);
and (n1489,n1377,n286);
nor (n1490,n1377,n286);
and (n1491,n1492,n75);
nand (n1492,n1493,n1494);
or (n1493,n69,n1470);
nand (n1494,n1495,n67);
not (n1495,n1496);
and (n1496,n1470,n69);
nor (n1497,n1498,n382);
nor (n1498,n1499,n1501);
and (n1499,n1500,n440);
nand (n1500,n1463,n442);
and (n1501,n1462,n444);
and (n1502,n1486,n1491);
xor (n1503,n1504,n1507);
xor (n1504,n1505,n1506);
and (n1505,n272,n1377);
and (n1506,n333,n1470);
nor (n1507,n522,n1462);
or (n1508,n1509,n1541);
and (n1509,n1510,n1531);
xor (n1510,n1511,n1521);
nand (n1511,n1512,n1517);
or (n1512,n1513,n1223);
not (n1513,n1514);
nand (n1514,n1515,n1516);
or (n1515,n133,n203);
or (n1516,n202,n134);
nand (n1517,n1238,n1518);
nand (n1518,n1519,n1520);
or (n1519,n348,n202);
nand (n1520,n348,n202);
nand (n1521,n1522,n1526);
or (n1522,n1523,n1173);
nor (n1523,n1524,n1525);
and (n1524,n341,n1181);
and (n1525,n340,n1175);
or (n1526,n1527,n1176);
not (n1527,n1528);
nor (n1528,n1529,n1530);
and (n1529,n1181,n485);
and (n1530,n483,n1175);
nand (n1531,n1532,n1537);
or (n1532,n171,n1533);
not (n1533,n1534);
nand (n1534,n1535,n1536);
or (n1535,n1130,n180);
or (n1536,n195,n1131);
or (n1537,n1538,n172);
nor (n1538,n1539,n1540);
and (n1539,n1305,n195);
and (n1540,n180,n1304);
and (n1541,n1511,n1521);
and (n1542,n1483,n1503);
xor (n1543,n1544,n1568);
xor (n1544,n1545,n1548);
or (n1545,n1546,n1547);
and (n1546,n1504,n1507);
and (n1547,n1505,n1506);
xor (n1548,n1549,n1562);
xor (n1549,n1550,n1556);
and (n1550,n1551,n48);
nand (n1551,n1552,n1553);
or (n1552,n259,n1377);
nand (n1553,n1554,n265);
not (n1554,n1555);
and (n1555,n1377,n259);
nor (n1556,n1557,n153);
not (n1557,n1558);
nand (n1558,n1559,n1560);
or (n1559,n1463,n378);
nand (n1560,n1561,n382);
nand (n1561,n1463,n378);
nor (n1562,n1563,n127);
nor (n1563,n1564,n1566);
and (n1564,n1565,n74);
nand (n1565,n1470,n335);
and (n1566,n1469,n1567);
not (n1567,n335);
or (n1568,n1569,n1614);
and (n1569,n1570,n1605);
xor (n1570,n1571,n1583);
nand (n1571,n1572,n1578);
or (n1572,n400,n1573);
not (n1573,n1574);
nor (n1574,n1575,n1577);
and (n1575,n395,n1576);
not (n1576,n1344);
and (n1577,n1344,n396);
or (n1578,n1579,n529);
not (n1579,n1580);
nand (n1580,n1581,n1582);
or (n1581,n935,n395);
nand (n1582,n935,n395);
nand (n1583,n1584,n1600);
or (n1584,n1585,n1590);
not (n1585,n1586);
nand (n1586,n1587,n1589);
or (n1587,n53,n1588);
not (n1588,n100);
nand (n1589,n53,n1588);
not (n1590,n1591);
and (n1591,n1592,n1597);
nand (n1592,n1593,n1596);
or (n1593,n1594,n100);
not (n1594,n1595);
nand (n1596,n100,n1594);
nor (n1597,n1598,n1599);
and (n1598,n1191,n1595);
and (n1599,n1192,n1594);
nand (n1600,n1601,n1602);
not (n1601,n1597);
nor (n1602,n1603,n1604);
and (n1603,n61,n1588);
and (n1604,n59,n100);
nand (n1605,n1606,n1610);
or (n1606,n315,n1607);
nor (n1607,n1608,n1609);
and (n1608,n1125,n290);
and (n1609,n291,n1124);
or (n1610,n1611,n316);
nor (n1611,n1612,n1613);
and (n1612,n290,n1131);
and (n1613,n1130,n291);
and (n1614,n1571,n1583);
and (n1615,n1366,n1480);
and (n1616,n1104,n1252);
xor (n1617,n1618,n1735);
xor (n1618,n1619,n1665);
xor (n1619,n1620,n1627);
xor (n1620,n1621,n1624);
or (n1621,n1622,n1623);
and (n1622,n1204,n1239);
and (n1623,n1205,n1217);
or (n1624,n1625,n1626);
and (n1625,n1156,n1187);
and (n1626,n1157,n1171);
or (n1627,n1628,n1664);
and (n1628,n1629,n1653);
xor (n1629,n1630,n1642);
nand (n1630,n1631,n1636);
or (n1631,n532,n1632);
not (n1632,n1633);
nor (n1633,n1634,n1635);
and (n1634,n1477,n127);
and (n1635,n1475,n128);
or (n1636,n332,n1637);
nor (n1637,n1638,n1640);
and (n1638,n127,n1639);
and (n1640,n1641,n128);
not (n1641,n1639);
nand (n1642,n1643,n1648);
or (n1643,n1590,n1644);
not (n1644,n1645);
nor (n1645,n1646,n1647);
and (n1646,n278,n1588);
and (n1647,n279,n100);
or (n1648,n1597,n1649);
not (n1649,n1650);
nand (n1650,n1651,n1652);
or (n1651,n100,n296);
nand (n1652,n100,n296);
nand (n1653,n1654,n1660);
or (n1654,n22,n1655);
not (n1655,n1656);
or (n1656,n1657,n1658);
and (n1657,n114,n32);
and (n1658,n1659,n33);
not (n1659,n114);
or (n1660,n1661,n23);
nor (n1661,n1662,n1663);
and (n1662,n134,n32);
and (n1663,n133,n33);
and (n1664,n1630,n1642);
xor (n1665,n1666,n1714);
xor (n1666,n1667,n1687);
xor (n1667,n1668,n1681);
xor (n1668,n1669,n1675);
nand (n1669,n1670,n1671);
nand (n1670,n1650,n1597,n1592);
nand (n1671,n1601,n1672);
nand (n1672,n1673,n1674);
or (n1673,n313,n1588);
nand (n1674,n313,n1588);
nand (n1675,n1676,n1677);
nand (n1676,n1213,n438,n445);
nand (n1677,n1678,n449);
nand (n1678,n1679,n1680);
or (n1679,n1344,n382);
nand (n1680,n1344,n382);
nand (n1681,n1682,n1683);
or (n1682,n1347,n470);
nand (n1683,n1684,n566);
nand (n1684,n1685,n1686);
or (n1685,n441,n158);
nand (n1686,n158,n441);
xor (n1687,n1688,n1707);
xor (n1688,n1689,n1696);
nand (n1689,n1690,n1695);
or (n1690,n424,n1691);
not (n1691,n1692);
nor (n1692,n1693,n1694);
and (n1693,n409,n521);
and (n1694,n434,n407);
nand (n1695,n1273,n421,n424);
nand (n1696,n1697,n1702);
or (n1697,n1698,n37);
not (n1698,n1699);
nor (n1699,n1700,n1701);
and (n1700,n41,n1379);
and (n1701,n1377,n42);
nand (n1702,n1703,n46);
nand (n1703,n1704,n1706);
or (n1704,n42,n1705);
not (n1705,n1244);
nand (n1706,n1705,n42);
nand (n1707,n1708,n1710);
or (n1708,n171,n1709);
not (n1709,n1263);
or (n1710,n1711,n172);
nor (n1711,n1712,n1713);
and (n1712,n195,n53);
and (n1713,n52,n180);
xor (n1714,n1715,n1729);
xor (n1715,n1716,n1722);
nand (n1716,n1717,n1718);
or (n1717,n532,n1637);
nand (n1718,n1719,n333);
nand (n1719,n1720,n1721);
or (n1720,n1163,n127);
nand (n1721,n1163,n127);
nand (n1722,n1723,n1725);
or (n1723,n1724,n1223);
not (n1724,n1235);
nand (n1725,n1726,n1238);
nand (n1726,n1727,n1728);
or (n1727,n79,n202);
nand (n1728,n202,n79);
nand (n1729,n1730,n1731);
or (n1730,n255,n1247);
or (n1731,n1732,n263);
nor (n1732,n1733,n1734);
and (n1733,n253,n1125);
and (n1734,n48,n1124);
xor (n1735,n1736,n1784);
xor (n1736,n1737,n1762);
xor (n1737,n1738,n1755);
xor (n1738,n1739,n1745);
nand (n1739,n1740,n1741);
or (n1740,n1313,n373);
nand (n1741,n1742,n380);
nor (n1742,n1743,n1744);
and (n1743,n1210,n151);
and (n1744,n153,n1399);
nand (n1745,n1746,n1751);
or (n1746,n1747,n118);
not (n1747,n1748);
nor (n1748,n1749,n1750);
and (n1749,n115,n1469);
and (n1750,n1470,n116);
nand (n1751,n1752,n125);
nor (n1752,n1753,n1754);
and (n1753,n115,n1477);
and (n1754,n1475,n116);
nand (n1755,n1756,n1758);
or (n1756,n1757,n281);
not (n1757,n1128);
nand (n1758,n288,n1759);
nand (n1759,n1760,n1761);
or (n1760,n1305,n265);
nand (n1761,n265,n1305);
xor (n1762,n1763,n1777);
xor (n1763,n1764,n1771);
nand (n1764,n1765,n1767);
or (n1765,n1766,n315);
not (n1766,n1308);
nand (n1767,n1768,n317);
nor (n1768,n1769,n1770);
and (n1769,n290,n217);
and (n1770,n215,n291);
nand (n1771,n1772,n1776);
nand (n1772,n1773,n1197);
nor (n1773,n1774,n1775);
and (n1774,n1191,n185);
and (n1775,n186,n1192);
nand (n1776,n1200,n1195);
nand (n1777,n1778,n1780);
or (n1778,n1779,n64);
not (n1779,n1166);
nand (n1780,n1781,n1006);
nor (n1781,n1782,n1783);
and (n1782,n74,n1356);
and (n1783,n1357,n75);
xor (n1784,n1785,n1799);
xor (n1785,n1786,n1792);
nand (n1786,n1787,n1788);
or (n1787,n1280,n103);
nand (n1788,n1789,n96);
nand (n1789,n1790,n1791);
or (n1790,n177,n279);
nand (n1791,n279,n177);
nand (n1792,n1793,n1798);
or (n1793,n1144,n1794);
not (n1794,n1795);
nand (n1795,n1796,n1797);
or (n1796,n416,n476);
or (n1797,n477,n415);
nand (n1798,n1139,n1151);
nand (n1799,n1800,n1801);
or (n1800,n234,n1360);
or (n1801,n235,n1802);
nor (n1802,n1803,n1804);
and (n1803,n1659,n68);
and (n1804,n114,n67);
xor (n1805,n1806,n1981);
xor (n1806,n1807,n1886);
xor (n1807,n1808,n1857);
xor (n1808,n1809,n1835);
xor (n1809,n1810,n1828);
xor (n1810,n1811,n1821);
nand (n1811,n1812,n1817);
or (n1812,n149,n1813);
not (n1813,n1814);
nand (n1814,n1815,n1816);
or (n1815,n147,n1323);
nand (n1816,n1323,n147);
or (n1817,n138,n1818);
nor (n1818,n1819,n1820);
and (n1819,n144,n1462);
and (n1820,n1463,n147);
nand (n1821,n1822,n1824);
or (n1822,n1823,n199);
not (n1823,n1115);
nand (n1824,n1825,n1118);
nand (n1825,n1826,n1827);
or (n1826,n28,n485);
nand (n1827,n28,n485);
nand (n1828,n1829,n1830);
or (n1829,n1290,n1424);
or (n1830,n1831,n1288);
not (n1831,n1832);
nor (n1832,n1833,n1834);
and (n1833,n1149,n399);
and (n1834,n397,n1146);
xor (n1835,n1836,n1850);
xor (n1836,n1837,n1844);
nand (n1837,n1838,n1840);
or (n1838,n1173,n1839);
not (n1839,n1184);
nand (n1840,n1841,n1177);
nor (n1841,n1842,n1843);
and (n1842,n1181,n360);
and (n1843,n358,n1175);
nand (n1844,n1845,n1846);
or (n1845,n1335,n400);
nand (n1846,n1847,n405);
nand (n1847,n1848,n1849);
or (n1848,n396,n370);
nand (n1849,n396,n370);
nand (n1850,n1851,n1856);
or (n1851,n23,n1852);
not (n1852,n1853);
nor (n1853,n1854,n1855);
and (n1854,n32,n347);
and (n1855,n348,n33);
or (n1856,n22,n1661);
xor (n1857,n1858,n1883);
xor (n1858,n1859,n1866);
or (n1859,n1860,n1865);
and (n1860,n1861,n1864);
xor (n1861,n1862,n1863);
and (n1862,n46,n1377);
and (n1863,n148,n1463);
nor (n1864,n664,n1469);
and (n1865,n1862,n1863);
xor (n1866,n1867,n1878);
xor (n1867,n1868,n1873);
nor (n1868,n1869,n41);
nor (n1869,n1870,n1871);
and (n1870,n1379,n45);
nor (n1871,n1872,n48);
and (n1872,n1377,n43);
and (n1873,n1874,n144);
nand (n1874,n1875,n1877);
or (n1875,n1876,n151);
and (n1876,n1463,n143);
or (n1877,n1463,n143);
nor (n1878,n1879,n115);
nor (n1879,n1880,n1882);
and (n1880,n1881,n127);
nand (n1881,n1470,n122);
and (n1882,n1469,n124);
or (n1883,n1884,n1885);
and (n1884,n1285,n1311);
and (n1885,n1286,n1299);
or (n1886,n1887,n1980);
and (n1887,n1888,n1977);
xor (n1888,n1889,n1890);
xor (n1889,n1629,n1653);
or (n1890,n1891,n1976);
and (n1891,n1892,n1942);
xor (n1892,n1893,n1918);
or (n1893,n1894,n1917);
and (n1894,n1895,n1910);
xor (n1895,n1896,n1903);
nand (n1896,n1897,n1899);
or (n1897,n1898,n1223);
not (n1898,n1518);
nand (n1899,n1900,n1238);
nor (n1900,n1901,n1902);
and (n1901,n202,n340);
and (n1902,n341,n203);
nand (n1903,n1904,n1909);
or (n1904,n1176,n1905);
not (n1905,n1906);
nor (n1906,n1907,n1908);
and (n1907,n1181,n491);
and (n1908,n489,n1175);
nand (n1909,n1528,n1174);
nand (n1910,n1911,n1916);
or (n1911,n172,n1912);
not (n1912,n1913);
nor (n1913,n1914,n1915);
and (n1914,n195,n955);
and (n1915,n956,n180);
or (n1916,n171,n1538);
and (n1917,n1896,n1903);
or (n1918,n1919,n1941);
and (n1919,n1920,n1934);
xor (n1920,n1921,n1928);
nand (n1921,n1922,n1927);
or (n1922,n1196,n1923);
not (n1923,n1924);
nor (n1924,n1925,n1926);
and (n1925,n296,n1191);
and (n1926,n297,n1192);
or (n1927,n1450,n1194);
nand (n1928,n1929,n1930);
or (n1929,n1455,n436);
nand (n1930,n449,n1931);
nand (n1931,n1932,n1933);
or (n1932,n1317,n382);
nand (n1933,n382,n1317);
nand (n1934,n1935,n1936);
or (n1935,n64,n1473);
or (n1936,n1937,n65);
not (n1937,n1938);
nand (n1938,n1939,n1940);
or (n1939,n75,n1641);
or (n1940,n1639,n74);
and (n1941,n1921,n1928);
or (n1942,n1943,n1975);
and (n1943,n1944,n1965);
xor (n1944,n1945,n1955);
nand (n1945,n1946,n1951);
or (n1946,n1947,n234);
not (n1947,n1948);
nand (n1948,n1949,n1950);
or (n1949,n1163,n67);
nand (n1950,n1163,n67);
nand (n1951,n1952,n247);
nor (n1952,n1953,n1954);
and (n1953,n67,n1168);
and (n1954,n1169,n68);
nand (n1955,n1956,n1961);
or (n1956,n1957,n103);
not (n1957,n1958);
nor (n1958,n1959,n1960);
and (n1959,n177,n217);
and (n1960,n215,n107);
nand (n1961,n1962,n96);
nor (n1962,n1963,n1964);
and (n1963,n222,n107);
and (n1964,n221,n177);
nand (n1965,n1966,n1971);
or (n1966,n1967,n199);
not (n1967,n1968);
nand (n1968,n1969,n1970);
or (n1969,n28,n1659);
or (n1970,n209,n114);
nand (n1971,n1118,n1972);
nand (n1972,n1973,n1974);
or (n1973,n134,n209);
or (n1974,n28,n133);
and (n1975,n1945,n1955);
and (n1976,n1893,n1918);
or (n1977,n1978,n1979);
and (n1978,n1544,n1568);
and (n1979,n1545,n1548);
and (n1980,n1889,n1890);
or (n1981,n1982,n2126);
and (n1982,n1983,n2067);
xor (n1983,n1984,n2009);
xor (n1984,n1985,n1990);
xor (n1985,n1986,n1989);
or (n1986,n1987,n1988);
and (n1987,n1549,n1562);
and (n1988,n1550,n1556);
xor (n1989,n1861,n1864);
or (n1990,n1991,n2008);
and (n1991,n1992,n2001);
xor (n1992,n1993,n1997);
nand (n1993,n1994,n1996);
or (n1994,n1995,n436);
not (n1995,n1931);
nand (n1996,n1208,n449);
nand (n1997,n1998,n2000);
or (n1998,n1999,n1223);
not (n1999,n1900);
nand (n2000,n1220,n1238);
nand (n2001,n2002,n2007);
or (n2002,n2003,n255);
not (n2003,n2004);
nand (n2004,n2005,n2006);
or (n2005,n1377,n253);
or (n2006,n1379,n48);
nand (n2007,n1242,n272);
and (n2008,n1993,n1997);
xor (n2009,n2010,n2054);
xor (n2010,n2011,n2032);
or (n2011,n2012,n2031);
and (n2012,n2013,n2025);
xor (n2013,n2014,n2021);
nand (n2014,n2015,n2020);
or (n2015,n2016,n532);
not (n2016,n2017);
nor (n2017,n2018,n2019);
and (n2018,n1469,n127);
and (n2019,n1470,n128);
nand (n2020,n1633,n333);
nand (n2021,n2022,n2024);
or (n2022,n2023,n1590);
not (n2023,n1602);
nand (n2024,n1645,n1601);
nand (n2025,n2026,n2030);
or (n2026,n22,n2027);
nor (n2027,n2028,n2029);
and (n2028,n32,n928);
and (n2029,n33,n927);
nand (n2030,n1656,n24);
and (n2031,n2014,n2021);
or (n2032,n2033,n2053);
and (n2033,n2034,n2046);
xor (n2034,n2035,n2039);
nand (n2035,n2036,n2038);
or (n2036,n2037,n199);
not (n2037,n1972);
nand (n2038,n1118,n1111);
nand (n2039,n2040,n2045);
or (n2040,n281,n2041);
not (n2041,n2042);
nor (n2042,n2043,n2044);
and (n2043,n1249,n265);
and (n2044,n1250,n266);
nand (n2045,n288,n1122);
nand (n2046,n2047,n2052);
or (n2047,n1138,n2048);
not (n2048,n2049);
nor (n2049,n2050,n2051);
and (n2050,n415,n388);
and (n2051,n389,n416);
or (n2052,n1135,n1144);
and (n2053,n2035,n2039);
or (n2054,n2055,n2066);
and (n2055,n2056,n2063);
xor (n2056,n2057,n2060);
nand (n2057,n2058,n2059);
or (n2058,n1937,n64);
nand (n2059,n1160,n1006);
nand (n2060,n2061,n2062);
or (n2061,n1176,n1178);
nand (n2062,n1906,n1174);
nand (n2063,n2064,n2065);
or (n2064,n1194,n1923);
or (n2065,n1189,n1196);
and (n2066,n2057,n2060);
or (n2067,n2068,n2125);
and (n2068,n2069,n2109);
xor (n2069,n2070,n2093);
or (n2070,n2071,n2092);
and (n2071,n2072,n2084);
xor (n2072,n2073,n2077);
nand (n2073,n2074,n2076);
or (n2074,n2075,n281);
not (n2075,n1381);
nand (n2076,n2042,n288);
nand (n2077,n2078,n2083);
or (n2078,n424,n2079);
not (n2079,n2080);
nor (n2080,n2081,n2082);
and (n2081,n162,n407);
and (n2082,n164,n409);
nand (n2083,n419,n1391);
nand (n2084,n2085,n2086);
or (n2085,n470,n1396);
or (n2086,n2087,n457);
not (n2087,n2088);
nor (n2088,n2089,n2091);
and (n2089,n440,n2090);
not (n2090,n1215);
and (n2091,n1215,n441);
and (n2092,n2073,n2077);
or (n2093,n2094,n2108);
and (n2094,n2095,n2105);
xor (n2095,n2096,n2099);
nand (n2096,n2097,n2098);
or (n2097,n1411,n1138);
nand (n2098,n2049,n1154);
nand (n2099,n2100,n2101);
or (n2100,n1426,n1424);
or (n2101,n2102,n1288);
nor (n2102,n2103,n2104);
and (n2103,n453,n1149);
and (n2104,n452,n1146);
nand (n2105,n2106,n2107);
or (n2106,n22,n1436);
or (n2107,n2027,n23);
and (n2108,n2096,n2099);
xor (n2109,n2110,n2119);
xor (n2110,n2111,n2115);
nand (n2111,n2112,n2114);
or (n2112,n1288,n2113);
not (n2113,n1295);
or (n2114,n2102,n1424);
nand (n2115,n2116,n2117);
or (n2116,n316,n1301);
nand (n2117,n2118,n656);
not (n2118,n1611);
nand (n2119,n2120,n2124);
or (n2120,n373,n2121);
nor (n2121,n2122,n2123);
and (n2122,n1462,n151);
and (n2123,n1463,n153);
or (n2124,n1321,n522);
and (n2125,n2070,n2093);
and (n2126,n1984,n2009);
xor (n2127,n2128,n2284);
xor (n2128,n2129,n2249);
or (n2129,n2130,n2248);
and (n2130,n2131,n2199);
xor (n2131,n2132,n2133);
xor (n2132,n1888,n1977);
or (n2133,n2134,n2198);
and (n2134,n2135,n2191);
xor (n2135,n2136,n2190);
or (n2136,n2137,n2189);
and (n2137,n2138,n2188);
xor (n2138,n2139,n2164);
or (n2139,n2140,n2163);
and (n2140,n2141,n2156);
xor (n2141,n2142,n2149);
nand (n2142,n2143,n2148);
or (n2143,n2144,n400);
not (n2144,n2145);
nor (n2145,n2146,n2147);
and (n2146,n395,n2090);
and (n2147,n1215,n396);
nand (n2148,n1574,n405);
nand (n2149,n2150,n2155);
or (n2150,n2151,n1590);
not (n2151,n2152);
nor (n2152,n2153,n2154);
and (n2153,n221,n1588);
and (n2154,n222,n100);
nand (n2155,n1586,n1601);
nand (n2156,n2157,n2162);
or (n2157,n315,n2158);
not (n2158,n2159);
nor (n2159,n2160,n2161);
and (n2160,n290,n1249);
and (n2161,n1250,n291);
or (n2162,n1607,n316);
and (n2163,n2142,n2149);
or (n2164,n2165,n2187);
and (n2165,n2166,n2181);
xor (n2166,n2167,n2174);
nand (n2167,n2168,n2173);
or (n2168,n2169,n234);
not (n2169,n2170);
nand (n2170,n2171,n2172);
or (n2171,n68,n1641);
nand (n2172,n68,n1641);
nand (n2173,n1948,n247);
nand (n2174,n2175,n2180);
or (n2175,n2176,n103);
not (n2176,n2177);
nand (n2177,n2178,n2179);
or (n2178,n107,n955);
nand (n2179,n955,n107);
nand (n2180,n1958,n96);
not (n2181,n2182);
nor (n2182,n2183,n2184);
and (n2183,n1118,n1968);
and (n2184,n2185,n2186);
not (n2185,n199);
xor (n2186,n928,n28);
and (n2187,n2167,n2174);
xor (n2188,n1944,n1965);
and (n2189,n2139,n2164);
xor (n2190,n2069,n2109);
or (n2191,n2192,n2197);
and (n2192,n2193,n2196);
xor (n2193,n2194,n2195);
xor (n2194,n1570,n1605);
xor (n2195,n2072,n2084);
xor (n2196,n1895,n1910);
and (n2197,n2194,n2195);
and (n2198,n2136,n2190);
xor (n2199,n2200,n2241);
xor (n2200,n2201,n2219);
or (n2201,n2202,n2218);
and (n2202,n2203,n2217);
xor (n2203,n2204,n2205);
xor (n2204,n1992,n2001);
xor (n2205,n2206,n2213);
xor (n2206,n2207,n2210);
nand (n2207,n2208,n2209);
or (n2208,n1579,n400);
nand (n2209,n1331,n405);
nand (n2210,n2211,n2212);
or (n2211,n2087,n470);
nand (n2212,n1342,n566);
nand (n2213,n2214,n2216);
or (n2214,n2215,n234);
not (n2215,n1952);
nand (n2216,n1354,n247);
xor (n2217,n2056,n2063);
and (n2218,n2204,n2205);
xor (n2219,n2220,n2238);
xor (n2220,n2221,n2235);
or (n2221,n2222,n2234);
and (n2222,n2223,n2230);
xor (n2223,n2224,n2227);
nand (n2224,n2225,n2226);
or (n2225,n1912,n171);
nand (n2226,n1259,n189);
nand (n2227,n2228,n2229);
or (n2228,n2079,n420);
nand (n2229,n1269,n413);
nand (n2230,n2231,n2233);
or (n2231,n103,n2232);
not (n2232,n1962);
or (n2233,n1276,n104);
and (n2234,n2224,n2227);
or (n2235,n2236,n2237);
and (n2236,n2206,n2213);
and (n2237,n2207,n2210);
or (n2238,n2239,n2240);
and (n2239,n2110,n2119);
and (n2240,n2111,n2115);
or (n2241,n2242,n2247);
and (n2242,n2243,n2246);
xor (n2243,n2244,n2245);
xor (n2244,n2013,n2025);
xor (n2245,n2034,n2046);
xor (n2246,n2223,n2230);
and (n2247,n2244,n2245);
and (n2248,n2132,n2133);
xor (n2249,n2250,n2265);
xor (n2250,n2251,n2254);
or (n2251,n2252,n2253);
and (n2252,n2200,n2241);
and (n2253,n2201,n2219);
xor (n2254,n2255,n2262);
xor (n2255,n2256,n2259);
or (n2256,n2257,n2258);
and (n2257,n2010,n2054);
and (n2258,n2011,n2032);
or (n2259,n2260,n2261);
and (n2260,n2220,n2238);
and (n2261,n2221,n2235);
or (n2262,n2263,n2264);
and (n2263,n1985,n1990);
and (n2264,n1986,n1989);
xor (n2265,n2266,n2273);
xor (n2266,n2267,n2270);
or (n2267,n2268,n2269);
and (n2268,n1105,n1203);
and (n2269,n1106,n1155);
or (n2270,n2271,n2272);
and (n2271,n1253,n1326);
and (n2272,n1254,n1284);
xor (n2273,n2274,n2281);
xor (n2274,n2275,n2278);
or (n2275,n2276,n2277);
and (n2276,n1255,n1274);
and (n2277,n1256,n1266);
or (n2278,n2279,n2280);
and (n2279,n1327,n1351);
and (n2280,n1328,n1339);
or (n2281,n2282,n2283);
and (n2282,n1107,n1133);
and (n2283,n1108,n1119);
or (n2284,n2285,n2296);
and (n2285,n2286,n2295);
xor (n2286,n2287,n2294);
or (n2287,n2288,n2293);
and (n2288,n2289,n2292);
xor (n2289,n2290,n2291);
xor (n2290,n1892,n1942);
xor (n2291,n2203,n2217);
xor (n2292,n2243,n2246);
and (n2293,n2290,n2291);
xor (n2294,n1983,n2067);
xor (n2295,n1103,n1363);
and (n2296,n2287,n2294);
or (n2297,n2298,n2479);
and (n2298,n2299,n2431);
xor (n2299,n2300,n2430);
or (n2300,n2301,n2429);
and (n2301,n2302,n2347);
xor (n2302,n2303,n2346);
or (n2303,n2304,n2345);
and (n2304,n2305,n2308);
xor (n2305,n2306,n2307);
xor (n2306,n2095,n2105);
xor (n2307,n1920,n1934);
or (n2308,n2309,n2344);
and (n2309,n2310,n2319);
xor (n2310,n2311,n2318);
or (n2311,n2312,n2317);
and (n2312,n2313,n2316);
xor (n2313,n2314,n2315);
nor (n2314,n730,n1379);
and (n2315,n1006,n1470);
nor (n2316,n438,n1462);
and (n2317,n2314,n2315);
xor (n2318,n1485,n1497);
or (n2319,n2320,n2343);
and (n2320,n2321,n2336);
xor (n2321,n2322,n2329);
nand (n2322,n2323,n2328);
or (n2323,n1194,n2324);
not (n2324,n2325);
nor (n2325,n2326,n2327);
and (n2326,n1191,n52);
and (n2327,n53,n1192);
nand (n2328,n1446,n1197);
nand (n2329,n2330,n2335);
or (n2330,n2331,n420);
not (n2331,n2332);
nor (n2332,n2333,n2334);
and (n2333,n1344,n407);
and (n2334,n1576,n409);
nand (n2335,n1387,n413);
nand (n2336,n2337,n2342);
or (n2337,n2338,n315);
not (n2338,n2339);
nor (n2339,n2340,n2341);
and (n2340,n1244,n291);
and (n2341,n1705,n290);
nand (n2342,n317,n2159);
and (n2343,n2322,n2329);
and (n2344,n2311,n2318);
and (n2345,n2306,n2307);
xor (n2346,n1365,n1543);
or (n2347,n2348,n2428);
and (n2348,n2349,n2427);
xor (n2349,n2350,n2351);
xor (n2350,n1482,n1508);
or (n2351,n2352,n2426);
and (n2352,n2353,n2402);
xor (n2353,n2354,n2378);
or (n2354,n2355,n2377);
and (n2355,n2356,n2371);
xor (n2356,n2357,n2364);
nand (n2357,n2358,n2363);
or (n2358,n2359,n22);
not (n2359,n2360);
nor (n2360,n2361,n2362);
and (n2361,n32,n1162);
and (n2362,n1163,n33);
nand (n2363,n1432,n24);
nand (n2364,n2365,n2370);
or (n2365,n2366,n470);
not (n2366,n2367);
nand (n2367,n2368,n2369);
or (n2368,n441,n1325);
nand (n2369,n441,n1325);
or (n2370,n1402,n457);
nand (n2371,n2372,n2376);
or (n2372,n2373,n1173);
nor (n2373,n2374,n2375);
and (n2374,n1181,n348);
and (n2375,n1175,n347);
or (n2376,n1523,n1176);
and (n2377,n2357,n2364);
or (n2378,n2379,n2401);
and (n2379,n2380,n2395);
xor (n2380,n2381,n2388);
nand (n2381,n2382,n2387);
or (n2382,n2383,n1590);
not (n2383,n2384);
nand (n2384,n2385,n2386);
or (n2385,n217,n100);
or (n2386,n1588,n215);
nand (n2387,n1601,n2152);
nand (n2388,n2389,n2394);
or (n2389,n2390,n171);
not (n2390,n2391);
nor (n2391,n2392,n2393);
and (n2392,n195,n1124);
and (n2393,n1125,n180);
nand (n2394,n1534,n189);
nand (n2395,n2396,n2400);
or (n2396,n1223,n2397);
nor (n2397,n2398,n2399);
and (n2398,n202,n114);
and (n2399,n203,n1659);
or (n2400,n1231,n1513);
and (n2401,n2381,n2388);
or (n2402,n2403,n2425);
and (n2403,n2404,n2419);
xor (n2404,n2405,n2412);
nand (n2405,n2406,n2411);
or (n2406,n2407,n103);
not (n2407,n2408);
nand (n2408,n2409,n2410);
or (n2409,n107,n1304);
nand (n2410,n1304,n107);
nand (n2411,n96,n2177);
nand (n2412,n2413,n2418);
or (n2413,n2414,n199);
not (n2414,n2415);
nor (n2415,n2416,n2417);
and (n2416,n1357,n28);
and (n2417,n1356,n209);
nand (n2418,n2186,n1118);
nand (n2419,n2420,n2424);
or (n2420,n400,n2421);
nor (n2421,n2422,n2423);
and (n2422,n395,n1210);
and (n2423,n396,n1399);
or (n2424,n2144,n529);
and (n2425,n2405,n2412);
and (n2426,n2354,n2378);
xor (n2427,n2138,n2188);
and (n2428,n2350,n2351);
and (n2429,n2303,n2346);
xor (n2430,n2131,n2199);
or (n2431,n2432,n2478);
and (n2432,n2433,n2477);
xor (n2433,n2434,n2476);
or (n2434,n2435,n2475);
and (n2435,n2436,n2468);
xor (n2436,n2437,n2467);
or (n2437,n2438,n2466);
and (n2438,n2439,n2465);
xor (n2439,n2440,n2464);
or (n2440,n2441,n2463);
and (n2441,n2442,n2457);
xor (n2442,n2443,n2450);
nand (n2443,n2444,n2449);
or (n2444,n2445,n234);
not (n2445,n2446);
nand (n2446,n2447,n2448);
or (n2447,n1475,n67);
nand (n2448,n1475,n67);
nand (n2449,n2170,n247);
nand (n2450,n2451,n2456);
or (n2451,n2452,n1138);
not (n2452,n2453);
nor (n2453,n2454,n2455);
and (n2454,n415,n158);
and (n2455,n156,n416);
or (n2456,n1416,n1144);
nand (n2457,n2458,n2462);
or (n2458,n2459,n1424);
nor (n2459,n2460,n2461);
and (n2460,n371,n1149);
and (n2461,n370,n1146);
or (n2462,n1421,n1288);
and (n2463,n2443,n2450);
xor (n2464,n2166,n2181);
xor (n2465,n2141,n2156);
and (n2466,n2440,n2464);
xor (n2467,n1368,n1440);
or (n2468,n2469,n2474);
and (n2469,n2470,n2473);
xor (n2470,n2471,n2472);
xor (n2471,n1371,n1394);
xor (n2472,n1510,n1531);
xor (n2473,n1442,n1465);
and (n2474,n2471,n2472);
and (n2475,n2437,n2467);
xor (n2476,n2135,n2191);
xor (n2477,n2289,n2292);
and (n2478,n2434,n2476);
and (n2479,n2300,n2430);
or (n2480,n2481,n2675);
and (n2481,n2482,n2674);
xor (n2482,n2483,n2484);
xor (n2483,n2286,n2295);
or (n2484,n2485,n2673);
and (n2485,n2486,n2624);
xor (n2486,n2487,n2623);
or (n2487,n2488,n2622);
and (n2488,n2489,n2621);
xor (n2489,n2490,n2491);
xor (n2490,n2193,n2196);
or (n2491,n2492,n2620);
and (n2492,n2493,n2568);
xor (n2493,n2494,n2495);
xor (n2494,n1408,n1429);
or (n2495,n2496,n2567);
and (n2496,n2497,n2544);
xor (n2497,n2498,n2521);
or (n2498,n2499,n2520);
and (n2499,n2500,n2514);
xor (n2500,n2501,n2508);
nand (n2501,n2502,n2507);
or (n2502,n2503,n22);
not (n2503,n2504);
nand (n2504,n2505,n2506);
or (n2505,n33,n1641);
nand (n2506,n1641,n33);
nand (n2507,n2360,n24);
nand (n2508,n2509,n2513);
or (n2509,n470,n2510);
nor (n2510,n2511,n2512);
and (n2511,n1462,n441);
and (n2512,n1463,n440);
nand (n2513,n566,n2367);
nand (n2514,n2515,n2519);
or (n2515,n2516,n1173);
nor (n2516,n2517,n2518);
and (n2517,n1181,n134);
and (n2518,n1175,n133);
or (n2519,n2373,n1176);
and (n2520,n2501,n2508);
or (n2521,n2522,n2543);
and (n2522,n2523,n2537);
xor (n2523,n2524,n2531);
nand (n2524,n2525,n2530);
or (n2525,n2526,n103);
not (n2526,n2527);
nand (n2527,n2528,n2529);
or (n2528,n1131,n177);
nand (n2529,n1131,n177);
nand (n2530,n2408,n96);
nand (n2531,n2532,n2533);
or (n2532,n200,n2414);
nand (n2533,n2185,n2534);
nand (n2534,n2535,n2536);
or (n2535,n28,n1168);
nand (n2536,n28,n1168);
nand (n2537,n2538,n2542);
or (n2538,n400,n2539);
nor (n2539,n2540,n2541);
and (n2540,n395,n1317);
and (n2541,n1316,n396);
or (n2542,n2421,n529);
and (n2543,n2524,n2531);
or (n2544,n2545,n2566);
and (n2545,n2546,n2560);
xor (n2546,n2547,n2553);
nand (n2547,n2548,n2552);
or (n2548,n2549,n1194);
nor (n2549,n2550,n2551);
and (n2550,n1191,n222);
and (n2551,n1192,n221);
or (n2552,n2324,n1196);
nand (n2553,n2554,n2555);
or (n2554,n424,n2331);
or (n2555,n420,n2556);
not (n2556,n2557);
nand (n2557,n2558,n2559);
or (n2558,n1215,n409);
nand (n2559,n409,n1215);
nand (n2560,n2561,n2565);
or (n2561,n315,n2562);
nor (n2562,n2563,n2564);
and (n2563,n1379,n291);
and (n2564,n1377,n290);
or (n2565,n2338,n316);
and (n2566,n2547,n2553);
and (n2567,n2498,n2521);
or (n2568,n2569,n2619);
and (n2569,n2570,n2595);
xor (n2570,n2571,n2594);
or (n2571,n2572,n2593);
and (n2572,n2573,n2586);
xor (n2573,n2574,n2581);
and (n2574,n2575,n291);
nand (n2575,n2576,n2579);
nand (n2576,n2577,n195);
not (n2577,n2578);
and (n2578,n1377,n319);
nand (n2579,n1379,n2580);
not (n2580,n319);
and (n2581,n2582,n68);
nand (n2582,n2583,n2584);
or (n2583,n1470,n237);
nand (n2584,n2585,n32);
nand (n2585,n1470,n237);
nor (n2586,n2587,n440);
and (n2587,n2588,n2591);
not (n2588,n2589);
nor (n2589,n2590,n396);
and (n2590,n1463,n459);
not (n2591,n2592);
nor (n2592,n1463,n459);
and (n2593,n2574,n2581);
xor (n2594,n2313,n2316);
or (n2595,n2596,n2618);
and (n2596,n2597,n2611);
xor (n2597,n2598,n2605);
nand (n2598,n2599,n2604);
or (n2599,n2600,n1590);
not (n2600,n2601);
nand (n2601,n2602,n2603);
or (n2602,n955,n100);
or (n2603,n1588,n956);
nand (n2604,n1601,n2384);
nand (n2605,n2606,n2610);
or (n2606,n171,n2607);
nor (n2607,n2608,n2609);
and (n2608,n1250,n195);
and (n2609,n1249,n180);
or (n2610,n172,n2390);
nand (n2611,n2612,n2617);
or (n2612,n1223,n2613);
not (n2613,n2614);
nor (n2614,n2615,n2616);
and (n2615,n928,n203);
and (n2616,n927,n202);
or (n2617,n2397,n1231);
and (n2618,n2598,n2605);
and (n2619,n2571,n2594);
and (n2620,n2494,n2495);
xor (n2621,n2305,n2308);
and (n2622,n2490,n2491);
xor (n2623,n2302,n2347);
or (n2624,n2625,n2672);
and (n2625,n2626,n2671);
xor (n2626,n2627,n2670);
or (n2627,n2628,n2669);
and (n2628,n2629,n2638);
xor (n2629,n2630,n2631);
xor (n2630,n2310,n2319);
or (n2631,n2632,n2637);
and (n2632,n2633,n2636);
xor (n2633,n2634,n2635);
xor (n2634,n2321,n2336);
xor (n2635,n2404,n2419);
xor (n2636,n2380,n2395);
and (n2637,n2634,n2635);
or (n2638,n2639,n2668);
and (n2639,n2640,n2667);
xor (n2640,n2641,n2666);
or (n2641,n2642,n2665);
and (n2642,n2643,n2658);
xor (n2643,n2644,n2651);
nand (n2644,n2645,n2650);
or (n2645,n2646,n234);
not (n2646,n2647);
nand (n2647,n2648,n2649);
or (n2648,n67,n1470);
or (n2649,n1469,n68);
nand (n2650,n2446,n247);
nand (n2651,n2652,n2657);
or (n2652,n2653,n1138);
not (n2653,n2654);
nand (n2654,n2655,n2656);
or (n2655,n937,n416);
or (n2656,n935,n415);
nand (n2657,n2453,n1154);
nand (n2658,n2659,n2664);
or (n2659,n1424,n2660);
not (n2660,n2661);
nand (n2661,n2662,n2663);
or (n2662,n164,n1146);
or (n2663,n162,n1149);
or (n2664,n2459,n1288);
and (n2665,n2644,n2651);
xor (n2666,n2356,n2371);
xor (n2667,n2442,n2457);
and (n2668,n2641,n2666);
and (n2669,n2630,n2631);
xor (n2670,n2349,n2427);
xor (n2671,n2436,n2468);
and (n2672,n2627,n2670);
and (n2673,n2487,n2623);
xor (n2674,n2299,n2431);
and (n2675,n2483,n2484);
nor (n2676,n2677,n2678);
xor (n2677,n2482,n2674);
or (n2678,n2679,n2696);
and (n2679,n2680,n2695);
xor (n2680,n2681,n2682);
xor (n2681,n2433,n2477);
or (n2682,n2683,n2694);
and (n2683,n2684,n2693);
xor (n2684,n2685,n2692);
or (n2685,n2686,n2691);
and (n2686,n2687,n2690);
xor (n2687,n2688,n2689);
xor (n2688,n2353,n2402);
xor (n2689,n2470,n2473);
xor (n2690,n2439,n2465);
and (n2691,n2688,n2689);
xor (n2692,n2489,n2621);
xor (n2693,n2626,n2671);
and (n2694,n2685,n2692);
xor (n2695,n2486,n2624);
and (n2696,n2681,n2682);
nor (n2697,n2698,n3577);
and (n2698,n2699,n3345);
nor (n2699,n2700,n3341);
and (n2700,n2701,n3239);
nor (n2701,n2702,n3119);
nor (n2702,n2703,n3001);
xor (n2703,n2704,n2988);
xor (n2704,n2705,n2834);
xor (n2705,n2706,n2821);
xor (n2706,n2707,n2820);
or (n2707,n2708,n2819);
and (n2708,n2709,n2818);
xor (n2709,n2710,n2783);
or (n2710,n2711,n2782);
and (n2711,n2712,n2760);
xor (n2712,n2713,n2737);
or (n2713,n2714,n2736);
and (n2714,n2715,n2730);
xor (n2715,n2716,n2723);
nand (n2716,n2717,n2722);
or (n2717,n2718,n199);
not (n2718,n2719);
nand (n2719,n2720,n2721);
or (n2720,n28,n1162);
nand (n2721,n28,n1162);
nand (n2722,n2534,n1118);
nand (n2723,n2724,n2729);
or (n2724,n2725,n103);
not (n2725,n2726);
nor (n2726,n2727,n2728);
and (n2727,n177,n1124);
and (n2728,n1125,n107);
nand (n2729,n2527,n96);
nand (n2730,n2731,n2732);
or (n2731,n1288,n2660);
or (n2732,n2733,n1424);
nor (n2733,n2734,n2735);
and (n2734,n156,n1149);
and (n2735,n1146,n158);
and (n2736,n2716,n2723);
or (n2737,n2738,n2759);
and (n2738,n2739,n2753);
xor (n2739,n2740,n2747);
nand (n2740,n2741,n2746);
or (n2741,n2742,n420);
not (n2742,n2743);
nor (n2743,n2744,n2745);
and (n2744,n409,n1399);
and (n2745,n1210,n407);
nand (n2746,n2557,n413);
nand (n2747,n2748,n2752);
or (n2748,n171,n2749);
nor (n2749,n2750,n2751);
and (n2750,n180,n1705);
and (n2751,n195,n1244);
or (n2752,n2607,n172);
nand (n2753,n2754,n2755);
or (n2754,n1144,n2653);
or (n2755,n1138,n2756);
nor (n2756,n2757,n2758);
and (n2757,n415,n1344);
and (n2758,n416,n1576);
and (n2759,n2740,n2747);
or (n2760,n2761,n2781);
and (n2761,n2762,n2775);
xor (n2762,n2763,n2769);
nand (n2763,n2764,n2768);
or (n2764,n400,n2765);
nor (n2765,n2766,n2767);
and (n2766,n1323,n395);
and (n2767,n1325,n396);
or (n2768,n2539,n529);
nand (n2769,n2770,n2774);
or (n2770,n2771,n1173);
nor (n2771,n2772,n2773);
and (n2772,n1175,n1659);
and (n2773,n1181,n114);
or (n2774,n2516,n1176);
nand (n2775,n2776,n2780);
or (n2776,n2777,n1194);
nor (n2777,n2778,n2779);
and (n2778,n215,n1191);
and (n2779,n217,n1192);
or (n2780,n2549,n1196);
and (n2781,n2763,n2769);
and (n2782,n2713,n2737);
or (n2783,n2784,n2817);
and (n2784,n2785,n2794);
xor (n2785,n2786,n2793);
or (n2786,n2787,n2792);
and (n2787,n2788,n2791);
xor (n2788,n2789,n2790);
and (n2789,n317,n1377);
and (n2790,n566,n1463);
and (n2791,n247,n1470);
and (n2792,n2789,n2790);
xor (n2793,n2573,n2586);
or (n2794,n2795,n2816);
and (n2795,n2796,n2810);
xor (n2796,n2797,n2804);
nand (n2797,n2798,n2803);
or (n2798,n2799,n1223);
not (n2799,n2800);
nor (n2800,n2801,n2802);
and (n2801,n1357,n203);
and (n2802,n1356,n202);
nand (n2803,n2614,n1238);
nand (n2804,n2805,n2806);
or (n2805,n1597,n2600);
nand (n2806,n1591,n2807);
nor (n2807,n2808,n2809);
and (n2808,n1304,n1588);
and (n2809,n1305,n100);
nand (n2810,n2811,n2812);
or (n2811,n2503,n23);
or (n2812,n22,n2813);
nor (n2813,n2814,n2815);
and (n2814,n1475,n32);
and (n2815,n1477,n33);
and (n2816,n2797,n2804);
and (n2817,n2786,n2793);
xor (n2818,n2570,n2595);
and (n2819,n2710,n2783);
xor (n2820,n2493,n2568);
or (n2821,n2822,n2833);
and (n2822,n2823,n2832);
xor (n2823,n2824,n2831);
or (n2824,n2825,n2830);
and (n2825,n2826,n2829);
xor (n2826,n2827,n2828);
xor (n2827,n2643,n2658);
xor (n2828,n2500,n2514);
xor (n2829,n2523,n2537);
and (n2830,n2827,n2828);
xor (n2831,n2497,n2544);
xor (n2832,n2640,n2667);
and (n2833,n2824,n2831);
or (n2834,n2835,n2987);
and (n2835,n2836,n2894);
xor (n2836,n2837,n2893);
or (n2837,n2838,n2892);
and (n2838,n2839,n2891);
xor (n2839,n2840,n2841);
xor (n2840,n2785,n2794);
or (n2841,n2842,n2890);
and (n2842,n2843,n2867);
xor (n2843,n2844,n2866);
or (n2844,n2845,n2865);
and (n2845,n2846,n2858);
xor (n2846,n2847,n2853);
and (n2847,n2848,n180);
nand (n2848,n2849,n2852);
nand (n2849,n2850,n177);
not (n2850,n2851);
and (n2851,n1377,n175);
nand (n2852,n1379,n174);
and (n2853,n2854,n396);
nand (n2854,n2855,n2856);
or (n2855,n1463,n404);
nand (n2856,n2857,n409);
nand (n2857,n1463,n404);
nor (n2858,n2859,n32);
and (n2859,n2860,n2863);
not (n2860,n2861);
nor (n2861,n2862,n28);
and (n2862,n1470,n27);
not (n2863,n2864);
nor (n2864,n1470,n27);
and (n2865,n2847,n2853);
xor (n2866,n2788,n2791);
or (n2867,n2868,n2889);
and (n2868,n2869,n2883);
xor (n2869,n2870,n2877);
nand (n2870,n2871,n2876);
or (n2871,n2872,n420);
not (n2872,n2873);
nor (n2873,n2874,n2875);
and (n2874,n1317,n407);
and (n2875,n1316,n409);
nand (n2876,n2743,n413);
nand (n2877,n2878,n2882);
or (n2878,n22,n2879);
nor (n2879,n2880,n2881);
and (n2880,n1469,n33);
and (n2881,n32,n1470);
or (n2882,n23,n2813);
nand (n2883,n2884,n2888);
or (n2884,n2885,n1194);
nor (n2885,n2886,n2887);
and (n2886,n956,n1191);
and (n2887,n955,n1192);
or (n2888,n2777,n1196);
and (n2889,n2870,n2877);
and (n2890,n2844,n2866);
xor (n2891,n2712,n2760);
and (n2892,n2840,n2841);
xor (n2893,n2823,n2832);
or (n2894,n2895,n2986);
and (n2895,n2896,n2905);
xor (n2896,n2897,n2904);
or (n2897,n2898,n2903);
and (n2898,n2899,n2902);
xor (n2899,n2900,n2901);
xor (n2900,n2796,n2810);
xor (n2901,n2762,n2775);
xor (n2902,n2715,n2730);
and (n2903,n2900,n2901);
xor (n2904,n2826,n2829);
xor (n2905,n2906,n2909);
xor (n2906,n2907,n2908);
xor (n2907,n2546,n2560);
xor (n2908,n2597,n2611);
or (n2909,n2910,n2985);
and (n2910,n2911,n2963);
xor (n2911,n2912,n2937);
or (n2912,n2913,n2936);
and (n2913,n2914,n2929);
xor (n2914,n2915,n2922);
nand (n2915,n2916,n2921);
or (n2916,n2917,n199);
not (n2917,n2918);
nor (n2918,n2919,n2920);
and (n2919,n1639,n28);
and (n2920,n1641,n209);
nand (n2921,n1118,n2719);
nand (n2922,n2923,n2928);
or (n2923,n103,n2924);
not (n2924,n2925);
nand (n2925,n2926,n2927);
or (n2926,n1250,n177);
nand (n2927,n1250,n177);
or (n2928,n104,n2725);
nand (n2929,n2930,n2935);
or (n2930,n2931,n1424);
not (n2931,n2932);
nor (n2932,n2933,n2934);
and (n2933,n1149,n937);
and (n2934,n935,n1146);
or (n2935,n2733,n1288);
and (n2936,n2915,n2922);
or (n2937,n2938,n2962);
and (n2938,n2939,n2954);
xor (n2939,n2940,n2947);
nand (n2940,n2941,n2946);
or (n2941,n2942,n1223);
not (n2942,n2943);
nor (n2943,n2944,n2945);
and (n2944,n202,n1168);
and (n2945,n1169,n203);
nand (n2946,n2800,n1238);
nand (n2947,n2948,n2953);
or (n2948,n2949,n171);
not (n2949,n2950);
nand (n2950,n2951,n2952);
or (n2951,n1377,n195);
or (n2952,n1379,n180);
or (n2953,n172,n2749);
nand (n2954,n2955,n2960);
or (n2955,n1590,n2956);
not (n2956,n2957);
nor (n2957,n2958,n2959);
and (n2958,n1130,n1588);
and (n2959,n1131,n100);
or (n2960,n2961,n1597);
not (n2961,n2807);
and (n2962,n2940,n2947);
or (n2963,n2964,n2984);
and (n2964,n2965,n2978);
xor (n2965,n2966,n2972);
nand (n2966,n2967,n2971);
or (n2967,n400,n2968);
nor (n2968,n2969,n2970);
and (n2969,n1462,n396);
and (n2970,n395,n1463);
or (n2971,n2765,n529);
nand (n2972,n2973,n2977);
or (n2973,n2974,n1173);
nor (n2974,n2975,n2976);
and (n2975,n1181,n928);
and (n2976,n1175,n927);
or (n2977,n2771,n1176);
nand (n2978,n2979,n2983);
or (n2979,n1138,n2980);
nor (n2980,n2981,n2982);
and (n2981,n415,n1215);
and (n2982,n416,n2090);
or (n2983,n2756,n1144);
and (n2984,n2966,n2972);
and (n2985,n2912,n2937);
and (n2986,n2897,n2904);
and (n2987,n2837,n2893);
xor (n2988,n2989,n2992);
xor (n2989,n2990,n2991);
xor (n2990,n2629,n2638);
xor (n2991,n2687,n2690);
or (n2992,n2993,n3000);
and (n2993,n2994,n2999);
xor (n2994,n2995,n2996);
xor (n2995,n2633,n2636);
or (n2996,n2997,n2998);
and (n2997,n2906,n2909);
and (n2998,n2907,n2908);
xor (n2999,n2709,n2818);
and (n3000,n2995,n2996);
or (n3001,n3002,n3118);
and (n3002,n3003,n3117);
xor (n3003,n3004,n3005);
xor (n3004,n2994,n2999);
or (n3005,n3006,n3116);
and (n3006,n3007,n3115);
xor (n3007,n3008,n3050);
or (n3008,n3009,n3049);
and (n3009,n3010,n3013);
xor (n3010,n3011,n3012);
xor (n3011,n2739,n2753);
xor (n3012,n2843,n2867);
or (n3013,n3014,n3048);
and (n3014,n3015,n3024);
xor (n3015,n3016,n3023);
or (n3016,n3017,n3022);
and (n3017,n3018,n3021);
xor (n3018,n3019,n3020);
and (n3019,n189,n1377);
and (n3020,n405,n1463);
nor (n3021,n23,n1469);
and (n3022,n3019,n3020);
xor (n3023,n2846,n2858);
or (n3024,n3025,n3047);
and (n3025,n3026,n3041);
xor (n3026,n3027,n3034);
nand (n3027,n3028,n3033);
or (n3028,n1424,n3029);
not (n3029,n3030);
nand (n3030,n3031,n3032);
or (n3031,n1344,n1149);
nand (n3032,n1344,n1149);
nand (n3033,n2932,n1289);
nand (n3034,n3035,n3040);
or (n3035,n3036,n420);
not (n3036,n3037);
nor (n3037,n3038,n3039);
and (n3038,n1323,n407);
and (n3039,n1325,n409);
nand (n3040,n2873,n413);
nand (n3041,n3042,n3046);
or (n3042,n3043,n1173);
nor (n3043,n3044,n3045);
and (n3044,n1181,n1357);
and (n3045,n1175,n1356);
or (n3046,n2974,n1176);
and (n3047,n3027,n3034);
and (n3048,n3016,n3023);
and (n3049,n3011,n3012);
or (n3050,n3051,n3114);
and (n3051,n3052,n3107);
xor (n3052,n3053,n3054);
xor (n3053,n2911,n2963);
or (n3054,n3055,n3106);
and (n3055,n3056,n3105);
xor (n3056,n3057,n3081);
or (n3057,n3058,n3080);
and (n3058,n3059,n3074);
xor (n3059,n3060,n3067);
nand (n3060,n3061,n3066);
or (n3061,n3062,n103);
not (n3062,n3063);
nand (n3063,n3064,n3065);
or (n3064,n1244,n177);
nand (n3065,n177,n1244);
nand (n3066,n96,n2925);
nand (n3067,n3068,n3073);
or (n3068,n3069,n1590);
not (n3069,n3070);
nand (n3070,n3071,n3072);
or (n3071,n1125,n1588);
nand (n3072,n1588,n1125);
nand (n3073,n1601,n2957);
nand (n3074,n3075,n3079);
or (n3075,n1138,n3076);
nor (n3076,n3077,n3078);
and (n3077,n415,n1210);
and (n3078,n1399,n416);
or (n3079,n2980,n1144);
and (n3080,n3060,n3067);
or (n3081,n3082,n3104);
and (n3082,n3083,n3098);
xor (n3083,n3084,n3091);
nand (n3084,n3085,n3090);
or (n3085,n3086,n1223);
not (n3086,n3087);
nor (n3087,n3088,n3089);
and (n3088,n202,n1162);
and (n3089,n1163,n203);
nand (n3090,n1238,n2943);
nand (n3091,n3092,n3097);
or (n3092,n3093,n1194);
not (n3093,n3094);
nand (n3094,n3095,n3096);
or (n3095,n1191,n1305);
nand (n3096,n1305,n1191);
or (n3097,n2885,n1196);
nand (n3098,n3099,n3103);
or (n3099,n199,n3100);
nor (n3100,n3101,n3102);
and (n3101,n209,n1475);
and (n3102,n28,n1477);
or (n3103,n200,n2917);
and (n3104,n3084,n3091);
xor (n3105,n2939,n2954);
and (n3106,n3057,n3081);
or (n3107,n3108,n3113);
and (n3108,n3109,n3112);
xor (n3109,n3110,n3111);
xor (n3110,n2914,n2929);
xor (n3111,n2965,n2978);
xor (n3112,n2869,n2883);
and (n3113,n3110,n3111);
and (n3114,n3053,n3054);
xor (n3115,n2839,n2891);
and (n3116,n3008,n3050);
xor (n3117,n2836,n2894);
and (n3118,n3004,n3005);
nor (n3119,n3120,n3121);
xor (n3120,n3003,n3117);
or (n3121,n3122,n3238);
and (n3122,n3123,n3237);
xor (n3123,n3124,n3125);
xor (n3124,n2896,n2905);
or (n3125,n3126,n3236);
and (n3126,n3127,n3235);
xor (n3127,n3128,n3129);
xor (n3128,n2899,n2902);
or (n3129,n3130,n3234);
and (n3130,n3131,n3183);
xor (n3131,n3132,n3182);
or (n3132,n3133,n3181);
and (n3133,n3134,n3157);
xor (n3134,n3135,n3156);
or (n3135,n3136,n3155);
and (n3136,n3137,n3150);
xor (n3137,n3138,n3143);
nor (n3138,n3139,n177);
nor (n3139,n3140,n3142);
and (n3140,n3141,n1588);
nand (n3141,n1377,n99);
nor (n3142,n1377,n99);
nor (n3143,n3144,n409);
and (n3144,n3145,n3148);
not (n3145,n3146);
nor (n3146,n3147,n416);
and (n3147,n1463,n417);
not (n3148,n3149);
nor (n3149,n1463,n417);
nor (n3150,n3151,n209);
nor (n3151,n3152,n3154);
and (n3152,n3153,n202);
nand (n3153,n1470,n204);
and (n3154,n1469,n206);
and (n3155,n3138,n3143);
xor (n3156,n3018,n3021);
or (n3157,n3158,n3180);
and (n3158,n3159,n3174);
xor (n3159,n3160,n3167);
nand (n3160,n3161,n3166);
or (n3161,n3162,n1223);
not (n3162,n3163);
nand (n3163,n3164,n3165);
or (n3164,n1639,n202);
nand (n3165,n1639,n202);
nand (n3166,n3087,n1238);
nand (n3167,n3168,n3173);
or (n3168,n1194,n3169);
not (n3169,n3170);
nor (n3170,n3171,n3172);
and (n3171,n1191,n1130);
and (n3172,n1131,n1192);
nand (n3173,n3094,n1197);
nand (n3174,n3175,n3179);
or (n3175,n199,n3176);
nor (n3176,n3177,n3178);
and (n3177,n1469,n28);
and (n3178,n209,n1470);
or (n3179,n3100,n200);
and (n3180,n3160,n3167);
and (n3181,n3135,n3156);
xor (n3182,n3015,n3024);
or (n3183,n3184,n3233);
and (n3184,n3185,n3232);
xor (n3185,n3186,n3209);
or (n3186,n3187,n3208);
and (n3187,n3188,n3202);
xor (n3188,n3189,n3196);
nand (n3189,n3190,n3195);
or (n3190,n3191,n103);
not (n3191,n3192);
nand (n3192,n3193,n3194);
or (n3193,n177,n1377);
or (n3194,n1379,n107);
nand (n3195,n96,n3063);
nand (n3196,n3197,n3201);
or (n3197,n1590,n3198);
nor (n3198,n3199,n3200);
and (n3199,n1250,n1588);
and (n3200,n1249,n100);
nand (n3201,n1601,n3070);
nand (n3202,n3203,n3207);
or (n3203,n1138,n3204);
nor (n3204,n3205,n3206);
and (n3205,n415,n1317);
and (n3206,n416,n1316);
or (n3207,n3076,n1144);
and (n3208,n3189,n3196);
or (n3209,n3210,n3231);
and (n3210,n3211,n3225);
xor (n3211,n3212,n3218);
nand (n3212,n3213,n3217);
or (n3213,n3214,n1424);
nor (n3214,n3215,n3216);
and (n3215,n1149,n1215);
and (n3216,n1146,n2090);
or (n3217,n3029,n1288);
nand (n3218,n3219,n3224);
or (n3219,n3220,n420);
not (n3220,n3221);
nand (n3221,n3222,n3223);
or (n3222,n409,n1463);
or (n3223,n1462,n407);
nand (n3224,n3037,n413);
nand (n3225,n3226,n3230);
or (n3226,n3227,n1173);
nor (n3227,n3228,n3229);
and (n3228,n1169,n1181);
and (n3229,n1168,n1175);
or (n3230,n3043,n1176);
and (n3231,n3212,n3218);
xor (n3232,n3083,n3098);
and (n3233,n3186,n3209);
and (n3234,n3132,n3182);
xor (n3235,n3010,n3013);
and (n3236,n3128,n3129);
xor (n3237,n3007,n3115);
and (n3238,n3124,n3125);
nand (n3239,n3240,n3340);
or (n3240,n3241,n3296);
nor (n3241,n3242,n3243);
xor (n3242,n3123,n3237);
or (n3243,n3244,n3295);
and (n3244,n3245,n3294);
xor (n3245,n3246,n3247);
xor (n3246,n3052,n3107);
or (n3247,n3248,n3293);
and (n3248,n3249,n3252);
xor (n3249,n3250,n3251);
xor (n3250,n3056,n3105);
xor (n3251,n3109,n3112);
or (n3252,n3253,n3292);
and (n3253,n3254,n3257);
xor (n3254,n3255,n3256);
xor (n3255,n3026,n3041);
xor (n3256,n3059,n3074);
or (n3257,n3258,n3291);
and (n3258,n3259,n3268);
xor (n3259,n3260,n3267);
or (n3260,n3261,n3266);
and (n3261,n3262,n3265);
xor (n3262,n3263,n3264);
and (n3263,n96,n1377);
and (n3264,n1118,n1470);
nor (n3265,n424,n1462);
and (n3266,n3263,n3264);
xor (n3267,n3137,n3150);
or (n3268,n3269,n3290);
and (n3269,n3270,n3284);
xor (n3270,n3271,n3278);
nand (n3271,n3272,n3277);
or (n3272,n3273,n1173);
not (n3273,n3274);
nor (n3274,n3275,n3276);
and (n3275,n1163,n1175);
and (n3276,n1181,n1162);
or (n3277,n3227,n1176);
nand (n3278,n3279,n3283);
or (n3279,n1138,n3280);
nor (n3280,n3281,n3282);
and (n3281,n415,n1323);
and (n3282,n1325,n416);
or (n3283,n3204,n1144);
nand (n3284,n3285,n3289);
or (n3285,n1590,n3286);
nor (n3286,n3287,n3288);
and (n3287,n1588,n1244);
and (n3288,n100,n1705);
or (n3289,n1597,n3198);
and (n3290,n3271,n3278);
and (n3291,n3260,n3267);
and (n3292,n3255,n3256);
and (n3293,n3250,n3251);
xor (n3294,n3127,n3235);
and (n3295,n3246,n3247);
nand (n3296,n3297,n3298);
xor (n3297,n3245,n3294);
or (n3298,n3299,n3339);
and (n3299,n3300,n3338);
xor (n3300,n3301,n3302);
xor (n3301,n3131,n3183);
or (n3302,n3303,n3337);
and (n3303,n3304,n3336);
xor (n3304,n3305,n3306);
xor (n3305,n3134,n3157);
or (n3306,n3307,n3335);
and (n3307,n3308,n3334);
xor (n3308,n3309,n3333);
or (n3309,n3310,n3332);
and (n3310,n3311,n3325);
xor (n3311,n3312,n3319);
nand (n3312,n3313,n3318);
or (n3313,n3314,n1223);
not (n3314,n3315);
nor (n3315,n3316,n3317);
and (n3316,n1475,n203);
and (n3317,n1477,n202);
nand (n3318,n3163,n1238);
nand (n3319,n3320,n3324);
or (n3320,n3321,n1424);
nor (n3321,n3322,n3323);
and (n3322,n1149,n1210);
and (n3323,n1399,n1146);
or (n3324,n3214,n1288);
nand (n3325,n3326,n3331);
or (n3326,n1194,n3327);
not (n3327,n3328);
nor (n3328,n3329,n3330);
and (n3329,n1125,n1192);
and (n3330,n1124,n1191);
or (n3331,n3169,n1196);
and (n3332,n3312,n3319);
xor (n3333,n3159,n3174);
xor (n3334,n3211,n3225);
and (n3335,n3309,n3333);
xor (n3336,n3185,n3232);
and (n3337,n3305,n3306);
xor (n3338,n3249,n3252);
and (n3339,n3301,n3302);
nand (n3340,n3242,n3243);
nor (n3341,n3342,n2702);
and (n3342,n3343,n3344);
nand (n3343,n2703,n3001);
nand (n3344,n3120,n3121);
nand (n3345,n2701,n3346);
nor (n3346,n3347,n3350);
nand (n3347,n3348,n3349);
or (n3348,n3298,n3297);
not (n3349,n3241);
nor (n3350,n3351,n3540,n3571);
and (n3351,n3352,n3456);
not (n3352,n3353);
nand (n3353,n3354,n3449);
or (n3354,n3355,n3442);
or (n3355,n3356,n3441);
and (n3356,n3357,n3389);
xor (n3357,n3358,n3388);
or (n3358,n3359,n3387);
and (n3359,n3360,n3386);
xor (n3360,n3361,n3385);
or (n3361,n3362,n3384);
and (n3362,n3363,n3377);
xor (n3363,n3364,n3371);
nand (n3364,n3365,n3370);
or (n3365,n1173,n3366);
not (n3366,n3367);
nor (n3367,n3368,n3369);
and (n3368,n1639,n1175);
and (n3369,n1641,n1181);
nand (n3370,n3274,n1177);
nand (n3371,n3372,n3373);
or (n3372,n1196,n3327);
nand (n3373,n3374,n1195);
nand (n3374,n3375,n3376);
or (n3375,n1250,n1191);
nand (n3376,n1191,n1250);
nand (n3377,n3378,n3383);
or (n3378,n3379,n1138);
not (n3379,n3380);
nand (n3380,n3381,n3382);
or (n3381,n415,n1463);
or (n3382,n1462,n416);
or (n3383,n3280,n1144);
and (n3384,n3364,n3371);
xor (n3385,n3311,n3325);
xor (n3386,n3270,n3284);
and (n3387,n3361,n3385);
xor (n3388,n3308,n3334);
xor (n3389,n3390,n3440);
xor (n3390,n3391,n3392);
xor (n3391,n3188,n3202);
or (n3392,n3393,n3439);
and (n3393,n3394,n3416);
xor (n3394,n3395,n3415);
or (n3395,n3396,n3414);
and (n3396,n3397,n3409);
xor (n3397,n3398,n3403);
nor (n3398,n3399,n1588);
nor (n3399,n3400,n3401);
and (n3400,n1379,n1594);
and (n3401,n3402,n1191);
nand (n3402,n1377,n1595);
and (n3403,n3404,n203);
nand (n3404,n3405,n3406);
or (n3405,n1470,n1227);
nand (n3406,n3407,n1181);
not (n3407,n3408);
and (n3408,n1470,n1227);
nor (n3409,n3410,n415);
nor (n3410,n3411,n3413);
and (n3411,n3412,n1149);
nand (n3412,n1463,n1142);
and (n3413,n1462,n1147);
and (n3414,n3398,n3403);
xor (n3415,n3262,n3265);
or (n3416,n3417,n3438);
and (n3417,n3418,n3432);
xor (n3418,n3419,n3425);
nand (n3419,n3420,n3424);
or (n3420,n1223,n3421);
nor (n3421,n3422,n3423);
and (n3422,n1469,n203);
and (n3423,n1470,n202);
or (n3424,n1231,n3314);
nand (n3425,n3426,n3431);
or (n3426,n1424,n3427);
not (n3427,n3428);
nor (n3428,n3429,n3430);
and (n3429,n1149,n1316);
and (n3430,n1317,n1146);
or (n3431,n3321,n1288);
nand (n3432,n3433,n3437);
or (n3433,n1590,n3434);
nor (n3434,n3435,n3436);
and (n3435,n1379,n100);
and (n3436,n1377,n1588);
or (n3437,n1597,n3286);
and (n3438,n3419,n3425);
and (n3439,n3395,n3415);
xor (n3440,n3259,n3268);
and (n3441,n3358,n3388);
xor (n3442,n3443,n3448);
xor (n3443,n3444,n3447);
or (n3444,n3445,n3446);
and (n3445,n3390,n3440);
and (n3446,n3391,n3392);
xor (n3447,n3254,n3257);
xor (n3448,n3304,n3336);
nand (n3449,n3450,n3452);
not (n3450,n3451);
xor (n3451,n3300,n3338);
not (n3452,n3453);
or (n3453,n3454,n3455);
and (n3454,n3443,n3448);
and (n3455,n3444,n3447);
nand (n3456,n3457,n3537);
or (n3457,n3458,n3501);
nor (n3458,n3459,n3500);
or (n3459,n3460,n3499);
and (n3460,n3461,n3498);
xor (n3461,n3462,n3497);
or (n3462,n3463,n3496);
and (n3463,n3464,n3473);
xor (n3464,n3465,n3472);
or (n3465,n3466,n3471);
and (n3466,n3467,n3470);
xor (n3467,n3468,n3469);
and (n3468,n1601,n1377);
and (n3469,n1154,n1463);
nor (n3470,n1231,n1469);
and (n3471,n3468,n3469);
xor (n3472,n3397,n3409);
or (n3473,n3474,n3495);
and (n3474,n3475,n3489);
xor (n3475,n3476,n3483);
nand (n3476,n3477,n3481);
or (n3477,n3478,n1194);
nor (n3478,n3479,n3480);
and (n3479,n1191,n1244);
and (n3480,n1192,n1705);
or (n3481,n3482,n1196);
not (n3482,n3374);
nand (n3483,n3484,n3485);
or (n3484,n1176,n3366);
or (n3485,n3486,n1173);
nor (n3486,n3487,n3488);
and (n3487,n1181,n1475);
and (n3488,n1477,n1175);
nand (n3489,n3490,n3491);
or (n3490,n1288,n3427);
or (n3491,n3492,n1424);
nor (n3492,n3493,n3494);
and (n3493,n1146,n1325);
and (n3494,n1149,n1323);
and (n3495,n3476,n3483);
and (n3496,n3465,n3472);
xor (n3497,n3394,n3416);
xor (n3498,n3360,n3386);
and (n3499,n3462,n3497);
xor (n3500,n3357,n3389);
nand (n3501,n3502,n3536);
or (n3502,n3503,n3535);
and (n3503,n3504,n3507);
xor (n3504,n3505,n3506);
xor (n3505,n3363,n3377);
xor (n3506,n3418,n3432);
or (n3507,n3508,n3534);
and (n3508,n3509,n3521);
xor (n3509,n3510,n3520);
or (n3510,n3511,n3519);
and (n3511,n3512,n3517);
xor (n3512,n3513,n3515);
and (n3513,n3514,n1192);
nand (n3514,n1377,n1197);
nor (n3515,n3516,n1149);
and (n3516,n1463,n1289);
nor (n3517,n3518,n1181);
and (n3518,n1470,n1177);
and (n3519,n3513,n3515);
xor (n3520,n3467,n3470);
or (n3521,n3522,n3533);
and (n3522,n3523,n3530);
xor (n3523,n3524,n3527);
nand (n3524,n3525,n3526);
or (n3525,n3478,n1196);
or (n3526,n1194,n1377);
nand (n3527,n3528,n3529);
or (n3528,n3492,n1288);
or (n3529,n1424,n1463);
nand (n3530,n3531,n3532);
or (n3531,n1470,n1173);
or (n3532,n3486,n1176);
and (n3533,n3524,n3527);
and (n3534,n3510,n3520);
and (n3535,n3505,n3506);
xor (n3536,n3461,n3498);
or (n3537,n3538,n3539);
not (n3538,n3500);
not (n3539,n3459);
nor (n3540,n3353,n3541);
nand (n3541,n3542,n3543);
not (n3542,n3458);
nor (n3543,n3544,n3568);
and (n3544,n3545,n3553);
nor (n3545,n3546,n3552);
and (n3546,n3547,n3550,n3551);
or (n3547,n3548,n3549);
xor (n3548,n3504,n3507);
xor (n3549,n3464,n3473);
xor (n3550,n3509,n3521);
xor (n3551,n3475,n3489);
and (n3552,n3548,n3549);
nand (n3553,n3547,n3554);
nor (n3554,n3555,n3560,n3561);
and (n3555,n3556,n3558);
not (n3556,n3557);
xor (n3557,n3523,n3530);
not (n3558,n3559);
xor (n3559,n3512,n3517);
nor (n3560,n3550,n3551);
nor (n3561,n3562,n3563,n3564);
and (n3562,n3516,n3518);
nor (n3563,n3556,n3558);
nor (n3564,n3565,n3514);
and (n3565,n3566,n3567);
not (n3566,n3518);
not (n3567,n3516);
and (n3568,n3569,n3570);
not (n3569,n3536);
not (n3570,n3502);
nand (n3571,n3572,n3576);
or (n3572,n3573,n3574,n3575);
not (n3573,n3449);
not (n3574,n3442);
not (n3575,n3355);
nand (n3576,n3451,n3453);
nand (n3577,n3578,n3591);
or (n3578,n3579,n3582);
or (n3579,n3580,n3581);
and (n3580,n2704,n2988);
and (n3581,n2705,n2834);
xor (n3582,n3583,n3590);
xor (n3583,n3584,n3587);
or (n3584,n3585,n3586);
and (n3585,n2706,n2821);
and (n3586,n2707,n2820);
or (n3587,n3588,n3589);
and (n3588,n2989,n2992);
and (n3589,n2990,n2991);
xor (n3590,n2684,n2693);
nand (n3591,n3592,n3594);
not (n3592,n3593);
xor (n3593,n2680,n2695);
not (n3594,n3595);
or (n3595,n3596,n3597);
and (n3596,n3583,n3590);
and (n3597,n3584,n3587);
nand (n3598,n1095,n3599);
nand (n3599,n3600,n3601);
or (n3600,n3594,n3592);
or (n3601,n3602,n3603);
not (n3602,n3591);
nand (n3603,n3582,n3579);
nand (n3604,n3605,n3606);
not (n3605,n1096);
nand (n3606,n3607,n3610);
or (n3607,n3608,n3609);
not (n3608,n2480);
not (n3609,n1097);
nand (n3610,n2677,n2678);
nor (n3611,n3612,n4140);
nor (n3612,n3613,n4131);
xor (n3613,n3614,n3883);
xor (n3614,n3615,n3874);
xor (n3615,n3616,n3803);
xor (n3616,n3617,n3758);
or (n3617,n3618,n3757);
and (n3618,n3619,n3754);
xor (n3619,n3620,n3688);
xor (n3620,n3621,n3664);
xor (n3621,n3622,n3640);
xor (n3622,n3623,n3634);
xor (n3623,n3624,n3627);
nand (n3624,n3625,n3626);
or (n3625,n1424,n1831);
nand (n3626,n1146,n1289);
nand (n3627,n3628,n3630);
or (n3628,n3629,n281);
not (n3629,n1759);
nand (n3630,n3631,n288);
nand (n3631,n3632,n3633);
or (n3632,n956,n265);
nand (n3633,n956,n265);
nand (n3634,n3635,n3636);
or (n3635,n1691,n420);
nand (n3636,n3637,n413);
nor (n3637,n3638,n3639);
and (n3638,n452,n409);
and (n3639,n453,n407);
xor (n3640,n3641,n3656);
xor (n3641,n3642,n3649);
nand (n3642,n3643,n3645);
or (n3643,n3644,n1223);
not (n3644,n1726);
nand (n3645,n3646,n1238);
nand (n3646,n3647,n3648);
or (n3647,n85,n202);
nand (n3648,n202,n85);
nand (n3649,n3650,n3652);
or (n3650,n3651,n37);
not (n3651,n1703);
nand (n3652,n46,n3653);
nand (n3653,n3654,n3655);
or (n3654,n1250,n41);
nand (n3655,n41,n1250);
nand (n3656,n3657,n3659);
or (n3657,n103,n3658);
not (n3658,n1789);
or (n3659,n3660,n104);
not (n3660,n3661);
nand (n3661,n3662,n3663);
or (n3662,n297,n177);
nand (n3663,n297,n177);
xor (n3664,n3665,n3680);
xor (n3665,n3666,n3673);
nand (n3666,n3667,n3669);
or (n3667,n3668,n199);
not (n3668,n1825);
nand (n3669,n1118,n3670);
nand (n3670,n3671,n3672);
or (n3671,n28,n491);
nand (n3672,n491,n28);
nand (n3673,n3674,n3676);
or (n3674,n400,n3675);
not (n3675,n1847);
nand (n3676,n3677,n405);
nand (n3677,n3678,n3679);
or (n3678,n396,n388);
nand (n3679,n388,n396);
nand (n3680,n3681,n3683);
or (n3681,n64,n3682);
not (n3682,n1781);
or (n3683,n65,n3684);
not (n3684,n3685);
nor (n3685,n3686,n3687);
and (n3686,n927,n74);
and (n3687,n928,n75);
xor (n3688,n3689,n3733);
xor (n3689,n3690,n3712);
xor (n3690,n3691,n3706);
xor (n3691,n3692,n3699);
nand (n3692,n3693,n3695);
or (n3693,n3694,n1590);
not (n3694,n1672);
nand (n3695,n3696,n1601);
nand (n3696,n3697,n3698);
or (n3697,n100,n327);
nand (n3698,n327,n100);
nand (n3699,n3700,n3702);
or (n3700,n3701,n470);
not (n3701,n1684);
nand (n3702,n3703,n566);
nor (n3703,n3704,n3705);
and (n3704,n440,n164);
and (n3705,n441,n162);
nand (n3706,n3707,n3708);
or (n3707,n1813,n138);
nand (n3708,n3709,n148);
nor (n3709,n3710,n3711);
and (n3710,n147,n1316);
and (n3711,n144,n1317);
xor (n3712,n3713,n3727);
xor (n3713,n3714,n3721);
nand (n3714,n3715,n3717);
or (n3715,n3716,n532);
not (n3716,n1719);
nand (n3717,n3718,n333);
nand (n3718,n3719,n3720);
or (n3719,n1169,n127);
nand (n3720,n127,n1169);
nand (n3721,n3722,n3723);
or (n3722,n1732,n255);
nand (n3723,n3724,n272);
nand (n3724,n3725,n3726);
or (n3725,n1131,n253);
nand (n3726,n253,n1131);
nand (n3727,n3728,n3729);
or (n3728,n1852,n22);
nand (n3729,n3730,n24);
nor (n3730,n3731,n3732);
and (n3731,n33,n341);
and (n3732,n32,n340);
xor (n3733,n3734,n3748);
xor (n3734,n3735,n3742);
nand (n3735,n3736,n3738);
or (n3736,n3737,n436);
not (n3737,n1678);
nand (n3738,n449,n3739);
nand (n3739,n3740,n3741);
or (n3740,n935,n382);
nand (n3741,n382,n935);
nand (n3742,n3743,n3744);
or (n3743,n1794,n1138);
nand (n3744,n3745,n1154);
nand (n3745,n3746,n3747);
or (n3746,n416,n465);
nand (n3747,n465,n416);
nand (n3748,n3749,n3750);
or (n3749,n234,n1802);
or (n3750,n235,n3751);
nor (n3751,n3752,n3753);
and (n3752,n134,n67);
and (n3753,n133,n68);
or (n3754,n3755,n3756);
and (n3755,n1808,n1857);
and (n3756,n1809,n1835);
and (n3757,n3620,n3688);
or (n3758,n3759,n3802);
and (n3759,n3760,n3767);
xor (n3760,n3761,n3764);
or (n3761,n3762,n3763);
and (n3762,n2255,n2262);
and (n3763,n2256,n2259);
or (n3764,n3765,n3766);
and (n3765,n2266,n2273);
and (n3766,n2267,n2270);
xor (n3767,n3768,n3799);
xor (n3768,n3769,n3796);
xor (n3769,n3770,n3780);
xor (n3770,n3771,n3777);
nand (n3771,n3772,n3773);
or (n3772,n171,n1711);
or (n3773,n172,n3774);
nor (n3774,n3775,n3776);
and (n3775,n195,n59);
and (n3776,n180,n61);
or (n3777,n3778,n3779);
and (n3778,n1867,n1878);
and (n3779,n1868,n1873);
xor (n3780,n3781,n3789);
nand (n3781,n3782,n3787);
or (n3782,n1196,n3783);
not (n3783,n3784);
nor (n3784,n3785,n3786);
and (n3785,n1191,n192);
and (n3786,n1192,n193);
or (n3787,n3788,n1194);
not (n3788,n1773);
nand (n3789,n3790,n3792);
or (n3790,n118,n3791);
not (n3791,n1752);
or (n3792,n3793,n664);
nor (n3793,n3794,n3795);
and (n3794,n115,n1639);
and (n3795,n1641,n116);
or (n3796,n3797,n3798);
and (n3797,n1858,n1883);
and (n3798,n1859,n1866);
or (n3799,n3800,n3801);
and (n3800,n2274,n2281);
and (n3801,n2275,n2278);
and (n3802,n3761,n3764);
or (n3803,n3804,n3873);
and (n3804,n3805,n3870);
xor (n3805,n3806,n3833);
xor (n3806,n3807,n3822);
xor (n3807,n3808,n3819);
xor (n3808,n3809,n3816);
xor (n3809,n3810,n3813);
or (n3810,n3811,n3812);
and (n3811,n1668,n1681);
and (n3812,n1669,n1675);
or (n3813,n3814,n3815);
and (n3814,n1688,n1707);
and (n3815,n1689,n1696);
or (n3816,n3817,n3818);
and (n3817,n1836,n1850);
and (n3818,n1837,n1844);
or (n3819,n3820,n3821);
and (n3820,n1736,n1784);
and (n3821,n1737,n1762);
xor (n3822,n3823,n3830);
xor (n3823,n3824,n3827);
or (n3824,n3825,n3826);
and (n3825,n1715,n1729);
and (n3826,n1716,n1722);
or (n3827,n3828,n3829);
and (n3828,n1810,n1828);
and (n3829,n1811,n1821);
or (n3830,n3831,n3832);
and (n3831,n1785,n1799);
and (n3832,n1786,n1792);
xor (n3833,n3834,n3867);
xor (n3834,n3835,n3838);
or (n3835,n3836,n3837);
and (n3836,n1620,n1627);
and (n3837,n1621,n1624);
xor (n3838,n3839,n3846);
xor (n3839,n3840,n3843);
or (n3840,n3841,n3842);
and (n3841,n1763,n1777);
and (n3842,n1764,n1771);
or (n3843,n3844,n3845);
and (n3844,n1738,n1755);
and (n3845,n1739,n1745);
xor (n3846,n3847,n3860);
xor (n3847,n3848,n3856);
nand (n3848,n3849,n3854);
or (n3849,n316,n3850);
not (n3850,n3851);
nand (n3851,n3852,n3853);
or (n3852,n290,n222);
nand (n3853,n290,n222);
or (n3854,n315,n3855);
not (n3855,n1768);
nand (n3856,n3857,n3859);
or (n3857,n3858,n1173);
not (n3858,n1841);
or (n3859,n1181,n1176);
nand (n3860,n3861,n3863);
or (n3861,n373,n3862);
not (n3862,n1742);
or (n3863,n3864,n522);
nor (n3864,n3865,n3866);
and (n3865,n153,n1215);
and (n3866,n151,n2090);
or (n3867,n3868,n3869);
and (n3868,n1666,n1714);
and (n3869,n1667,n1687);
or (n3870,n3871,n3872);
and (n3871,n1618,n1735);
and (n3872,n1619,n1665);
and (n3873,n3806,n3833);
or (n3874,n3875,n3882);
and (n3875,n3876,n3879);
xor (n3876,n3877,n3878);
xor (n3877,n3760,n3767);
xor (n3878,n3805,n3870);
or (n3879,n3880,n3881);
and (n3880,n1100,n1805);
and (n3881,n1101,n1617);
and (n3882,n3877,n3878);
xor (n3883,n3884,n4120);
xor (n3884,n3885,n3921);
xor (n3885,n3886,n3918);
xor (n3886,n3887,n3890);
or (n3887,n3888,n3889);
and (n3888,n3807,n3822);
and (n3889,n3808,n3819);
xor (n3890,n3891,n3898);
xor (n3891,n3892,n3895);
or (n3892,n3893,n3894);
and (n3893,n3823,n3830);
and (n3894,n3824,n3827);
or (n3895,n3896,n3897);
and (n3896,n3809,n3816);
and (n3897,n3810,n3813);
xor (n3898,n3899,n3917);
xor (n3899,n3900,n3906);
nand (n3900,n3901,n3902);
or (n3901,n171,n3774);
or (n3902,n172,n3903);
nor (n3903,n3904,n3905);
and (n3904,n195,n279);
and (n3905,n180,n278);
xor (n3906,n3907,n3910);
nor (n3907,n3908,n3909);
and (n3908,n1192,n1197);
and (n3909,n3784,n1195);
not (n3910,n3911);
nand (n3911,n3912,n3913);
or (n3912,n3793,n118);
nand (n3913,n3914,n125);
nor (n3914,n3915,n3916);
and (n3915,n116,n1163);
and (n3916,n115,n1162);
and (n3917,n3781,n3789);
or (n3918,n3919,n3920);
and (n3919,n3834,n3867);
and (n3920,n3835,n3838);
xor (n3921,n3922,n3994);
xor (n3922,n3923,n3942);
xor (n3923,n3924,n3939);
xor (n3924,n3925,n3928);
or (n3925,n3926,n3927);
and (n3926,n3689,n3733);
and (n3927,n3690,n3712);
xor (n3928,n3929,n3936);
xor (n3929,n3930,n3933);
or (n3930,n3931,n3932);
and (n3931,n3623,n3634);
and (n3932,n3624,n3627);
or (n3933,n3934,n3935);
and (n3934,n3691,n3706);
and (n3935,n3692,n3699);
or (n3936,n3937,n3938);
and (n3937,n3665,n3680);
and (n3938,n3666,n3673);
or (n3939,n3940,n3941);
and (n3940,n3621,n3664);
and (n3941,n3622,n3640);
xor (n3942,n3943,n3958);
xor (n3943,n3944,n3947);
or (n3944,n3945,n3946);
and (n3945,n3839,n3846);
and (n3946,n3840,n3843);
xor (n3947,n3948,n3955);
xor (n3948,n3949,n3952);
or (n3949,n3950,n3951);
and (n3950,n3713,n3727);
and (n3951,n3714,n3721);
or (n3952,n3953,n3954);
and (n3953,n3734,n3748);
and (n3954,n3735,n3742);
or (n3955,n3956,n3957);
and (n3956,n3847,n3860);
and (n3957,n3848,n3856);
xor (n3958,n3959,n3980);
xor (n3959,n3960,n3963);
or (n3960,n3961,n3962);
and (n3961,n3641,n3656);
and (n3962,n3642,n3649);
xor (n3963,n3964,n3972);
xor (n3964,n1146,n3965);
nand (n3965,n3966,n3968);
or (n3966,n3967,n281);
not (n3967,n3631);
nand (n3968,n288,n3969);
nand (n3969,n3970,n3971);
or (n3970,n217,n266);
nand (n3971,n217,n266);
nand (n3972,n3973,n3975);
or (n3973,n420,n3974);
not (n3974,n3637);
or (n3975,n3976,n424);
not (n3976,n3977);
nand (n3977,n3978,n3979);
or (n3978,n477,n409);
nand (n3979,n409,n477);
xor (n3980,n3981,n3988);
xor (n3981,n3982,n1175);
nand (n3982,n3983,n3984);
or (n3983,n3850,n315);
nand (n3984,n317,n3985);
nand (n3985,n3986,n3987);
or (n3986,n53,n290);
nand (n3987,n290,n53);
nand (n3988,n3989,n3990);
or (n3989,n373,n3864);
or (n3990,n522,n3991);
nor (n3991,n3992,n3993);
and (n3992,n153,n1344);
and (n3993,n151,n1576);
xor (n3994,n3995,n4117);
xor (n3995,n3996,n4065);
xor (n3996,n3997,n4041);
xor (n3997,n3998,n4020);
xor (n3998,n3999,n4014);
xor (n3999,n4000,n4007);
nand (n4000,n4001,n4003);
or (n4001,n4002,n1223);
not (n4002,n3646);
nand (n4003,n4004,n1238);
nand (n4004,n4005,n4006);
or (n4005,n358,n202);
nand (n4006,n202,n358);
nand (n4007,n4008,n4010);
or (n4008,n4009,n37);
not (n4009,n3653);
nand (n4010,n4011,n46);
nand (n4011,n4012,n4013);
or (n4012,n42,n1124);
nand (n4013,n42,n1124);
nand (n4014,n4015,n4016);
or (n4015,n3660,n103);
nand (n4016,n96,n4017);
nand (n4017,n4018,n4019);
or (n4018,n107,n312);
nand (n4019,n312,n107);
xor (n4020,n4021,n4035);
xor (n4021,n4022,n4028);
nand (n4022,n4023,n4024);
nand (n4023,n3670,n200,n207);
nand (n4024,n4025,n1118);
nand (n4025,n4026,n4027);
or (n4026,n79,n209);
nand (n4027,n209,n79);
nand (n4028,n4029,n4031);
or (n4029,n4030,n400);
not (n4030,n3677);
nand (n4031,n4032,n405);
nand (n4032,n4033,n4034);
or (n4033,n434,n395);
nand (n4034,n395,n434);
nand (n4035,n4036,n4037);
or (n4036,n3684,n64);
nand (n4037,n4038,n1006);
nor (n4038,n4039,n4040);
and (n4039,n1659,n74);
and (n4040,n114,n75);
xor (n4041,n4042,n4057);
xor (n4042,n4043,n4050);
nand (n4043,n4044,n4046);
or (n4044,n4045,n1590);
not (n4045,n3696);
nand (n4046,n4047,n1601);
nand (n4047,n4048,n4049);
or (n4048,n186,n1588);
nand (n4049,n1588,n186);
nand (n4050,n4051,n4053);
or (n4051,n4052,n470);
not (n4052,n3703);
nand (n4053,n566,n4054);
nand (n4054,n4055,n4056);
or (n4055,n371,n440);
nand (n4056,n440,n371);
nand (n4057,n4058,n4063);
or (n4058,n149,n4059);
not (n4059,n4060);
nor (n4060,n4061,n4062);
and (n4061,n147,n1399);
and (n4062,n144,n1210);
or (n4063,n138,n4064);
not (n4064,n3709);
xor (n4065,n4066,n4114);
xor (n4066,n4067,n4091);
xor (n4067,n4068,n4083);
xor (n4068,n4069,n4076);
nand (n4069,n4070,n4072);
or (n4070,n4071,n532);
not (n4071,n3718);
nand (n4072,n4073,n333);
nand (n4073,n4074,n4075);
or (n4074,n1357,n127);
nand (n4075,n127,n1357);
nand (n4076,n4077,n4079);
or (n4077,n4078,n255);
not (n4078,n3724);
nand (n4079,n4080,n272);
nand (n4080,n4081,n4082);
or (n4081,n1305,n253);
nand (n4082,n1305,n253);
nand (n4083,n4084,n4086);
or (n4084,n22,n4085);
not (n4085,n3730);
or (n4086,n4087,n23);
not (n4087,n4088);
nor (n4088,n4089,n4090);
and (n4089,n33,n483);
and (n4090,n32,n485);
xor (n4091,n4092,n4107);
xor (n4092,n4093,n4100);
nand (n4093,n4094,n4096);
or (n4094,n4095,n436);
not (n4095,n3739);
nand (n4096,n4097,n449);
nand (n4097,n4098,n4099);
or (n4098,n156,n382);
nand (n4099,n382,n156);
nand (n4100,n4101,n4103);
or (n4101,n4102,n1138);
not (n4102,n3745);
nand (n4103,n4104,n1154);
nand (n4104,n4105,n4106);
or (n4105,n397,n415);
nand (n4106,n397,n415);
nand (n4107,n4108,n4113);
or (n4108,n4109,n235);
not (n4109,n4110);
nand (n4110,n4111,n4112);
or (n4111,n348,n67);
or (n4112,n347,n68);
or (n4113,n234,n3751);
or (n4114,n4115,n4116);
and (n4115,n3770,n3780);
and (n4116,n3771,n3777);
or (n4117,n4118,n4119);
and (n4118,n3768,n3799);
and (n4119,n3769,n3796);
or (n4120,n4121,n4130);
and (n4121,n4122,n4127);
xor (n4122,n4123,n4124);
xor (n4123,n3619,n3754);
or (n4124,n4125,n4126);
and (n4125,n1806,n1981);
and (n4126,n1807,n1886);
or (n4127,n4128,n4129);
and (n4128,n2250,n2265);
and (n4129,n2251,n2254);
and (n4130,n4123,n4124);
or (n4131,n4132,n4139);
and (n4132,n4133,n4138);
xor (n4133,n4134,n4135);
xor (n4134,n4122,n4127);
or (n4135,n4136,n4137);
and (n4136,n2128,n2284);
and (n4137,n2129,n2249);
xor (n4138,n3876,n3879);
and (n4139,n4134,n4135);
nor (n4140,n4141,n4142);
xor (n4141,n4133,n4138);
or (n4142,n4143,n4144);
and (n4143,n1098,n2297);
and (n4144,n1099,n2127);
nor (n4145,n4146,n4928);
nor (n4146,n4147,n4897);
xor (n4147,n4148,n4862);
xor (n4148,n4149,n4669);
xor (n4149,n4150,n4607);
xor (n4150,n4151,n4275);
xor (n4151,n4152,n4268);
xor (n4152,n4153,n4239);
or (n4153,n4154,n4238);
and (n4154,n4155,n4209);
xor (n4155,n4156,n4182);
xor (n4156,n4157,n4172);
xor (n4157,n4158,n4162);
not (n4158,n4159);
nor (n4159,n4160,n415);
and (n4160,n4161,n1144);
not (n4161,n1140);
nand (n4162,n4163,n4168);
or (n4163,n4164,n373);
not (n4164,n4165);
nor (n4165,n4166,n4167);
and (n4166,n153,n158);
and (n4167,n151,n156);
nand (n4168,n4169,n380);
nor (n4169,n4170,n4171);
and (n4170,n153,n164);
and (n4171,n151,n162);
nand (n4172,n4173,n4178);
or (n4173,n4174,n64);
not (n4174,n4175);
nor (n4175,n4176,n4177);
and (n4176,n75,n348);
and (n4177,n74,n347);
nand (n4178,n4179,n1006);
nand (n4179,n4180,n4181);
or (n4180,n340,n75);
or (n4181,n74,n341);
xor (n4182,n4183,n4200);
xor (n4183,n4184,n4191);
nand (n4184,n4185,n4190);
or (n4185,n4186,n281);
not (n4186,n4187);
nand (n4187,n4188,n4189);
or (n4188,n53,n265);
nand (n4189,n53,n265);
nand (n4190,n980,n288);
nand (n4191,n4192,n4196);
or (n4192,n4193,n22);
nor (n4193,n4194,n4195);
and (n4194,n32,n79);
and (n4195,n33,n81);
nand (n4196,n4197,n24);
nor (n4197,n4198,n4199);
and (n4198,n32,n87);
and (n4199,n33,n85);
nand (n4200,n4201,n4205);
or (n4201,n470,n4202);
nor (n4202,n4203,n4204);
and (n4203,n440,n434);
and (n4204,n441,n521);
or (n4205,n4206,n457);
nor (n4206,n4207,n4208);
and (n4207,n453,n440);
and (n4208,n452,n441);
xor (n4209,n4210,n4232);
xor (n4210,n4211,n4222);
nand (n4211,n4212,n4217);
or (n4212,n316,n4213);
not (n4213,n4214);
nor (n4214,n4215,n4216);
and (n4215,n290,n296);
and (n4216,n291,n297);
or (n4217,n315,n4218);
not (n4218,n4219);
nand (n4219,n4220,n4221);
or (n4220,n291,n278);
nand (n4221,n291,n278);
nand (n4222,n4223,n4228);
or (n4223,n4224,n400);
not (n4224,n4225);
nor (n4225,n4226,n4227);
and (n4226,n476,n395);
and (n4227,n477,n396);
or (n4228,n4229,n529);
nor (n4229,n4230,n4231);
and (n4230,n395,n466);
and (n4231,n465,n396);
nand (n4232,n4233,n4237);
or (n4233,n4234,n199);
nor (n4234,n4235,n4236);
and (n4235,n360,n28);
and (n4236,n358,n209);
nand (n4237,n1118,n28);
and (n4238,n4156,n4182);
xor (n4239,n4240,n4258);
xor (n4240,n4241,n4242);
xor (n4241,n915,n931);
xor (n4242,n4243,n4254);
xor (n4243,n4244,n4251);
nand (n4244,n4245,n4250);
or (n4245,n4246,n436);
not (n4246,n4247);
nor (n4247,n4248,n4249);
and (n4248,n388,n382);
and (n4249,n389,n383);
nand (n4250,n432,n449);
nand (n4251,n4252,n4253);
or (n4252,n4206,n470);
nand (n4253,n566,n474);
nand (n4254,n4255,n4257);
or (n4255,n64,n4256);
not (n4256,n4179);
or (n4257,n481,n65);
xor (n4258,n4259,n4267);
xor (n4259,n4260,n4264);
nand (n4260,n4261,n4263);
or (n4261,n373,n4262);
not (n4262,n4169);
or (n4263,n368,n522);
nand (n4264,n4265,n4266);
or (n4265,n400,n4229);
or (n4266,n393,n529);
not (n4267,n411);
xor (n4268,n4269,n4274);
xor (n4269,n4270,n4273);
or (n4270,n4271,n4272);
and (n4271,n4157,n4172);
and (n4272,n4158,n4162);
xor (n4273,n942,n950);
xor (n4274,n962,n977);
or (n4275,n4276,n4606);
and (n4276,n4277,n4477);
xor (n4277,n4278,n4380);
xor (n4278,n4279,n4328);
xor (n4279,n4280,n4304);
xor (n4280,n4281,n4295);
xor (n4281,n4282,n4288);
nand (n4282,n4283,n4287);
or (n4283,n138,n4284);
nor (n4284,n4285,n4286);
and (n4285,n147,n1344);
and (n4286,n144,n1576);
or (n4287,n933,n149);
nand (n4288,n4289,n4294);
or (n4289,n436,n4290);
not (n4290,n4291);
nor (n4291,n4292,n4293);
and (n4292,n371,n383);
and (n4293,n370,n382);
or (n4294,n438,n4246);
nand (n4295,n4296,n4300);
or (n4296,n532,n4297);
nor (n4297,n4298,n4299);
and (n4298,n127,n114);
and (n4299,n128,n1659);
or (n4300,n4301,n332);
nor (n4301,n4302,n4303);
and (n4302,n127,n134);
and (n4303,n133,n128);
xor (n4304,n4305,n4320);
xor (n4305,n4306,n4313);
nand (n4306,n4307,n4308);
or (n4307,n263,n972);
or (n4308,n255,n4309);
not (n4309,n4310);
nand (n4310,n4311,n4312);
or (n4311,n48,n217);
nand (n4312,n217,n48);
nand (n4313,n4314,n4319);
or (n4314,n4315,n171);
not (n4315,n4316);
nor (n4316,n4317,n4318);
and (n4317,n312,n195);
and (n4318,n313,n180);
nand (n4319,n189,n946);
nand (n4320,n4321,n4326);
or (n4321,n103,n4322);
not (n4322,n4323);
nand (n4323,n4324,n4325);
or (n4324,n107,n185);
or (n4325,n177,n186);
or (n4326,n104,n4327);
not (n4327,n918);
or (n4328,n4329,n4379);
and (n4329,n4330,n4371);
xor (n4330,n4331,n4347);
or (n4331,n4332,n4340);
nand (n4332,n4333,n4335);
or (n4333,n281,n4334);
not (n4334,n3969);
nand (n4335,n4336,n288);
not (n4336,n4337);
nor (n4337,n4338,n4339);
and (n4338,n222,n265);
and (n4339,n221,n266);
nand (n4340,n4341,n4343);
or (n4341,n4342,n532);
not (n4342,n4073);
nand (n4343,n4344,n333);
nand (n4344,n4345,n4346);
or (n4345,n927,n128);
or (n4346,n127,n928);
or (n4347,n4348,n4370);
and (n4348,n4349,n4363);
xor (n4349,n4350,n4356);
nand (n4350,n4351,n4352);
or (n4351,n3976,n420);
nand (n4352,n4353,n413);
nand (n4353,n4354,n4355);
or (n4354,n466,n409);
nand (n4355,n409,n466);
nand (n4356,n4357,n4359);
or (n4357,n4358,n37);
not (n4358,n4011);
nand (n4359,n46,n4360);
nor (n4360,n4361,n4362);
and (n4361,n1130,n41);
and (n4362,n1131,n42);
nand (n4363,n4364,n4366);
or (n4364,n4365,n118);
not (n4365,n3914);
nand (n4366,n125,n4367);
nor (n4367,n4368,n4369);
and (n4368,n115,n1168);
and (n4369,n116,n1169);
and (n4370,n4350,n4356);
or (n4371,n4372,n4378);
and (n4372,n4373,n1181);
xor (n4373,n1191,n4374);
nand (n4374,n4375,n4377);
or (n4375,n4376,n1138);
not (n4376,n4104);
nand (n4377,n1154,n416);
and (n4378,n1191,n4374);
and (n4379,n4331,n4347);
or (n4380,n4381,n4476);
and (n4381,n4382,n4475);
xor (n4382,n4383,n4434);
or (n4383,n4384,n4433);
and (n4384,n4385,n4409);
xor (n4385,n4386,n4387);
xor (n4386,n4349,n4363);
xor (n4387,n4388,n4402);
xor (n4388,n4389,n4395);
nand (n4389,n4390,n4391);
or (n4390,n4087,n22);
nand (n4391,n24,n4392);
nand (n4392,n4393,n4394);
or (n4393,n489,n32);
nand (n4394,n489,n32);
nand (n4395,n4396,n4398);
or (n4396,n4397,n470);
not (n4397,n4054);
nand (n4398,n566,n4399);
nand (n4399,n4400,n4401);
or (n4400,n389,n440);
nand (n4401,n440,n389);
nand (n4402,n4403,n4405);
or (n4403,n400,n4404);
not (n4404,n4032);
or (n4405,n4406,n529);
nor (n4406,n4407,n4408);
and (n4407,n453,n395);
and (n4408,n452,n396);
xor (n4409,n4410,n4425);
xor (n4410,n4411,n4418);
nand (n4411,n4412,n4414);
or (n4412,n4413,n1590);
not (n4413,n4047);
nand (n4414,n1601,n4415);
nor (n4415,n4416,n4417);
and (n4416,n192,n1588);
and (n4417,n193,n100);
nand (n4418,n4419,n4421);
or (n4419,n436,n4420);
not (n4420,n4097);
nand (n4421,n449,n4422);
nand (n4422,n4423,n4424);
or (n4423,n164,n383);
or (n4424,n382,n162);
nand (n4425,n4426,n4428);
or (n4426,n255,n4427);
not (n4427,n4080);
or (n4428,n263,n4429);
not (n4429,n4430);
nand (n4430,n4431,n4432);
or (n4431,n48,n955);
nand (n4432,n955,n48);
and (n4433,n4386,n4387);
xor (n4434,n4435,n4462);
xor (n4435,n4436,n4459);
or (n4436,n4437,n4458);
and (n4437,n4438,n4450);
xor (n4438,n4439,n4446);
nand (n4439,n4440,n4442);
or (n4440,n4441,n199);
not (n4441,n4025);
nand (n4442,n1118,n4443);
nand (n4443,n4444,n4445);
or (n4444,n85,n209);
or (n4445,n87,n28);
nand (n4446,n4447,n4449);
or (n4447,n4448,n1223);
not (n4448,n4004);
nand (n4449,n1238,n203);
nand (n4450,n4451,n4456);
or (n4451,n4452,n104);
not (n4452,n4453);
nand (n4453,n4454,n4455);
or (n4454,n327,n107);
or (n4455,n177,n328);
or (n4456,n103,n4457);
not (n4457,n4017);
and (n4458,n4439,n4446);
or (n4459,n4460,n4461);
and (n4460,n4388,n4402);
and (n4461,n4389,n4395);
xor (n4462,n4463,n4471);
xor (n4463,n4464,n4467);
nand (n4464,n4465,n4466);
or (n4465,n281,n4337);
nand (n4466,n288,n4187);
nand (n4467,n4468,n4470);
or (n4468,n22,n4469);
not (n4469,n4392);
or (n4470,n4193,n23);
nand (n4471,n4472,n4474);
or (n4472,n470,n4473);
not (n4473,n4399);
or (n4474,n4202,n457);
xor (n4475,n4330,n4371);
and (n4476,n4383,n4434);
xor (n4477,n4478,n4577);
xor (n4478,n4479,n4527);
or (n4479,n4480,n4526);
and (n4480,n4481,n4523);
xor (n4481,n4482,n4499);
or (n4482,n4483,n4498);
and (n4483,n4484,n4491);
xor (n4484,n4485,n1149);
nand (n4485,n4486,n4487);
or (n4486,n4059,n138);
nand (n4487,n4488,n148);
nor (n4488,n4489,n4490);
and (n4489,n147,n2090);
and (n4490,n144,n1215);
nand (n4491,n4492,n4494);
or (n4492,n315,n4493);
not (n4493,n3985);
or (n4494,n4495,n316);
nor (n4495,n4496,n4497);
and (n4496,n290,n59);
and (n4497,n291,n61);
and (n4498,n4485,n1149);
or (n4499,n4500,n4522);
and (n4500,n4501,n4515);
xor (n4501,n4502,n4508);
nand (n4502,n4503,n4504);
or (n4503,n4109,n234);
nand (n4504,n4505,n247);
nand (n4505,n4506,n4507);
or (n4506,n341,n67);
nand (n4507,n341,n67);
nand (n4508,n4509,n4511);
or (n4509,n4510,n64);
not (n4510,n4038);
nand (n4511,n4512,n1006);
nor (n4512,n4513,n4514);
and (n4513,n74,n133);
and (n4514,n75,n134);
nand (n4515,n4516,n4517);
or (n4516,n373,n3991);
or (n4517,n4518,n522);
not (n4518,n4519);
nor (n4519,n4520,n4521);
and (n4520,n153,n937);
and (n4521,n151,n935);
and (n4522,n4502,n4508);
or (n4523,n4524,n4525);
and (n4524,n4410,n4425);
and (n4525,n4411,n4418);
and (n4526,n4482,n4499);
xor (n4527,n4528,n4560);
xor (n4528,n4529,n4546);
or (n4529,n4530,n4545);
and (n4530,n4531,n4542);
xor (n4531,n4532,n4535);
nand (n4532,n4533,n4534);
or (n4533,n4429,n255);
nand (n4534,n4310,n272);
nand (n4535,n4536,n4541);
or (n4536,n4537,n171);
not (n4537,n4538);
nor (n4538,n4539,n4540);
and (n4539,n195,n296);
and (n4540,n180,n297);
nand (n4541,n4316,n189);
nand (n4542,n4543,n4544);
or (n4543,n4452,n103);
nand (n4544,n96,n4323);
and (n4545,n4532,n4535);
or (n4546,n4547,n4559);
and (n4547,n4548,n4555);
xor (n4548,n4549,n4552);
nand (n4549,n4550,n4551);
or (n4550,n4495,n315);
nand (n4551,n4219,n317);
nand (n4552,n4553,n4554);
or (n4553,n4406,n400);
nand (n4554,n4225,n405);
nand (n4555,n4556,n4558);
or (n4556,n199,n4557);
not (n4557,n4443);
or (n4558,n4234,n200);
and (n4559,n4549,n4552);
or (n4560,n4561,n4576);
and (n4561,n4562,n4572);
xor (n4562,n4563,n4568);
nand (n4563,n4564,n4566);
or (n4564,n4565,n138);
not (n4565,n4488);
nand (n4566,n4567,n148);
not (n4567,n4284);
nand (n4568,n4569,n4571);
or (n4569,n4570,n436);
not (n4570,n4422);
nand (n4571,n449,n4291);
nand (n4572,n4573,n4575);
or (n4573,n532,n4574);
not (n4574,n4344);
or (n4575,n4297,n332);
and (n4576,n4563,n4568);
or (n4577,n4578,n4605);
and (n4578,n4579,n4604);
xor (n4579,n4580,n4603);
xor (n4580,n4581,n4596);
xor (n4581,n4582,n4589);
nand (n4582,n4583,n4585);
or (n4583,n4584,n37);
not (n4584,n4360);
nand (n4585,n46,n4586);
nor (n4586,n4587,n4588);
and (n4587,n41,n1304);
and (n4588,n42,n1305);
nand (n4589,n4590,n4592);
or (n4590,n4591,n234);
not (n4591,n4505);
nand (n4592,n4593,n247);
nor (n4593,n4594,n4595);
and (n4594,n67,n485);
and (n4595,n68,n483);
nand (n4596,n4597,n4599);
or (n4597,n420,n4598);
not (n4598,n4353);
or (n4599,n4600,n424);
nor (n4600,n4601,n4602);
and (n4601,n409,n397);
and (n4602,n407,n399);
xor (n4603,n4548,n4555);
xor (n4604,n4562,n4572);
and (n4605,n4580,n4603);
and (n4606,n4278,n4380);
xor (n4607,n4608,n4615);
xor (n4608,n4609,n4612);
or (n4609,n4610,n4611);
and (n4610,n4279,n4328);
and (n4611,n4280,n4304);
or (n4612,n4613,n4614);
and (n4613,n4478,n4577);
and (n4614,n4479,n4527);
xor (n4615,n4616,n4666);
xor (n4616,n4617,n4629);
xor (n4617,n4618,n4625);
xor (n4618,n4619,n4622);
nand (n4619,n4620,n4621);
or (n4620,n315,n4213);
or (n4621,n309,n316);
nand (n4622,n4623,n4624);
or (n4623,n532,n4301);
or (n4624,n345,n332);
nand (n4625,n4626,n4627);
or (n4626,n356,n23);
or (n4627,n22,n4628);
not (n4628,n4197);
or (n4629,n4630,n4665);
and (n4630,n4631,n4654);
xor (n4631,n4632,n4651);
or (n4632,n4633,n4650);
and (n4633,n4634,n4646);
xor (n4634,n4635,n4639);
nand (n4635,n4636,n4638);
or (n4636,n4637,n1590);
not (n4637,n4415);
nand (n4638,n1601,n100);
nand (n4639,n4640,n4642);
or (n4640,n4641,n118);
not (n4641,n4367);
nand (n4642,n4643,n125);
nor (n4643,n4644,n4645);
and (n4644,n115,n1356);
and (n4645,n116,n1357);
not (n4646,n4647);
nand (n4647,n4648,n203);
or (n4648,n1238,n4649);
not (n4649,n1223);
and (n4650,n4635,n4639);
or (n4651,n4652,n4653);
and (n4652,n4463,n4471);
and (n4653,n4464,n4467);
or (n4654,n4655,n4664);
and (n4655,n4656,n4660);
xor (n4656,n4159,n4657);
nand (n4657,n4658,n4659);
or (n4658,n4518,n373);
nand (n4659,n4165,n380);
nand (n4660,n4661,n4663);
or (n4661,n4662,n64);
not (n4662,n4512);
nand (n4663,n4175,n1006);
and (n4664,n4159,n4657);
and (n4665,n4632,n4651);
or (n4666,n4667,n4668);
and (n4667,n4528,n4560);
and (n4668,n4529,n4546);
xor (n4669,n4670,n4815);
xor (n4670,n4671,n4787);
xor (n4671,n4672,n4740);
xor (n4672,n4673,n4688);
or (n4673,n4674,n4687);
and (n4674,n4675,n4686);
xor (n4675,n4676,n4683);
or (n4676,n4677,n4682);
and (n4677,n4678,n4681);
xor (n4678,n4679,n4680);
xor (n4679,n4656,n4660);
xor (n4680,n4531,n4542);
xor (n4681,n4634,n4646);
and (n4682,n4679,n4680);
or (n4683,n4684,n4685);
and (n4684,n4435,n4462);
and (n4685,n4436,n4459);
xor (n4686,n4631,n4654);
and (n4687,n4676,n4683);
xor (n4688,n4689,n4731);
xor (n4689,n4690,n4708);
xor (n4690,n4691,n4705);
xor (n4691,n4692,n4702);
or (n4692,n4693,n4701);
and (n4693,n4694,n4647);
xor (n4694,n4695,n4697);
nand (n4695,n4696,n100);
or (n4696,n1594,n1191);
nand (n4697,n4698,n4700);
or (n4698,n4699,n118);
not (n4699,n4643);
nand (n4700,n925,n125);
and (n4701,n4695,n4697);
or (n4702,n4703,n4704);
and (n4703,n4183,n4200);
and (n4704,n4184,n4191);
or (n4705,n4706,n4707);
and (n4706,n4210,n4232);
and (n4707,n4211,n4222);
xor (n4708,n4709,n4728);
xor (n4709,n4710,n4725);
or (n4710,n4711,n4724);
and (n4711,n4712,n4721);
xor (n4712,n4713,n4717);
nand (n4713,n4714,n4716);
or (n4714,n4715,n37);
not (n4715,n4586);
nand (n4716,n953,n46);
nand (n4717,n4718,n4720);
or (n4718,n4719,n234);
not (n4719,n4593);
nand (n4720,n966,n247);
nand (n4721,n4722,n4723);
or (n4722,n420,n4600);
or (n4723,n424,n409);
and (n4724,n4713,n4717);
or (n4725,n4726,n4727);
and (n4726,n4305,n4320);
and (n4727,n4306,n4313);
or (n4728,n4729,n4730);
and (n4729,n4281,n4295);
and (n4730,n4282,n4288);
or (n4731,n4732,n4739);
and (n4732,n4733,n4738);
xor (n4733,n4734,n4737);
or (n4734,n4735,n4736);
and (n4735,n4581,n4596);
and (n4736,n4582,n4589);
xor (n4737,n4694,n4647);
xor (n4738,n4712,n4721);
and (n4739,n4734,n4737);
or (n4740,n4741,n4786);
and (n4741,n4742,n4745);
xor (n4742,n4743,n4744);
xor (n4743,n4155,n4209);
xor (n4744,n4733,n4738);
or (n4745,n4746,n4785);
and (n4746,n4747,n4772);
xor (n4747,n4748,n4761);
or (n4748,n4749,n4760);
and (n4749,n4750,n4757);
xor (n4750,n4751,n4754);
or (n4751,n4752,n4753);
and (n4752,n4021,n4035);
and (n4753,n4022,n4028);
or (n4754,n4755,n4756);
and (n4755,n4092,n4107);
and (n4756,n4093,n4100);
or (n4757,n4758,n4759);
and (n4758,n4042,n4057);
and (n4759,n4043,n4050);
and (n4760,n4751,n4754);
or (n4761,n4762,n4771);
and (n4762,n4763,n4768);
xor (n4763,n4764,n4767);
nand (n4764,n4765,n4766);
or (n4765,n171,n3903);
or (n4766,n172,n4537);
nor (n4767,n3910,n3907);
or (n4768,n4769,n4770);
and (n4769,n4068,n4083);
and (n4770,n4069,n4076);
and (n4771,n4764,n4767);
or (n4772,n4773,n4784);
and (n4773,n4774,n4781);
xor (n4774,n4775,n4778);
or (n4775,n4776,n4777);
and (n4776,n3999,n4014);
and (n4777,n4000,n4007);
or (n4778,n4779,n4780);
and (n4779,n3964,n3972);
and (n4780,n1146,n3965);
or (n4781,n4782,n4783);
and (n4782,n3981,n3988);
and (n4783,n3982,n1175);
and (n4784,n4775,n4778);
and (n4785,n4748,n4761);
and (n4786,n4743,n4744);
or (n4787,n4788,n4814);
and (n4788,n4789,n4813);
xor (n4789,n4790,n4812);
or (n4790,n4791,n4811);
and (n4791,n4792,n4802);
xor (n4792,n4793,n4801);
or (n4793,n4794,n4800);
and (n4794,n4795,n4799);
xor (n4795,n4796,n4798);
nand (n4796,n4331,n4797);
nand (n4797,n4332,n4340);
xor (n4798,n4438,n4450);
xor (n4799,n4484,n4491);
and (n4800,n4796,n4798);
xor (n4801,n4481,n4523);
or (n4802,n4803,n4810);
and (n4803,n4804,n4807);
xor (n4804,n4805,n4806);
xor (n4805,n4501,n4515);
xor (n4806,n4373,n1181);
or (n4807,n4808,n4809);
and (n4808,n3899,n3917);
and (n4809,n3900,n3906);
and (n4810,n4805,n4806);
and (n4811,n4793,n4801);
xor (n4812,n4675,n4686);
xor (n4813,n4742,n4745);
and (n4814,n4790,n4812);
or (n4815,n4816,n4861);
and (n4816,n4817,n4860);
xor (n4817,n4818,n4835);
or (n4818,n4819,n4834);
and (n4819,n4820,n4823);
xor (n4820,n4821,n4822);
xor (n4821,n4678,n4681);
xor (n4822,n4579,n4604);
or (n4823,n4824,n4833);
and (n4824,n4825,n4830);
xor (n4825,n4826,n4829);
or (n4826,n4827,n4828);
and (n4827,n3929,n3936);
and (n4828,n3930,n3933);
xor (n4829,n4763,n4768);
or (n4830,n4831,n4832);
and (n4831,n3948,n3955);
and (n4832,n3949,n3952);
and (n4833,n4826,n4829);
and (n4834,n4821,n4822);
or (n4835,n4836,n4859);
and (n4836,n4837,n4850);
xor (n4837,n4838,n4849);
or (n4838,n4839,n4848);
and (n4839,n4840,n4845);
xor (n4840,n4841,n4842);
xor (n4841,n4750,n4757);
or (n4842,n4843,n4844);
and (n4843,n3997,n4041);
and (n4844,n3998,n4020);
or (n4845,n4846,n4847);
and (n4846,n3959,n3980);
and (n4847,n3960,n3963);
and (n4848,n4841,n4842);
xor (n4849,n4747,n4772);
or (n4850,n4851,n4858);
and (n4851,n4852,n4855);
xor (n4852,n4853,n4854);
xor (n4853,n4774,n4781);
xor (n4854,n4795,n4799);
or (n4855,n4856,n4857);
and (n4856,n4066,n4114);
and (n4857,n4067,n4091);
and (n4858,n4853,n4854);
and (n4859,n4838,n4849);
xor (n4860,n4277,n4477);
and (n4861,n4818,n4835);
or (n4862,n4863,n4896);
and (n4863,n4864,n4881);
xor (n4864,n4865,n4866);
xor (n4865,n4789,n4813);
or (n4866,n4867,n4880);
and (n4867,n4868,n4871);
xor (n4868,n4869,n4870);
xor (n4869,n4382,n4475);
xor (n4870,n4792,n4802);
or (n4871,n4872,n4879);
and (n4872,n4873,n4876);
xor (n4873,n4874,n4875);
xor (n4874,n4385,n4409);
xor (n4875,n4804,n4807);
or (n4876,n4877,n4878);
and (n4877,n3891,n3898);
and (n4878,n3892,n3895);
and (n4879,n4874,n4875);
and (n4880,n4869,n4870);
or (n4881,n4882,n4895);
and (n4882,n4883,n4894);
xor (n4883,n4884,n4885);
xor (n4884,n4820,n4823);
or (n4885,n4886,n4893);
and (n4886,n4887,n4892);
xor (n4887,n4888,n4889);
xor (n4888,n4825,n4830);
or (n4889,n4890,n4891);
and (n4890,n3924,n3939);
and (n4891,n3925,n3928);
xor (n4892,n4840,n4845);
and (n4893,n4888,n4889);
xor (n4894,n4837,n4850);
and (n4895,n4884,n4885);
and (n4896,n4865,n4866);
or (n4897,n4898,n4927);
and (n4898,n4899,n4902);
xor (n4899,n4900,n4901);
xor (n4900,n4817,n4860);
xor (n4901,n4864,n4881);
or (n4902,n4903,n4926);
and (n4903,n4904,n4917);
xor (n4904,n4905,n4916);
or (n4905,n4906,n4915);
and (n4906,n4907,n4914);
xor (n4907,n4908,n4911);
or (n4908,n4909,n4910);
and (n4909,n3943,n3958);
and (n4910,n3944,n3947);
or (n4911,n4912,n4913);
and (n4912,n3995,n4117);
and (n4913,n3996,n4065);
xor (n4914,n4873,n4876);
and (n4915,n4908,n4911);
xor (n4916,n4868,n4871);
or (n4917,n4918,n4925);
and (n4918,n4919,n4924);
xor (n4919,n4920,n4921);
xor (n4920,n4852,n4855);
or (n4921,n4922,n4923);
and (n4922,n3886,n3918);
and (n4923,n3887,n3890);
xor (n4924,n4887,n4892);
and (n4925,n4920,n4921);
and (n4926,n4905,n4916);
and (n4927,n4900,n4901);
nor (n4928,n4929,n4930);
xor (n4929,n4899,n4902);
or (n4930,n4931,n4944);
and (n4931,n4932,n4935);
xor (n4932,n4933,n4934);
xor (n4933,n4883,n4894);
xor (n4934,n4904,n4917);
or (n4935,n4936,n4943);
and (n4936,n4937,n4942);
xor (n4937,n4938,n4941);
or (n4938,n4939,n4940);
and (n4939,n3922,n3994);
and (n4940,n3923,n3942);
xor (n4941,n4907,n4914);
xor (n4942,n4919,n4924);
and (n4943,n4938,n4941);
and (n4944,n4933,n4934);
nor (n4945,n4946,n4959);
nor (n4946,n4947,n4956);
xor (n4947,n4948,n4953);
xor (n4948,n4949,n4952);
or (n4949,n4950,n4951);
and (n4950,n3616,n3803);
and (n4951,n3617,n3758);
xor (n4952,n4937,n4942);
or (n4953,n4954,n4955);
and (n4954,n3884,n4120);
and (n4955,n3885,n3921);
or (n4956,n4957,n4958);
and (n4957,n3614,n3883);
and (n4958,n3615,n3874);
nor (n4959,n4960,n4961);
xor (n4960,n4932,n4935);
or (n4961,n4962,n4963);
and (n4962,n4948,n4953);
and (n4963,n4949,n4952);
nor (n4964,n4965,n5038);
nor (n4965,n4966,n4969);
or (n4966,n4967,n4968);
and (n4967,n4148,n4862);
and (n4968,n4149,n4669);
xor (n4969,n4970,n5035);
xor (n4970,n4971,n4974);
or (n4971,n4972,n4973);
and (n4972,n4150,n4607);
and (n4973,n4151,n4275);
xor (n4974,n4975,n5006);
xor (n4975,n4976,n5003);
xor (n4976,n4977,n5000);
xor (n4977,n4978,n4981);
or (n4978,n4979,n4980);
and (n4979,n4689,n4731);
and (n4980,n4690,n4708);
xor (n4981,n4982,n4989);
xor (n4982,n4983,n4986);
or (n4983,n4984,n4985);
and (n4984,n4709,n4728);
and (n4985,n4710,n4725);
or (n4986,n4987,n4988);
and (n4987,n4691,n4705);
and (n4988,n4692,n4702);
xor (n4989,n4990,n4997);
xor (n4990,n4991,n4994);
or (n4991,n4992,n4993);
and (n4992,n4243,n4254);
and (n4993,n4244,n4251);
or (n4994,n4995,n4996);
and (n4995,n4259,n4267);
and (n4996,n4260,n4264);
or (n4997,n4998,n4999);
and (n4998,n4618,n4625);
and (n4999,n4619,n4622);
or (n5000,n5001,n5002);
and (n5001,n4152,n4268);
and (n5002,n4153,n4239);
or (n5003,n5004,n5005);
and (n5004,n4672,n4740);
and (n5005,n4673,n4688);
xor (n5006,n5007,n5032);
xor (n5007,n5008,n5017);
xor (n5008,n5009,n5014);
xor (n5009,n5010,n5011);
xor (n5010,n912,n960);
or (n5011,n5012,n5013);
and (n5012,n4269,n4274);
and (n5013,n4270,n4273);
or (n5014,n5015,n5016);
and (n5015,n4240,n4258);
and (n5016,n4241,n4242);
xor (n5017,n5018,n5029);
xor (n5018,n5019,n5024);
xor (n5019,n5020,n5023);
xor (n5020,n5021,n5022);
xor (n5021,n227,n273);
xor (n5022,n93,n136);
xor (n5023,n168,n211);
xor (n5024,n5025,n5028);
xor (n5025,n5026,n5027);
xor (n5026,n428,n479);
xor (n5027,n365,n411);
xor (n5028,n306,n354);
or (n5029,n5030,n5031);
and (n5030,n4616,n4666);
and (n5031,n4617,n4629);
or (n5032,n5033,n5034);
and (n5033,n4608,n4615);
and (n5034,n4609,n4612);
or (n5035,n5036,n5037);
and (n5036,n4670,n4815);
and (n5037,n4671,n4787);
nor (n5038,n5039,n5042);
or (n5039,n5040,n5041);
and (n5040,n4970,n5035);
and (n5041,n4971,n4974);
xor (n5042,n5043,n5082);
xor (n5043,n5044,n5047);
or (n5044,n5045,n5046);
and (n5045,n5007,n5032);
and (n5046,n5008,n5017);
xor (n5047,n5048,n5061);
xor (n5048,n5049,n5058);
xor (n5049,n5050,n5055);
xor (n5050,n5051,n5052);
xor (n5051,n907,n910);
or (n5052,n5053,n5054);
and (n5053,n5009,n5014);
and (n5054,n5010,n5011);
or (n5055,n5056,n5057);
and (n5056,n4982,n4989);
and (n5057,n4983,n4986);
or (n5058,n5059,n5060);
and (n5059,n4977,n5000);
and (n5060,n4978,n4981);
xor (n5061,n5062,n5079);
xor (n5062,n5063,n5072);
xor (n5063,n5064,n5071);
xor (n5064,n5065,n5068);
or (n5065,n5066,n5067);
and (n5066,n5020,n5023);
and (n5067,n5021,n5022);
or (n5068,n5069,n5070);
and (n5069,n5025,n5028);
and (n5070,n5026,n5027);
xor (n5071,n624,n627);
xor (n5072,n5073,n5078);
xor (n5073,n5074,n5077);
or (n5074,n5075,n5076);
and (n5075,n4990,n4997);
and (n5076,n4991,n4994);
xor (n5077,n303,n426);
xor (n5078,n90,n225);
or (n5079,n5080,n5081);
and (n5080,n5018,n5029);
and (n5081,n5019,n5024);
or (n5082,n5083,n5084);
and (n5083,n4975,n5006);
and (n5084,n4976,n5003);
not (n5085,n5086);
nand (n5086,n5087,n5128);
nor (n5087,n5088,n5115);
nor (n5088,n5089,n5112);
xor (n5089,n5090,n5109);
xor (n5090,n5091,n5100);
xor (n5091,n5092,n5099);
xor (n5092,n5093,n5096);
or (n5093,n5094,n5095);
and (n5094,n5073,n5078);
and (n5095,n5074,n5077);
or (n5096,n5097,n5098);
and (n5097,n5064,n5071);
and (n5098,n5065,n5068);
xor (n5099,n497,n622);
xor (n5100,n5101,n5106);
xor (n5101,n5102,n5103);
xor (n5102,n903,n987);
or (n5103,n5104,n5105);
and (n5104,n5050,n5055);
and (n5105,n5051,n5052);
or (n5106,n5107,n5108);
and (n5107,n5062,n5079);
and (n5108,n5063,n5072);
or (n5109,n5110,n5111);
and (n5110,n5048,n5061);
and (n5111,n5049,n5058);
or (n5112,n5113,n5114);
and (n5113,n5043,n5082);
and (n5114,n5044,n5047);
nor (n5115,n5116,n5119);
or (n5116,n5117,n5118);
and (n5117,n5090,n5109);
and (n5118,n5091,n5100);
xor (n5119,n5120,n5125);
xor (n5120,n5121,n5124);
or (n5121,n5122,n5123);
and (n5122,n5092,n5099);
and (n5123,n5093,n5096);
xor (n5124,n899,n989);
or (n5125,n5126,n5127);
and (n5126,n5101,n5106);
and (n5127,n5102,n5103);
or (n5128,n5129,n5132);
or (n5129,n5130,n5131);
and (n5130,n5120,n5125);
and (n5131,n5121,n5124);
xor (n5132,n10,n897);
nand (n5133,n5134,n5085);
nand (n5134,n5135,n5154);
or (n5135,n5136,n5152);
not (n5136,n5137);
nand (n5137,n5138,n5145);
or (n5138,n5139,n5144);
not (n5139,n5140);
nand (n5140,n5141,n5143);
or (n5141,n3612,n5142);
nand (n5142,n4141,n4142);
nand (n5143,n3613,n4131);
not (n5144,n4945);
nand (n5145,n5146,n5151);
or (n5146,n5147,n5149);
not (n5147,n5148);
nand (n5148,n4960,n4961);
not (n5149,n5150);
nand (n5150,n4947,n4956);
not (n5151,n4959);
not (n5152,n5153);
and (n5153,n4145,n4964);
nor (n5154,n5155,n5164);
and (n5155,n5156,n4964);
not (n5156,n5157);
nand (n5157,n5158,n5163);
or (n5158,n5159,n5161);
not (n5159,n5160);
nand (n5160,n4929,n4930);
not (n5161,n5162);
nand (n5162,n4147,n4897);
not (n5163,n4146);
nand (n5164,n5165,n5167);
or (n5165,n5166,n5038);
nand (n5166,n4966,n4969);
nand (n5167,n5039,n5042);
nand (n5168,n5169,n5128);
or (n5169,n5170,n5174);
nand (n5170,n5171,n5173);
or (n5171,n5172,n5115);
nand (n5172,n5089,n5112);
nand (n5173,n5116,n5119);
and (n5174,n5129,n5132);
nand (n5175,n1087,n5);
not (n5176,n5177);
nor (n5177,n5178,n5180);
not (n5178,n5179);
or (n5181,n5177,n5182);
not (n5182,n5183);
or (n5184,n5185,n10415);
and (n5185,n5186,n5177);
xor (n5186,n5187,n10230);
xor (n5187,n5188,n8563);
xor (n5188,n5189,n8407);
xor (n5189,n5190,n6803);
xor (n5190,n5191,n6505);
xor (n5191,n5192,n6801);
xor (n5192,n5193,n6500);
xor (n5193,n5194,n6794);
xor (n5194,n5195,n3711);
xor (n5195,n5196,n6782);
xor (n5196,n5197,n4062);
xor (n5197,n5198,n6765);
xor (n5198,n5199,n4490);
xor (n5199,n5200,n6743);
xor (n5200,n5201,n6479);
xor (n5201,n5202,n6716);
xor (n5202,n5203,n6473);
xor (n5203,n5204,n6684);
xor (n5204,n5205,n6467);
xor (n5205,n5206,n6647);
xor (n5206,n5207,n6461);
xor (n5207,n5208,n6605);
xor (n5208,n5209,n6455);
xor (n5209,n5210,n6558);
xor (n5210,n5211,n6449);
xor (n5211,n5212,n6506);
xor (n5212,n5213,n6443);
xor (n5213,n5214,n6440);
xor (n5214,n5215,n6439);
xor (n5215,n5216,n6365);
xor (n5216,n5217,n6364);
xor (n5217,n5218,n6288);
xor (n5218,n5219,n6287);
xor (n5219,n5220,n6200);
xor (n5220,n5221,n6199);
or (n5221,n5222,n6113);
and (n5222,n5223,n6112);
or (n5223,n5224,n6023);
and (n5224,n5225,n6022);
or (n5225,n5226,n5938);
and (n5226,n5227,n565);
or (n5227,n5228,n5850);
and (n5228,n5229,n5849);
or (n5229,n5230,n5763);
and (n5230,n5231,n5762);
or (n5231,n5232,n5673);
and (n5232,n5233,n5672);
or (n5233,n5234,n5592);
and (n5234,n5235,n5591);
or (n5235,n5236,n5503);
and (n5236,n5237,n5502);
or (n5237,n5238,n5416);
and (n5238,n5239,n5415);
or (n5239,n5240,n5326);
and (n5240,n5241,n5325);
and (n5241,n1834,n5242);
or (n5242,n5243,n5245);
and (n5243,n5244,n1293);
and (n5244,n397,n1289);
and (n5245,n5246,n5247);
xor (n5246,n5244,n1293);
or (n5247,n5248,n5250);
and (n5248,n5249,n1297);
and (n5249,n466,n1289);
and (n5250,n5251,n5252);
xor (n5251,n5249,n1297);
or (n5252,n5253,n5256);
and (n5253,n5254,n5255);
and (n5254,n477,n1289);
and (n5255,n453,n1146);
and (n5256,n5257,n5258);
xor (n5257,n5254,n5255);
or (n5258,n5259,n5262);
and (n5259,n5260,n5261);
and (n5260,n453,n1289);
and (n5261,n434,n1146);
and (n5262,n5263,n5264);
xor (n5263,n5260,n5261);
or (n5264,n5265,n5268);
and (n5265,n5266,n5267);
and (n5266,n434,n1289);
and (n5267,n389,n1146);
and (n5268,n5269,n5270);
xor (n5269,n5266,n5267);
or (n5270,n5271,n5274);
and (n5271,n5272,n5273);
and (n5272,n389,n1289);
and (n5273,n371,n1146);
and (n5274,n5275,n5276);
xor (n5275,n5272,n5273);
or (n5276,n5277,n5280);
and (n5277,n5278,n5279);
and (n5278,n371,n1289);
and (n5279,n162,n1146);
and (n5280,n5281,n5282);
xor (n5281,n5278,n5279);
or (n5282,n5283,n5286);
and (n5283,n5284,n5285);
and (n5284,n162,n1289);
and (n5285,n156,n1146);
and (n5286,n5287,n5288);
xor (n5287,n5284,n5285);
or (n5288,n5289,n5291);
and (n5289,n5290,n2934);
and (n5290,n156,n1289);
and (n5291,n5292,n5293);
xor (n5292,n5290,n2934);
or (n5293,n5294,n5297);
and (n5294,n5295,n5296);
and (n5295,n935,n1289);
and (n5296,n1344,n1146);
and (n5297,n5298,n5299);
xor (n5298,n5295,n5296);
or (n5299,n5300,n5303);
and (n5300,n5301,n5302);
and (n5301,n1344,n1289);
and (n5302,n1215,n1146);
and (n5303,n5304,n5305);
xor (n5304,n5301,n5302);
or (n5305,n5306,n5309);
and (n5306,n5307,n5308);
and (n5307,n1215,n1289);
and (n5308,n1210,n1146);
and (n5309,n5310,n5311);
xor (n5310,n5307,n5308);
or (n5311,n5312,n5314);
and (n5312,n5313,n3430);
and (n5313,n1210,n1289);
and (n5314,n5315,n5316);
xor (n5315,n5313,n3430);
or (n5316,n5317,n5320);
and (n5317,n5318,n5319);
and (n5318,n1317,n1289);
and (n5319,n1323,n1146);
and (n5320,n5321,n5322);
xor (n5321,n5318,n5319);
and (n5322,n5323,n5324);
and (n5323,n1323,n1289);
and (n5324,n1463,n1146);
and (n5325,n397,n1142);
and (n5326,n5327,n5328);
xor (n5327,n5241,n5325);
or (n5328,n5329,n5332);
and (n5329,n5330,n5331);
xor (n5330,n1834,n5242);
and (n5331,n466,n1142);
and (n5332,n5333,n5334);
xor (n5333,n5330,n5331);
or (n5334,n5335,n5338);
and (n5335,n5336,n5337);
xor (n5336,n5246,n5247);
and (n5337,n477,n1142);
and (n5338,n5339,n5340);
xor (n5339,n5336,n5337);
or (n5340,n5341,n5344);
and (n5341,n5342,n5343);
xor (n5342,n5251,n5252);
and (n5343,n453,n1142);
and (n5344,n5345,n5346);
xor (n5345,n5342,n5343);
or (n5346,n5347,n5350);
and (n5347,n5348,n5349);
xor (n5348,n5257,n5258);
and (n5349,n434,n1142);
and (n5350,n5351,n5352);
xor (n5351,n5348,n5349);
or (n5352,n5353,n5356);
and (n5353,n5354,n5355);
xor (n5354,n5263,n5264);
and (n5355,n389,n1142);
and (n5356,n5357,n5358);
xor (n5357,n5354,n5355);
or (n5358,n5359,n5362);
and (n5359,n5360,n5361);
xor (n5360,n5269,n5270);
and (n5361,n371,n1142);
and (n5362,n5363,n5364);
xor (n5363,n5360,n5361);
or (n5364,n5365,n5368);
and (n5365,n5366,n5367);
xor (n5366,n5275,n5276);
and (n5367,n162,n1142);
and (n5368,n5369,n5370);
xor (n5369,n5366,n5367);
or (n5370,n5371,n5374);
and (n5371,n5372,n5373);
xor (n5372,n5281,n5282);
and (n5373,n156,n1142);
and (n5374,n5375,n5376);
xor (n5375,n5372,n5373);
or (n5376,n5377,n5380);
and (n5377,n5378,n5379);
xor (n5378,n5287,n5288);
and (n5379,n935,n1142);
and (n5380,n5381,n5382);
xor (n5381,n5378,n5379);
or (n5382,n5383,n5386);
and (n5383,n5384,n5385);
xor (n5384,n5292,n5293);
and (n5385,n1344,n1142);
and (n5386,n5387,n5388);
xor (n5387,n5384,n5385);
or (n5388,n5389,n5392);
and (n5389,n5390,n5391);
xor (n5390,n5298,n5299);
and (n5391,n1215,n1142);
and (n5392,n5393,n5394);
xor (n5393,n5390,n5391);
or (n5394,n5395,n5398);
and (n5395,n5396,n5397);
xor (n5396,n5304,n5305);
and (n5397,n1210,n1142);
and (n5398,n5399,n5400);
xor (n5399,n5396,n5397);
or (n5400,n5401,n5404);
and (n5401,n5402,n5403);
xor (n5402,n5310,n5311);
and (n5403,n1317,n1142);
and (n5404,n5405,n5406);
xor (n5405,n5402,n5403);
or (n5406,n5407,n5410);
and (n5407,n5408,n5409);
xor (n5408,n5315,n5316);
and (n5409,n1323,n1142);
and (n5410,n5411,n5412);
xor (n5411,n5408,n5409);
and (n5412,n5413,n5414);
xor (n5413,n5321,n5322);
not (n5414,n3412);
and (n5415,n397,n416);
and (n5416,n5417,n5418);
xor (n5417,n5239,n5415);
or (n5418,n5419,n5422);
and (n5419,n5420,n5421);
xor (n5420,n5327,n5328);
and (n5421,n466,n416);
and (n5422,n5423,n5424);
xor (n5423,n5420,n5421);
or (n5424,n5425,n5428);
and (n5425,n5426,n5427);
xor (n5426,n5333,n5334);
and (n5427,n477,n416);
and (n5428,n5429,n5430);
xor (n5429,n5426,n5427);
or (n5430,n5431,n5433);
and (n5431,n5432,n1152);
xor (n5432,n5339,n5340);
and (n5433,n5434,n5435);
xor (n5434,n5432,n1152);
or (n5435,n5436,n5439);
and (n5436,n5437,n5438);
xor (n5437,n5345,n5346);
and (n5438,n434,n416);
and (n5439,n5440,n5441);
xor (n5440,n5437,n5438);
or (n5441,n5442,n5444);
and (n5442,n5443,n2051);
xor (n5443,n5351,n5352);
and (n5444,n5445,n5446);
xor (n5445,n5443,n2051);
or (n5446,n5447,n5450);
and (n5447,n5448,n5449);
xor (n5448,n5357,n5358);
and (n5449,n371,n416);
and (n5450,n5451,n5452);
xor (n5451,n5448,n5449);
or (n5452,n5453,n5456);
and (n5453,n5454,n5455);
xor (n5454,n5363,n5364);
and (n5455,n162,n416);
and (n5456,n5457,n5458);
xor (n5457,n5454,n5455);
or (n5458,n5459,n5461);
and (n5459,n5460,n2455);
xor (n5460,n5369,n5370);
and (n5461,n5462,n5463);
xor (n5462,n5460,n2455);
or (n5463,n5464,n5467);
and (n5464,n5465,n5466);
xor (n5465,n5375,n5376);
and (n5466,n935,n416);
and (n5467,n5468,n5469);
xor (n5468,n5465,n5466);
or (n5469,n5470,n5473);
and (n5470,n5471,n5472);
xor (n5471,n5381,n5382);
and (n5472,n1344,n416);
and (n5473,n5474,n5475);
xor (n5474,n5471,n5472);
or (n5475,n5476,n5479);
and (n5476,n5477,n5478);
xor (n5477,n5387,n5388);
and (n5478,n1215,n416);
and (n5479,n5480,n5481);
xor (n5480,n5477,n5478);
or (n5481,n5482,n5485);
and (n5482,n5483,n5484);
xor (n5483,n5393,n5394);
and (n5484,n1210,n416);
and (n5485,n5486,n5487);
xor (n5486,n5483,n5484);
or (n5487,n5488,n5491);
and (n5488,n5489,n5490);
xor (n5489,n5399,n5400);
and (n5490,n1317,n416);
and (n5491,n5492,n5493);
xor (n5492,n5489,n5490);
or (n5493,n5494,n5497);
and (n5494,n5495,n5496);
xor (n5495,n5405,n5406);
and (n5496,n1323,n416);
and (n5497,n5498,n5499);
xor (n5498,n5495,n5496);
and (n5499,n5500,n5501);
xor (n5500,n5411,n5412);
and (n5501,n1463,n416);
and (n5502,n397,n417);
and (n5503,n5504,n5505);
xor (n5504,n5237,n5502);
or (n5505,n5506,n5509);
and (n5506,n5507,n5508);
xor (n5507,n5417,n5418);
and (n5508,n466,n417);
and (n5509,n5510,n5511);
xor (n5510,n5507,n5508);
or (n5511,n5512,n5515);
and (n5512,n5513,n5514);
xor (n5513,n5423,n5424);
and (n5514,n477,n417);
and (n5515,n5516,n5517);
xor (n5516,n5513,n5514);
or (n5517,n5518,n5521);
and (n5518,n5519,n5520);
xor (n5519,n5429,n5430);
and (n5520,n453,n417);
and (n5521,n5522,n5523);
xor (n5522,n5519,n5520);
or (n5523,n5524,n5527);
and (n5524,n5525,n5526);
xor (n5525,n5434,n5435);
and (n5526,n434,n417);
and (n5527,n5528,n5529);
xor (n5528,n5525,n5526);
or (n5529,n5530,n5533);
and (n5530,n5531,n5532);
xor (n5531,n5440,n5441);
and (n5532,n389,n417);
and (n5533,n5534,n5535);
xor (n5534,n5531,n5532);
or (n5535,n5536,n5539);
and (n5536,n5537,n5538);
xor (n5537,n5445,n5446);
and (n5538,n371,n417);
and (n5539,n5540,n5541);
xor (n5540,n5537,n5538);
or (n5541,n5542,n5545);
and (n5542,n5543,n5544);
xor (n5543,n5451,n5452);
and (n5544,n162,n417);
and (n5545,n5546,n5547);
xor (n5546,n5543,n5544);
or (n5547,n5548,n5551);
and (n5548,n5549,n5550);
xor (n5549,n5457,n5458);
and (n5550,n156,n417);
and (n5551,n5552,n5553);
xor (n5552,n5549,n5550);
or (n5553,n5554,n5557);
and (n5554,n5555,n5556);
xor (n5555,n5462,n5463);
and (n5556,n935,n417);
and (n5557,n5558,n5559);
xor (n5558,n5555,n5556);
or (n5559,n5560,n5563);
and (n5560,n5561,n5562);
xor (n5561,n5468,n5469);
and (n5562,n1344,n417);
and (n5563,n5564,n5565);
xor (n5564,n5561,n5562);
or (n5565,n5566,n5569);
and (n5566,n5567,n5568);
xor (n5567,n5474,n5475);
and (n5568,n1215,n417);
and (n5569,n5570,n5571);
xor (n5570,n5567,n5568);
or (n5571,n5572,n5575);
and (n5572,n5573,n5574);
xor (n5573,n5480,n5481);
and (n5574,n1210,n417);
and (n5575,n5576,n5577);
xor (n5576,n5573,n5574);
or (n5577,n5578,n5581);
and (n5578,n5579,n5580);
xor (n5579,n5486,n5487);
and (n5580,n1317,n417);
and (n5581,n5582,n5583);
xor (n5582,n5579,n5580);
or (n5583,n5584,n5587);
and (n5584,n5585,n5586);
xor (n5585,n5492,n5493);
and (n5586,n1323,n417);
and (n5587,n5588,n5589);
xor (n5588,n5585,n5586);
and (n5589,n5590,n3147);
xor (n5590,n5498,n5499);
and (n5591,n397,n407);
and (n5592,n5593,n5594);
xor (n5593,n5235,n5591);
or (n5594,n5595,n5598);
and (n5595,n5596,n5597);
xor (n5596,n5504,n5505);
and (n5597,n466,n407);
and (n5598,n5599,n5600);
xor (n5599,n5596,n5597);
or (n5600,n5601,n5604);
and (n5601,n5602,n5603);
xor (n5602,n5510,n5511);
and (n5603,n477,n407);
and (n5604,n5605,n5606);
xor (n5605,n5602,n5603);
or (n5606,n5607,n5609);
and (n5607,n5608,n3639);
xor (n5608,n5516,n5517);
and (n5609,n5610,n5611);
xor (n5610,n5608,n3639);
or (n5611,n5612,n5614);
and (n5612,n5613,n1694);
xor (n5613,n5522,n5523);
and (n5614,n5615,n5616);
xor (n5615,n5613,n1694);
or (n5616,n5617,n5620);
and (n5617,n5618,n5619);
xor (n5618,n5528,n5529);
and (n5619,n389,n407);
and (n5620,n5621,n5622);
xor (n5621,n5618,n5619);
or (n5622,n5623,n5625);
and (n5623,n5624,n1271);
xor (n5624,n5534,n5535);
and (n5625,n5626,n5627);
xor (n5626,n5624,n1271);
or (n5627,n5628,n5630);
and (n5628,n5629,n2081);
xor (n5629,n5540,n5541);
and (n5630,n5631,n5632);
xor (n5631,n5629,n2081);
or (n5632,n5633,n5636);
and (n5633,n5634,n5635);
xor (n5634,n5546,n5547);
and (n5635,n156,n407);
and (n5636,n5637,n5638);
xor (n5637,n5634,n5635);
or (n5638,n5639,n5641);
and (n5639,n5640,n1389);
xor (n5640,n5552,n5553);
and (n5641,n5642,n5643);
xor (n5642,n5640,n1389);
or (n5643,n5644,n5646);
and (n5644,n5645,n2333);
xor (n5645,n5558,n5559);
and (n5646,n5647,n5648);
xor (n5647,n5645,n2333);
or (n5648,n5649,n5652);
and (n5649,n5650,n5651);
xor (n5650,n5564,n5565);
and (n5651,n1215,n407);
and (n5652,n5653,n5654);
xor (n5653,n5650,n5651);
or (n5654,n5655,n5657);
and (n5655,n5656,n2745);
xor (n5656,n5570,n5571);
and (n5657,n5658,n5659);
xor (n5658,n5656,n2745);
or (n5659,n5660,n5662);
and (n5660,n5661,n2874);
xor (n5661,n5576,n5577);
and (n5662,n5663,n5664);
xor (n5663,n5661,n2874);
or (n5664,n5665,n5667);
and (n5665,n5666,n3038);
xor (n5666,n5582,n5583);
and (n5667,n5668,n5669);
xor (n5668,n5666,n3038);
and (n5669,n5670,n5671);
xor (n5670,n5588,n5589);
and (n5671,n1463,n407);
and (n5672,n397,n404);
and (n5673,n5674,n5675);
xor (n5674,n5233,n5672);
or (n5675,n5676,n5679);
and (n5676,n5677,n5678);
xor (n5677,n5593,n5594);
and (n5678,n466,n404);
and (n5679,n5680,n5681);
xor (n5680,n5677,n5678);
or (n5681,n5682,n5685);
and (n5682,n5683,n5684);
xor (n5683,n5599,n5600);
and (n5684,n477,n404);
and (n5685,n5686,n5687);
xor (n5686,n5683,n5684);
or (n5687,n5688,n5691);
and (n5688,n5689,n5690);
xor (n5689,n5605,n5606);
and (n5690,n453,n404);
and (n5691,n5692,n5693);
xor (n5692,n5689,n5690);
or (n5693,n5694,n5697);
and (n5694,n5695,n5696);
xor (n5695,n5610,n5611);
and (n5696,n434,n404);
and (n5697,n5698,n5699);
xor (n5698,n5695,n5696);
or (n5699,n5700,n5703);
and (n5700,n5701,n5702);
xor (n5701,n5615,n5616);
and (n5702,n389,n404);
and (n5703,n5704,n5705);
xor (n5704,n5701,n5702);
or (n5705,n5706,n5709);
and (n5706,n5707,n5708);
xor (n5707,n5621,n5622);
and (n5708,n371,n404);
and (n5709,n5710,n5711);
xor (n5710,n5707,n5708);
or (n5711,n5712,n5715);
and (n5712,n5713,n5714);
xor (n5713,n5626,n5627);
and (n5714,n162,n404);
and (n5715,n5716,n5717);
xor (n5716,n5713,n5714);
or (n5717,n5718,n5721);
and (n5718,n5719,n5720);
xor (n5719,n5631,n5632);
and (n5720,n156,n404);
and (n5721,n5722,n5723);
xor (n5722,n5719,n5720);
or (n5723,n5724,n5727);
and (n5724,n5725,n5726);
xor (n5725,n5637,n5638);
and (n5726,n935,n404);
and (n5727,n5728,n5729);
xor (n5728,n5725,n5726);
or (n5729,n5730,n5733);
and (n5730,n5731,n5732);
xor (n5731,n5642,n5643);
and (n5732,n1344,n404);
and (n5733,n5734,n5735);
xor (n5734,n5731,n5732);
or (n5735,n5736,n5739);
and (n5736,n5737,n5738);
xor (n5737,n5647,n5648);
and (n5738,n1215,n404);
and (n5739,n5740,n5741);
xor (n5740,n5737,n5738);
or (n5741,n5742,n5745);
and (n5742,n5743,n5744);
xor (n5743,n5653,n5654);
and (n5744,n1210,n404);
and (n5745,n5746,n5747);
xor (n5746,n5743,n5744);
or (n5747,n5748,n5751);
and (n5748,n5749,n5750);
xor (n5749,n5658,n5659);
and (n5750,n1317,n404);
and (n5751,n5752,n5753);
xor (n5752,n5749,n5750);
or (n5753,n5754,n5757);
and (n5754,n5755,n5756);
xor (n5755,n5663,n5664);
and (n5756,n1323,n404);
and (n5757,n5758,n5759);
xor (n5758,n5755,n5756);
and (n5759,n5760,n5761);
xor (n5760,n5668,n5669);
not (n5761,n2857);
and (n5762,n397,n396);
and (n5763,n5764,n5765);
xor (n5764,n5231,n5762);
or (n5765,n5766,n5769);
and (n5766,n5767,n5768);
xor (n5767,n5674,n5675);
and (n5768,n466,n396);
and (n5769,n5770,n5771);
xor (n5770,n5767,n5768);
or (n5771,n5772,n5774);
and (n5772,n5773,n4227);
xor (n5773,n5680,n5681);
and (n5774,n5775,n5776);
xor (n5775,n5773,n4227);
or (n5776,n5777,n5780);
and (n5777,n5778,n5779);
xor (n5778,n5686,n5687);
and (n5779,n453,n396);
and (n5780,n5781,n5782);
xor (n5781,n5778,n5779);
or (n5782,n5783,n5786);
and (n5783,n5784,n5785);
xor (n5784,n5692,n5693);
and (n5785,n434,n396);
and (n5786,n5787,n5788);
xor (n5787,n5784,n5785);
or (n5788,n5789,n5792);
and (n5789,n5790,n5791);
xor (n5790,n5698,n5699);
and (n5791,n389,n396);
and (n5792,n5793,n5794);
xor (n5793,n5790,n5791);
or (n5794,n5795,n5798);
and (n5795,n5796,n5797);
xor (n5796,n5704,n5705);
and (n5797,n371,n396);
and (n5798,n5799,n5800);
xor (n5799,n5796,n5797);
or (n5800,n5801,n5804);
and (n5801,n5802,n5803);
xor (n5802,n5710,n5711);
and (n5803,n162,n396);
and (n5804,n5805,n5806);
xor (n5805,n5802,n5803);
or (n5806,n5807,n5810);
and (n5807,n5808,n5809);
xor (n5808,n5716,n5717);
and (n5809,n156,n396);
and (n5810,n5811,n5812);
xor (n5811,n5808,n5809);
or (n5812,n5813,n5816);
and (n5813,n5814,n5815);
xor (n5814,n5722,n5723);
and (n5815,n935,n396);
and (n5816,n5817,n5818);
xor (n5817,n5814,n5815);
or (n5818,n5819,n5821);
and (n5819,n5820,n1577);
xor (n5820,n5728,n5729);
and (n5821,n5822,n5823);
xor (n5822,n5820,n1577);
or (n5823,n5824,n5826);
and (n5824,n5825,n2147);
xor (n5825,n5734,n5735);
and (n5826,n5827,n5828);
xor (n5827,n5825,n2147);
or (n5828,n5829,n5832);
and (n5829,n5830,n5831);
xor (n5830,n5740,n5741);
and (n5831,n1210,n396);
and (n5832,n5833,n5834);
xor (n5833,n5830,n5831);
or (n5834,n5835,n5838);
and (n5835,n5836,n5837);
xor (n5836,n5746,n5747);
and (n5837,n1317,n396);
and (n5838,n5839,n5840);
xor (n5839,n5836,n5837);
or (n5840,n5841,n5844);
and (n5841,n5842,n5843);
xor (n5842,n5752,n5753);
and (n5843,n1323,n396);
and (n5844,n5845,n5846);
xor (n5845,n5842,n5843);
and (n5846,n5847,n5848);
xor (n5847,n5758,n5759);
and (n5848,n1463,n396);
and (n5849,n397,n459);
and (n5850,n5851,n5852);
xor (n5851,n5229,n5849);
or (n5852,n5853,n5856);
and (n5853,n5854,n5855);
xor (n5854,n5764,n5765);
and (n5855,n466,n459);
and (n5856,n5857,n5858);
xor (n5857,n5854,n5855);
or (n5858,n5859,n5862);
and (n5859,n5860,n5861);
xor (n5860,n5770,n5771);
and (n5861,n477,n459);
and (n5862,n5863,n5864);
xor (n5863,n5860,n5861);
or (n5864,n5865,n5868);
and (n5865,n5866,n5867);
xor (n5866,n5775,n5776);
and (n5867,n453,n459);
and (n5868,n5869,n5870);
xor (n5869,n5866,n5867);
or (n5870,n5871,n5874);
and (n5871,n5872,n5873);
xor (n5872,n5781,n5782);
and (n5873,n434,n459);
and (n5874,n5875,n5876);
xor (n5875,n5872,n5873);
or (n5876,n5877,n5880);
and (n5877,n5878,n5879);
xor (n5878,n5787,n5788);
and (n5879,n389,n459);
and (n5880,n5881,n5882);
xor (n5881,n5878,n5879);
or (n5882,n5883,n5886);
and (n5883,n5884,n5885);
xor (n5884,n5793,n5794);
and (n5885,n371,n459);
and (n5886,n5887,n5888);
xor (n5887,n5884,n5885);
or (n5888,n5889,n5892);
and (n5889,n5890,n5891);
xor (n5890,n5799,n5800);
and (n5891,n162,n459);
and (n5892,n5893,n5894);
xor (n5893,n5890,n5891);
or (n5894,n5895,n5898);
and (n5895,n5896,n5897);
xor (n5896,n5805,n5806);
and (n5897,n156,n459);
and (n5898,n5899,n5900);
xor (n5899,n5896,n5897);
or (n5900,n5901,n5904);
and (n5901,n5902,n5903);
xor (n5902,n5811,n5812);
and (n5903,n935,n459);
and (n5904,n5905,n5906);
xor (n5905,n5902,n5903);
or (n5906,n5907,n5910);
and (n5907,n5908,n5909);
xor (n5908,n5817,n5818);
and (n5909,n1344,n459);
and (n5910,n5911,n5912);
xor (n5911,n5908,n5909);
or (n5912,n5913,n5916);
and (n5913,n5914,n5915);
xor (n5914,n5822,n5823);
and (n5915,n1215,n459);
and (n5916,n5917,n5918);
xor (n5917,n5914,n5915);
or (n5918,n5919,n5922);
and (n5919,n5920,n5921);
xor (n5920,n5827,n5828);
and (n5921,n1210,n459);
and (n5922,n5923,n5924);
xor (n5923,n5920,n5921);
or (n5924,n5925,n5928);
and (n5925,n5926,n5927);
xor (n5926,n5833,n5834);
and (n5927,n1317,n459);
and (n5928,n5929,n5930);
xor (n5929,n5926,n5927);
or (n5930,n5931,n5934);
and (n5931,n5932,n5933);
xor (n5932,n5839,n5840);
and (n5933,n1323,n459);
and (n5934,n5935,n5936);
xor (n5935,n5932,n5933);
and (n5936,n5937,n2590);
xor (n5937,n5845,n5846);
and (n5938,n5939,n5940);
xor (n5939,n5227,n565);
or (n5940,n5941,n5943);
and (n5941,n5942,n467);
xor (n5942,n5851,n5852);
and (n5943,n5944,n5945);
xor (n5944,n5942,n467);
or (n5945,n5946,n5948);
and (n5946,n5947,n478);
xor (n5947,n5857,n5858);
and (n5948,n5949,n5950);
xor (n5949,n5947,n478);
or (n5950,n5951,n5954);
and (n5951,n5952,n5953);
xor (n5952,n5863,n5864);
and (n5953,n453,n441);
and (n5954,n5955,n5956);
xor (n5955,n5952,n5953);
or (n5956,n5957,n5960);
and (n5957,n5958,n5959);
xor (n5958,n5869,n5870);
and (n5959,n434,n441);
and (n5960,n5961,n5962);
xor (n5961,n5958,n5959);
or (n5962,n5963,n5966);
and (n5963,n5964,n5965);
xor (n5964,n5875,n5876);
and (n5965,n389,n441);
and (n5966,n5967,n5968);
xor (n5967,n5964,n5965);
or (n5968,n5969,n5972);
and (n5969,n5970,n5971);
xor (n5970,n5881,n5882);
and (n5971,n371,n441);
and (n5972,n5973,n5974);
xor (n5973,n5970,n5971);
or (n5974,n5975,n5977);
and (n5975,n5976,n3705);
xor (n5976,n5887,n5888);
and (n5977,n5978,n5979);
xor (n5978,n5976,n3705);
or (n5979,n5980,n5983);
and (n5980,n5981,n5982);
xor (n5981,n5893,n5894);
and (n5982,n156,n441);
and (n5983,n5984,n5985);
xor (n5984,n5981,n5982);
or (n5985,n5986,n5988);
and (n5986,n5987,n1350);
xor (n5987,n5899,n5900);
and (n5988,n5989,n5990);
xor (n5989,n5987,n1350);
or (n5990,n5991,n5994);
and (n5991,n5992,n5993);
xor (n5992,n5905,n5906);
and (n5993,n1344,n441);
and (n5994,n5995,n5996);
xor (n5995,n5992,n5993);
or (n5996,n5997,n5999);
and (n5997,n5998,n2091);
xor (n5998,n5911,n5912);
and (n5999,n6000,n6001);
xor (n6000,n5998,n2091);
or (n6001,n6002,n6005);
and (n6002,n6003,n6004);
xor (n6003,n5917,n5918);
and (n6004,n1210,n441);
and (n6005,n6006,n6007);
xor (n6006,n6003,n6004);
or (n6007,n6008,n6011);
and (n6008,n6009,n6010);
xor (n6009,n5923,n5924);
and (n6010,n1317,n441);
and (n6011,n6012,n6013);
xor (n6012,n6009,n6010);
or (n6013,n6014,n6017);
and (n6014,n6015,n6016);
xor (n6015,n5929,n5930);
and (n6016,n1323,n441);
and (n6017,n6018,n6019);
xor (n6018,n6015,n6016);
and (n6019,n6020,n6021);
xor (n6020,n5935,n5936);
and (n6021,n1463,n441);
and (n6022,n397,n442);
and (n6023,n6024,n6025);
xor (n6024,n5225,n6022);
or (n6025,n6026,n6029);
and (n6026,n6027,n6028);
xor (n6027,n5939,n5940);
and (n6028,n466,n442);
and (n6029,n6030,n6031);
xor (n6030,n6027,n6028);
or (n6031,n6032,n6035);
and (n6032,n6033,n6034);
xor (n6033,n5944,n5945);
and (n6034,n477,n442);
and (n6035,n6036,n6037);
xor (n6036,n6033,n6034);
or (n6037,n6038,n6041);
and (n6038,n6039,n6040);
xor (n6039,n5949,n5950);
and (n6040,n453,n442);
and (n6041,n6042,n6043);
xor (n6042,n6039,n6040);
or (n6043,n6044,n6047);
and (n6044,n6045,n6046);
xor (n6045,n5955,n5956);
and (n6046,n434,n442);
and (n6047,n6048,n6049);
xor (n6048,n6045,n6046);
or (n6049,n6050,n6053);
and (n6050,n6051,n6052);
xor (n6051,n5961,n5962);
and (n6052,n389,n442);
and (n6053,n6054,n6055);
xor (n6054,n6051,n6052);
or (n6055,n6056,n6059);
and (n6056,n6057,n6058);
xor (n6057,n5967,n5968);
and (n6058,n371,n442);
and (n6059,n6060,n6061);
xor (n6060,n6057,n6058);
or (n6061,n6062,n6065);
and (n6062,n6063,n6064);
xor (n6063,n5973,n5974);
and (n6064,n162,n442);
and (n6065,n6066,n6067);
xor (n6066,n6063,n6064);
or (n6067,n6068,n6071);
and (n6068,n6069,n6070);
xor (n6069,n5978,n5979);
and (n6070,n156,n442);
and (n6071,n6072,n6073);
xor (n6072,n6069,n6070);
or (n6073,n6074,n6077);
and (n6074,n6075,n6076);
xor (n6075,n5984,n5985);
and (n6076,n935,n442);
and (n6077,n6078,n6079);
xor (n6078,n6075,n6076);
or (n6079,n6080,n6083);
and (n6080,n6081,n6082);
xor (n6081,n5989,n5990);
and (n6082,n1344,n442);
and (n6083,n6084,n6085);
xor (n6084,n6081,n6082);
or (n6085,n6086,n6089);
and (n6086,n6087,n6088);
xor (n6087,n5995,n5996);
and (n6088,n1215,n442);
and (n6089,n6090,n6091);
xor (n6090,n6087,n6088);
or (n6091,n6092,n6095);
and (n6092,n6093,n6094);
xor (n6093,n6000,n6001);
and (n6094,n1210,n442);
and (n6095,n6096,n6097);
xor (n6096,n6093,n6094);
or (n6097,n6098,n6101);
and (n6098,n6099,n6100);
xor (n6099,n6006,n6007);
and (n6100,n1317,n442);
and (n6101,n6102,n6103);
xor (n6102,n6099,n6100);
or (n6103,n6104,n6107);
and (n6104,n6105,n6106);
xor (n6105,n6012,n6013);
and (n6106,n1323,n442);
and (n6107,n6108,n6109);
xor (n6108,n6105,n6106);
and (n6109,n6110,n6111);
xor (n6110,n6018,n6019);
not (n6111,n1500);
and (n6112,n397,n383);
and (n6113,n6114,n6115);
xor (n6114,n5223,n6112);
or (n6115,n6116,n6119);
and (n6116,n6117,n6118);
xor (n6117,n6024,n6025);
and (n6118,n466,n383);
and (n6119,n6120,n6121);
xor (n6120,n6117,n6118);
or (n6121,n6122,n6125);
and (n6122,n6123,n6124);
xor (n6123,n6030,n6031);
and (n6124,n477,n383);
and (n6125,n6126,n6127);
xor (n6126,n6123,n6124);
or (n6127,n6128,n6130);
and (n6128,n6129,n454);
xor (n6129,n6036,n6037);
and (n6130,n6131,n6132);
xor (n6131,n6129,n454);
or (n6132,n6133,n6136);
and (n6133,n6134,n6135);
xor (n6134,n6042,n6043);
and (n6135,n434,n383);
and (n6136,n6137,n6138);
xor (n6137,n6134,n6135);
or (n6138,n6139,n6141);
and (n6139,n6140,n4249);
xor (n6140,n6048,n6049);
and (n6141,n6142,n6143);
xor (n6142,n6140,n4249);
or (n6143,n6144,n6146);
and (n6144,n6145,n4292);
xor (n6145,n6054,n6055);
and (n6146,n6147,n6148);
xor (n6147,n6145,n4292);
or (n6148,n6149,n6152);
and (n6149,n6150,n6151);
xor (n6150,n6060,n6061);
and (n6151,n162,n383);
and (n6152,n6153,n6154);
xor (n6153,n6150,n6151);
or (n6154,n6155,n6158);
and (n6155,n6156,n6157);
xor (n6156,n6066,n6067);
and (n6157,n156,n383);
and (n6158,n6159,n6160);
xor (n6159,n6156,n6157);
or (n6160,n6161,n6164);
and (n6161,n6162,n6163);
xor (n6162,n6072,n6073);
and (n6163,n935,n383);
and (n6164,n6165,n6166);
xor (n6165,n6162,n6163);
or (n6166,n6167,n6170);
and (n6167,n6168,n6169);
xor (n6168,n6078,n6079);
and (n6169,n1344,n383);
and (n6170,n6171,n6172);
xor (n6171,n6168,n6169);
or (n6172,n6173,n6176);
and (n6173,n6174,n6175);
xor (n6174,n6084,n6085);
and (n6175,n1215,n383);
and (n6176,n6177,n6178);
xor (n6177,n6174,n6175);
or (n6178,n6179,n6182);
and (n6179,n6180,n6181);
xor (n6180,n6090,n6091);
and (n6181,n1210,n383);
and (n6182,n6183,n6184);
xor (n6183,n6180,n6181);
or (n6184,n6185,n6188);
and (n6185,n6186,n6187);
xor (n6186,n6096,n6097);
and (n6187,n1317,n383);
and (n6188,n6189,n6190);
xor (n6189,n6186,n6187);
or (n6190,n6191,n6194);
and (n6191,n6192,n6193);
xor (n6192,n6102,n6103);
and (n6193,n1323,n383);
and (n6194,n6195,n6196);
xor (n6195,n6192,n6193);
and (n6196,n6197,n6198);
xor (n6197,n6108,n6109);
and (n6198,n1463,n383);
and (n6199,n397,n378);
or (n6200,n6201,n6204);
and (n6201,n6202,n6203);
xor (n6202,n6114,n6115);
and (n6203,n466,n378);
and (n6204,n6205,n6206);
xor (n6205,n6202,n6203);
or (n6206,n6207,n6210);
and (n6207,n6208,n6209);
xor (n6208,n6120,n6121);
and (n6209,n477,n378);
and (n6210,n6211,n6212);
xor (n6211,n6208,n6209);
or (n6212,n6213,n6216);
and (n6213,n6214,n6215);
xor (n6214,n6126,n6127);
and (n6215,n453,n378);
and (n6216,n6217,n6218);
xor (n6217,n6214,n6215);
or (n6218,n6219,n6222);
and (n6219,n6220,n6221);
xor (n6220,n6131,n6132);
and (n6221,n434,n378);
and (n6222,n6223,n6224);
xor (n6223,n6220,n6221);
or (n6224,n6225,n6228);
and (n6225,n6226,n6227);
xor (n6226,n6137,n6138);
and (n6227,n389,n378);
and (n6228,n6229,n6230);
xor (n6229,n6226,n6227);
or (n6230,n6231,n6234);
and (n6231,n6232,n6233);
xor (n6232,n6142,n6143);
and (n6233,n371,n378);
and (n6234,n6235,n6236);
xor (n6235,n6232,n6233);
or (n6236,n6237,n6240);
and (n6237,n6238,n6239);
xor (n6238,n6147,n6148);
and (n6239,n162,n378);
and (n6240,n6241,n6242);
xor (n6241,n6238,n6239);
or (n6242,n6243,n6246);
and (n6243,n6244,n6245);
xor (n6244,n6153,n6154);
and (n6245,n156,n378);
and (n6246,n6247,n6248);
xor (n6247,n6244,n6245);
or (n6248,n6249,n6252);
and (n6249,n6250,n6251);
xor (n6250,n6159,n6160);
and (n6251,n935,n378);
and (n6252,n6253,n6254);
xor (n6253,n6250,n6251);
or (n6254,n6255,n6258);
and (n6255,n6256,n6257);
xor (n6256,n6165,n6166);
and (n6257,n1344,n378);
and (n6258,n6259,n6260);
xor (n6259,n6256,n6257);
or (n6260,n6261,n6264);
and (n6261,n6262,n6263);
xor (n6262,n6171,n6172);
and (n6263,n1215,n378);
and (n6264,n6265,n6266);
xor (n6265,n6262,n6263);
or (n6266,n6267,n6270);
and (n6267,n6268,n6269);
xor (n6268,n6177,n6178);
and (n6269,n1210,n378);
and (n6270,n6271,n6272);
xor (n6271,n6268,n6269);
or (n6272,n6273,n6276);
and (n6273,n6274,n6275);
xor (n6274,n6183,n6184);
and (n6275,n1317,n378);
and (n6276,n6277,n6278);
xor (n6277,n6274,n6275);
or (n6278,n6279,n6282);
and (n6279,n6280,n6281);
xor (n6280,n6189,n6190);
and (n6281,n1323,n378);
and (n6282,n6283,n6284);
xor (n6283,n6280,n6281);
and (n6284,n6285,n6286);
xor (n6285,n6195,n6196);
not (n6286,n1561);
and (n6287,n466,n151);
or (n6288,n6289,n6292);
and (n6289,n6290,n6291);
xor (n6290,n6205,n6206);
and (n6291,n477,n151);
and (n6292,n6293,n6294);
xor (n6293,n6290,n6291);
or (n6294,n6295,n6298);
and (n6295,n6296,n6297);
xor (n6296,n6211,n6212);
and (n6297,n453,n151);
and (n6298,n6299,n6300);
xor (n6299,n6296,n6297);
or (n6300,n6301,n6304);
and (n6301,n6302,n6303);
xor (n6302,n6217,n6218);
and (n6303,n434,n151);
and (n6304,n6305,n6306);
xor (n6305,n6302,n6303);
or (n6306,n6307,n6309);
and (n6307,n6308,n390);
xor (n6308,n6223,n6224);
and (n6309,n6310,n6311);
xor (n6310,n6308,n390);
or (n6311,n6312,n6315);
and (n6312,n6313,n6314);
xor (n6313,n6229,n6230);
and (n6314,n371,n151);
and (n6315,n6316,n6317);
xor (n6316,n6313,n6314);
or (n6317,n6318,n6320);
and (n6318,n6319,n4171);
xor (n6319,n6235,n6236);
and (n6320,n6321,n6322);
xor (n6321,n6319,n4171);
or (n6322,n6323,n6325);
and (n6323,n6324,n4167);
xor (n6324,n6241,n6242);
and (n6325,n6326,n6327);
xor (n6326,n6324,n4167);
or (n6327,n6328,n6330);
and (n6328,n6329,n4521);
xor (n6329,n6247,n6248);
and (n6330,n6331,n6332);
xor (n6331,n6329,n4521);
or (n6332,n6333,n6336);
and (n6333,n6334,n6335);
xor (n6334,n6253,n6254);
and (n6335,n1344,n151);
and (n6336,n6337,n6338);
xor (n6337,n6334,n6335);
or (n6338,n6339,n6342);
and (n6339,n6340,n6341);
xor (n6340,n6259,n6260);
and (n6341,n1215,n151);
and (n6342,n6343,n6344);
xor (n6343,n6340,n6341);
or (n6344,n6345,n6347);
and (n6345,n6346,n1743);
xor (n6346,n6265,n6266);
and (n6347,n6348,n6349);
xor (n6348,n6346,n1743);
or (n6349,n6350,n6353);
and (n6350,n6351,n6352);
xor (n6351,n6271,n6272);
and (n6352,n1317,n151);
and (n6353,n6354,n6355);
xor (n6354,n6351,n6352);
or (n6355,n6356,n6359);
and (n6356,n6357,n6358);
xor (n6357,n6277,n6278);
and (n6358,n1323,n151);
and (n6359,n6360,n6361);
xor (n6360,n6357,n6358);
and (n6361,n6362,n6363);
xor (n6362,n6283,n6284);
and (n6363,n1463,n151);
and (n6364,n477,n143);
or (n6365,n6366,n6369);
and (n6366,n6367,n6368);
xor (n6367,n6293,n6294);
and (n6368,n453,n143);
and (n6369,n6370,n6371);
xor (n6370,n6367,n6368);
or (n6371,n6372,n6375);
and (n6372,n6373,n6374);
xor (n6373,n6299,n6300);
and (n6374,n434,n143);
and (n6375,n6376,n6377);
xor (n6376,n6373,n6374);
or (n6377,n6378,n6381);
and (n6378,n6379,n6380);
xor (n6379,n6305,n6306);
and (n6380,n389,n143);
and (n6381,n6382,n6383);
xor (n6382,n6379,n6380);
or (n6383,n6384,n6387);
and (n6384,n6385,n6386);
xor (n6385,n6310,n6311);
and (n6386,n371,n143);
and (n6387,n6388,n6389);
xor (n6388,n6385,n6386);
or (n6389,n6390,n6393);
and (n6390,n6391,n6392);
xor (n6391,n6316,n6317);
and (n6392,n162,n143);
and (n6393,n6394,n6395);
xor (n6394,n6391,n6392);
or (n6395,n6396,n6399);
and (n6396,n6397,n6398);
xor (n6397,n6321,n6322);
and (n6398,n156,n143);
and (n6399,n6400,n6401);
xor (n6400,n6397,n6398);
or (n6401,n6402,n6405);
and (n6402,n6403,n6404);
xor (n6403,n6326,n6327);
and (n6404,n935,n143);
and (n6405,n6406,n6407);
xor (n6406,n6403,n6404);
or (n6407,n6408,n6411);
and (n6408,n6409,n6410);
xor (n6409,n6331,n6332);
and (n6410,n1344,n143);
and (n6411,n6412,n6413);
xor (n6412,n6409,n6410);
or (n6413,n6414,n6417);
and (n6414,n6415,n6416);
xor (n6415,n6337,n6338);
and (n6416,n1215,n143);
and (n6417,n6418,n6419);
xor (n6418,n6415,n6416);
or (n6419,n6420,n6423);
and (n6420,n6421,n6422);
xor (n6421,n6343,n6344);
and (n6422,n1210,n143);
and (n6423,n6424,n6425);
xor (n6424,n6421,n6422);
or (n6425,n6426,n6429);
and (n6426,n6427,n6428);
xor (n6427,n6348,n6349);
and (n6428,n1317,n143);
and (n6429,n6430,n6431);
xor (n6430,n6427,n6428);
or (n6431,n6432,n6435);
and (n6432,n6433,n6434);
xor (n6433,n6354,n6355);
and (n6434,n1323,n143);
and (n6435,n6436,n6437);
xor (n6436,n6433,n6434);
and (n6437,n6438,n1876);
xor (n6438,n6360,n6361);
and (n6439,n453,n144);
or (n6440,n6441,n6444);
and (n6441,n6442,n6443);
xor (n6442,n6370,n6371);
and (n6443,n434,n144);
and (n6444,n6445,n6446);
xor (n6445,n6442,n6443);
or (n6446,n6447,n6450);
and (n6447,n6448,n6449);
xor (n6448,n6376,n6377);
and (n6449,n389,n144);
and (n6450,n6451,n6452);
xor (n6451,n6448,n6449);
or (n6452,n6453,n6456);
and (n6453,n6454,n6455);
xor (n6454,n6382,n6383);
and (n6455,n371,n144);
and (n6456,n6457,n6458);
xor (n6457,n6454,n6455);
or (n6458,n6459,n6462);
and (n6459,n6460,n6461);
xor (n6460,n6388,n6389);
and (n6461,n162,n144);
and (n6462,n6463,n6464);
xor (n6463,n6460,n6461);
or (n6464,n6465,n6468);
and (n6465,n6466,n6467);
xor (n6466,n6394,n6395);
and (n6467,n156,n144);
and (n6468,n6469,n6470);
xor (n6469,n6466,n6467);
or (n6470,n6471,n6474);
and (n6471,n6472,n6473);
xor (n6472,n6400,n6401);
and (n6473,n935,n144);
and (n6474,n6475,n6476);
xor (n6475,n6472,n6473);
or (n6476,n6477,n6480);
and (n6477,n6478,n6479);
xor (n6478,n6406,n6407);
and (n6479,n1344,n144);
and (n6480,n6481,n6482);
xor (n6481,n6478,n6479);
or (n6482,n6483,n6485);
and (n6483,n6484,n4490);
xor (n6484,n6412,n6413);
and (n6485,n6486,n6487);
xor (n6486,n6484,n4490);
or (n6487,n6488,n6490);
and (n6488,n6489,n4062);
xor (n6489,n6418,n6419);
and (n6490,n6491,n6492);
xor (n6491,n6489,n4062);
or (n6492,n6493,n6495);
and (n6493,n6494,n3711);
xor (n6494,n6424,n6425);
and (n6495,n6496,n6497);
xor (n6496,n6494,n3711);
or (n6497,n6498,n6501);
and (n6498,n6499,n6500);
xor (n6499,n6430,n6431);
and (n6500,n1323,n144);
and (n6501,n6502,n6503);
xor (n6502,n6499,n6500);
and (n6503,n6504,n6505);
xor (n6504,n6436,n6437);
and (n6505,n1463,n144);
or (n6506,n6507,n6509);
and (n6507,n6508,n6449);
xor (n6508,n6445,n6446);
and (n6509,n6510,n6511);
xor (n6510,n6508,n6449);
or (n6511,n6512,n6514);
and (n6512,n6513,n6455);
xor (n6513,n6451,n6452);
and (n6514,n6515,n6516);
xor (n6515,n6513,n6455);
or (n6516,n6517,n6519);
and (n6517,n6518,n6461);
xor (n6518,n6457,n6458);
and (n6519,n6520,n6521);
xor (n6520,n6518,n6461);
or (n6521,n6522,n6524);
and (n6522,n6523,n6467);
xor (n6523,n6463,n6464);
and (n6524,n6525,n6526);
xor (n6525,n6523,n6467);
or (n6526,n6527,n6529);
and (n6527,n6528,n6473);
xor (n6528,n6469,n6470);
and (n6529,n6530,n6531);
xor (n6530,n6528,n6473);
or (n6531,n6532,n6534);
and (n6532,n6533,n6479);
xor (n6533,n6475,n6476);
and (n6534,n6535,n6536);
xor (n6535,n6533,n6479);
or (n6536,n6537,n6539);
and (n6537,n6538,n4490);
xor (n6538,n6481,n6482);
and (n6539,n6540,n6541);
xor (n6540,n6538,n4490);
or (n6541,n6542,n6544);
and (n6542,n6543,n4062);
xor (n6543,n6486,n6487);
and (n6544,n6545,n6546);
xor (n6545,n6543,n4062);
or (n6546,n6547,n6549);
and (n6547,n6548,n3711);
xor (n6548,n6491,n6492);
and (n6549,n6550,n6551);
xor (n6550,n6548,n3711);
or (n6551,n6552,n6554);
and (n6552,n6553,n6500);
xor (n6553,n6496,n6497);
and (n6554,n6555,n6556);
xor (n6555,n6553,n6500);
and (n6556,n6557,n6505);
xor (n6557,n6502,n6503);
or (n6558,n6559,n6561);
and (n6559,n6560,n6455);
xor (n6560,n6510,n6511);
and (n6561,n6562,n6563);
xor (n6562,n6560,n6455);
or (n6563,n6564,n6566);
and (n6564,n6565,n6461);
xor (n6565,n6515,n6516);
and (n6566,n6567,n6568);
xor (n6567,n6565,n6461);
or (n6568,n6569,n6571);
and (n6569,n6570,n6467);
xor (n6570,n6520,n6521);
and (n6571,n6572,n6573);
xor (n6572,n6570,n6467);
or (n6573,n6574,n6576);
and (n6574,n6575,n6473);
xor (n6575,n6525,n6526);
and (n6576,n6577,n6578);
xor (n6577,n6575,n6473);
or (n6578,n6579,n6581);
and (n6579,n6580,n6479);
xor (n6580,n6530,n6531);
and (n6581,n6582,n6583);
xor (n6582,n6580,n6479);
or (n6583,n6584,n6586);
and (n6584,n6585,n4490);
xor (n6585,n6535,n6536);
and (n6586,n6587,n6588);
xor (n6587,n6585,n4490);
or (n6588,n6589,n6591);
and (n6589,n6590,n4062);
xor (n6590,n6540,n6541);
and (n6591,n6592,n6593);
xor (n6592,n6590,n4062);
or (n6593,n6594,n6596);
and (n6594,n6595,n3711);
xor (n6595,n6545,n6546);
and (n6596,n6597,n6598);
xor (n6597,n6595,n3711);
or (n6598,n6599,n6601);
and (n6599,n6600,n6500);
xor (n6600,n6550,n6551);
and (n6601,n6602,n6603);
xor (n6602,n6600,n6500);
and (n6603,n6604,n6505);
xor (n6604,n6555,n6556);
or (n6605,n6606,n6608);
and (n6606,n6607,n6461);
xor (n6607,n6562,n6563);
and (n6608,n6609,n6610);
xor (n6609,n6607,n6461);
or (n6610,n6611,n6613);
and (n6611,n6612,n6467);
xor (n6612,n6567,n6568);
and (n6613,n6614,n6615);
xor (n6614,n6612,n6467);
or (n6615,n6616,n6618);
and (n6616,n6617,n6473);
xor (n6617,n6572,n6573);
and (n6618,n6619,n6620);
xor (n6619,n6617,n6473);
or (n6620,n6621,n6623);
and (n6621,n6622,n6479);
xor (n6622,n6577,n6578);
and (n6623,n6624,n6625);
xor (n6624,n6622,n6479);
or (n6625,n6626,n6628);
and (n6626,n6627,n4490);
xor (n6627,n6582,n6583);
and (n6628,n6629,n6630);
xor (n6629,n6627,n4490);
or (n6630,n6631,n6633);
and (n6631,n6632,n4062);
xor (n6632,n6587,n6588);
and (n6633,n6634,n6635);
xor (n6634,n6632,n4062);
or (n6635,n6636,n6638);
and (n6636,n6637,n3711);
xor (n6637,n6592,n6593);
and (n6638,n6639,n6640);
xor (n6639,n6637,n3711);
or (n6640,n6641,n6643);
and (n6641,n6642,n6500);
xor (n6642,n6597,n6598);
and (n6643,n6644,n6645);
xor (n6644,n6642,n6500);
and (n6645,n6646,n6505);
xor (n6646,n6602,n6603);
or (n6647,n6648,n6650);
and (n6648,n6649,n6467);
xor (n6649,n6609,n6610);
and (n6650,n6651,n6652);
xor (n6651,n6649,n6467);
or (n6652,n6653,n6655);
and (n6653,n6654,n6473);
xor (n6654,n6614,n6615);
and (n6655,n6656,n6657);
xor (n6656,n6654,n6473);
or (n6657,n6658,n6660);
and (n6658,n6659,n6479);
xor (n6659,n6619,n6620);
and (n6660,n6661,n6662);
xor (n6661,n6659,n6479);
or (n6662,n6663,n6665);
and (n6663,n6664,n4490);
xor (n6664,n6624,n6625);
and (n6665,n6666,n6667);
xor (n6666,n6664,n4490);
or (n6667,n6668,n6670);
and (n6668,n6669,n4062);
xor (n6669,n6629,n6630);
and (n6670,n6671,n6672);
xor (n6671,n6669,n4062);
or (n6672,n6673,n6675);
and (n6673,n6674,n3711);
xor (n6674,n6634,n6635);
and (n6675,n6676,n6677);
xor (n6676,n6674,n3711);
or (n6677,n6678,n6680);
and (n6678,n6679,n6500);
xor (n6679,n6639,n6640);
and (n6680,n6681,n6682);
xor (n6681,n6679,n6500);
and (n6682,n6683,n6505);
xor (n6683,n6644,n6645);
or (n6684,n6685,n6687);
and (n6685,n6686,n6473);
xor (n6686,n6651,n6652);
and (n6687,n6688,n6689);
xor (n6688,n6686,n6473);
or (n6689,n6690,n6692);
and (n6690,n6691,n6479);
xor (n6691,n6656,n6657);
and (n6692,n6693,n6694);
xor (n6693,n6691,n6479);
or (n6694,n6695,n6697);
and (n6695,n6696,n4490);
xor (n6696,n6661,n6662);
and (n6697,n6698,n6699);
xor (n6698,n6696,n4490);
or (n6699,n6700,n6702);
and (n6700,n6701,n4062);
xor (n6701,n6666,n6667);
and (n6702,n6703,n6704);
xor (n6703,n6701,n4062);
or (n6704,n6705,n6707);
and (n6705,n6706,n3711);
xor (n6706,n6671,n6672);
and (n6707,n6708,n6709);
xor (n6708,n6706,n3711);
or (n6709,n6710,n6712);
and (n6710,n6711,n6500);
xor (n6711,n6676,n6677);
and (n6712,n6713,n6714);
xor (n6713,n6711,n6500);
and (n6714,n6715,n6505);
xor (n6715,n6681,n6682);
or (n6716,n6717,n6719);
and (n6717,n6718,n6479);
xor (n6718,n6688,n6689);
and (n6719,n6720,n6721);
xor (n6720,n6718,n6479);
or (n6721,n6722,n6724);
and (n6722,n6723,n4490);
xor (n6723,n6693,n6694);
and (n6724,n6725,n6726);
xor (n6725,n6723,n4490);
or (n6726,n6727,n6729);
and (n6727,n6728,n4062);
xor (n6728,n6698,n6699);
and (n6729,n6730,n6731);
xor (n6730,n6728,n4062);
or (n6731,n6732,n6734);
and (n6732,n6733,n3711);
xor (n6733,n6703,n6704);
and (n6734,n6735,n6736);
xor (n6735,n6733,n3711);
or (n6736,n6737,n6739);
and (n6737,n6738,n6500);
xor (n6738,n6708,n6709);
and (n6739,n6740,n6741);
xor (n6740,n6738,n6500);
and (n6741,n6742,n6505);
xor (n6742,n6713,n6714);
or (n6743,n6744,n6746);
and (n6744,n6745,n4490);
xor (n6745,n6720,n6721);
and (n6746,n6747,n6748);
xor (n6747,n6745,n4490);
or (n6748,n6749,n6751);
and (n6749,n6750,n4062);
xor (n6750,n6725,n6726);
and (n6751,n6752,n6753);
xor (n6752,n6750,n4062);
or (n6753,n6754,n6756);
and (n6754,n6755,n3711);
xor (n6755,n6730,n6731);
and (n6756,n6757,n6758);
xor (n6757,n6755,n3711);
or (n6758,n6759,n6761);
and (n6759,n6760,n6500);
xor (n6760,n6735,n6736);
and (n6761,n6762,n6763);
xor (n6762,n6760,n6500);
and (n6763,n6764,n6505);
xor (n6764,n6740,n6741);
or (n6765,n6766,n6768);
and (n6766,n6767,n4062);
xor (n6767,n6747,n6748);
and (n6768,n6769,n6770);
xor (n6769,n6767,n4062);
or (n6770,n6771,n6773);
and (n6771,n6772,n3711);
xor (n6772,n6752,n6753);
and (n6773,n6774,n6775);
xor (n6774,n6772,n3711);
or (n6775,n6776,n6778);
and (n6776,n6777,n6500);
xor (n6777,n6757,n6758);
and (n6778,n6779,n6780);
xor (n6779,n6777,n6500);
and (n6780,n6781,n6505);
xor (n6781,n6762,n6763);
or (n6782,n6783,n6785);
and (n6783,n6784,n3711);
xor (n6784,n6769,n6770);
and (n6785,n6786,n6787);
xor (n6786,n6784,n3711);
or (n6787,n6788,n6790);
and (n6788,n6789,n6500);
xor (n6789,n6774,n6775);
and (n6790,n6791,n6792);
xor (n6791,n6789,n6500);
and (n6792,n6793,n6505);
xor (n6793,n6779,n6780);
or (n6794,n6795,n6797);
and (n6795,n6796,n6500);
xor (n6796,n6786,n6787);
and (n6797,n6798,n6799);
xor (n6798,n6796,n6500);
and (n6799,n6800,n6505);
xor (n6800,n6791,n6792);
and (n6801,n6802,n6505);
xor (n6802,n6798,n6799);
xor (n6803,n6804,n1750);
xor (n6804,n6805,n8405);
xor (n6805,n6806,n1754);
xor (n6806,n6807,n8398);
xor (n6807,n6808,n8100);
xor (n6808,n6809,n8386);
xor (n6809,n6810,n3915);
xor (n6810,n6811,n8369);
xor (n6811,n6812,n4369);
xor (n6812,n6813,n8347);
xor (n6813,n6814,n4645);
xor (n6814,n6815,n8320);
xor (n6815,n6816,n929);
xor (n6816,n6817,n8288);
xor (n6817,n6818,n8074);
xor (n6818,n6819,n8251);
xor (n6819,n6820,n135);
xor (n6820,n6821,n8209);
xor (n6821,n6822,n513);
xor (n6822,n6823,n8162);
xor (n6823,n6824,n8058);
xor (n6824,n6825,n8110);
xor (n6825,n6826,n8052);
xor (n6826,n6827,n8049);
xor (n6827,n6828,n8048);
xor (n6828,n6829,n7973);
xor (n6829,n6830,n7972);
xor (n6830,n6831,n7895);
xor (n6831,n6832,n7894);
xor (n6832,n6833,n7807);
xor (n6833,n6834,n7806);
or (n6834,n6835,n7723);
and (n6835,n6836,n7722);
or (n6836,n6837,n7634);
and (n6837,n6838,n7633);
or (n6838,n6839,n7550);
and (n6839,n6840,n591);
or (n6840,n6841,n7461);
and (n6841,n6842,n7460);
or (n6842,n6843,n7377);
and (n6843,n6844,n7376);
or (n6844,n6845,n7288);
and (n6845,n6846,n7287);
or (n6846,n6847,n7200);
and (n6847,n6848,n7199);
or (n6848,n6849,n7110);
and (n6849,n6850,n7109);
or (n6850,n6851,n7026);
and (n6851,n6852,n7025);
or (n6852,n6853,n6937);
and (n6853,n6854,n6936);
and (n6854,n1843,n6855);
or (n6855,n6856,n6858);
and (n6856,n6857,n1186);
and (n6857,n358,n1177);
and (n6858,n6859,n6860);
xor (n6859,n6857,n1186);
or (n6860,n6861,n6863);
and (n6861,n6862,n1182);
and (n6862,n85,n1177);
and (n6863,n6864,n6865);
xor (n6864,n6862,n1182);
or (n6865,n6866,n6868);
and (n6866,n6867,n1908);
and (n6867,n79,n1177);
and (n6868,n6869,n6870);
xor (n6869,n6867,n1908);
or (n6870,n6871,n6873);
and (n6871,n6872,n1530);
and (n6872,n489,n1177);
and (n6873,n6874,n6875);
xor (n6874,n6872,n1530);
or (n6875,n6876,n6879);
and (n6876,n6877,n6878);
and (n6877,n483,n1177);
and (n6878,n341,n1175);
and (n6879,n6880,n6881);
xor (n6880,n6877,n6878);
or (n6881,n6882,n6885);
and (n6882,n6883,n6884);
and (n6883,n341,n1177);
and (n6884,n348,n1175);
and (n6885,n6886,n6887);
xor (n6886,n6883,n6884);
or (n6887,n6888,n6891);
and (n6888,n6889,n6890);
and (n6889,n348,n1177);
and (n6890,n134,n1175);
and (n6891,n6892,n6893);
xor (n6892,n6889,n6890);
or (n6893,n6894,n6897);
and (n6894,n6895,n6896);
and (n6895,n134,n1177);
and (n6896,n114,n1175);
and (n6897,n6898,n6899);
xor (n6898,n6895,n6896);
or (n6899,n6900,n6903);
and (n6900,n6901,n6902);
and (n6901,n114,n1177);
and (n6902,n928,n1175);
and (n6903,n6904,n6905);
xor (n6904,n6901,n6902);
or (n6905,n6906,n6909);
and (n6906,n6907,n6908);
and (n6907,n928,n1177);
and (n6908,n1357,n1175);
and (n6909,n6910,n6911);
xor (n6910,n6907,n6908);
or (n6911,n6912,n6915);
and (n6912,n6913,n6914);
and (n6913,n1357,n1177);
and (n6914,n1169,n1175);
and (n6915,n6916,n6917);
xor (n6916,n6913,n6914);
or (n6917,n6918,n6920);
and (n6918,n6919,n3275);
and (n6919,n1169,n1177);
and (n6920,n6921,n6922);
xor (n6921,n6919,n3275);
or (n6922,n6923,n6925);
and (n6923,n6924,n3368);
and (n6924,n1163,n1177);
and (n6925,n6926,n6927);
xor (n6926,n6924,n3368);
or (n6927,n6928,n6931);
and (n6928,n6929,n6930);
and (n6929,n1639,n1177);
and (n6930,n1475,n1175);
and (n6931,n6932,n6933);
xor (n6932,n6929,n6930);
and (n6933,n6934,n6935);
and (n6934,n1475,n1177);
and (n6935,n1470,n1175);
and (n6936,n358,n1227);
and (n6937,n6938,n6939);
xor (n6938,n6854,n6936);
or (n6939,n6940,n6943);
and (n6940,n6941,n6942);
xor (n6941,n1843,n6855);
and (n6942,n85,n1227);
and (n6943,n6944,n6945);
xor (n6944,n6941,n6942);
or (n6945,n6946,n6949);
and (n6946,n6947,n6948);
xor (n6947,n6859,n6860);
and (n6948,n79,n1227);
and (n6949,n6950,n6951);
xor (n6950,n6947,n6948);
or (n6951,n6952,n6955);
and (n6952,n6953,n6954);
xor (n6953,n6864,n6865);
and (n6954,n489,n1227);
and (n6955,n6956,n6957);
xor (n6956,n6953,n6954);
or (n6957,n6958,n6961);
and (n6958,n6959,n6960);
xor (n6959,n6869,n6870);
and (n6960,n483,n1227);
and (n6961,n6962,n6963);
xor (n6962,n6959,n6960);
or (n6963,n6964,n6967);
and (n6964,n6965,n6966);
xor (n6965,n6874,n6875);
and (n6966,n341,n1227);
and (n6967,n6968,n6969);
xor (n6968,n6965,n6966);
or (n6969,n6970,n6973);
and (n6970,n6971,n6972);
xor (n6971,n6880,n6881);
and (n6972,n348,n1227);
and (n6973,n6974,n6975);
xor (n6974,n6971,n6972);
or (n6975,n6976,n6979);
and (n6976,n6977,n6978);
xor (n6977,n6886,n6887);
and (n6978,n134,n1227);
and (n6979,n6980,n6981);
xor (n6980,n6977,n6978);
or (n6981,n6982,n6985);
and (n6982,n6983,n6984);
xor (n6983,n6892,n6893);
and (n6984,n114,n1227);
and (n6985,n6986,n6987);
xor (n6986,n6983,n6984);
or (n6987,n6988,n6991);
and (n6988,n6989,n6990);
xor (n6989,n6898,n6899);
and (n6990,n928,n1227);
and (n6991,n6992,n6993);
xor (n6992,n6989,n6990);
or (n6993,n6994,n6997);
and (n6994,n6995,n6996);
xor (n6995,n6904,n6905);
and (n6996,n1357,n1227);
and (n6997,n6998,n6999);
xor (n6998,n6995,n6996);
or (n6999,n7000,n7003);
and (n7000,n7001,n7002);
xor (n7001,n6910,n6911);
and (n7002,n1169,n1227);
and (n7003,n7004,n7005);
xor (n7004,n7001,n7002);
or (n7005,n7006,n7009);
and (n7006,n7007,n7008);
xor (n7007,n6916,n6917);
and (n7008,n1163,n1227);
and (n7009,n7010,n7011);
xor (n7010,n7007,n7008);
or (n7011,n7012,n7015);
and (n7012,n7013,n7014);
xor (n7013,n6921,n6922);
and (n7014,n1639,n1227);
and (n7015,n7016,n7017);
xor (n7016,n7013,n7014);
or (n7017,n7018,n7021);
and (n7018,n7019,n7020);
xor (n7019,n6926,n6927);
and (n7020,n1475,n1227);
and (n7021,n7022,n7023);
xor (n7022,n7019,n7020);
and (n7023,n7024,n3408);
xor (n7024,n6932,n6933);
and (n7025,n358,n203);
and (n7026,n7027,n7028);
xor (n7027,n6852,n7025);
or (n7028,n7029,n7032);
and (n7029,n7030,n7031);
xor (n7030,n6938,n6939);
and (n7031,n85,n203);
and (n7032,n7033,n7034);
xor (n7033,n7030,n7031);
or (n7034,n7035,n7038);
and (n7035,n7036,n7037);
xor (n7036,n6944,n6945);
and (n7037,n79,n203);
and (n7038,n7039,n7040);
xor (n7039,n7036,n7037);
or (n7040,n7041,n7044);
and (n7041,n7042,n7043);
xor (n7042,n6950,n6951);
and (n7043,n489,n203);
and (n7044,n7045,n7046);
xor (n7045,n7042,n7043);
or (n7046,n7047,n7050);
and (n7047,n7048,n7049);
xor (n7048,n6956,n6957);
and (n7049,n483,n203);
and (n7050,n7051,n7052);
xor (n7051,n7048,n7049);
or (n7052,n7053,n7055);
and (n7053,n7054,n1902);
xor (n7054,n6962,n6963);
and (n7055,n7056,n7057);
xor (n7056,n7054,n1902);
or (n7057,n7058,n7061);
and (n7058,n7059,n7060);
xor (n7059,n6968,n6969);
and (n7060,n348,n203);
and (n7061,n7062,n7063);
xor (n7062,n7059,n7060);
or (n7063,n7064,n7067);
and (n7064,n7065,n7066);
xor (n7065,n6974,n6975);
and (n7066,n134,n203);
and (n7067,n7068,n7069);
xor (n7068,n7065,n7066);
or (n7069,n7070,n7073);
and (n7070,n7071,n7072);
xor (n7071,n6980,n6981);
and (n7072,n114,n203);
and (n7073,n7074,n7075);
xor (n7074,n7071,n7072);
or (n7075,n7076,n7078);
and (n7076,n7077,n2615);
xor (n7077,n6986,n6987);
and (n7078,n7079,n7080);
xor (n7079,n7077,n2615);
or (n7080,n7081,n7083);
and (n7081,n7082,n2801);
xor (n7082,n6992,n6993);
and (n7083,n7084,n7085);
xor (n7084,n7082,n2801);
or (n7085,n7086,n7088);
and (n7086,n7087,n2945);
xor (n7087,n6998,n6999);
and (n7088,n7089,n7090);
xor (n7089,n7087,n2945);
or (n7090,n7091,n7093);
and (n7091,n7092,n3089);
xor (n7092,n7004,n7005);
and (n7093,n7094,n7095);
xor (n7094,n7092,n3089);
or (n7095,n7096,n7099);
and (n7096,n7097,n7098);
xor (n7097,n7010,n7011);
and (n7098,n1639,n203);
and (n7099,n7100,n7101);
xor (n7100,n7097,n7098);
or (n7101,n7102,n7104);
and (n7102,n7103,n3316);
xor (n7103,n7016,n7017);
and (n7104,n7105,n7106);
xor (n7105,n7103,n3316);
and (n7106,n7107,n7108);
xor (n7107,n7022,n7023);
and (n7108,n1470,n203);
and (n7109,n358,n204);
and (n7110,n7111,n7112);
xor (n7111,n6850,n7109);
or (n7112,n7113,n7116);
and (n7113,n7114,n7115);
xor (n7114,n7027,n7028);
and (n7115,n85,n204);
and (n7116,n7117,n7118);
xor (n7117,n7114,n7115);
or (n7118,n7119,n7122);
and (n7119,n7120,n7121);
xor (n7120,n7033,n7034);
and (n7121,n79,n204);
and (n7122,n7123,n7124);
xor (n7123,n7120,n7121);
or (n7124,n7125,n7128);
and (n7125,n7126,n7127);
xor (n7126,n7039,n7040);
and (n7127,n489,n204);
and (n7128,n7129,n7130);
xor (n7129,n7126,n7127);
or (n7130,n7131,n7134);
and (n7131,n7132,n7133);
xor (n7132,n7045,n7046);
and (n7133,n483,n204);
and (n7134,n7135,n7136);
xor (n7135,n7132,n7133);
or (n7136,n7137,n7140);
and (n7137,n7138,n7139);
xor (n7138,n7051,n7052);
and (n7139,n341,n204);
and (n7140,n7141,n7142);
xor (n7141,n7138,n7139);
or (n7142,n7143,n7146);
and (n7143,n7144,n7145);
xor (n7144,n7056,n7057);
and (n7145,n348,n204);
and (n7146,n7147,n7148);
xor (n7147,n7144,n7145);
or (n7148,n7149,n7152);
and (n7149,n7150,n7151);
xor (n7150,n7062,n7063);
and (n7151,n134,n204);
and (n7152,n7153,n7154);
xor (n7153,n7150,n7151);
or (n7154,n7155,n7158);
and (n7155,n7156,n7157);
xor (n7156,n7068,n7069);
and (n7157,n114,n204);
and (n7158,n7159,n7160);
xor (n7159,n7156,n7157);
or (n7160,n7161,n7164);
and (n7161,n7162,n7163);
xor (n7162,n7074,n7075);
and (n7163,n928,n204);
and (n7164,n7165,n7166);
xor (n7165,n7162,n7163);
or (n7166,n7167,n7170);
and (n7167,n7168,n7169);
xor (n7168,n7079,n7080);
and (n7169,n1357,n204);
and (n7170,n7171,n7172);
xor (n7171,n7168,n7169);
or (n7172,n7173,n7176);
and (n7173,n7174,n7175);
xor (n7174,n7084,n7085);
and (n7175,n1169,n204);
and (n7176,n7177,n7178);
xor (n7177,n7174,n7175);
or (n7178,n7179,n7182);
and (n7179,n7180,n7181);
xor (n7180,n7089,n7090);
and (n7181,n1163,n204);
and (n7182,n7183,n7184);
xor (n7183,n7180,n7181);
or (n7184,n7185,n7188);
and (n7185,n7186,n7187);
xor (n7186,n7094,n7095);
and (n7187,n1639,n204);
and (n7188,n7189,n7190);
xor (n7189,n7186,n7187);
or (n7190,n7191,n7194);
and (n7191,n7192,n7193);
xor (n7192,n7100,n7101);
and (n7193,n1475,n204);
and (n7194,n7195,n7196);
xor (n7195,n7192,n7193);
and (n7196,n7197,n7198);
xor (n7197,n7105,n7106);
not (n7198,n3153);
and (n7199,n358,n28);
and (n7200,n7201,n7202);
xor (n7201,n6848,n7199);
or (n7202,n7203,n7206);
and (n7203,n7204,n7205);
xor (n7204,n7111,n7112);
and (n7205,n85,n28);
and (n7206,n7207,n7208);
xor (n7207,n7204,n7205);
or (n7208,n7209,n7212);
and (n7209,n7210,n7211);
xor (n7210,n7117,n7118);
and (n7211,n79,n28);
and (n7212,n7213,n7214);
xor (n7213,n7210,n7211);
or (n7214,n7215,n7218);
and (n7215,n7216,n7217);
xor (n7216,n7123,n7124);
and (n7217,n489,n28);
and (n7218,n7219,n7220);
xor (n7219,n7216,n7217);
or (n7220,n7221,n7224);
and (n7221,n7222,n7223);
xor (n7222,n7129,n7130);
and (n7223,n483,n28);
and (n7224,n7225,n7226);
xor (n7225,n7222,n7223);
or (n7226,n7227,n7230);
and (n7227,n7228,n7229);
xor (n7228,n7135,n7136);
and (n7229,n341,n28);
and (n7230,n7231,n7232);
xor (n7231,n7228,n7229);
or (n7232,n7233,n7236);
and (n7233,n7234,n7235);
xor (n7234,n7141,n7142);
and (n7235,n348,n28);
and (n7236,n7237,n7238);
xor (n7237,n7234,n7235);
or (n7238,n7239,n7242);
and (n7239,n7240,n7241);
xor (n7240,n7147,n7148);
and (n7241,n134,n28);
and (n7242,n7243,n7244);
xor (n7243,n7240,n7241);
or (n7244,n7245,n7248);
and (n7245,n7246,n7247);
xor (n7246,n7153,n7154);
and (n7247,n114,n28);
and (n7248,n7249,n7250);
xor (n7249,n7246,n7247);
or (n7250,n7251,n7254);
and (n7251,n7252,n7253);
xor (n7252,n7159,n7160);
and (n7253,n928,n28);
and (n7254,n7255,n7256);
xor (n7255,n7252,n7253);
or (n7256,n7257,n7259);
and (n7257,n7258,n2416);
xor (n7258,n7165,n7166);
and (n7259,n7260,n7261);
xor (n7260,n7258,n2416);
or (n7261,n7262,n7265);
and (n7262,n7263,n7264);
xor (n7263,n7171,n7172);
and (n7264,n1169,n28);
and (n7265,n7266,n7267);
xor (n7266,n7263,n7264);
or (n7267,n7268,n7271);
and (n7268,n7269,n7270);
xor (n7269,n7177,n7178);
and (n7270,n1163,n28);
and (n7271,n7272,n7273);
xor (n7272,n7269,n7270);
or (n7273,n7274,n7276);
and (n7274,n7275,n2919);
xor (n7275,n7183,n7184);
and (n7276,n7277,n7278);
xor (n7277,n7275,n2919);
or (n7278,n7279,n7282);
and (n7279,n7280,n7281);
xor (n7280,n7189,n7190);
and (n7281,n1475,n28);
and (n7282,n7283,n7284);
xor (n7283,n7280,n7281);
and (n7284,n7285,n7286);
xor (n7285,n7195,n7196);
and (n7286,n1470,n28);
and (n7287,n358,n27);
and (n7288,n7289,n7290);
xor (n7289,n6846,n7287);
or (n7290,n7291,n7294);
and (n7291,n7292,n7293);
xor (n7292,n7201,n7202);
and (n7293,n85,n27);
and (n7294,n7295,n7296);
xor (n7295,n7292,n7293);
or (n7296,n7297,n7300);
and (n7297,n7298,n7299);
xor (n7298,n7207,n7208);
and (n7299,n79,n27);
and (n7300,n7301,n7302);
xor (n7301,n7298,n7299);
or (n7302,n7303,n7306);
and (n7303,n7304,n7305);
xor (n7304,n7213,n7214);
and (n7305,n489,n27);
and (n7306,n7307,n7308);
xor (n7307,n7304,n7305);
or (n7308,n7309,n7312);
and (n7309,n7310,n7311);
xor (n7310,n7219,n7220);
and (n7311,n483,n27);
and (n7312,n7313,n7314);
xor (n7313,n7310,n7311);
or (n7314,n7315,n7318);
and (n7315,n7316,n7317);
xor (n7316,n7225,n7226);
and (n7317,n341,n27);
and (n7318,n7319,n7320);
xor (n7319,n7316,n7317);
or (n7320,n7321,n7324);
and (n7321,n7322,n7323);
xor (n7322,n7231,n7232);
and (n7323,n348,n27);
and (n7324,n7325,n7326);
xor (n7325,n7322,n7323);
or (n7326,n7327,n7330);
and (n7327,n7328,n7329);
xor (n7328,n7237,n7238);
and (n7329,n134,n27);
and (n7330,n7331,n7332);
xor (n7331,n7328,n7329);
or (n7332,n7333,n7336);
and (n7333,n7334,n7335);
xor (n7334,n7243,n7244);
and (n7335,n114,n27);
and (n7336,n7337,n7338);
xor (n7337,n7334,n7335);
or (n7338,n7339,n7342);
and (n7339,n7340,n7341);
xor (n7340,n7249,n7250);
and (n7341,n928,n27);
and (n7342,n7343,n7344);
xor (n7343,n7340,n7341);
or (n7344,n7345,n7348);
and (n7345,n7346,n7347);
xor (n7346,n7255,n7256);
and (n7347,n1357,n27);
and (n7348,n7349,n7350);
xor (n7349,n7346,n7347);
or (n7350,n7351,n7354);
and (n7351,n7352,n7353);
xor (n7352,n7260,n7261);
and (n7353,n1169,n27);
and (n7354,n7355,n7356);
xor (n7355,n7352,n7353);
or (n7356,n7357,n7360);
and (n7357,n7358,n7359);
xor (n7358,n7266,n7267);
and (n7359,n1163,n27);
and (n7360,n7361,n7362);
xor (n7361,n7358,n7359);
or (n7362,n7363,n7366);
and (n7363,n7364,n7365);
xor (n7364,n7272,n7273);
and (n7365,n1639,n27);
and (n7366,n7367,n7368);
xor (n7367,n7364,n7365);
or (n7368,n7369,n7372);
and (n7369,n7370,n7371);
xor (n7370,n7277,n7278);
and (n7371,n1475,n27);
and (n7372,n7373,n7374);
xor (n7373,n7370,n7371);
and (n7374,n7375,n2862);
xor (n7375,n7283,n7284);
and (n7376,n358,n33);
and (n7377,n7378,n7379);
xor (n7378,n6844,n7376);
or (n7379,n7380,n7382);
and (n7380,n7381,n4199);
xor (n7381,n7289,n7290);
and (n7382,n7383,n7384);
xor (n7383,n7381,n4199);
or (n7384,n7385,n7388);
and (n7385,n7386,n7387);
xor (n7386,n7295,n7296);
and (n7387,n79,n33);
and (n7388,n7389,n7390);
xor (n7389,n7386,n7387);
or (n7390,n7391,n7394);
and (n7391,n7392,n7393);
xor (n7392,n7301,n7302);
and (n7393,n489,n33);
and (n7394,n7395,n7396);
xor (n7395,n7392,n7393);
or (n7396,n7397,n7399);
and (n7397,n7398,n4089);
xor (n7398,n7307,n7308);
and (n7399,n7400,n7401);
xor (n7400,n7398,n4089);
or (n7401,n7402,n7404);
and (n7402,n7403,n3731);
xor (n7403,n7313,n7314);
and (n7404,n7405,n7406);
xor (n7405,n7403,n3731);
or (n7406,n7407,n7409);
and (n7407,n7408,n1855);
xor (n7408,n7319,n7320);
and (n7409,n7410,n7411);
xor (n7410,n7408,n1855);
or (n7411,n7412,n7415);
and (n7412,n7413,n7414);
xor (n7413,n7325,n7326);
and (n7414,n134,n33);
and (n7415,n7416,n7417);
xor (n7416,n7413,n7414);
or (n7417,n7418,n7421);
and (n7418,n7419,n7420);
xor (n7419,n7331,n7332);
and (n7420,n114,n33);
and (n7421,n7422,n7423);
xor (n7422,n7419,n7420);
or (n7423,n7424,n7427);
and (n7424,n7425,n7426);
xor (n7425,n7337,n7338);
and (n7426,n928,n33);
and (n7427,n7428,n7429);
xor (n7428,n7425,n7426);
or (n7429,n7430,n7433);
and (n7430,n7431,n7432);
xor (n7431,n7343,n7344);
and (n7432,n1357,n33);
and (n7433,n7434,n7435);
xor (n7434,n7431,n7432);
or (n7435,n7436,n7438);
and (n7436,n7437,n1434);
xor (n7437,n7349,n7350);
and (n7438,n7439,n7440);
xor (n7439,n7437,n1434);
or (n7440,n7441,n7443);
and (n7441,n7442,n2362);
xor (n7442,n7355,n7356);
and (n7443,n7444,n7445);
xor (n7444,n7442,n2362);
or (n7445,n7446,n7449);
and (n7446,n7447,n7448);
xor (n7447,n7361,n7362);
and (n7448,n1639,n33);
and (n7449,n7450,n7451);
xor (n7450,n7447,n7448);
or (n7451,n7452,n7455);
and (n7452,n7453,n7454);
xor (n7453,n7367,n7368);
and (n7454,n1475,n33);
and (n7455,n7456,n7457);
xor (n7456,n7453,n7454);
and (n7457,n7458,n7459);
xor (n7458,n7373,n7374);
and (n7459,n1470,n33);
and (n7460,n358,n237);
and (n7461,n7462,n7463);
xor (n7462,n6842,n7460);
or (n7463,n7464,n7467);
and (n7464,n7465,n7466);
xor (n7465,n7378,n7379);
and (n7466,n85,n237);
and (n7467,n7468,n7469);
xor (n7468,n7465,n7466);
or (n7469,n7470,n7473);
and (n7470,n7471,n7472);
xor (n7471,n7383,n7384);
and (n7472,n79,n237);
and (n7473,n7474,n7475);
xor (n7474,n7471,n7472);
or (n7475,n7476,n7479);
and (n7476,n7477,n7478);
xor (n7477,n7389,n7390);
and (n7478,n489,n237);
and (n7479,n7480,n7481);
xor (n7480,n7477,n7478);
or (n7481,n7482,n7485);
and (n7482,n7483,n7484);
xor (n7483,n7395,n7396);
and (n7484,n483,n237);
and (n7485,n7486,n7487);
xor (n7486,n7483,n7484);
or (n7487,n7488,n7491);
and (n7488,n7489,n7490);
xor (n7489,n7400,n7401);
and (n7490,n341,n237);
and (n7491,n7492,n7493);
xor (n7492,n7489,n7490);
or (n7493,n7494,n7497);
and (n7494,n7495,n7496);
xor (n7495,n7405,n7406);
and (n7496,n348,n237);
and (n7497,n7498,n7499);
xor (n7498,n7495,n7496);
or (n7499,n7500,n7503);
and (n7500,n7501,n7502);
xor (n7501,n7410,n7411);
and (n7502,n134,n237);
and (n7503,n7504,n7505);
xor (n7504,n7501,n7502);
or (n7505,n7506,n7509);
and (n7506,n7507,n7508);
xor (n7507,n7416,n7417);
and (n7508,n114,n237);
and (n7509,n7510,n7511);
xor (n7510,n7507,n7508);
or (n7511,n7512,n7515);
and (n7512,n7513,n7514);
xor (n7513,n7422,n7423);
and (n7514,n928,n237);
and (n7515,n7516,n7517);
xor (n7516,n7513,n7514);
or (n7517,n7518,n7521);
and (n7518,n7519,n7520);
xor (n7519,n7428,n7429);
and (n7520,n1357,n237);
and (n7521,n7522,n7523);
xor (n7522,n7519,n7520);
or (n7523,n7524,n7527);
and (n7524,n7525,n7526);
xor (n7525,n7434,n7435);
and (n7526,n1169,n237);
and (n7527,n7528,n7529);
xor (n7528,n7525,n7526);
or (n7529,n7530,n7533);
and (n7530,n7531,n7532);
xor (n7531,n7439,n7440);
and (n7532,n1163,n237);
and (n7533,n7534,n7535);
xor (n7534,n7531,n7532);
or (n7535,n7536,n7539);
and (n7536,n7537,n7538);
xor (n7537,n7444,n7445);
and (n7538,n1639,n237);
and (n7539,n7540,n7541);
xor (n7540,n7537,n7538);
or (n7541,n7542,n7545);
and (n7542,n7543,n7544);
xor (n7543,n7450,n7451);
and (n7544,n1475,n237);
and (n7545,n7546,n7547);
xor (n7546,n7543,n7544);
and (n7547,n7548,n7549);
xor (n7548,n7456,n7457);
not (n7549,n2585);
and (n7550,n7551,n7552);
xor (n7551,n6840,n591);
or (n7552,n7553,n7555);
and (n7553,n7554,n246);
xor (n7554,n7462,n7463);
and (n7555,n7556,n7557);
xor (n7556,n7554,n246);
or (n7557,n7558,n7560);
and (n7558,n7559,n233);
xor (n7559,n7468,n7469);
and (n7560,n7561,n7562);
xor (n7561,n7559,n233);
or (n7562,n7563,n7565);
and (n7563,n7564,n968);
xor (n7564,n7474,n7475);
and (n7565,n7566,n7567);
xor (n7566,n7564,n968);
or (n7567,n7568,n7570);
and (n7568,n7569,n4595);
xor (n7569,n7480,n7481);
and (n7570,n7571,n7572);
xor (n7571,n7569,n4595);
or (n7572,n7573,n7576);
and (n7573,n7574,n7575);
xor (n7574,n7486,n7487);
and (n7575,n341,n68);
and (n7576,n7577,n7578);
xor (n7577,n7574,n7575);
or (n7578,n7579,n7582);
and (n7579,n7580,n7581);
xor (n7580,n7492,n7493);
and (n7581,n348,n68);
and (n7582,n7583,n7584);
xor (n7583,n7580,n7581);
or (n7584,n7585,n7588);
and (n7585,n7586,n7587);
xor (n7586,n7498,n7499);
and (n7587,n134,n68);
and (n7588,n7589,n7590);
xor (n7589,n7586,n7587);
or (n7590,n7591,n7594);
and (n7591,n7592,n7593);
xor (n7592,n7504,n7505);
and (n7593,n114,n68);
and (n7594,n7595,n7596);
xor (n7595,n7592,n7593);
or (n7596,n7597,n7600);
and (n7597,n7598,n7599);
xor (n7598,n7510,n7511);
and (n7599,n928,n68);
and (n7600,n7601,n7602);
xor (n7601,n7598,n7599);
or (n7602,n7603,n7605);
and (n7603,n7604,n1358);
xor (n7604,n7516,n7517);
and (n7605,n7606,n7607);
xor (n7606,n7604,n1358);
or (n7607,n7608,n7610);
and (n7608,n7609,n1954);
xor (n7609,n7522,n7523);
and (n7610,n7611,n7612);
xor (n7611,n7609,n1954);
or (n7612,n7613,n7616);
and (n7613,n7614,n7615);
xor (n7614,n7528,n7529);
and (n7615,n1163,n68);
and (n7616,n7617,n7618);
xor (n7617,n7614,n7615);
or (n7618,n7619,n7622);
and (n7619,n7620,n7621);
xor (n7620,n7534,n7535);
and (n7621,n1639,n68);
and (n7622,n7623,n7624);
xor (n7623,n7620,n7621);
or (n7624,n7625,n7628);
and (n7625,n7626,n7627);
xor (n7626,n7540,n7541);
and (n7627,n1475,n68);
and (n7628,n7629,n7630);
xor (n7629,n7626,n7627);
and (n7630,n7631,n7632);
xor (n7631,n7546,n7547);
and (n7632,n1470,n68);
and (n7633,n358,n69);
and (n7634,n7635,n7636);
xor (n7635,n6838,n7633);
or (n7636,n7637,n7640);
and (n7637,n7638,n7639);
xor (n7638,n7551,n7552);
and (n7639,n85,n69);
and (n7640,n7641,n7642);
xor (n7641,n7638,n7639);
or (n7642,n7643,n7646);
and (n7643,n7644,n7645);
xor (n7644,n7556,n7557);
and (n7645,n79,n69);
and (n7646,n7647,n7648);
xor (n7647,n7644,n7645);
or (n7648,n7649,n7652);
and (n7649,n7650,n7651);
xor (n7650,n7561,n7562);
and (n7651,n489,n69);
and (n7652,n7653,n7654);
xor (n7653,n7650,n7651);
or (n7654,n7655,n7658);
and (n7655,n7656,n7657);
xor (n7656,n7566,n7567);
and (n7657,n483,n69);
and (n7658,n7659,n7660);
xor (n7659,n7656,n7657);
or (n7660,n7661,n7664);
and (n7661,n7662,n7663);
xor (n7662,n7571,n7572);
and (n7663,n341,n69);
and (n7664,n7665,n7666);
xor (n7665,n7662,n7663);
or (n7666,n7667,n7670);
and (n7667,n7668,n7669);
xor (n7668,n7577,n7578);
and (n7669,n348,n69);
and (n7670,n7671,n7672);
xor (n7671,n7668,n7669);
or (n7672,n7673,n7676);
and (n7673,n7674,n7675);
xor (n7674,n7583,n7584);
and (n7675,n134,n69);
and (n7676,n7677,n7678);
xor (n7677,n7674,n7675);
or (n7678,n7679,n7682);
and (n7679,n7680,n7681);
xor (n7680,n7589,n7590);
and (n7681,n114,n69);
and (n7682,n7683,n7684);
xor (n7683,n7680,n7681);
or (n7684,n7685,n7688);
and (n7685,n7686,n7687);
xor (n7686,n7595,n7596);
and (n7687,n928,n69);
and (n7688,n7689,n7690);
xor (n7689,n7686,n7687);
or (n7690,n7691,n7694);
and (n7691,n7692,n7693);
xor (n7692,n7601,n7602);
and (n7693,n1357,n69);
and (n7694,n7695,n7696);
xor (n7695,n7692,n7693);
or (n7696,n7697,n7700);
and (n7697,n7698,n7699);
xor (n7698,n7606,n7607);
and (n7699,n1169,n69);
and (n7700,n7701,n7702);
xor (n7701,n7698,n7699);
or (n7702,n7703,n7706);
and (n7703,n7704,n7705);
xor (n7704,n7611,n7612);
and (n7705,n1163,n69);
and (n7706,n7707,n7708);
xor (n7707,n7704,n7705);
or (n7708,n7709,n7712);
and (n7709,n7710,n7711);
xor (n7710,n7617,n7618);
and (n7711,n1639,n69);
and (n7712,n7713,n7714);
xor (n7713,n7710,n7711);
or (n7714,n7715,n7718);
and (n7715,n7716,n7717);
xor (n7716,n7623,n7624);
and (n7717,n1475,n69);
and (n7718,n7719,n7720);
xor (n7719,n7716,n7717);
and (n7720,n7721,n1496);
xor (n7721,n7629,n7630);
and (n7722,n358,n75);
and (n7723,n7724,n7725);
xor (n7724,n6836,n7722);
or (n7725,n7726,n7729);
and (n7726,n7727,n7728);
xor (n7727,n7635,n7636);
and (n7728,n85,n75);
and (n7729,n7730,n7731);
xor (n7730,n7727,n7728);
or (n7731,n7732,n7735);
and (n7732,n7733,n7734);
xor (n7733,n7641,n7642);
and (n7734,n79,n75);
and (n7735,n7736,n7737);
xor (n7736,n7733,n7734);
or (n7737,n7738,n7741);
and (n7738,n7739,n7740);
xor (n7739,n7647,n7648);
and (n7740,n489,n75);
and (n7741,n7742,n7743);
xor (n7742,n7739,n7740);
or (n7743,n7744,n7747);
and (n7744,n7745,n7746);
xor (n7745,n7653,n7654);
and (n7746,n483,n75);
and (n7747,n7748,n7749);
xor (n7748,n7745,n7746);
or (n7749,n7750,n7753);
and (n7750,n7751,n7752);
xor (n7751,n7659,n7660);
and (n7752,n341,n75);
and (n7753,n7754,n7755);
xor (n7754,n7751,n7752);
or (n7755,n7756,n7758);
and (n7756,n7757,n4176);
xor (n7757,n7665,n7666);
and (n7758,n7759,n7760);
xor (n7759,n7757,n4176);
or (n7760,n7761,n7763);
and (n7761,n7762,n4514);
xor (n7762,n7671,n7672);
and (n7763,n7764,n7765);
xor (n7764,n7762,n4514);
or (n7765,n7766,n7768);
and (n7766,n7767,n4040);
xor (n7767,n7677,n7678);
and (n7768,n7769,n7770);
xor (n7769,n7767,n4040);
or (n7770,n7771,n7773);
and (n7771,n7772,n3687);
xor (n7772,n7683,n7684);
and (n7773,n7774,n7775);
xor (n7774,n7772,n3687);
or (n7775,n7776,n7778);
and (n7776,n7777,n1783);
xor (n7777,n7689,n7690);
and (n7778,n7779,n7780);
xor (n7779,n7777,n1783);
or (n7780,n7781,n7784);
and (n7781,n7782,n7783);
xor (n7782,n7695,n7696);
and (n7783,n1169,n75);
and (n7784,n7785,n7786);
xor (n7785,n7782,n7783);
or (n7786,n7787,n7789);
and (n7787,n7788,n1164);
xor (n7788,n7701,n7702);
and (n7789,n7790,n7791);
xor (n7790,n7788,n1164);
or (n7791,n7792,n7795);
and (n7792,n7793,n7794);
xor (n7793,n7707,n7708);
and (n7794,n1639,n75);
and (n7795,n7796,n7797);
xor (n7796,n7793,n7794);
or (n7797,n7798,n7801);
and (n7798,n7799,n7800);
xor (n7799,n7713,n7714);
and (n7800,n1475,n75);
and (n7801,n7802,n7803);
xor (n7802,n7799,n7800);
and (n7803,n7804,n7805);
xor (n7804,n7719,n7720);
and (n7805,n1470,n75);
and (n7806,n358,n335);
or (n7807,n7808,n7811);
and (n7808,n7809,n7810);
xor (n7809,n7724,n7725);
and (n7810,n85,n335);
and (n7811,n7812,n7813);
xor (n7812,n7809,n7810);
or (n7813,n7814,n7817);
and (n7814,n7815,n7816);
xor (n7815,n7730,n7731);
and (n7816,n79,n335);
and (n7817,n7818,n7819);
xor (n7818,n7815,n7816);
or (n7819,n7820,n7823);
and (n7820,n7821,n7822);
xor (n7821,n7736,n7737);
and (n7822,n489,n335);
and (n7823,n7824,n7825);
xor (n7824,n7821,n7822);
or (n7825,n7826,n7829);
and (n7826,n7827,n7828);
xor (n7827,n7742,n7743);
and (n7828,n483,n335);
and (n7829,n7830,n7831);
xor (n7830,n7827,n7828);
or (n7831,n7832,n7835);
and (n7832,n7833,n7834);
xor (n7833,n7748,n7749);
and (n7834,n341,n335);
and (n7835,n7836,n7837);
xor (n7836,n7833,n7834);
or (n7837,n7838,n7841);
and (n7838,n7839,n7840);
xor (n7839,n7754,n7755);
and (n7840,n348,n335);
and (n7841,n7842,n7843);
xor (n7842,n7839,n7840);
or (n7843,n7844,n7847);
and (n7844,n7845,n7846);
xor (n7845,n7759,n7760);
and (n7846,n134,n335);
and (n7847,n7848,n7849);
xor (n7848,n7845,n7846);
or (n7849,n7850,n7853);
and (n7850,n7851,n7852);
xor (n7851,n7764,n7765);
and (n7852,n114,n335);
and (n7853,n7854,n7855);
xor (n7854,n7851,n7852);
or (n7855,n7856,n7859);
and (n7856,n7857,n7858);
xor (n7857,n7769,n7770);
and (n7858,n928,n335);
and (n7859,n7860,n7861);
xor (n7860,n7857,n7858);
or (n7861,n7862,n7865);
and (n7862,n7863,n7864);
xor (n7863,n7774,n7775);
and (n7864,n1357,n335);
and (n7865,n7866,n7867);
xor (n7866,n7863,n7864);
or (n7867,n7868,n7871);
and (n7868,n7869,n7870);
xor (n7869,n7779,n7780);
and (n7870,n1169,n335);
and (n7871,n7872,n7873);
xor (n7872,n7869,n7870);
or (n7873,n7874,n7877);
and (n7874,n7875,n7876);
xor (n7875,n7785,n7786);
and (n7876,n1163,n335);
and (n7877,n7878,n7879);
xor (n7878,n7875,n7876);
or (n7879,n7880,n7883);
and (n7880,n7881,n7882);
xor (n7881,n7790,n7791);
and (n7882,n1639,n335);
and (n7883,n7884,n7885);
xor (n7884,n7881,n7882);
or (n7885,n7886,n7889);
and (n7886,n7887,n7888);
xor (n7887,n7796,n7797);
and (n7888,n1475,n335);
and (n7889,n7890,n7891);
xor (n7890,n7887,n7888);
and (n7891,n7892,n7893);
xor (n7892,n7802,n7803);
not (n7893,n1565);
and (n7894,n85,n128);
or (n7895,n7896,n7898);
and (n7896,n7897,n752);
xor (n7897,n7812,n7813);
and (n7898,n7899,n7900);
xor (n7899,n7897,n752);
or (n7900,n7901,n7904);
and (n7901,n7902,n7903);
xor (n7902,n7818,n7819);
and (n7903,n489,n128);
and (n7904,n7905,n7906);
xor (n7905,n7902,n7903);
or (n7906,n7907,n7909);
and (n7907,n7908,n536);
xor (n7908,n7824,n7825);
and (n7909,n7910,n7911);
xor (n7910,n7908,n536);
or (n7911,n7912,n7915);
and (n7912,n7913,n7914);
xor (n7913,n7830,n7831);
and (n7914,n341,n128);
and (n7915,n7916,n7917);
xor (n7916,n7913,n7914);
or (n7917,n7918,n7921);
and (n7918,n7919,n7920);
xor (n7919,n7836,n7837);
and (n7920,n348,n128);
and (n7921,n7922,n7923);
xor (n7922,n7919,n7920);
or (n7923,n7924,n7927);
and (n7924,n7925,n7926);
xor (n7925,n7842,n7843);
and (n7926,n134,n128);
and (n7927,n7928,n7929);
xor (n7928,n7925,n7926);
or (n7929,n7930,n7933);
and (n7930,n7931,n7932);
xor (n7931,n7848,n7849);
and (n7932,n114,n128);
and (n7933,n7934,n7935);
xor (n7934,n7931,n7932);
or (n7935,n7936,n7939);
and (n7936,n7937,n7938);
xor (n7937,n7854,n7855);
and (n7938,n928,n128);
and (n7939,n7940,n7941);
xor (n7940,n7937,n7938);
or (n7941,n7942,n7945);
and (n7942,n7943,n7944);
xor (n7943,n7860,n7861);
and (n7944,n1357,n128);
and (n7945,n7946,n7947);
xor (n7946,n7943,n7944);
or (n7947,n7948,n7951);
and (n7948,n7949,n7950);
xor (n7949,n7866,n7867);
and (n7950,n1169,n128);
and (n7951,n7952,n7953);
xor (n7952,n7949,n7950);
or (n7953,n7954,n7957);
and (n7954,n7955,n7956);
xor (n7955,n7872,n7873);
and (n7956,n1163,n128);
and (n7957,n7958,n7959);
xor (n7958,n7955,n7956);
or (n7959,n7960,n7963);
and (n7960,n7961,n7962);
xor (n7961,n7878,n7879);
and (n7962,n1639,n128);
and (n7963,n7964,n7965);
xor (n7964,n7961,n7962);
or (n7965,n7966,n7968);
and (n7966,n7967,n1635);
xor (n7967,n7884,n7885);
and (n7968,n7969,n7970);
xor (n7969,n7967,n1635);
and (n7970,n7971,n2019);
xor (n7971,n7890,n7891);
and (n7972,n79,n122);
or (n7973,n7974,n7977);
and (n7974,n7975,n7976);
xor (n7975,n7899,n7900);
and (n7976,n489,n122);
and (n7977,n7978,n7979);
xor (n7978,n7975,n7976);
or (n7979,n7980,n7983);
and (n7980,n7981,n7982);
xor (n7981,n7905,n7906);
and (n7982,n483,n122);
and (n7983,n7984,n7985);
xor (n7984,n7981,n7982);
or (n7985,n7986,n7989);
and (n7986,n7987,n7988);
xor (n7987,n7910,n7911);
and (n7988,n341,n122);
and (n7989,n7990,n7991);
xor (n7990,n7987,n7988);
or (n7991,n7992,n7995);
and (n7992,n7993,n7994);
xor (n7993,n7916,n7917);
and (n7994,n348,n122);
and (n7995,n7996,n7997);
xor (n7996,n7993,n7994);
or (n7997,n7998,n8001);
and (n7998,n7999,n8000);
xor (n7999,n7922,n7923);
and (n8000,n134,n122);
and (n8001,n8002,n8003);
xor (n8002,n7999,n8000);
or (n8003,n8004,n8007);
and (n8004,n8005,n8006);
xor (n8005,n7928,n7929);
and (n8006,n114,n122);
and (n8007,n8008,n8009);
xor (n8008,n8005,n8006);
or (n8009,n8010,n8013);
and (n8010,n8011,n8012);
xor (n8011,n7934,n7935);
and (n8012,n928,n122);
and (n8013,n8014,n8015);
xor (n8014,n8011,n8012);
or (n8015,n8016,n8019);
and (n8016,n8017,n8018);
xor (n8017,n7940,n7941);
and (n8018,n1357,n122);
and (n8019,n8020,n8021);
xor (n8020,n8017,n8018);
or (n8021,n8022,n8025);
and (n8022,n8023,n8024);
xor (n8023,n7946,n7947);
and (n8024,n1169,n122);
and (n8025,n8026,n8027);
xor (n8026,n8023,n8024);
or (n8027,n8028,n8031);
and (n8028,n8029,n8030);
xor (n8029,n7952,n7953);
and (n8030,n1163,n122);
and (n8031,n8032,n8033);
xor (n8032,n8029,n8030);
or (n8033,n8034,n8037);
and (n8034,n8035,n8036);
xor (n8035,n7958,n7959);
and (n8036,n1639,n122);
and (n8037,n8038,n8039);
xor (n8038,n8035,n8036);
or (n8039,n8040,n8043);
and (n8040,n8041,n8042);
xor (n8041,n7964,n7965);
and (n8042,n1475,n122);
and (n8043,n8044,n8045);
xor (n8044,n8041,n8042);
and (n8045,n8046,n8047);
xor (n8046,n7969,n7970);
not (n8047,n1881);
and (n8048,n489,n116);
or (n8049,n8050,n8053);
and (n8050,n8051,n8052);
xor (n8051,n7978,n7979);
and (n8052,n483,n116);
and (n8053,n8054,n8055);
xor (n8054,n8051,n8052);
or (n8055,n8056,n8059);
and (n8056,n8057,n8058);
xor (n8057,n7984,n7985);
and (n8058,n341,n116);
and (n8059,n8060,n8061);
xor (n8060,n8057,n8058);
or (n8061,n8062,n8064);
and (n8062,n8063,n513);
xor (n8063,n7990,n7991);
and (n8064,n8065,n8066);
xor (n8065,n8063,n513);
or (n8066,n8067,n8069);
and (n8067,n8068,n135);
xor (n8068,n7996,n7997);
and (n8069,n8070,n8071);
xor (n8070,n8068,n135);
or (n8071,n8072,n8075);
and (n8072,n8073,n8074);
xor (n8073,n8002,n8003);
and (n8074,n114,n116);
and (n8075,n8076,n8077);
xor (n8076,n8073,n8074);
or (n8077,n8078,n8080);
and (n8078,n8079,n929);
xor (n8079,n8008,n8009);
and (n8080,n8081,n8082);
xor (n8081,n8079,n929);
or (n8082,n8083,n8085);
and (n8083,n8084,n4645);
xor (n8084,n8014,n8015);
and (n8085,n8086,n8087);
xor (n8086,n8084,n4645);
or (n8087,n8088,n8090);
and (n8088,n8089,n4369);
xor (n8089,n8020,n8021);
and (n8090,n8091,n8092);
xor (n8091,n8089,n4369);
or (n8092,n8093,n8095);
and (n8093,n8094,n3915);
xor (n8094,n8026,n8027);
and (n8095,n8096,n8097);
xor (n8096,n8094,n3915);
or (n8097,n8098,n8101);
and (n8098,n8099,n8100);
xor (n8099,n8032,n8033);
and (n8100,n1639,n116);
and (n8101,n8102,n8103);
xor (n8102,n8099,n8100);
or (n8103,n8104,n8106);
and (n8104,n8105,n1754);
xor (n8105,n8038,n8039);
and (n8106,n8107,n8108);
xor (n8107,n8105,n1754);
and (n8108,n8109,n1750);
xor (n8109,n8044,n8045);
or (n8110,n8111,n8113);
and (n8111,n8112,n8058);
xor (n8112,n8054,n8055);
and (n8113,n8114,n8115);
xor (n8114,n8112,n8058);
or (n8115,n8116,n8118);
and (n8116,n8117,n513);
xor (n8117,n8060,n8061);
and (n8118,n8119,n8120);
xor (n8119,n8117,n513);
or (n8120,n8121,n8123);
and (n8121,n8122,n135);
xor (n8122,n8065,n8066);
and (n8123,n8124,n8125);
xor (n8124,n8122,n135);
or (n8125,n8126,n8128);
and (n8126,n8127,n8074);
xor (n8127,n8070,n8071);
and (n8128,n8129,n8130);
xor (n8129,n8127,n8074);
or (n8130,n8131,n8133);
and (n8131,n8132,n929);
xor (n8132,n8076,n8077);
and (n8133,n8134,n8135);
xor (n8134,n8132,n929);
or (n8135,n8136,n8138);
and (n8136,n8137,n4645);
xor (n8137,n8081,n8082);
and (n8138,n8139,n8140);
xor (n8139,n8137,n4645);
or (n8140,n8141,n8143);
and (n8141,n8142,n4369);
xor (n8142,n8086,n8087);
and (n8143,n8144,n8145);
xor (n8144,n8142,n4369);
or (n8145,n8146,n8148);
and (n8146,n8147,n3915);
xor (n8147,n8091,n8092);
and (n8148,n8149,n8150);
xor (n8149,n8147,n3915);
or (n8150,n8151,n8153);
and (n8151,n8152,n8100);
xor (n8152,n8096,n8097);
and (n8153,n8154,n8155);
xor (n8154,n8152,n8100);
or (n8155,n8156,n8158);
and (n8156,n8157,n1754);
xor (n8157,n8102,n8103);
and (n8158,n8159,n8160);
xor (n8159,n8157,n1754);
and (n8160,n8161,n1750);
xor (n8161,n8107,n8108);
or (n8162,n8163,n8165);
and (n8163,n8164,n513);
xor (n8164,n8114,n8115);
and (n8165,n8166,n8167);
xor (n8166,n8164,n513);
or (n8167,n8168,n8170);
and (n8168,n8169,n135);
xor (n8169,n8119,n8120);
and (n8170,n8171,n8172);
xor (n8171,n8169,n135);
or (n8172,n8173,n8175);
and (n8173,n8174,n8074);
xor (n8174,n8124,n8125);
and (n8175,n8176,n8177);
xor (n8176,n8174,n8074);
or (n8177,n8178,n8180);
and (n8178,n8179,n929);
xor (n8179,n8129,n8130);
and (n8180,n8181,n8182);
xor (n8181,n8179,n929);
or (n8182,n8183,n8185);
and (n8183,n8184,n4645);
xor (n8184,n8134,n8135);
and (n8185,n8186,n8187);
xor (n8186,n8184,n4645);
or (n8187,n8188,n8190);
and (n8188,n8189,n4369);
xor (n8189,n8139,n8140);
and (n8190,n8191,n8192);
xor (n8191,n8189,n4369);
or (n8192,n8193,n8195);
and (n8193,n8194,n3915);
xor (n8194,n8144,n8145);
and (n8195,n8196,n8197);
xor (n8196,n8194,n3915);
or (n8197,n8198,n8200);
and (n8198,n8199,n8100);
xor (n8199,n8149,n8150);
and (n8200,n8201,n8202);
xor (n8201,n8199,n8100);
or (n8202,n8203,n8205);
and (n8203,n8204,n1754);
xor (n8204,n8154,n8155);
and (n8205,n8206,n8207);
xor (n8206,n8204,n1754);
and (n8207,n8208,n1750);
xor (n8208,n8159,n8160);
or (n8209,n8210,n8212);
and (n8210,n8211,n135);
xor (n8211,n8166,n8167);
and (n8212,n8213,n8214);
xor (n8213,n8211,n135);
or (n8214,n8215,n8217);
and (n8215,n8216,n8074);
xor (n8216,n8171,n8172);
and (n8217,n8218,n8219);
xor (n8218,n8216,n8074);
or (n8219,n8220,n8222);
and (n8220,n8221,n929);
xor (n8221,n8176,n8177);
and (n8222,n8223,n8224);
xor (n8223,n8221,n929);
or (n8224,n8225,n8227);
and (n8225,n8226,n4645);
xor (n8226,n8181,n8182);
and (n8227,n8228,n8229);
xor (n8228,n8226,n4645);
or (n8229,n8230,n8232);
and (n8230,n8231,n4369);
xor (n8231,n8186,n8187);
and (n8232,n8233,n8234);
xor (n8233,n8231,n4369);
or (n8234,n8235,n8237);
and (n8235,n8236,n3915);
xor (n8236,n8191,n8192);
and (n8237,n8238,n8239);
xor (n8238,n8236,n3915);
or (n8239,n8240,n8242);
and (n8240,n8241,n8100);
xor (n8241,n8196,n8197);
and (n8242,n8243,n8244);
xor (n8243,n8241,n8100);
or (n8244,n8245,n8247);
and (n8245,n8246,n1754);
xor (n8246,n8201,n8202);
and (n8247,n8248,n8249);
xor (n8248,n8246,n1754);
and (n8249,n8250,n1750);
xor (n8250,n8206,n8207);
or (n8251,n8252,n8254);
and (n8252,n8253,n8074);
xor (n8253,n8213,n8214);
and (n8254,n8255,n8256);
xor (n8255,n8253,n8074);
or (n8256,n8257,n8259);
and (n8257,n8258,n929);
xor (n8258,n8218,n8219);
and (n8259,n8260,n8261);
xor (n8260,n8258,n929);
or (n8261,n8262,n8264);
and (n8262,n8263,n4645);
xor (n8263,n8223,n8224);
and (n8264,n8265,n8266);
xor (n8265,n8263,n4645);
or (n8266,n8267,n8269);
and (n8267,n8268,n4369);
xor (n8268,n8228,n8229);
and (n8269,n8270,n8271);
xor (n8270,n8268,n4369);
or (n8271,n8272,n8274);
and (n8272,n8273,n3915);
xor (n8273,n8233,n8234);
and (n8274,n8275,n8276);
xor (n8275,n8273,n3915);
or (n8276,n8277,n8279);
and (n8277,n8278,n8100);
xor (n8278,n8238,n8239);
and (n8279,n8280,n8281);
xor (n8280,n8278,n8100);
or (n8281,n8282,n8284);
and (n8282,n8283,n1754);
xor (n8283,n8243,n8244);
and (n8284,n8285,n8286);
xor (n8285,n8283,n1754);
and (n8286,n8287,n1750);
xor (n8287,n8248,n8249);
or (n8288,n8289,n8291);
and (n8289,n8290,n929);
xor (n8290,n8255,n8256);
and (n8291,n8292,n8293);
xor (n8292,n8290,n929);
or (n8293,n8294,n8296);
and (n8294,n8295,n4645);
xor (n8295,n8260,n8261);
and (n8296,n8297,n8298);
xor (n8297,n8295,n4645);
or (n8298,n8299,n8301);
and (n8299,n8300,n4369);
xor (n8300,n8265,n8266);
and (n8301,n8302,n8303);
xor (n8302,n8300,n4369);
or (n8303,n8304,n8306);
and (n8304,n8305,n3915);
xor (n8305,n8270,n8271);
and (n8306,n8307,n8308);
xor (n8307,n8305,n3915);
or (n8308,n8309,n8311);
and (n8309,n8310,n8100);
xor (n8310,n8275,n8276);
and (n8311,n8312,n8313);
xor (n8312,n8310,n8100);
or (n8313,n8314,n8316);
and (n8314,n8315,n1754);
xor (n8315,n8280,n8281);
and (n8316,n8317,n8318);
xor (n8317,n8315,n1754);
and (n8318,n8319,n1750);
xor (n8319,n8285,n8286);
or (n8320,n8321,n8323);
and (n8321,n8322,n4645);
xor (n8322,n8292,n8293);
and (n8323,n8324,n8325);
xor (n8324,n8322,n4645);
or (n8325,n8326,n8328);
and (n8326,n8327,n4369);
xor (n8327,n8297,n8298);
and (n8328,n8329,n8330);
xor (n8329,n8327,n4369);
or (n8330,n8331,n8333);
and (n8331,n8332,n3915);
xor (n8332,n8302,n8303);
and (n8333,n8334,n8335);
xor (n8334,n8332,n3915);
or (n8335,n8336,n8338);
and (n8336,n8337,n8100);
xor (n8337,n8307,n8308);
and (n8338,n8339,n8340);
xor (n8339,n8337,n8100);
or (n8340,n8341,n8343);
and (n8341,n8342,n1754);
xor (n8342,n8312,n8313);
and (n8343,n8344,n8345);
xor (n8344,n8342,n1754);
and (n8345,n8346,n1750);
xor (n8346,n8317,n8318);
or (n8347,n8348,n8350);
and (n8348,n8349,n4369);
xor (n8349,n8324,n8325);
and (n8350,n8351,n8352);
xor (n8351,n8349,n4369);
or (n8352,n8353,n8355);
and (n8353,n8354,n3915);
xor (n8354,n8329,n8330);
and (n8355,n8356,n8357);
xor (n8356,n8354,n3915);
or (n8357,n8358,n8360);
and (n8358,n8359,n8100);
xor (n8359,n8334,n8335);
and (n8360,n8361,n8362);
xor (n8361,n8359,n8100);
or (n8362,n8363,n8365);
and (n8363,n8364,n1754);
xor (n8364,n8339,n8340);
and (n8365,n8366,n8367);
xor (n8366,n8364,n1754);
and (n8367,n8368,n1750);
xor (n8368,n8344,n8345);
or (n8369,n8370,n8372);
and (n8370,n8371,n3915);
xor (n8371,n8351,n8352);
and (n8372,n8373,n8374);
xor (n8373,n8371,n3915);
or (n8374,n8375,n8377);
and (n8375,n8376,n8100);
xor (n8376,n8356,n8357);
and (n8377,n8378,n8379);
xor (n8378,n8376,n8100);
or (n8379,n8380,n8382);
and (n8380,n8381,n1754);
xor (n8381,n8361,n8362);
and (n8382,n8383,n8384);
xor (n8383,n8381,n1754);
and (n8384,n8385,n1750);
xor (n8385,n8366,n8367);
or (n8386,n8387,n8389);
and (n8387,n8388,n8100);
xor (n8388,n8373,n8374);
and (n8389,n8390,n8391);
xor (n8390,n8388,n8100);
or (n8391,n8392,n8394);
and (n8392,n8393,n1754);
xor (n8393,n8378,n8379);
and (n8394,n8395,n8396);
xor (n8395,n8393,n1754);
and (n8396,n8397,n1750);
xor (n8397,n8383,n8384);
or (n8398,n8399,n8401);
and (n8399,n8400,n1754);
xor (n8400,n8390,n8391);
and (n8401,n8402,n8403);
xor (n8402,n8400,n1754);
and (n8403,n8404,n1750);
xor (n8404,n8395,n8396);
and (n8405,n8406,n1750);
xor (n8406,n8402,n8403);
or (n8407,n8408,n8411,n8562);
and (n8408,n8409,n8410);
xor (n8409,n6802,n6505);
xor (n8410,n8406,n1750);
and (n8411,n8410,n8412);
or (n8412,n8413,n8416,n8561);
and (n8413,n8414,n8415);
xor (n8414,n6800,n6505);
xor (n8415,n8404,n1750);
and (n8416,n8415,n8417);
or (n8417,n8418,n8421,n8560);
and (n8418,n8419,n8420);
xor (n8419,n6793,n6505);
xor (n8420,n8397,n1750);
and (n8421,n8420,n8422);
or (n8422,n8423,n8426,n8559);
and (n8423,n8424,n8425);
xor (n8424,n6781,n6505);
xor (n8425,n8385,n1750);
and (n8426,n8425,n8427);
or (n8427,n8428,n8431,n8558);
and (n8428,n8429,n8430);
xor (n8429,n6764,n6505);
xor (n8430,n8368,n1750);
and (n8431,n8430,n8432);
or (n8432,n8433,n8436,n8557);
and (n8433,n8434,n8435);
xor (n8434,n6742,n6505);
xor (n8435,n8346,n1750);
and (n8436,n8435,n8437);
or (n8437,n8438,n8441,n8556);
and (n8438,n8439,n8440);
xor (n8439,n6715,n6505);
xor (n8440,n8319,n1750);
and (n8441,n8440,n8442);
or (n8442,n8443,n8446,n8555);
and (n8443,n8444,n8445);
xor (n8444,n6683,n6505);
xor (n8445,n8287,n1750);
and (n8446,n8445,n8447);
or (n8447,n8448,n8451,n8554);
and (n8448,n8449,n8450);
xor (n8449,n6646,n6505);
xor (n8450,n8250,n1750);
and (n8451,n8450,n8452);
or (n8452,n8453,n8456,n8553);
and (n8453,n8454,n8455);
xor (n8454,n6604,n6505);
xor (n8455,n8208,n1750);
and (n8456,n8455,n8457);
or (n8457,n8458,n8461,n8552);
and (n8458,n8459,n8460);
xor (n8459,n6557,n6505);
xor (n8460,n8161,n1750);
and (n8461,n8460,n8462);
or (n8462,n8463,n8466,n8551);
and (n8463,n8464,n8465);
xor (n8464,n6504,n6505);
xor (n8465,n8109,n1750);
and (n8466,n8465,n8467);
or (n8467,n8468,n8471,n8550);
and (n8468,n8469,n8470);
xor (n8469,n6438,n1876);
xor (n8470,n8046,n8047);
and (n8471,n8470,n8472);
or (n8472,n8473,n8476,n8549);
and (n8473,n8474,n8475);
xor (n8474,n6362,n6363);
xor (n8475,n7971,n2019);
and (n8476,n8475,n8477);
or (n8477,n8478,n8481,n8548);
and (n8478,n8479,n8480);
xor (n8479,n6285,n6286);
xor (n8480,n7892,n7893);
and (n8481,n8480,n8482);
or (n8482,n8483,n8486,n8547);
and (n8483,n8484,n8485);
xor (n8484,n6197,n6198);
xor (n8485,n7804,n7805);
and (n8486,n8485,n8487);
or (n8487,n8488,n8491,n8546);
and (n8488,n8489,n8490);
xor (n8489,n6110,n6111);
xor (n8490,n7721,n1496);
and (n8491,n8490,n8492);
or (n8492,n8493,n8496,n8545);
and (n8493,n8494,n8495);
xor (n8494,n6020,n6021);
xor (n8495,n7631,n7632);
and (n8496,n8495,n8497);
or (n8497,n8498,n8501,n8544);
and (n8498,n8499,n8500);
xor (n8499,n5937,n2590);
xor (n8500,n7548,n7549);
and (n8501,n8500,n8502);
or (n8502,n8503,n8506,n8543);
and (n8503,n8504,n8505);
xor (n8504,n5847,n5848);
xor (n8505,n7458,n7459);
and (n8506,n8505,n8507);
or (n8507,n8508,n8511,n8542);
and (n8508,n8509,n8510);
xor (n8509,n5760,n5761);
xor (n8510,n7375,n2862);
and (n8511,n8510,n8512);
or (n8512,n8513,n8516,n8541);
and (n8513,n8514,n8515);
xor (n8514,n5670,n5671);
xor (n8515,n7285,n7286);
and (n8516,n8515,n8517);
or (n8517,n8518,n8521,n8540);
and (n8518,n8519,n8520);
xor (n8519,n5590,n3147);
xor (n8520,n7197,n7198);
and (n8521,n8520,n8522);
or (n8522,n8523,n8526,n8539);
and (n8523,n8524,n8525);
xor (n8524,n5500,n5501);
xor (n8525,n7107,n7108);
and (n8526,n8525,n8527);
or (n8527,n8528,n8531,n8538);
and (n8528,n8529,n8530);
xor (n8529,n5413,n5414);
xor (n8530,n7024,n3408);
and (n8531,n8530,n8532);
or (n8532,n8533,n8536,n8537);
and (n8533,n8534,n8535);
xor (n8534,n5323,n5324);
xor (n8535,n6934,n6935);
and (n8536,n8535,n3562);
and (n8537,n8534,n3562);
and (n8538,n8529,n8532);
and (n8539,n8524,n8527);
and (n8540,n8519,n8522);
and (n8541,n8514,n8517);
and (n8542,n8509,n8512);
and (n8543,n8504,n8507);
and (n8544,n8499,n8502);
and (n8545,n8494,n8497);
and (n8546,n8489,n8492);
and (n8547,n8484,n8487);
and (n8548,n8479,n8482);
and (n8549,n8474,n8477);
and (n8550,n8469,n8472);
and (n8551,n8464,n8467);
and (n8552,n8459,n8462);
and (n8553,n8454,n8457);
and (n8554,n8449,n8452);
and (n8555,n8444,n8447);
and (n8556,n8439,n8442);
and (n8557,n8434,n8437);
and (n8558,n8429,n8432);
and (n8559,n8424,n8427);
and (n8560,n8419,n8422);
and (n8561,n8414,n8417);
and (n8562,n8409,n8412);
xor (n8563,n8564,n1701);
xor (n8564,n8565,n10228);
xor (n8565,n8566,n9928);
xor (n8566,n8567,n10221);
xor (n8567,n8568,n9922);
xor (n8568,n8569,n10209);
xor (n8569,n8570,n9916);
xor (n8570,n8571,n10192);
xor (n8571,n8572,n4362);
xor (n8572,n8573,n10170);
xor (n8573,n8574,n4588);
xor (n8574,n8575,n10143);
xor (n8575,n8576,n957);
xor (n8576,n8577,n10111);
xor (n8577,n8578,n9895);
xor (n8578,n8579,n10074);
xor (n8579,n8580,n9889);
xor (n8580,n8581,n10032);
xor (n8581,n8582,n9883);
xor (n8582,n8583,n9985);
xor (n8583,n8584,n9877);
xor (n8584,n8585,n9933);
xor (n8585,n8586,n9871);
xor (n8586,n8587,n9868);
xor (n8587,n8588,n9867);
xor (n8588,n8589,n9793);
xor (n8589,n8590,n9792);
xor (n8590,n8591,n9715);
xor (n8591,n8592,n9714);
xor (n8592,n8593,n9628);
xor (n8593,n8594,n9627);
xor (n8594,n8595,n9540);
xor (n8595,n8596,n9539);
or (n8596,n8597,n9445);
and (n8597,n8598,n9444);
or (n8598,n8599,n9356);
and (n8599,n8600,n653);
or (n8600,n8601,n9262);
and (n8601,n8602,n9261);
or (n8602,n8603,n9172);
and (n8603,n8604,n9171);
or (n8604,n8605,n9077);
and (n8605,n8606,n9076);
or (n8606,n8607,n8985);
and (n8607,n8608,n8984);
or (n8608,n8609,n8889);
and (n8609,n8610,n8888);
or (n8610,n8611,n8798);
and (n8611,n8612,n4417);
or (n8612,n8613,n8703);
and (n8613,n8614,n8702);
and (n8614,n3786,n8615);
or (n8615,n8616,n8618);
and (n8616,n8617,n1775);
and (n8617,n193,n1197);
and (n8618,n8619,n8620);
xor (n8619,n8617,n1775);
or (n8620,n8621,n8623);
and (n8621,n8622,n1202);
and (n8622,n186,n1197);
and (n8623,n8624,n8625);
xor (n8624,n8622,n1202);
or (n8625,n8626,n8629);
and (n8626,n8627,n8628);
and (n8627,n328,n1197);
and (n8628,n313,n1192);
and (n8629,n8630,n8631);
xor (n8630,n8627,n8628);
or (n8631,n8632,n8634);
and (n8632,n8633,n1926);
and (n8633,n313,n1197);
and (n8634,n8635,n8636);
xor (n8635,n8633,n1926);
or (n8636,n8637,n8640);
and (n8637,n8638,n8639);
and (n8638,n297,n1197);
and (n8639,n279,n1192);
and (n8640,n8641,n8642);
xor (n8641,n8638,n8639);
or (n8642,n8643,n8646);
and (n8643,n8644,n8645);
and (n8644,n279,n1197);
and (n8645,n59,n1192);
and (n8646,n8647,n8648);
xor (n8647,n8644,n8645);
or (n8648,n8649,n8651);
and (n8649,n8650,n2327);
and (n8650,n59,n1197);
and (n8651,n8652,n8653);
xor (n8652,n8650,n2327);
or (n8653,n8654,n8657);
and (n8654,n8655,n8656);
and (n8655,n53,n1197);
and (n8656,n222,n1192);
and (n8657,n8658,n8659);
xor (n8658,n8655,n8656);
or (n8659,n8660,n8663);
and (n8660,n8661,n8662);
and (n8661,n222,n1197);
and (n8662,n215,n1192);
and (n8663,n8664,n8665);
xor (n8664,n8661,n8662);
or (n8665,n8666,n8669);
and (n8666,n8667,n8668);
and (n8667,n215,n1197);
and (n8668,n956,n1192);
and (n8669,n8670,n8671);
xor (n8670,n8667,n8668);
or (n8671,n8672,n8675);
and (n8672,n8673,n8674);
and (n8673,n956,n1197);
and (n8674,n1305,n1192);
and (n8675,n8676,n8677);
xor (n8676,n8673,n8674);
or (n8677,n8678,n8680);
and (n8678,n8679,n3172);
and (n8679,n1305,n1197);
and (n8680,n8681,n8682);
xor (n8681,n8679,n3172);
or (n8682,n8683,n8685);
and (n8683,n8684,n3329);
and (n8684,n1131,n1197);
and (n8685,n8686,n8687);
xor (n8686,n8684,n3329);
or (n8687,n8688,n8691);
and (n8688,n8689,n8690);
and (n8689,n1125,n1197);
and (n8690,n1250,n1192);
and (n8691,n8692,n8693);
xor (n8692,n8689,n8690);
or (n8693,n8694,n8697);
and (n8694,n8695,n8696);
and (n8695,n1250,n1197);
and (n8696,n1244,n1192);
and (n8697,n8698,n8699);
xor (n8698,n8695,n8696);
and (n8699,n8700,n8701);
and (n8700,n1244,n1197);
and (n8701,n1377,n1192);
and (n8702,n193,n1595);
and (n8703,n8704,n8705);
xor (n8704,n8614,n8702);
or (n8705,n8706,n8709);
and (n8706,n8707,n8708);
xor (n8707,n3786,n8615);
and (n8708,n186,n1595);
and (n8709,n8710,n8711);
xor (n8710,n8707,n8708);
or (n8711,n8712,n8715);
and (n8712,n8713,n8714);
xor (n8713,n8619,n8620);
and (n8714,n328,n1595);
and (n8715,n8716,n8717);
xor (n8716,n8713,n8714);
or (n8717,n8718,n8721);
and (n8718,n8719,n8720);
xor (n8719,n8624,n8625);
and (n8720,n313,n1595);
and (n8721,n8722,n8723);
xor (n8722,n8719,n8720);
or (n8723,n8724,n8727);
and (n8724,n8725,n8726);
xor (n8725,n8630,n8631);
and (n8726,n297,n1595);
and (n8727,n8728,n8729);
xor (n8728,n8725,n8726);
or (n8729,n8730,n8733);
and (n8730,n8731,n8732);
xor (n8731,n8635,n8636);
and (n8732,n279,n1595);
and (n8733,n8734,n8735);
xor (n8734,n8731,n8732);
or (n8735,n8736,n8739);
and (n8736,n8737,n8738);
xor (n8737,n8641,n8642);
and (n8738,n59,n1595);
and (n8739,n8740,n8741);
xor (n8740,n8737,n8738);
or (n8741,n8742,n8745);
and (n8742,n8743,n8744);
xor (n8743,n8647,n8648);
and (n8744,n53,n1595);
and (n8745,n8746,n8747);
xor (n8746,n8743,n8744);
or (n8747,n8748,n8751);
and (n8748,n8749,n8750);
xor (n8749,n8652,n8653);
and (n8750,n222,n1595);
and (n8751,n8752,n8753);
xor (n8752,n8749,n8750);
or (n8753,n8754,n8757);
and (n8754,n8755,n8756);
xor (n8755,n8658,n8659);
and (n8756,n215,n1595);
and (n8757,n8758,n8759);
xor (n8758,n8755,n8756);
or (n8759,n8760,n8763);
and (n8760,n8761,n8762);
xor (n8761,n8664,n8665);
and (n8762,n956,n1595);
and (n8763,n8764,n8765);
xor (n8764,n8761,n8762);
or (n8765,n8766,n8769);
and (n8766,n8767,n8768);
xor (n8767,n8670,n8671);
and (n8768,n1305,n1595);
and (n8769,n8770,n8771);
xor (n8770,n8767,n8768);
or (n8771,n8772,n8775);
and (n8772,n8773,n8774);
xor (n8773,n8676,n8677);
and (n8774,n1131,n1595);
and (n8775,n8776,n8777);
xor (n8776,n8773,n8774);
or (n8777,n8778,n8781);
and (n8778,n8779,n8780);
xor (n8779,n8681,n8682);
and (n8780,n1125,n1595);
and (n8781,n8782,n8783);
xor (n8782,n8779,n8780);
or (n8783,n8784,n8787);
and (n8784,n8785,n8786);
xor (n8785,n8686,n8687);
and (n8786,n1250,n1595);
and (n8787,n8788,n8789);
xor (n8788,n8785,n8786);
or (n8789,n8790,n8793);
and (n8790,n8791,n8792);
xor (n8791,n8692,n8693);
and (n8792,n1244,n1595);
and (n8793,n8794,n8795);
xor (n8794,n8791,n8792);
and (n8795,n8796,n8797);
xor (n8796,n8698,n8699);
not (n8797,n3402);
and (n8798,n8799,n8800);
xor (n8799,n8612,n4417);
or (n8800,n8801,n8804);
and (n8801,n8802,n8803);
xor (n8802,n8704,n8705);
and (n8803,n186,n100);
and (n8804,n8805,n8806);
xor (n8805,n8802,n8803);
or (n8806,n8807,n8810);
and (n8807,n8808,n8809);
xor (n8808,n8710,n8711);
and (n8809,n328,n100);
and (n8810,n8811,n8812);
xor (n8811,n8808,n8809);
or (n8812,n8813,n8816);
and (n8813,n8814,n8815);
xor (n8814,n8716,n8717);
and (n8815,n313,n100);
and (n8816,n8817,n8818);
xor (n8817,n8814,n8815);
or (n8818,n8819,n8822);
and (n8819,n8820,n8821);
xor (n8820,n8722,n8723);
and (n8821,n297,n100);
and (n8822,n8823,n8824);
xor (n8823,n8820,n8821);
or (n8824,n8825,n8827);
and (n8825,n8826,n1647);
xor (n8826,n8728,n8729);
and (n8827,n8828,n8829);
xor (n8828,n8826,n1647);
or (n8829,n8830,n8832);
and (n8830,n8831,n1604);
xor (n8831,n8734,n8735);
and (n8832,n8833,n8834);
xor (n8833,n8831,n1604);
or (n8834,n8835,n8838);
and (n8835,n8836,n8837);
xor (n8836,n8740,n8741);
and (n8837,n53,n100);
and (n8838,n8839,n8840);
xor (n8839,n8836,n8837);
or (n8840,n8841,n8843);
and (n8841,n8842,n2154);
xor (n8842,n8746,n8747);
and (n8843,n8844,n8845);
xor (n8844,n8842,n2154);
or (n8845,n8846,n8849);
and (n8846,n8847,n8848);
xor (n8847,n8752,n8753);
and (n8848,n215,n100);
and (n8849,n8850,n8851);
xor (n8850,n8847,n8848);
or (n8851,n8852,n8855);
and (n8852,n8853,n8854);
xor (n8853,n8758,n8759);
and (n8854,n956,n100);
and (n8855,n8856,n8857);
xor (n8856,n8853,n8854);
or (n8857,n8858,n8860);
and (n8858,n8859,n2809);
xor (n8859,n8764,n8765);
and (n8860,n8861,n8862);
xor (n8861,n8859,n2809);
or (n8862,n8863,n8865);
and (n8863,n8864,n2959);
xor (n8864,n8770,n8771);
and (n8865,n8866,n8867);
xor (n8866,n8864,n2959);
or (n8867,n8868,n8871);
and (n8868,n8869,n8870);
xor (n8869,n8776,n8777);
and (n8870,n1125,n100);
and (n8871,n8872,n8873);
xor (n8872,n8869,n8870);
or (n8873,n8874,n8877);
and (n8874,n8875,n8876);
xor (n8875,n8782,n8783);
and (n8876,n1250,n100);
and (n8877,n8878,n8879);
xor (n8878,n8875,n8876);
or (n8879,n8880,n8883);
and (n8880,n8881,n8882);
xor (n8881,n8788,n8789);
and (n8882,n1244,n100);
and (n8883,n8884,n8885);
xor (n8884,n8881,n8882);
and (n8885,n8886,n8887);
xor (n8886,n8794,n8795);
and (n8887,n1377,n100);
and (n8888,n193,n99);
and (n8889,n8890,n8891);
xor (n8890,n8610,n8888);
or (n8891,n8892,n8895);
and (n8892,n8893,n8894);
xor (n8893,n8799,n8800);
and (n8894,n186,n99);
and (n8895,n8896,n8897);
xor (n8896,n8893,n8894);
or (n8897,n8898,n8901);
and (n8898,n8899,n8900);
xor (n8899,n8805,n8806);
and (n8900,n328,n99);
and (n8901,n8902,n8903);
xor (n8902,n8899,n8900);
or (n8903,n8904,n8907);
and (n8904,n8905,n8906);
xor (n8905,n8811,n8812);
and (n8906,n313,n99);
and (n8907,n8908,n8909);
xor (n8908,n8905,n8906);
or (n8909,n8910,n8913);
and (n8910,n8911,n8912);
xor (n8911,n8817,n8818);
and (n8912,n297,n99);
and (n8913,n8914,n8915);
xor (n8914,n8911,n8912);
or (n8915,n8916,n8919);
and (n8916,n8917,n8918);
xor (n8917,n8823,n8824);
and (n8918,n279,n99);
and (n8919,n8920,n8921);
xor (n8920,n8917,n8918);
or (n8921,n8922,n8925);
and (n8922,n8923,n8924);
xor (n8923,n8828,n8829);
and (n8924,n59,n99);
and (n8925,n8926,n8927);
xor (n8926,n8923,n8924);
or (n8927,n8928,n8931);
and (n8928,n8929,n8930);
xor (n8929,n8833,n8834);
and (n8930,n53,n99);
and (n8931,n8932,n8933);
xor (n8932,n8929,n8930);
or (n8933,n8934,n8937);
and (n8934,n8935,n8936);
xor (n8935,n8839,n8840);
and (n8936,n222,n99);
and (n8937,n8938,n8939);
xor (n8938,n8935,n8936);
or (n8939,n8940,n8943);
and (n8940,n8941,n8942);
xor (n8941,n8844,n8845);
and (n8942,n215,n99);
and (n8943,n8944,n8945);
xor (n8944,n8941,n8942);
or (n8945,n8946,n8949);
and (n8946,n8947,n8948);
xor (n8947,n8850,n8851);
and (n8948,n956,n99);
and (n8949,n8950,n8951);
xor (n8950,n8947,n8948);
or (n8951,n8952,n8955);
and (n8952,n8953,n8954);
xor (n8953,n8856,n8857);
and (n8954,n1305,n99);
and (n8955,n8956,n8957);
xor (n8956,n8953,n8954);
or (n8957,n8958,n8961);
and (n8958,n8959,n8960);
xor (n8959,n8861,n8862);
and (n8960,n1131,n99);
and (n8961,n8962,n8963);
xor (n8962,n8959,n8960);
or (n8963,n8964,n8967);
and (n8964,n8965,n8966);
xor (n8965,n8866,n8867);
and (n8966,n1125,n99);
and (n8967,n8968,n8969);
xor (n8968,n8965,n8966);
or (n8969,n8970,n8973);
and (n8970,n8971,n8972);
xor (n8971,n8872,n8873);
and (n8972,n1250,n99);
and (n8973,n8974,n8975);
xor (n8974,n8971,n8972);
or (n8975,n8976,n8979);
and (n8976,n8977,n8978);
xor (n8977,n8878,n8879);
and (n8978,n1244,n99);
and (n8979,n8980,n8981);
xor (n8980,n8977,n8978);
and (n8981,n8982,n8983);
xor (n8982,n8884,n8885);
not (n8983,n3141);
and (n8984,n193,n107);
and (n8985,n8986,n8987);
xor (n8986,n8608,n8984);
or (n8987,n8988,n8991);
and (n8988,n8989,n8990);
xor (n8989,n8890,n8891);
and (n8990,n186,n107);
and (n8991,n8992,n8993);
xor (n8992,n8989,n8990);
or (n8993,n8994,n8997);
and (n8994,n8995,n8996);
xor (n8995,n8896,n8897);
and (n8996,n328,n107);
and (n8997,n8998,n8999);
xor (n8998,n8995,n8996);
or (n8999,n9000,n9003);
and (n9000,n9001,n9002);
xor (n9001,n8902,n8903);
and (n9002,n313,n107);
and (n9003,n9004,n9005);
xor (n9004,n9001,n9002);
or (n9005,n9006,n9009);
and (n9006,n9007,n9008);
xor (n9007,n8908,n8909);
and (n9008,n297,n107);
and (n9009,n9010,n9011);
xor (n9010,n9007,n9008);
or (n9011,n9012,n9015);
and (n9012,n9013,n9014);
xor (n9013,n8914,n8915);
and (n9014,n279,n107);
and (n9015,n9016,n9017);
xor (n9016,n9013,n9014);
or (n9017,n9018,n9020);
and (n9018,n9019,n1283);
xor (n9019,n8920,n8921);
and (n9020,n9021,n9022);
xor (n9021,n9019,n1283);
or (n9022,n9023,n9026);
and (n9023,n9024,n9025);
xor (n9024,n8926,n8927);
and (n9025,n53,n107);
and (n9026,n9027,n9028);
xor (n9027,n9024,n9025);
or (n9028,n9029,n9031);
and (n9029,n9030,n1963);
xor (n9030,n8932,n8933);
and (n9031,n9032,n9033);
xor (n9032,n9030,n1963);
or (n9033,n9034,n9036);
and (n9034,n9035,n1960);
xor (n9035,n8938,n8939);
and (n9036,n9037,n9038);
xor (n9037,n9035,n1960);
or (n9038,n9039,n9042);
and (n9039,n9040,n9041);
xor (n9040,n8944,n8945);
and (n9041,n956,n107);
and (n9042,n9043,n9044);
xor (n9043,n9040,n9041);
or (n9044,n9045,n9048);
and (n9045,n9046,n9047);
xor (n9046,n8950,n8951);
and (n9047,n1305,n107);
and (n9048,n9049,n9050);
xor (n9049,n9046,n9047);
or (n9050,n9051,n9054);
and (n9051,n9052,n9053);
xor (n9052,n8956,n8957);
and (n9053,n1131,n107);
and (n9054,n9055,n9056);
xor (n9055,n9052,n9053);
or (n9056,n9057,n9059);
and (n9057,n9058,n2728);
xor (n9058,n8962,n8963);
and (n9059,n9060,n9061);
xor (n9060,n9058,n2728);
or (n9061,n9062,n9065);
and (n9062,n9063,n9064);
xor (n9063,n8968,n8969);
and (n9064,n1250,n107);
and (n9065,n9066,n9067);
xor (n9066,n9063,n9064);
or (n9067,n9068,n9071);
and (n9068,n9069,n9070);
xor (n9069,n8974,n8975);
and (n9070,n1244,n107);
and (n9071,n9072,n9073);
xor (n9072,n9069,n9070);
and (n9073,n9074,n9075);
xor (n9074,n8980,n8981);
and (n9075,n1377,n107);
and (n9076,n193,n175);
and (n9077,n9078,n9079);
xor (n9078,n8606,n9076);
or (n9079,n9080,n9083);
and (n9080,n9081,n9082);
xor (n9081,n8986,n8987);
and (n9082,n186,n175);
and (n9083,n9084,n9085);
xor (n9084,n9081,n9082);
or (n9085,n9086,n9089);
and (n9086,n9087,n9088);
xor (n9087,n8992,n8993);
and (n9088,n328,n175);
and (n9089,n9090,n9091);
xor (n9090,n9087,n9088);
or (n9091,n9092,n9095);
and (n9092,n9093,n9094);
xor (n9093,n8998,n8999);
and (n9094,n313,n175);
and (n9095,n9096,n9097);
xor (n9096,n9093,n9094);
or (n9097,n9098,n9101);
and (n9098,n9099,n9100);
xor (n9099,n9004,n9005);
and (n9100,n297,n175);
and (n9101,n9102,n9103);
xor (n9102,n9099,n9100);
or (n9103,n9104,n9107);
and (n9104,n9105,n9106);
xor (n9105,n9010,n9011);
and (n9106,n279,n175);
and (n9107,n9108,n9109);
xor (n9108,n9105,n9106);
or (n9109,n9110,n9113);
and (n9110,n9111,n9112);
xor (n9111,n9016,n9017);
and (n9112,n59,n175);
and (n9113,n9114,n9115);
xor (n9114,n9111,n9112);
or (n9115,n9116,n9119);
and (n9116,n9117,n9118);
xor (n9117,n9021,n9022);
and (n9118,n53,n175);
and (n9119,n9120,n9121);
xor (n9120,n9117,n9118);
or (n9121,n9122,n9125);
and (n9122,n9123,n9124);
xor (n9123,n9027,n9028);
and (n9124,n222,n175);
and (n9125,n9126,n9127);
xor (n9126,n9123,n9124);
or (n9127,n9128,n9131);
and (n9128,n9129,n9130);
xor (n9129,n9032,n9033);
and (n9130,n215,n175);
and (n9131,n9132,n9133);
xor (n9132,n9129,n9130);
or (n9133,n9134,n9137);
and (n9134,n9135,n9136);
xor (n9135,n9037,n9038);
and (n9136,n956,n175);
and (n9137,n9138,n9139);
xor (n9138,n9135,n9136);
or (n9139,n9140,n9143);
and (n9140,n9141,n9142);
xor (n9141,n9043,n9044);
and (n9142,n1305,n175);
and (n9143,n9144,n9145);
xor (n9144,n9141,n9142);
or (n9145,n9146,n9149);
and (n9146,n9147,n9148);
xor (n9147,n9049,n9050);
and (n9148,n1131,n175);
and (n9149,n9150,n9151);
xor (n9150,n9147,n9148);
or (n9151,n9152,n9155);
and (n9152,n9153,n9154);
xor (n9153,n9055,n9056);
and (n9154,n1125,n175);
and (n9155,n9156,n9157);
xor (n9156,n9153,n9154);
or (n9157,n9158,n9161);
and (n9158,n9159,n9160);
xor (n9159,n9060,n9061);
and (n9160,n1250,n175);
and (n9161,n9162,n9163);
xor (n9162,n9159,n9160);
or (n9163,n9164,n9167);
and (n9164,n9165,n9166);
xor (n9165,n9066,n9067);
and (n9166,n1244,n175);
and (n9167,n9168,n9169);
xor (n9168,n9165,n9166);
and (n9169,n9170,n2851);
xor (n9170,n9072,n9073);
and (n9171,n193,n180);
and (n9172,n9173,n9174);
xor (n9173,n8604,n9171);
or (n9174,n9175,n9178);
and (n9175,n9176,n9177);
xor (n9176,n9078,n9079);
and (n9177,n186,n180);
and (n9178,n9179,n9180);
xor (n9179,n9176,n9177);
or (n9180,n9181,n9183);
and (n9181,n9182,n948);
xor (n9182,n9084,n9085);
and (n9183,n9184,n9185);
xor (n9184,n9182,n948);
or (n9185,n9186,n9188);
and (n9186,n9187,n4318);
xor (n9187,n9090,n9091);
and (n9188,n9189,n9190);
xor (n9189,n9187,n4318);
or (n9190,n9191,n9193);
and (n9191,n9192,n4540);
xor (n9192,n9096,n9097);
and (n9193,n9194,n9195);
xor (n9194,n9192,n4540);
or (n9195,n9196,n9199);
and (n9196,n9197,n9198);
xor (n9197,n9102,n9103);
and (n9198,n279,n180);
and (n9199,n9200,n9201);
xor (n9200,n9197,n9198);
or (n9201,n9202,n9205);
and (n9202,n9203,n9204);
xor (n9203,n9108,n9109);
and (n9204,n59,n180);
and (n9205,n9206,n9207);
xor (n9206,n9203,n9204);
or (n9207,n9208,n9211);
and (n9208,n9209,n9210);
xor (n9209,n9114,n9115);
and (n9210,n53,n180);
and (n9211,n9212,n9213);
xor (n9212,n9209,n9210);
or (n9213,n9214,n9217);
and (n9214,n9215,n9216);
xor (n9215,n9120,n9121);
and (n9216,n222,n180);
and (n9217,n9218,n9219);
xor (n9218,n9215,n9216);
or (n9219,n9220,n9222);
and (n9220,n9221,n1261);
xor (n9221,n9126,n9127);
and (n9222,n9223,n9224);
xor (n9223,n9221,n1261);
or (n9224,n9225,n9227);
and (n9225,n9226,n1915);
xor (n9226,n9132,n9133);
and (n9227,n9228,n9229);
xor (n9228,n9226,n1915);
or (n9229,n9230,n9233);
and (n9230,n9231,n9232);
xor (n9231,n9138,n9139);
and (n9232,n1305,n180);
and (n9233,n9234,n9235);
xor (n9234,n9231,n9232);
or (n9235,n9236,n9239);
and (n9236,n9237,n9238);
xor (n9237,n9144,n9145);
and (n9238,n1131,n180);
and (n9239,n9240,n9241);
xor (n9240,n9237,n9238);
or (n9241,n9242,n9244);
and (n9242,n9243,n2393);
xor (n9243,n9150,n9151);
and (n9244,n9245,n9246);
xor (n9245,n9243,n2393);
or (n9246,n9247,n9250);
and (n9247,n9248,n9249);
xor (n9248,n9156,n9157);
and (n9249,n1250,n180);
and (n9250,n9251,n9252);
xor (n9251,n9248,n9249);
or (n9252,n9253,n9256);
and (n9253,n9254,n9255);
xor (n9254,n9162,n9163);
and (n9255,n1244,n180);
and (n9256,n9257,n9258);
xor (n9257,n9254,n9255);
and (n9258,n9259,n9260);
xor (n9259,n9168,n9169);
and (n9260,n1377,n180);
and (n9261,n193,n319);
and (n9262,n9263,n9264);
xor (n9263,n8602,n9261);
or (n9264,n9265,n9268);
and (n9265,n9266,n9267);
xor (n9266,n9173,n9174);
and (n9267,n186,n319);
and (n9268,n9269,n9270);
xor (n9269,n9266,n9267);
or (n9270,n9271,n9274);
and (n9271,n9272,n9273);
xor (n9272,n9179,n9180);
and (n9273,n328,n319);
and (n9274,n9275,n9276);
xor (n9275,n9272,n9273);
or (n9276,n9277,n9280);
and (n9277,n9278,n9279);
xor (n9278,n9184,n9185);
and (n9279,n313,n319);
and (n9280,n9281,n9282);
xor (n9281,n9278,n9279);
or (n9282,n9283,n9286);
and (n9283,n9284,n9285);
xor (n9284,n9189,n9190);
and (n9285,n297,n319);
and (n9286,n9287,n9288);
xor (n9287,n9284,n9285);
or (n9288,n9289,n9292);
and (n9289,n9290,n9291);
xor (n9290,n9194,n9195);
and (n9291,n279,n319);
and (n9292,n9293,n9294);
xor (n9293,n9290,n9291);
or (n9294,n9295,n9298);
and (n9295,n9296,n9297);
xor (n9296,n9200,n9201);
and (n9297,n59,n319);
and (n9298,n9299,n9300);
xor (n9299,n9296,n9297);
or (n9300,n9301,n9304);
and (n9301,n9302,n9303);
xor (n9302,n9206,n9207);
and (n9303,n53,n319);
and (n9304,n9305,n9306);
xor (n9305,n9302,n9303);
or (n9306,n9307,n9310);
and (n9307,n9308,n9309);
xor (n9308,n9212,n9213);
and (n9309,n222,n319);
and (n9310,n9311,n9312);
xor (n9311,n9308,n9309);
or (n9312,n9313,n9316);
and (n9313,n9314,n9315);
xor (n9314,n9218,n9219);
and (n9315,n215,n319);
and (n9316,n9317,n9318);
xor (n9317,n9314,n9315);
or (n9318,n9319,n9322);
and (n9319,n9320,n9321);
xor (n9320,n9223,n9224);
and (n9321,n956,n319);
and (n9322,n9323,n9324);
xor (n9323,n9320,n9321);
or (n9324,n9325,n9328);
and (n9325,n9326,n9327);
xor (n9326,n9228,n9229);
and (n9327,n1305,n319);
and (n9328,n9329,n9330);
xor (n9329,n9326,n9327);
or (n9330,n9331,n9334);
and (n9331,n9332,n9333);
xor (n9332,n9234,n9235);
and (n9333,n1131,n319);
and (n9334,n9335,n9336);
xor (n9335,n9332,n9333);
or (n9336,n9337,n9340);
and (n9337,n9338,n9339);
xor (n9338,n9240,n9241);
and (n9339,n1125,n319);
and (n9340,n9341,n9342);
xor (n9341,n9338,n9339);
or (n9342,n9343,n9346);
and (n9343,n9344,n9345);
xor (n9344,n9245,n9246);
and (n9345,n1250,n319);
and (n9346,n9347,n9348);
xor (n9347,n9344,n9345);
or (n9348,n9349,n9352);
and (n9349,n9350,n9351);
xor (n9350,n9251,n9252);
and (n9351,n1244,n319);
and (n9352,n9353,n9354);
xor (n9353,n9350,n9351);
and (n9354,n9355,n2578);
xor (n9355,n9257,n9258);
and (n9356,n9357,n9358);
xor (n9357,n8600,n653);
or (n9358,n9359,n9362);
and (n9359,n9360,n9361);
xor (n9360,n9263,n9264);
and (n9361,n186,n291);
and (n9362,n9363,n9364);
xor (n9363,n9360,n9361);
or (n9364,n9365,n9367);
and (n9365,n9366,n329);
xor (n9366,n9269,n9270);
and (n9367,n9368,n9369);
xor (n9368,n9366,n329);
or (n9369,n9370,n9372);
and (n9370,n9371,n314);
xor (n9371,n9275,n9276);
and (n9372,n9373,n9374);
xor (n9373,n9371,n314);
or (n9374,n9375,n9377);
and (n9375,n9376,n4216);
xor (n9376,n9281,n9282);
and (n9377,n9378,n9379);
xor (n9378,n9376,n4216);
or (n9379,n9380,n9383);
and (n9380,n9381,n9382);
xor (n9381,n9287,n9288);
and (n9382,n279,n291);
and (n9383,n9384,n9385);
xor (n9384,n9381,n9382);
or (n9385,n9386,n9389);
and (n9386,n9387,n9388);
xor (n9387,n9293,n9294);
and (n9388,n59,n291);
and (n9389,n9390,n9391);
xor (n9390,n9387,n9388);
or (n9391,n9392,n9395);
and (n9392,n9393,n9394);
xor (n9393,n9299,n9300);
and (n9394,n53,n291);
and (n9395,n9396,n9397);
xor (n9396,n9393,n9394);
or (n9397,n9398,n9401);
and (n9398,n9399,n9400);
xor (n9399,n9305,n9306);
and (n9400,n222,n291);
and (n9401,n9402,n9403);
xor (n9402,n9399,n9400);
or (n9403,n9404,n9406);
and (n9404,n9405,n1770);
xor (n9405,n9311,n9312);
and (n9406,n9407,n9408);
xor (n9407,n9405,n1770);
or (n9408,n9409,n9412);
and (n9409,n9410,n9411);
xor (n9410,n9317,n9318);
and (n9411,n956,n291);
and (n9412,n9413,n9414);
xor (n9413,n9410,n9411);
or (n9414,n9415,n9417);
and (n9415,n9416,n1306);
xor (n9416,n9323,n9324);
and (n9417,n9418,n9419);
xor (n9418,n9416,n1306);
or (n9419,n9420,n9423);
and (n9420,n9421,n9422);
xor (n9421,n9329,n9330);
and (n9422,n1131,n291);
and (n9423,n9424,n9425);
xor (n9424,n9421,n9422);
or (n9425,n9426,n9429);
and (n9426,n9427,n9428);
xor (n9427,n9335,n9336);
and (n9428,n1125,n291);
and (n9429,n9430,n9431);
xor (n9430,n9427,n9428);
or (n9431,n9432,n9434);
and (n9432,n9433,n2161);
xor (n9433,n9341,n9342);
and (n9434,n9435,n9436);
xor (n9435,n9433,n2161);
or (n9436,n9437,n9439);
and (n9437,n9438,n2340);
xor (n9438,n9347,n9348);
and (n9439,n9440,n9441);
xor (n9440,n9438,n2340);
and (n9441,n9442,n9443);
xor (n9442,n9353,n9354);
and (n9443,n1377,n291);
and (n9444,n193,n286);
and (n9445,n9446,n9447);
xor (n9446,n8598,n9444);
or (n9447,n9448,n9451);
and (n9448,n9449,n9450);
xor (n9449,n9357,n9358);
and (n9450,n186,n286);
and (n9451,n9452,n9453);
xor (n9452,n9449,n9450);
or (n9453,n9454,n9457);
and (n9454,n9455,n9456);
xor (n9455,n9363,n9364);
and (n9456,n328,n286);
and (n9457,n9458,n9459);
xor (n9458,n9455,n9456);
or (n9459,n9460,n9463);
and (n9460,n9461,n9462);
xor (n9461,n9368,n9369);
and (n9462,n313,n286);
and (n9463,n9464,n9465);
xor (n9464,n9461,n9462);
or (n9465,n9466,n9469);
and (n9466,n9467,n9468);
xor (n9467,n9373,n9374);
and (n9468,n297,n286);
and (n9469,n9470,n9471);
xor (n9470,n9467,n9468);
or (n9471,n9472,n9475);
and (n9472,n9473,n9474);
xor (n9473,n9378,n9379);
and (n9474,n279,n286);
and (n9475,n9476,n9477);
xor (n9476,n9473,n9474);
or (n9477,n9478,n9481);
and (n9478,n9479,n9480);
xor (n9479,n9384,n9385);
and (n9480,n59,n286);
and (n9481,n9482,n9483);
xor (n9482,n9479,n9480);
or (n9483,n9484,n9487);
and (n9484,n9485,n9486);
xor (n9485,n9390,n9391);
and (n9486,n53,n286);
and (n9487,n9488,n9489);
xor (n9488,n9485,n9486);
or (n9489,n9490,n9493);
and (n9490,n9491,n9492);
xor (n9491,n9396,n9397);
and (n9492,n222,n286);
and (n9493,n9494,n9495);
xor (n9494,n9491,n9492);
or (n9495,n9496,n9499);
and (n9496,n9497,n9498);
xor (n9497,n9402,n9403);
and (n9498,n215,n286);
and (n9499,n9500,n9501);
xor (n9500,n9497,n9498);
or (n9501,n9502,n9505);
and (n9502,n9503,n9504);
xor (n9503,n9407,n9408);
and (n9504,n956,n286);
and (n9505,n9506,n9507);
xor (n9506,n9503,n9504);
or (n9507,n9508,n9511);
and (n9508,n9509,n9510);
xor (n9509,n9413,n9414);
and (n9510,n1305,n286);
and (n9511,n9512,n9513);
xor (n9512,n9509,n9510);
or (n9513,n9514,n9517);
and (n9514,n9515,n9516);
xor (n9515,n9418,n9419);
and (n9516,n1131,n286);
and (n9517,n9518,n9519);
xor (n9518,n9515,n9516);
or (n9519,n9520,n9523);
and (n9520,n9521,n9522);
xor (n9521,n9424,n9425);
and (n9522,n1125,n286);
and (n9523,n9524,n9525);
xor (n9524,n9521,n9522);
or (n9525,n9526,n9529);
and (n9526,n9527,n9528);
xor (n9527,n9430,n9431);
and (n9528,n1250,n286);
and (n9529,n9530,n9531);
xor (n9530,n9527,n9528);
or (n9531,n9532,n9535);
and (n9532,n9533,n9534);
xor (n9533,n9435,n9436);
and (n9534,n1244,n286);
and (n9535,n9536,n9537);
xor (n9536,n9533,n9534);
and (n9537,n9538,n1489);
xor (n9538,n9440,n9441);
and (n9539,n193,n266);
or (n9540,n9541,n9544);
and (n9541,n9542,n9543);
xor (n9542,n9446,n9447);
and (n9543,n186,n266);
and (n9544,n9545,n9546);
xor (n9545,n9542,n9543);
or (n9546,n9547,n9549);
and (n9547,n9548,n646);
xor (n9548,n9452,n9453);
and (n9549,n9550,n9551);
xor (n9550,n9548,n646);
or (n9551,n9552,n9555);
and (n9552,n9553,n9554);
xor (n9553,n9458,n9459);
and (n9554,n313,n266);
and (n9555,n9556,n9557);
xor (n9556,n9553,n9554);
or (n9557,n9558,n9560);
and (n9558,n9559,n298);
xor (n9559,n9464,n9465);
and (n9560,n9561,n9562);
xor (n9561,n9559,n298);
or (n9562,n9563,n9565);
and (n9563,n9564,n280);
xor (n9564,n9470,n9471);
and (n9565,n9566,n9567);
xor (n9566,n9564,n280);
or (n9567,n9568,n9570);
and (n9568,n9569,n982);
xor (n9569,n9476,n9477);
and (n9570,n9571,n9572);
xor (n9571,n9569,n982);
or (n9572,n9573,n9576);
and (n9573,n9574,n9575);
xor (n9574,n9482,n9483);
and (n9575,n53,n266);
and (n9576,n9577,n9578);
xor (n9577,n9574,n9575);
or (n9578,n9579,n9582);
and (n9579,n9580,n9581);
xor (n9580,n9488,n9489);
and (n9581,n222,n266);
and (n9582,n9583,n9584);
xor (n9583,n9580,n9581);
or (n9584,n9585,n9588);
and (n9585,n9586,n9587);
xor (n9586,n9494,n9495);
and (n9587,n215,n266);
and (n9588,n9589,n9590);
xor (n9589,n9586,n9587);
or (n9590,n9591,n9594);
and (n9591,n9592,n9593);
xor (n9592,n9500,n9501);
and (n9593,n956,n266);
and (n9594,n9595,n9596);
xor (n9595,n9592,n9593);
or (n9596,n9597,n9600);
and (n9597,n9598,n9599);
xor (n9598,n9506,n9507);
and (n9599,n1305,n266);
and (n9600,n9601,n9602);
xor (n9601,n9598,n9599);
or (n9602,n9603,n9606);
and (n9603,n9604,n9605);
xor (n9604,n9512,n9513);
and (n9605,n1131,n266);
and (n9606,n9607,n9608);
xor (n9607,n9604,n9605);
or (n9608,n9609,n9611);
and (n9609,n9610,n1126);
xor (n9610,n9518,n9519);
and (n9611,n9612,n9613);
xor (n9612,n9610,n1126);
or (n9613,n9614,n9616);
and (n9614,n9615,n2044);
xor (n9615,n9524,n9525);
and (n9616,n9617,n9618);
xor (n9617,n9615,n2044);
or (n9618,n9619,n9622);
and (n9619,n9620,n9621);
xor (n9620,n9530,n9531);
and (n9621,n1244,n266);
and (n9622,n9623,n9624);
xor (n9623,n9620,n9621);
and (n9624,n9625,n9626);
xor (n9625,n9536,n9537);
and (n9626,n1377,n266);
and (n9627,n186,n259);
or (n9628,n9629,n9632);
and (n9629,n9630,n9631);
xor (n9630,n9545,n9546);
and (n9631,n328,n259);
and (n9632,n9633,n9634);
xor (n9633,n9630,n9631);
or (n9634,n9635,n9638);
and (n9635,n9636,n9637);
xor (n9636,n9550,n9551);
and (n9637,n313,n259);
and (n9638,n9639,n9640);
xor (n9639,n9636,n9637);
or (n9640,n9641,n9644);
and (n9641,n9642,n9643);
xor (n9642,n9556,n9557);
and (n9643,n297,n259);
and (n9644,n9645,n9646);
xor (n9645,n9642,n9643);
or (n9646,n9647,n9650);
and (n9647,n9648,n9649);
xor (n9648,n9561,n9562);
and (n9649,n279,n259);
and (n9650,n9651,n9652);
xor (n9651,n9648,n9649);
or (n9652,n9653,n9656);
and (n9653,n9654,n9655);
xor (n9654,n9566,n9567);
and (n9655,n59,n259);
and (n9656,n9657,n9658);
xor (n9657,n9654,n9655);
or (n9658,n9659,n9662);
and (n9659,n9660,n9661);
xor (n9660,n9571,n9572);
and (n9661,n53,n259);
and (n9662,n9663,n9664);
xor (n9663,n9660,n9661);
or (n9664,n9665,n9668);
and (n9665,n9666,n9667);
xor (n9666,n9577,n9578);
and (n9667,n222,n259);
and (n9668,n9669,n9670);
xor (n9669,n9666,n9667);
or (n9670,n9671,n9674);
and (n9671,n9672,n9673);
xor (n9672,n9583,n9584);
and (n9673,n215,n259);
and (n9674,n9675,n9676);
xor (n9675,n9672,n9673);
or (n9676,n9677,n9680);
and (n9677,n9678,n9679);
xor (n9678,n9589,n9590);
and (n9679,n956,n259);
and (n9680,n9681,n9682);
xor (n9681,n9678,n9679);
or (n9682,n9683,n9686);
and (n9683,n9684,n9685);
xor (n9684,n9595,n9596);
and (n9685,n1305,n259);
and (n9686,n9687,n9688);
xor (n9687,n9684,n9685);
or (n9688,n9689,n9692);
and (n9689,n9690,n9691);
xor (n9690,n9601,n9602);
and (n9691,n1131,n259);
and (n9692,n9693,n9694);
xor (n9693,n9690,n9691);
or (n9694,n9695,n9698);
and (n9695,n9696,n9697);
xor (n9696,n9607,n9608);
and (n9697,n1125,n259);
and (n9698,n9699,n9700);
xor (n9699,n9696,n9697);
or (n9700,n9701,n9704);
and (n9701,n9702,n9703);
xor (n9702,n9612,n9613);
and (n9703,n1250,n259);
and (n9704,n9705,n9706);
xor (n9705,n9702,n9703);
or (n9706,n9707,n9710);
and (n9707,n9708,n9709);
xor (n9708,n9617,n9618);
and (n9709,n1244,n259);
and (n9710,n9711,n9712);
xor (n9711,n9708,n9709);
and (n9712,n9713,n1555);
xor (n9713,n9623,n9624);
and (n9714,n328,n48);
or (n9715,n9716,n9719);
and (n9716,n9717,n9718);
xor (n9717,n9633,n9634);
and (n9718,n313,n48);
and (n9719,n9720,n9721);
xor (n9720,n9717,n9718);
or (n9721,n9722,n9725);
and (n9722,n9723,n9724);
xor (n9723,n9639,n9640);
and (n9724,n297,n48);
and (n9725,n9726,n9727);
xor (n9726,n9723,n9724);
or (n9727,n9728,n9730);
and (n9728,n9729,n598);
xor (n9729,n9645,n9646);
and (n9730,n9731,n9732);
xor (n9731,n9729,n598);
or (n9732,n9733,n9735);
and (n9733,n9734,n271);
xor (n9734,n9651,n9652);
and (n9735,n9736,n9737);
xor (n9736,n9734,n271);
or (n9737,n9738,n9740);
and (n9738,n9739,n254);
xor (n9739,n9657,n9658);
and (n9740,n9741,n9742);
xor (n9741,n9739,n254);
or (n9742,n9743,n9745);
and (n9743,n9744,n975);
xor (n9744,n9663,n9664);
and (n9745,n9746,n9747);
xor (n9746,n9744,n975);
or (n9747,n9748,n9751);
and (n9748,n9749,n9750);
xor (n9749,n9669,n9670);
and (n9750,n215,n48);
and (n9751,n9752,n9753);
xor (n9752,n9749,n9750);
or (n9753,n9754,n9757);
and (n9754,n9755,n9756);
xor (n9755,n9675,n9676);
and (n9756,n956,n48);
and (n9757,n9758,n9759);
xor (n9758,n9755,n9756);
or (n9759,n9760,n9763);
and (n9760,n9761,n9762);
xor (n9761,n9681,n9682);
and (n9762,n1305,n48);
and (n9763,n9764,n9765);
xor (n9764,n9761,n9762);
or (n9765,n9766,n9769);
and (n9766,n9767,n9768);
xor (n9767,n9687,n9688);
and (n9768,n1131,n48);
and (n9769,n9770,n9771);
xor (n9770,n9767,n9768);
or (n9771,n9772,n9775);
and (n9772,n9773,n9774);
xor (n9773,n9693,n9694);
and (n9774,n1125,n48);
and (n9775,n9776,n9777);
xor (n9776,n9773,n9774);
or (n9777,n9778,n9781);
and (n9778,n9779,n9780);
xor (n9779,n9699,n9700);
and (n9780,n1250,n48);
and (n9781,n9782,n9783);
xor (n9782,n9779,n9780);
or (n9783,n9784,n9787);
and (n9784,n9785,n9786);
xor (n9785,n9705,n9706);
and (n9786,n1244,n48);
and (n9787,n9788,n9789);
xor (n9788,n9785,n9786);
and (n9789,n9790,n9791);
xor (n9790,n9711,n9712);
and (n9791,n1377,n48);
and (n9792,n313,n43);
or (n9793,n9794,n9797);
and (n9794,n9795,n9796);
xor (n9795,n9720,n9721);
and (n9796,n297,n43);
and (n9797,n9798,n9799);
xor (n9798,n9795,n9796);
or (n9799,n9800,n9803);
and (n9800,n9801,n9802);
xor (n9801,n9726,n9727);
and (n9802,n279,n43);
and (n9803,n9804,n9805);
xor (n9804,n9801,n9802);
or (n9805,n9806,n9809);
and (n9806,n9807,n9808);
xor (n9807,n9731,n9732);
and (n9808,n59,n43);
and (n9809,n9810,n9811);
xor (n9810,n9807,n9808);
or (n9811,n9812,n9815);
and (n9812,n9813,n9814);
xor (n9813,n9736,n9737);
and (n9814,n53,n43);
and (n9815,n9816,n9817);
xor (n9816,n9813,n9814);
or (n9817,n9818,n9821);
and (n9818,n9819,n9820);
xor (n9819,n9741,n9742);
and (n9820,n222,n43);
and (n9821,n9822,n9823);
xor (n9822,n9819,n9820);
or (n9823,n9824,n9827);
and (n9824,n9825,n9826);
xor (n9825,n9746,n9747);
and (n9826,n215,n43);
and (n9827,n9828,n9829);
xor (n9828,n9825,n9826);
or (n9829,n9830,n9833);
and (n9830,n9831,n9832);
xor (n9831,n9752,n9753);
and (n9832,n956,n43);
and (n9833,n9834,n9835);
xor (n9834,n9831,n9832);
or (n9835,n9836,n9839);
and (n9836,n9837,n9838);
xor (n9837,n9758,n9759);
and (n9838,n1305,n43);
and (n9839,n9840,n9841);
xor (n9840,n9837,n9838);
or (n9841,n9842,n9845);
and (n9842,n9843,n9844);
xor (n9843,n9764,n9765);
and (n9844,n1131,n43);
and (n9845,n9846,n9847);
xor (n9846,n9843,n9844);
or (n9847,n9848,n9851);
and (n9848,n9849,n9850);
xor (n9849,n9770,n9771);
and (n9850,n1125,n43);
and (n9851,n9852,n9853);
xor (n9852,n9849,n9850);
or (n9853,n9854,n9857);
and (n9854,n9855,n9856);
xor (n9855,n9776,n9777);
and (n9856,n1250,n43);
and (n9857,n9858,n9859);
xor (n9858,n9855,n9856);
or (n9859,n9860,n9863);
and (n9860,n9861,n9862);
xor (n9861,n9782,n9783);
and (n9862,n1244,n43);
and (n9863,n9864,n9865);
xor (n9864,n9861,n9862);
and (n9865,n9866,n1872);
xor (n9866,n9788,n9789);
and (n9867,n297,n42);
or (n9868,n9869,n9872);
and (n9869,n9870,n9871);
xor (n9870,n9798,n9799);
and (n9871,n279,n42);
and (n9872,n9873,n9874);
xor (n9873,n9870,n9871);
or (n9874,n9875,n9878);
and (n9875,n9876,n9877);
xor (n9876,n9804,n9805);
and (n9877,n59,n42);
and (n9878,n9879,n9880);
xor (n9879,n9876,n9877);
or (n9880,n9881,n9884);
and (n9881,n9882,n9883);
xor (n9882,n9810,n9811);
and (n9883,n53,n42);
and (n9884,n9885,n9886);
xor (n9885,n9882,n9883);
or (n9886,n9887,n9890);
and (n9887,n9888,n9889);
xor (n9888,n9816,n9817);
and (n9889,n222,n42);
and (n9890,n9891,n9892);
xor (n9891,n9888,n9889);
or (n9892,n9893,n9896);
and (n9893,n9894,n9895);
xor (n9894,n9822,n9823);
and (n9895,n215,n42);
and (n9896,n9897,n9898);
xor (n9897,n9894,n9895);
or (n9898,n9899,n9901);
and (n9899,n9900,n957);
xor (n9900,n9828,n9829);
and (n9901,n9902,n9903);
xor (n9902,n9900,n957);
or (n9903,n9904,n9906);
and (n9904,n9905,n4588);
xor (n9905,n9834,n9835);
and (n9906,n9907,n9908);
xor (n9907,n9905,n4588);
or (n9908,n9909,n9911);
and (n9909,n9910,n4362);
xor (n9910,n9840,n9841);
and (n9911,n9912,n9913);
xor (n9912,n9910,n4362);
or (n9913,n9914,n9917);
and (n9914,n9915,n9916);
xor (n9915,n9846,n9847);
and (n9916,n1125,n42);
and (n9917,n9918,n9919);
xor (n9918,n9915,n9916);
or (n9919,n9920,n9923);
and (n9920,n9921,n9922);
xor (n9921,n9852,n9853);
and (n9922,n1250,n42);
and (n9923,n9924,n9925);
xor (n9924,n9921,n9922);
or (n9925,n9926,n9929);
and (n9926,n9927,n9928);
xor (n9927,n9858,n9859);
and (n9928,n1244,n42);
and (n9929,n9930,n9931);
xor (n9930,n9927,n9928);
and (n9931,n9932,n1701);
xor (n9932,n9864,n9865);
or (n9933,n9934,n9936);
and (n9934,n9935,n9877);
xor (n9935,n9873,n9874);
and (n9936,n9937,n9938);
xor (n9937,n9935,n9877);
or (n9938,n9939,n9941);
and (n9939,n9940,n9883);
xor (n9940,n9879,n9880);
and (n9941,n9942,n9943);
xor (n9942,n9940,n9883);
or (n9943,n9944,n9946);
and (n9944,n9945,n9889);
xor (n9945,n9885,n9886);
and (n9946,n9947,n9948);
xor (n9947,n9945,n9889);
or (n9948,n9949,n9951);
and (n9949,n9950,n9895);
xor (n9950,n9891,n9892);
and (n9951,n9952,n9953);
xor (n9952,n9950,n9895);
or (n9953,n9954,n9956);
and (n9954,n9955,n957);
xor (n9955,n9897,n9898);
and (n9956,n9957,n9958);
xor (n9957,n9955,n957);
or (n9958,n9959,n9961);
and (n9959,n9960,n4588);
xor (n9960,n9902,n9903);
and (n9961,n9962,n9963);
xor (n9962,n9960,n4588);
or (n9963,n9964,n9966);
and (n9964,n9965,n4362);
xor (n9965,n9907,n9908);
and (n9966,n9967,n9968);
xor (n9967,n9965,n4362);
or (n9968,n9969,n9971);
and (n9969,n9970,n9916);
xor (n9970,n9912,n9913);
and (n9971,n9972,n9973);
xor (n9972,n9970,n9916);
or (n9973,n9974,n9976);
and (n9974,n9975,n9922);
xor (n9975,n9918,n9919);
and (n9976,n9977,n9978);
xor (n9977,n9975,n9922);
or (n9978,n9979,n9981);
and (n9979,n9980,n9928);
xor (n9980,n9924,n9925);
and (n9981,n9982,n9983);
xor (n9982,n9980,n9928);
and (n9983,n9984,n1701);
xor (n9984,n9930,n9931);
or (n9985,n9986,n9988);
and (n9986,n9987,n9883);
xor (n9987,n9937,n9938);
and (n9988,n9989,n9990);
xor (n9989,n9987,n9883);
or (n9990,n9991,n9993);
and (n9991,n9992,n9889);
xor (n9992,n9942,n9943);
and (n9993,n9994,n9995);
xor (n9994,n9992,n9889);
or (n9995,n9996,n9998);
and (n9996,n9997,n9895);
xor (n9997,n9947,n9948);
and (n9998,n9999,n10000);
xor (n9999,n9997,n9895);
or (n10000,n10001,n10003);
and (n10001,n10002,n957);
xor (n10002,n9952,n9953);
and (n10003,n10004,n10005);
xor (n10004,n10002,n957);
or (n10005,n10006,n10008);
and (n10006,n10007,n4588);
xor (n10007,n9957,n9958);
and (n10008,n10009,n10010);
xor (n10009,n10007,n4588);
or (n10010,n10011,n10013);
and (n10011,n10012,n4362);
xor (n10012,n9962,n9963);
and (n10013,n10014,n10015);
xor (n10014,n10012,n4362);
or (n10015,n10016,n10018);
and (n10016,n10017,n9916);
xor (n10017,n9967,n9968);
and (n10018,n10019,n10020);
xor (n10019,n10017,n9916);
or (n10020,n10021,n10023);
and (n10021,n10022,n9922);
xor (n10022,n9972,n9973);
and (n10023,n10024,n10025);
xor (n10024,n10022,n9922);
or (n10025,n10026,n10028);
and (n10026,n10027,n9928);
xor (n10027,n9977,n9978);
and (n10028,n10029,n10030);
xor (n10029,n10027,n9928);
and (n10030,n10031,n1701);
xor (n10031,n9982,n9983);
or (n10032,n10033,n10035);
and (n10033,n10034,n9889);
xor (n10034,n9989,n9990);
and (n10035,n10036,n10037);
xor (n10036,n10034,n9889);
or (n10037,n10038,n10040);
and (n10038,n10039,n9895);
xor (n10039,n9994,n9995);
and (n10040,n10041,n10042);
xor (n10041,n10039,n9895);
or (n10042,n10043,n10045);
and (n10043,n10044,n957);
xor (n10044,n9999,n10000);
and (n10045,n10046,n10047);
xor (n10046,n10044,n957);
or (n10047,n10048,n10050);
and (n10048,n10049,n4588);
xor (n10049,n10004,n10005);
and (n10050,n10051,n10052);
xor (n10051,n10049,n4588);
or (n10052,n10053,n10055);
and (n10053,n10054,n4362);
xor (n10054,n10009,n10010);
and (n10055,n10056,n10057);
xor (n10056,n10054,n4362);
or (n10057,n10058,n10060);
and (n10058,n10059,n9916);
xor (n10059,n10014,n10015);
and (n10060,n10061,n10062);
xor (n10061,n10059,n9916);
or (n10062,n10063,n10065);
and (n10063,n10064,n9922);
xor (n10064,n10019,n10020);
and (n10065,n10066,n10067);
xor (n10066,n10064,n9922);
or (n10067,n10068,n10070);
and (n10068,n10069,n9928);
xor (n10069,n10024,n10025);
and (n10070,n10071,n10072);
xor (n10071,n10069,n9928);
and (n10072,n10073,n1701);
xor (n10073,n10029,n10030);
or (n10074,n10075,n10077);
and (n10075,n10076,n9895);
xor (n10076,n10036,n10037);
and (n10077,n10078,n10079);
xor (n10078,n10076,n9895);
or (n10079,n10080,n10082);
and (n10080,n10081,n957);
xor (n10081,n10041,n10042);
and (n10082,n10083,n10084);
xor (n10083,n10081,n957);
or (n10084,n10085,n10087);
and (n10085,n10086,n4588);
xor (n10086,n10046,n10047);
and (n10087,n10088,n10089);
xor (n10088,n10086,n4588);
or (n10089,n10090,n10092);
and (n10090,n10091,n4362);
xor (n10091,n10051,n10052);
and (n10092,n10093,n10094);
xor (n10093,n10091,n4362);
or (n10094,n10095,n10097);
and (n10095,n10096,n9916);
xor (n10096,n10056,n10057);
and (n10097,n10098,n10099);
xor (n10098,n10096,n9916);
or (n10099,n10100,n10102);
and (n10100,n10101,n9922);
xor (n10101,n10061,n10062);
and (n10102,n10103,n10104);
xor (n10103,n10101,n9922);
or (n10104,n10105,n10107);
and (n10105,n10106,n9928);
xor (n10106,n10066,n10067);
and (n10107,n10108,n10109);
xor (n10108,n10106,n9928);
and (n10109,n10110,n1701);
xor (n10110,n10071,n10072);
or (n10111,n10112,n10114);
and (n10112,n10113,n957);
xor (n10113,n10078,n10079);
and (n10114,n10115,n10116);
xor (n10115,n10113,n957);
or (n10116,n10117,n10119);
and (n10117,n10118,n4588);
xor (n10118,n10083,n10084);
and (n10119,n10120,n10121);
xor (n10120,n10118,n4588);
or (n10121,n10122,n10124);
and (n10122,n10123,n4362);
xor (n10123,n10088,n10089);
and (n10124,n10125,n10126);
xor (n10125,n10123,n4362);
or (n10126,n10127,n10129);
and (n10127,n10128,n9916);
xor (n10128,n10093,n10094);
and (n10129,n10130,n10131);
xor (n10130,n10128,n9916);
or (n10131,n10132,n10134);
and (n10132,n10133,n9922);
xor (n10133,n10098,n10099);
and (n10134,n10135,n10136);
xor (n10135,n10133,n9922);
or (n10136,n10137,n10139);
and (n10137,n10138,n9928);
xor (n10138,n10103,n10104);
and (n10139,n10140,n10141);
xor (n10140,n10138,n9928);
and (n10141,n10142,n1701);
xor (n10142,n10108,n10109);
or (n10143,n10144,n10146);
and (n10144,n10145,n4588);
xor (n10145,n10115,n10116);
and (n10146,n10147,n10148);
xor (n10147,n10145,n4588);
or (n10148,n10149,n10151);
and (n10149,n10150,n4362);
xor (n10150,n10120,n10121);
and (n10151,n10152,n10153);
xor (n10152,n10150,n4362);
or (n10153,n10154,n10156);
and (n10154,n10155,n9916);
xor (n10155,n10125,n10126);
and (n10156,n10157,n10158);
xor (n10157,n10155,n9916);
or (n10158,n10159,n10161);
and (n10159,n10160,n9922);
xor (n10160,n10130,n10131);
and (n10161,n10162,n10163);
xor (n10162,n10160,n9922);
or (n10163,n10164,n10166);
and (n10164,n10165,n9928);
xor (n10165,n10135,n10136);
and (n10166,n10167,n10168);
xor (n10167,n10165,n9928);
and (n10168,n10169,n1701);
xor (n10169,n10140,n10141);
or (n10170,n10171,n10173);
and (n10171,n10172,n4362);
xor (n10172,n10147,n10148);
and (n10173,n10174,n10175);
xor (n10174,n10172,n4362);
or (n10175,n10176,n10178);
and (n10176,n10177,n9916);
xor (n10177,n10152,n10153);
and (n10178,n10179,n10180);
xor (n10179,n10177,n9916);
or (n10180,n10181,n10183);
and (n10181,n10182,n9922);
xor (n10182,n10157,n10158);
and (n10183,n10184,n10185);
xor (n10184,n10182,n9922);
or (n10185,n10186,n10188);
and (n10186,n10187,n9928);
xor (n10187,n10162,n10163);
and (n10188,n10189,n10190);
xor (n10189,n10187,n9928);
and (n10190,n10191,n1701);
xor (n10191,n10167,n10168);
or (n10192,n10193,n10195);
and (n10193,n10194,n9916);
xor (n10194,n10174,n10175);
and (n10195,n10196,n10197);
xor (n10196,n10194,n9916);
or (n10197,n10198,n10200);
and (n10198,n10199,n9922);
xor (n10199,n10179,n10180);
and (n10200,n10201,n10202);
xor (n10201,n10199,n9922);
or (n10202,n10203,n10205);
and (n10203,n10204,n9928);
xor (n10204,n10184,n10185);
and (n10205,n10206,n10207);
xor (n10206,n10204,n9928);
and (n10207,n10208,n1701);
xor (n10208,n10189,n10190);
or (n10209,n10210,n10212);
and (n10210,n10211,n9922);
xor (n10211,n10196,n10197);
and (n10212,n10213,n10214);
xor (n10213,n10211,n9922);
or (n10214,n10215,n10217);
and (n10215,n10216,n9928);
xor (n10216,n10201,n10202);
and (n10217,n10218,n10219);
xor (n10218,n10216,n9928);
and (n10219,n10220,n1701);
xor (n10220,n10206,n10207);
or (n10221,n10222,n10224);
and (n10222,n10223,n9928);
xor (n10223,n10213,n10214);
and (n10224,n10225,n10226);
xor (n10225,n10223,n9928);
and (n10226,n10227,n1701);
xor (n10227,n10218,n10219);
and (n10228,n10229,n1701);
xor (n10229,n10225,n10226);
or (n10230,n10231,n10235,n10414);
and (n10231,n10232,n10234);
xor (n10232,n10233,n8412);
xor (n10233,n8409,n8410);
xor (n10234,n10229,n1701);
and (n10235,n10234,n10236);
or (n10236,n10237,n10241,n10413);
and (n10237,n10238,n10240);
xor (n10238,n10239,n8417);
xor (n10239,n8414,n8415);
xor (n10240,n10227,n1701);
and (n10241,n10240,n10242);
or (n10242,n10243,n10247,n10412);
and (n10243,n10244,n10246);
xor (n10244,n10245,n8422);
xor (n10245,n8419,n8420);
xor (n10246,n10220,n1701);
and (n10247,n10246,n10248);
or (n10248,n10249,n10253,n10411);
and (n10249,n10250,n10252);
xor (n10250,n10251,n8427);
xor (n10251,n8424,n8425);
xor (n10252,n10208,n1701);
and (n10253,n10252,n10254);
or (n10254,n10255,n10259,n10410);
and (n10255,n10256,n10258);
xor (n10256,n10257,n8432);
xor (n10257,n8429,n8430);
xor (n10258,n10191,n1701);
and (n10259,n10258,n10260);
or (n10260,n10261,n10265,n10409);
and (n10261,n10262,n10264);
xor (n10262,n10263,n8437);
xor (n10263,n8434,n8435);
xor (n10264,n10169,n1701);
and (n10265,n10264,n10266);
or (n10266,n10267,n10271,n10408);
and (n10267,n10268,n10270);
xor (n10268,n10269,n8442);
xor (n10269,n8439,n8440);
xor (n10270,n10142,n1701);
and (n10271,n10270,n10272);
or (n10272,n10273,n10277,n10407);
and (n10273,n10274,n10276);
xor (n10274,n10275,n8447);
xor (n10275,n8444,n8445);
xor (n10276,n10110,n1701);
and (n10277,n10276,n10278);
or (n10278,n10279,n10283,n10406);
and (n10279,n10280,n10282);
xor (n10280,n10281,n8452);
xor (n10281,n8449,n8450);
xor (n10282,n10073,n1701);
and (n10283,n10282,n10284);
or (n10284,n10285,n10289,n10405);
and (n10285,n10286,n10288);
xor (n10286,n10287,n8457);
xor (n10287,n8454,n8455);
xor (n10288,n10031,n1701);
and (n10289,n10288,n10290);
or (n10290,n10291,n10295,n10404);
and (n10291,n10292,n10294);
xor (n10292,n10293,n8462);
xor (n10293,n8459,n8460);
xor (n10294,n9984,n1701);
and (n10295,n10294,n10296);
or (n10296,n10297,n10301,n10403);
and (n10297,n10298,n10300);
xor (n10298,n10299,n8467);
xor (n10299,n8464,n8465);
xor (n10300,n9932,n1701);
and (n10301,n10300,n10302);
or (n10302,n10303,n10307,n10402);
and (n10303,n10304,n10306);
xor (n10304,n10305,n8472);
xor (n10305,n8469,n8470);
xor (n10306,n9866,n1872);
and (n10307,n10306,n10308);
or (n10308,n10309,n10313,n10401);
and (n10309,n10310,n10312);
xor (n10310,n10311,n8477);
xor (n10311,n8474,n8475);
xor (n10312,n9790,n9791);
and (n10313,n10312,n10314);
or (n10314,n10315,n10319,n10400);
and (n10315,n10316,n10318);
xor (n10316,n10317,n8482);
xor (n10317,n8479,n8480);
xor (n10318,n9713,n1555);
and (n10319,n10318,n10320);
or (n10320,n10321,n10325,n10399);
and (n10321,n10322,n10324);
xor (n10322,n10323,n8487);
xor (n10323,n8484,n8485);
xor (n10324,n9625,n9626);
and (n10325,n10324,n10326);
or (n10326,n10327,n10331,n10398);
and (n10327,n10328,n10330);
xor (n10328,n10329,n8492);
xor (n10329,n8489,n8490);
xor (n10330,n9538,n1489);
and (n10331,n10330,n10332);
or (n10332,n10333,n10337,n10397);
and (n10333,n10334,n10336);
xor (n10334,n10335,n8497);
xor (n10335,n8494,n8495);
xor (n10336,n9442,n9443);
and (n10337,n10336,n10338);
or (n10338,n10339,n10343,n10396);
and (n10339,n10340,n10342);
xor (n10340,n10341,n8502);
xor (n10341,n8499,n8500);
xor (n10342,n9355,n2578);
and (n10343,n10342,n10344);
or (n10344,n10345,n10349,n10395);
and (n10345,n10346,n10348);
xor (n10346,n10347,n8507);
xor (n10347,n8504,n8505);
xor (n10348,n9259,n9260);
and (n10349,n10348,n10350);
or (n10350,n10351,n10355,n10394);
and (n10351,n10352,n10354);
xor (n10352,n10353,n8512);
xor (n10353,n8509,n8510);
xor (n10354,n9170,n2851);
and (n10355,n10354,n10356);
or (n10356,n10357,n10361,n10393);
and (n10357,n10358,n10360);
xor (n10358,n10359,n8517);
xor (n10359,n8514,n8515);
xor (n10360,n9074,n9075);
and (n10361,n10360,n10362);
or (n10362,n10363,n10367,n10392);
and (n10363,n10364,n10366);
xor (n10364,n10365,n8522);
xor (n10365,n8519,n8520);
xor (n10366,n8982,n8983);
and (n10367,n10366,n10368);
or (n10368,n10369,n10373,n10391);
and (n10369,n10370,n10372);
xor (n10370,n10371,n8527);
xor (n10371,n8524,n8525);
xor (n10372,n8886,n8887);
and (n10373,n10372,n10374);
or (n10374,n10375,n10379,n10390);
and (n10375,n10376,n10378);
xor (n10376,n10377,n8532);
xor (n10377,n8529,n8530);
xor (n10378,n8796,n8797);
and (n10379,n10378,n10380);
or (n10380,n10381,n10385,n10389);
and (n10381,n10382,n10384);
xor (n10382,n10383,n3562);
xor (n10383,n8534,n8535);
xor (n10384,n8700,n8701);
and (n10385,n10384,n10386);
and (n10386,n10387,n10388);
xor (n10387,n3516,n3518);
not (n10388,n3514);
and (n10389,n10382,n10386);
and (n10390,n10376,n10380);
and (n10391,n10370,n10374);
and (n10392,n10364,n10368);
and (n10393,n10358,n10362);
and (n10394,n10352,n10356);
and (n10395,n10346,n10350);
and (n10396,n10340,n10344);
and (n10397,n10334,n10338);
and (n10398,n10328,n10332);
and (n10399,n10322,n10326);
and (n10400,n10316,n10320);
and (n10401,n10310,n10314);
and (n10402,n10304,n10308);
and (n10403,n10298,n10302);
and (n10404,n10292,n10296);
and (n10405,n10286,n10290);
and (n10406,n10280,n10284);
and (n10407,n10274,n10278);
and (n10408,n10268,n10272);
and (n10409,n10262,n10266);
and (n10410,n10256,n10260);
and (n10411,n10250,n10254);
and (n10412,n10244,n10248);
and (n10413,n10238,n10242);
and (n10414,n10232,n10236);
not (n10415,n5181);
endmodule
