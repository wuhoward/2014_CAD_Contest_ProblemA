module top (out,n18,n20,n26,n28,n38,n46,n47,n53,n54
        ,n62,n74,n79,n83,n89,n98,n99,n101,n106,n107
        ,n111,n118,n126,n132,n141,n152,n158,n167,n175,n177
        ,n182,n188,n202,n213,n220);
output out;
input n18;
input n20;
input n26;
input n28;
input n38;
input n46;
input n47;
input n53;
input n54;
input n62;
input n74;
input n79;
input n83;
input n89;
input n98;
input n99;
input n101;
input n106;
input n107;
input n111;
input n118;
input n126;
input n132;
input n141;
input n152;
input n158;
input n167;
input n175;
input n177;
input n182;
input n188;
input n202;
input n213;
input n220;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n19;
wire n21;
wire n22;
wire n23;
wire n24;
wire n25;
wire n27;
wire n29;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n75;
wire n76;
wire n77;
wire n78;
wire n80;
wire n81;
wire n82;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n100;
wire n102;
wire n103;
wire n104;
wire n105;
wire n108;
wire n109;
wire n110;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n176;
wire n178;
wire n179;
wire n180;
wire n181;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
xor (out,n0,n1006);
nand (n0,n1,n1005);
or (n1,n2,n494);
not (n2,n3);
nand (n3,n4,n493);
not (n4,n5);
nor (n5,n6,n434);
xor (n6,n7,n364);
xor (n7,n8,n222);
xor (n8,n9,n144);
xor (n9,n10,n92);
xor (n10,n11,n68);
xor (n11,n12,n40);
nand (n12,n13,n34);
or (n13,n14,n22);
not (n14,n15);
nor (n15,n16,n21);
and (n16,n17,n19);
not (n17,n18);
not (n19,n20);
and (n21,n18,n20);
not (n22,n23);
nor (n23,n24,n30);
nand (n24,n25,n29);
or (n25,n26,n27);
not (n27,n28);
nand (n29,n26,n27);
nor (n30,n31,n33);
and (n31,n32,n20);
not (n32,n26);
and (n33,n26,n19);
nand (n34,n24,n35);
nand (n35,n36,n39);
or (n36,n37,n20);
not (n37,n38);
or (n39,n19,n38);
nand (n40,n41,n57);
or (n41,n42,n49);
not (n42,n43);
nand (n43,n44,n48);
or (n44,n45,n47);
not (n45,n46);
nand (n48,n47,n45);
not (n49,n50);
nand (n50,n51,n55);
or (n51,n52,n54);
not (n52,n53);
or (n55,n56,n53);
not (n56,n54);
nand (n57,n58,n64);
not (n58,n59);
nor (n59,n60,n63);
and (n60,n54,n61);
not (n61,n62);
and (n63,n56,n62);
and (n64,n42,n65);
nand (n65,n66,n67);
nand (n66,n54,n45);
nand (n67,n46,n56);
nand (n68,n69,n86);
or (n69,n70,n81);
nand (n70,n71,n76);
nor (n71,n72,n75);
and (n72,n73,n54);
not (n73,n74);
and (n75,n74,n56);
nor (n76,n77,n80);
and (n77,n73,n78);
not (n78,n79);
and (n80,n74,n79);
nor (n81,n82,n84);
and (n82,n83,n78);
and (n84,n79,n85);
not (n85,n83);
or (n86,n87,n71);
nor (n87,n88,n90);
and (n88,n89,n78);
and (n90,n79,n91);
not (n91,n89);
xor (n92,n93,n120);
xor (n93,n94,n102);
and (n94,n95,n101);
nand (n95,n96,n100);
or (n96,n97,n99);
not (n97,n98);
nand (n100,n99,n97);
nand (n102,n103,n114);
or (n103,n104,n108);
nand (n104,n105,n107);
not (n105,n106);
nor (n108,n109,n112);
and (n109,n110,n111);
not (n110,n107);
and (n112,n107,n113);
not (n113,n111);
nand (n114,n115,n106);
nor (n115,n116,n119);
and (n116,n117,n110);
not (n117,n118);
and (n119,n118,n107);
nand (n120,n121,n134);
or (n121,n122,n128);
not (n122,n123);
nor (n123,n124,n127);
and (n124,n125,n27);
not (n125,n126);
and (n127,n126,n28);
not (n128,n129);
nand (n129,n130,n133);
or (n130,n131,n107);
not (n131,n132);
nand (n133,n107,n131);
or (n134,n135,n139);
nand (n135,n128,n136);
nand (n136,n137,n138);
or (n137,n131,n28);
nand (n138,n131,n28);
nor (n139,n140,n142);
and (n140,n27,n141);
and (n142,n28,n143);
not (n143,n141);
xor (n144,n145,n196);
xor (n145,n146,n169);
nand (n146,n147,n163);
or (n147,n148,n154);
not (n148,n149);
nor (n149,n150,n153);
and (n150,n151,n97);
not (n151,n152);
and (n153,n152,n98);
nand (n154,n155,n160);
not (n155,n156);
nand (n156,n157,n159);
or (n157,n78,n158);
nand (n159,n158,n78);
nand (n160,n161,n162);
or (n161,n158,n97);
nand (n162,n97,n158);
nand (n163,n156,n164);
nor (n164,n165,n168);
and (n165,n166,n97);
not (n166,n167);
and (n168,n167,n98);
nand (n169,n170,n184);
or (n170,n171,n179);
not (n171,n172);
nor (n172,n173,n178);
and (n173,n174,n176);
not (n174,n175);
not (n176,n177);
and (n178,n175,n177);
not (n179,n180);
nand (n180,n181,n183);
or (n181,n19,n182);
nand (n183,n182,n19);
nand (n184,n185,n191);
not (n185,n186);
nor (n186,n187,n189);
and (n187,n176,n188);
and (n189,n177,n190);
not (n190,n188);
not (n191,n192);
nand (n192,n193,n179);
nand (n193,n194,n195);
or (n194,n182,n176);
nand (n195,n176,n182);
nand (n196,n197,n215);
or (n197,n198,n209);
not (n198,n199);
nor (n199,n200,n204);
nand (n200,n201,n203);
or (n201,n176,n202);
nand (n203,n176,n202);
nor (n204,n205,n207);
and (n205,n206,n202);
not (n206,n47);
and (n207,n47,n208);
not (n208,n202);
not (n209,n210);
nor (n210,n211,n214);
and (n211,n212,n206);
not (n212,n213);
and (n214,n213,n47);
or (n215,n216,n217);
not (n216,n200);
nor (n217,n218,n221);
and (n218,n219,n47);
not (n219,n220);
and (n221,n220,n206);
or (n222,n223,n363);
and (n223,n224,n302);
xor (n224,n225,n265);
or (n225,n226,n264);
and (n226,n227,n247);
xor (n227,n228,n238);
nand (n228,n229,n234);
or (n229,n230,n231);
not (n230,n64);
nor (n231,n232,n233);
and (n232,n56,n83);
and (n233,n54,n85);
or (n234,n42,n235);
nor (n235,n236,n237);
and (n236,n56,n89);
and (n237,n54,n91);
nand (n238,n239,n243);
or (n239,n70,n240);
nor (n240,n241,n242);
and (n241,n78,n152);
and (n242,n79,n151);
or (n243,n71,n244);
nor (n244,n245,n246);
and (n245,n78,n167);
and (n246,n79,n166);
and (n247,n248,n254);
nor (n248,n249,n78);
nor (n249,n250,n252);
and (n250,n251,n56);
nand (n251,n101,n74);
and (n252,n253,n73);
not (n253,n101);
nand (n254,n255,n260);
or (n255,n104,n256);
not (n256,n257);
nor (n257,n258,n259);
and (n258,n37,n110);
and (n259,n38,n107);
or (n260,n261,n105);
nor (n261,n262,n263);
and (n262,n110,n141);
and (n263,n107,n143);
and (n264,n228,n238);
xor (n265,n266,n284);
xor (n266,n267,n270);
nand (n267,n268,n269);
or (n268,n70,n244);
or (n269,n71,n81);
xor (n270,n271,n277);
nor (n271,n272,n97);
nor (n272,n273,n275);
and (n273,n274,n78);
nand (n274,n101,n158);
and (n275,n253,n276);
not (n276,n158);
nand (n277,n278,n283);
or (n278,n104,n279);
not (n279,n280);
nor (n280,n281,n282);
and (n281,n126,n107);
and (n282,n125,n110);
or (n283,n108,n105);
or (n284,n285,n301);
and (n285,n286,n291);
xor (n286,n287,n288);
nor (n287,n155,n253);
nand (n288,n289,n290);
or (n289,n105,n279);
or (n290,n261,n104);
nand (n291,n292,n296);
or (n292,n135,n293);
nor (n293,n294,n295);
and (n294,n18,n27);
and (n295,n17,n28);
or (n296,n128,n297);
not (n297,n298);
nor (n298,n299,n300);
and (n299,n38,n28);
and (n300,n37,n27);
and (n301,n287,n288);
or (n302,n303,n362);
and (n303,n304,n361);
xor (n304,n305,n335);
or (n305,n306,n334);
and (n306,n307,n325);
xor (n307,n308,n315);
nand (n308,n309,n313);
or (n309,n135,n310);
nor (n310,n311,n312);
and (n311,n175,n27);
and (n312,n174,n28);
nand (n313,n314,n129);
not (n314,n293);
nand (n315,n316,n321);
or (n316,n317,n179);
not (n317,n318);
nor (n318,n319,n320);
and (n319,n213,n177);
and (n320,n212,n176);
or (n321,n192,n322);
nor (n322,n323,n324);
and (n323,n52,n177);
and (n324,n53,n176);
nand (n325,n326,n330);
or (n326,n198,n327);
nor (n327,n328,n329);
and (n328,n206,n89);
and (n329,n91,n47);
or (n330,n216,n331);
nor (n331,n332,n333);
and (n332,n206,n62);
and (n333,n47,n61);
and (n334,n308,n315);
or (n335,n336,n360);
and (n336,n337,n354);
xor (n337,n338,n348);
nand (n338,n339,n343);
or (n339,n340,n22);
nor (n340,n341,n342);
and (n341,n19,n220);
and (n342,n20,n219);
nand (n343,n344,n24);
not (n344,n345);
nor (n345,n346,n347);
and (n346,n19,n188);
and (n347,n20,n190);
nand (n348,n349,n353);
or (n349,n230,n350);
nor (n350,n351,n352);
and (n351,n56,n167);
and (n352,n54,n166);
or (n353,n42,n231);
nand (n354,n355,n359);
or (n355,n70,n356);
nor (n356,n357,n358);
and (n357,n253,n79);
and (n358,n101,n78);
or (n359,n240,n71);
and (n360,n338,n348);
xor (n361,n286,n291);
and (n362,n305,n335);
and (n363,n225,n265);
xor (n364,n365,n415);
xor (n365,n366,n369);
or (n366,n367,n368);
and (n367,n266,n284);
and (n368,n267,n270);
xor (n369,n370,n394);
xor (n370,n371,n372);
and (n371,n271,n277);
or (n372,n373,n393);
and (n373,n374,n386);
xor (n374,n375,n379);
nand (n375,n376,n377);
or (n376,n297,n135);
nand (n377,n378,n129);
not (n378,n139);
nand (n379,n380,n385);
or (n380,n381,n154);
not (n381,n382);
nand (n382,n383,n384);
or (n383,n97,n101);
or (n384,n253,n98);
nand (n385,n156,n149);
nand (n386,n387,n392);
or (n387,n192,n388);
not (n388,n389);
nor (n389,n390,n391);
and (n390,n220,n177);
and (n391,n219,n176);
or (n392,n179,n186);
and (n393,n375,n379);
or (n394,n395,n414);
and (n395,n396,n411);
xor (n396,n397,n404);
nand (n397,n398,n403);
or (n398,n399,n198);
not (n399,n400);
nor (n400,n401,n402);
and (n401,n52,n206);
and (n402,n53,n47);
nand (n403,n200,n210);
nand (n404,n405,n407);
or (n405,n14,n406);
not (n406,n24);
or (n407,n22,n408);
nor (n408,n409,n410);
and (n409,n19,n175);
and (n410,n20,n174);
nand (n411,n412,n413);
or (n412,n230,n235);
or (n413,n42,n59);
and (n414,n397,n404);
or (n415,n416,n433);
and (n416,n417,n432);
xor (n417,n418,n431);
or (n418,n419,n430);
and (n419,n420,n427);
xor (n420,n421,n424);
nand (n421,n422,n423);
or (n422,n317,n192);
nand (n423,n180,n389);
nand (n424,n425,n426);
or (n425,n198,n331);
nand (n426,n200,n400);
nand (n427,n428,n429);
or (n428,n22,n345);
or (n429,n406,n408);
and (n430,n421,n424);
xor (n431,n396,n411);
xor (n432,n374,n386);
and (n433,n418,n431);
or (n434,n435,n492);
and (n435,n436,n491);
xor (n436,n437,n438);
xor (n437,n417,n432);
or (n438,n439,n490);
and (n439,n440,n443);
xor (n440,n441,n442);
xor (n441,n420,n427);
xor (n442,n227,n247);
or (n443,n444,n489);
and (n444,n445,n464);
xor (n445,n446,n447);
xor (n446,n248,n254);
or (n447,n448,n463);
and (n448,n449,n456);
xor (n449,n450,n451);
nor (n450,n71,n253);
nand (n451,n452,n454);
or (n452,n135,n453);
xor (n453,n188,n27);
nand (n454,n455,n129);
not (n455,n310);
nand (n456,n457,n462);
or (n457,n192,n458);
not (n458,n459);
nor (n459,n460,n461);
and (n460,n61,n176);
and (n461,n62,n177);
or (n462,n179,n322);
and (n463,n450,n451);
or (n464,n465,n488);
and (n465,n466,n482);
xor (n466,n467,n475);
nand (n467,n468,n473);
or (n468,n469,n198);
not (n469,n470);
nand (n470,n471,n472);
or (n471,n47,n85);
or (n472,n83,n206);
nand (n473,n474,n200);
not (n474,n327);
nand (n475,n476,n481);
or (n476,n104,n477);
not (n477,n478);
nor (n478,n479,n480);
and (n479,n17,n110);
and (n480,n18,n107);
nand (n481,n257,n106);
nand (n482,n483,n487);
or (n483,n230,n484);
nor (n484,n485,n486);
and (n485,n56,n152);
and (n486,n54,n151);
or (n487,n42,n350);
and (n488,n467,n475);
and (n489,n446,n447);
and (n490,n441,n442);
xor (n491,n224,n302);
and (n492,n437,n438);
nand (n493,n6,n434);
not (n494,n495);
nand (n495,n496,n711);
nor (n496,n497,n710);
and (n497,n498,n562);
nand (n498,n499,n501);
not (n499,n500);
xor (n500,n436,n491);
not (n501,n502);
or (n502,n503,n561);
and (n503,n504,n507);
xor (n504,n505,n506);
xor (n505,n304,n361);
xor (n506,n440,n443);
or (n507,n508,n560);
and (n508,n509,n512);
xor (n509,n510,n511);
xor (n510,n337,n354);
xor (n511,n307,n325);
or (n512,n513,n559);
and (n513,n514,n535);
xor (n514,n515,n521);
nand (n515,n516,n520);
or (n516,n22,n517);
nor (n517,n518,n519);
and (n518,n19,n213);
and (n519,n20,n212);
or (n520,n406,n340);
and (n521,n522,n528);
nand (n522,n523,n524);
or (n523,n453,n128);
or (n524,n135,n525);
nor (n525,n526,n527);
and (n526,n220,n27);
and (n527,n219,n28);
not (n528,n529);
nand (n529,n530,n54);
nand (n530,n531,n532);
or (n531,n101,n46);
nand (n532,n533,n206);
not (n533,n534);
and (n534,n101,n46);
or (n535,n536,n558);
and (n536,n537,n552);
xor (n537,n538,n545);
nand (n538,n539,n544);
or (n539,n540,n192);
not (n540,n541);
nand (n541,n542,n543);
or (n542,n177,n91);
or (n543,n176,n89);
nand (n544,n180,n459);
nand (n545,n546,n551);
or (n546,n547,n198);
not (n547,n548);
nand (n548,n549,n550);
or (n549,n47,n166);
or (n550,n206,n167);
nand (n551,n200,n470);
nand (n552,n553,n554);
or (n553,n105,n477);
or (n554,n555,n104);
nor (n555,n556,n557);
and (n556,n110,n175);
and (n557,n107,n174);
and (n558,n538,n545);
and (n559,n515,n521);
and (n560,n510,n511);
and (n561,n505,n506);
nand (n562,n563,n709);
or (n563,n564,n701);
not (n564,n565);
nand (n565,n566,n700);
or (n566,n567,n650);
nor (n567,n568,n598);
xor (n568,n569,n597);
xor (n569,n570,n571);
xor (n570,n445,n464);
or (n571,n572,n596);
and (n572,n573,n576);
xor (n573,n574,n575);
xor (n574,n466,n482);
xor (n575,n449,n456);
or (n576,n577,n595);
and (n577,n578,n591);
xor (n578,n579,n585);
nand (n579,n580,n584);
or (n580,n230,n581);
nor (n581,n582,n583);
and (n582,n253,n54);
and (n583,n101,n56);
or (n584,n42,n484);
nand (n585,n586,n590);
or (n586,n22,n587);
nor (n587,n588,n589);
and (n588,n19,n53);
and (n589,n20,n52);
or (n590,n406,n517);
nand (n591,n592,n594);
or (n592,n528,n593);
not (n593,n522);
or (n594,n522,n529);
and (n595,n579,n585);
and (n596,n574,n575);
xor (n597,n509,n512);
or (n598,n599,n649);
and (n599,n600,n648);
xor (n600,n601,n602);
xor (n601,n514,n535);
or (n602,n603,n647);
and (n603,n604,n646);
xor (n604,n605,n623);
or (n605,n606,n622);
and (n606,n607,n616);
xor (n607,n608,n609);
nor (n608,n42,n253);
nand (n609,n610,n614);
or (n610,n611,n135);
nor (n611,n612,n613);
and (n612,n27,n213);
and (n613,n28,n212);
nand (n614,n615,n129);
not (n615,n525);
nand (n616,n617,n618);
or (n617,n540,n179);
or (n618,n192,n619);
nor (n619,n620,n621);
and (n620,n176,n83);
and (n621,n177,n85);
and (n622,n608,n609);
or (n623,n624,n645);
and (n624,n625,n639);
xor (n625,n626,n633);
nand (n626,n627,n632);
or (n627,n628,n198);
not (n628,n629);
nand (n629,n630,n631);
or (n630,n47,n151);
or (n631,n206,n152);
nand (n632,n200,n548);
nand (n633,n634,n638);
or (n634,n635,n104);
nor (n635,n636,n637);
and (n636,n110,n188);
and (n637,n107,n190);
or (n638,n555,n105);
nand (n639,n640,n644);
or (n640,n22,n641);
nor (n641,n642,n643);
and (n642,n19,n62);
and (n643,n20,n61);
or (n644,n406,n587);
and (n645,n626,n633);
xor (n646,n537,n552);
and (n647,n605,n623);
xor (n648,n573,n576);
and (n649,n601,n602);
nand (n650,n651,n699);
or (n651,n652,n698);
and (n652,n653,n656);
xor (n653,n654,n655);
xor (n654,n578,n591);
xor (n655,n604,n646);
or (n656,n657,n697);
and (n657,n658,n696);
xor (n658,n659,n672);
and (n659,n660,n666);
and (n660,n661,n47);
nand (n661,n662,n663);
or (n662,n101,n202);
nand (n663,n664,n176);
not (n664,n665);
and (n665,n101,n202);
nand (n666,n667,n671);
or (n667,n135,n668);
nor (n668,n669,n670);
and (n669,n27,n53);
and (n670,n28,n52);
or (n671,n128,n611);
or (n672,n673,n695);
and (n673,n674,n689);
xor (n674,n675,n682);
nand (n675,n676,n680);
or (n676,n677,n192);
nor (n677,n678,n679);
and (n678,n176,n167);
and (n679,n177,n166);
nand (n680,n681,n180);
not (n681,n619);
nand (n682,n683,n684);
or (n683,n628,n216);
nand (n684,n685,n199);
not (n685,n686);
nor (n686,n687,n688);
and (n687,n253,n47);
and (n688,n206,n101);
nand (n689,n690,n694);
or (n690,n104,n691);
nor (n691,n692,n693);
and (n692,n110,n220);
and (n693,n107,n219);
or (n694,n635,n105);
and (n695,n675,n682);
xor (n696,n607,n616);
and (n697,n659,n672);
and (n698,n654,n655);
xor (n699,n600,n648);
nand (n700,n568,n598);
not (n701,n702);
nand (n702,n703,n705);
not (n703,n704);
xor (n704,n504,n507);
not (n705,n706);
or (n706,n707,n708);
and (n707,n569,n597);
and (n708,n570,n571);
nand (n709,n704,n706);
nor (n710,n499,n501);
nand (n711,n712,n498,n1001);
nand (n712,n713,n1000);
or (n713,n714,n751);
not (n714,n715);
or (n715,n716,n717);
xor (n716,n653,n656);
or (n717,n718,n750);
and (n718,n719,n749);
xor (n719,n720,n721);
xor (n720,n625,n639);
or (n721,n722,n748);
and (n722,n723,n731);
xor (n723,n724,n730);
nand (n724,n725,n729);
or (n725,n22,n726);
nor (n726,n727,n728);
and (n727,n19,n89);
and (n728,n20,n91);
or (n729,n406,n641);
xor (n730,n660,n666);
or (n731,n732,n747);
and (n732,n733,n741);
xor (n733,n734,n735);
nor (n734,n216,n253);
nand (n735,n736,n740);
or (n736,n737,n104);
nor (n737,n738,n739);
and (n738,n212,n107);
and (n739,n213,n110);
or (n740,n691,n105);
nand (n741,n742,n746);
or (n742,n192,n743);
nor (n743,n744,n745);
and (n744,n176,n152);
and (n745,n177,n151);
or (n746,n179,n677);
and (n747,n734,n735);
and (n748,n724,n730);
xor (n749,n658,n696);
and (n750,n720,n721);
not (n751,n752);
or (n752,n753,n999);
and (n753,n754,n794);
xor (n754,n755,n793);
or (n755,n756,n792);
and (n756,n757,n791);
xor (n757,n758,n759);
xor (n758,n674,n689);
or (n759,n760,n790);
and (n760,n761,n776);
xor (n761,n762,n770);
nand (n762,n763,n768);
or (n763,n764,n135);
not (n764,n765);
nand (n765,n766,n767);
or (n766,n28,n61);
or (n767,n27,n62);
nand (n768,n769,n129);
not (n769,n668);
nand (n770,n771,n775);
or (n771,n22,n772);
nor (n772,n773,n774);
and (n773,n19,n83);
and (n774,n20,n85);
or (n775,n406,n726);
and (n776,n777,n783);
nor (n777,n778,n176);
nor (n778,n779,n781);
and (n779,n253,n780);
not (n780,n182);
nor (n781,n782,n20);
and (n782,n101,n182);
nand (n783,n784,n789);
or (n784,n104,n785);
not (n785,n786);
nor (n786,n787,n788);
and (n787,n52,n110);
and (n788,n53,n107);
or (n789,n737,n105);
and (n790,n762,n770);
xor (n791,n723,n731);
and (n792,n758,n759);
xor (n793,n719,n749);
nand (n794,n795,n996,n998);
nand (n795,n796,n831,n991);
nand (n796,n797,n799);
not (n797,n798);
xor (n798,n757,n791);
not (n799,n800);
or (n800,n801,n830);
and (n801,n802,n829);
xor (n802,n803,n828);
or (n803,n804,n827);
and (n804,n805,n821);
xor (n805,n806,n814);
nand (n806,n807,n812);
or (n807,n808,n192);
not (n808,n809);
nand (n809,n810,n811);
or (n810,n176,n101);
or (n811,n253,n177);
nand (n812,n813,n180);
not (n813,n743);
nand (n814,n815,n820);
or (n815,n816,n135);
not (n816,n817);
nand (n817,n818,n819);
or (n818,n28,n91);
or (n819,n27,n89);
nand (n820,n129,n765);
nand (n821,n822,n826);
or (n822,n22,n823);
nor (n823,n824,n825);
and (n824,n19,n167);
and (n825,n20,n166);
or (n826,n406,n772);
and (n827,n806,n814);
xor (n828,n733,n741);
xor (n829,n761,n776);
and (n830,n803,n828);
nand (n831,n832,n990);
or (n832,n833,n883);
not (n833,n834);
nand (n834,n835,n859);
not (n835,n836);
xor (n836,n837,n858);
xor (n837,n838,n839);
xor (n838,n777,n783);
or (n839,n840,n857);
and (n840,n841,n850);
xor (n841,n842,n843);
and (n842,n180,n101);
nand (n843,n844,n849);
or (n844,n104,n845);
not (n845,n846);
nor (n846,n847,n848);
and (n847,n61,n110);
and (n848,n62,n107);
nand (n849,n786,n106);
nand (n850,n851,n856);
or (n851,n852,n135);
not (n852,n853);
nor (n853,n854,n855);
and (n854,n85,n27);
and (n855,n83,n28);
nand (n856,n129,n817);
and (n857,n842,n843);
xor (n858,n805,n821);
not (n859,n860);
or (n860,n861,n882);
and (n861,n862,n881);
xor (n862,n863,n869);
nand (n863,n864,n868);
or (n864,n22,n865);
nor (n865,n866,n867);
and (n866,n151,n20);
and (n867,n152,n19);
or (n868,n406,n823);
and (n869,n870,n875);
and (n870,n871,n20);
nand (n871,n872,n874);
or (n872,n873,n28);
and (n873,n101,n26);
or (n874,n101,n26);
nand (n875,n876,n877);
or (n876,n105,n845);
or (n877,n878,n104);
nor (n878,n879,n880);
and (n879,n110,n89);
and (n880,n107,n91);
xor (n881,n841,n850);
and (n882,n863,n869);
not (n883,n884);
nand (n884,n885,n989);
or (n885,n886,n909);
not (n886,n887);
nand (n887,n888,n890);
not (n888,n889);
xor (n889,n862,n881);
not (n890,n891);
or (n891,n892,n908);
and (n892,n893,n907);
xor (n893,n894,n901);
nand (n894,n895,n900);
or (n895,n896,n135);
not (n896,n897);
nor (n897,n898,n899);
and (n898,n166,n27);
and (n899,n167,n28);
nand (n900,n853,n129);
nand (n901,n902,n903);
or (n902,n406,n865);
nand (n903,n23,n904);
nand (n904,n905,n906);
or (n905,n101,n19);
or (n906,n253,n20);
xor (n907,n870,n875);
and (n908,n894,n901);
not (n909,n910);
or (n910,n911,n988);
and (n911,n912,n933);
xor (n912,n913,n932);
or (n913,n914,n931);
and (n914,n915,n924);
xor (n915,n916,n917);
and (n916,n24,n101);
nand (n917,n918,n923);
or (n918,n919,n135);
not (n919,n920);
nor (n920,n921,n922);
and (n921,n151,n27);
and (n922,n152,n28);
nand (n923,n897,n129);
nand (n924,n925,n930);
or (n925,n104,n926);
not (n926,n927);
nor (n927,n928,n929);
and (n928,n85,n110);
and (n929,n83,n107);
or (n930,n878,n105);
and (n931,n916,n917);
xor (n932,n893,n907);
nand (n933,n934,n987);
or (n934,n935,n951);
nor (n935,n936,n937);
xor (n936,n915,n924);
nor (n937,n938,n946);
not (n938,n939);
nand (n939,n940,n941);
or (n940,n105,n926);
nand (n941,n942,n945);
nand (n942,n943,n944);
or (n943,n167,n110);
nand (n944,n110,n167);
not (n945,n104);
nand (n946,n947,n28);
nand (n947,n948,n950);
or (n948,n949,n107);
and (n949,n101,n132);
or (n950,n101,n132);
nor (n951,n952,n986);
and (n952,n953,n965);
nand (n953,n954,n961);
not (n954,n955);
nand (n955,n956,n960);
or (n956,n135,n957);
nor (n957,n958,n959);
and (n958,n28,n253);
and (n959,n101,n27);
or (n960,n128,n919);
nor (n961,n962,n963);
and (n962,n946,n939);
and (n963,n964,n938);
not (n964,n946);
or (n965,n966,n985);
and (n966,n967,n976);
xor (n967,n968,n969);
nor (n968,n128,n253);
nand (n969,n970,n975);
or (n970,n104,n971);
not (n971,n972);
nand (n972,n973,n974);
or (n973,n151,n107);
nand (n974,n107,n151);
nand (n975,n942,n106);
nor (n976,n977,n983);
nor (n977,n978,n979);
and (n978,n972,n106);
nor (n979,n980,n104);
nor (n980,n981,n982);
and (n981,n253,n107);
and (n982,n101,n110);
or (n983,n984,n110);
and (n984,n101,n106);
and (n985,n968,n969);
nor (n986,n954,n961);
nand (n987,n936,n937);
and (n988,n913,n932);
nand (n989,n889,n891);
nand (n990,n836,n860);
or (n991,n992,n995);
or (n992,n993,n994);
and (n993,n837,n858);
and (n994,n838,n839);
xor (n995,n802,n829);
nand (n996,n796,n997);
and (n997,n995,n992);
nand (n998,n800,n798);
and (n999,n755,n793);
nand (n1000,n716,n717);
nor (n1001,n701,n1002);
nand (n1002,n1003,n1004);
not (n1003,n567);
or (n1004,n651,n699);
or (n1005,n495,n3);
xor (n1006,n1007,n1706);
xor (n1007,n1008,n1703);
xor (n1008,n1009,n153);
xor (n1009,n1010,n1694);
xor (n1010,n1011,n1693);
xor (n1011,n1012,n1678);
xor (n1012,n1013,n1677);
xor (n1013,n1014,n1656);
xor (n1014,n1015,n1655);
xor (n1015,n1016,n1628);
xor (n1016,n1017,n1627);
xor (n1017,n1018,n1595);
xor (n1018,n1019,n1594);
xor (n1019,n1020,n1556);
xor (n1020,n1021,n214);
xor (n1021,n1022,n1512);
xor (n1022,n1023,n1511);
xor (n1023,n1024,n1463);
xor (n1024,n1025,n1462);
xor (n1025,n1026,n1406);
xor (n1026,n1027,n1405);
xor (n1027,n1028,n1342);
xor (n1028,n1029,n21);
xor (n1029,n1030,n1274);
xor (n1030,n1031,n1273);
xor (n1031,n1032,n1202);
xor (n1032,n1033,n1201);
xor (n1033,n1034,n1121);
xor (n1034,n1035,n1120);
xor (n1035,n1036,n1039);
xor (n1036,n1037,n1038);
and (n1037,n118,n106);
and (n1038,n111,n107);
or (n1039,n1040,n1042);
and (n1040,n1041,n281);
and (n1041,n111,n106);
and (n1042,n1043,n1044);
xor (n1043,n1041,n281);
or (n1044,n1045,n1048);
and (n1045,n1046,n1047);
and (n1046,n126,n106);
and (n1047,n141,n107);
and (n1048,n1049,n1050);
xor (n1049,n1046,n1047);
or (n1050,n1051,n1053);
and (n1051,n1052,n259);
and (n1052,n141,n106);
and (n1053,n1054,n1055);
xor (n1054,n1052,n259);
or (n1055,n1056,n1058);
and (n1056,n1057,n480);
and (n1057,n38,n106);
and (n1058,n1059,n1060);
xor (n1059,n1057,n480);
or (n1060,n1061,n1064);
and (n1061,n1062,n1063);
and (n1062,n18,n106);
and (n1063,n175,n107);
and (n1064,n1065,n1066);
xor (n1065,n1062,n1063);
or (n1066,n1067,n1070);
and (n1067,n1068,n1069);
and (n1068,n175,n106);
and (n1069,n188,n107);
and (n1070,n1071,n1072);
xor (n1071,n1068,n1069);
or (n1072,n1073,n1076);
and (n1073,n1074,n1075);
and (n1074,n188,n106);
and (n1075,n220,n107);
and (n1076,n1077,n1078);
xor (n1077,n1074,n1075);
or (n1078,n1079,n1082);
and (n1079,n1080,n1081);
and (n1080,n220,n106);
and (n1081,n213,n107);
and (n1082,n1083,n1084);
xor (n1083,n1080,n1081);
or (n1084,n1085,n1087);
and (n1085,n1086,n788);
and (n1086,n213,n106);
and (n1087,n1088,n1089);
xor (n1088,n1086,n788);
or (n1089,n1090,n1092);
and (n1090,n1091,n848);
and (n1091,n53,n106);
and (n1092,n1093,n1094);
xor (n1093,n1091,n848);
or (n1094,n1095,n1098);
and (n1095,n1096,n1097);
and (n1096,n62,n106);
and (n1097,n89,n107);
and (n1098,n1099,n1100);
xor (n1099,n1096,n1097);
or (n1100,n1101,n1103);
and (n1101,n1102,n929);
and (n1102,n89,n106);
and (n1103,n1104,n1105);
xor (n1104,n1102,n929);
or (n1105,n1106,n1109);
and (n1106,n1107,n1108);
and (n1107,n83,n106);
and (n1108,n167,n107);
and (n1109,n1110,n1111);
xor (n1110,n1107,n1108);
or (n1111,n1112,n1115);
and (n1112,n1113,n1114);
and (n1113,n167,n106);
and (n1114,n152,n107);
and (n1115,n1116,n1117);
xor (n1116,n1113,n1114);
and (n1117,n1118,n1119);
and (n1118,n152,n106);
and (n1119,n101,n107);
and (n1120,n126,n132);
or (n1121,n1122,n1125);
and (n1122,n1123,n1124);
xor (n1123,n1043,n1044);
and (n1124,n141,n132);
and (n1125,n1126,n1127);
xor (n1126,n1123,n1124);
or (n1127,n1128,n1131);
and (n1128,n1129,n1130);
xor (n1129,n1049,n1050);
and (n1130,n38,n132);
and (n1131,n1132,n1133);
xor (n1132,n1129,n1130);
or (n1133,n1134,n1137);
and (n1134,n1135,n1136);
xor (n1135,n1054,n1055);
and (n1136,n18,n132);
and (n1137,n1138,n1139);
xor (n1138,n1135,n1136);
or (n1139,n1140,n1143);
and (n1140,n1141,n1142);
xor (n1141,n1059,n1060);
and (n1142,n175,n132);
and (n1143,n1144,n1145);
xor (n1144,n1141,n1142);
or (n1145,n1146,n1149);
and (n1146,n1147,n1148);
xor (n1147,n1065,n1066);
and (n1148,n188,n132);
and (n1149,n1150,n1151);
xor (n1150,n1147,n1148);
or (n1151,n1152,n1155);
and (n1152,n1153,n1154);
xor (n1153,n1071,n1072);
and (n1154,n220,n132);
and (n1155,n1156,n1157);
xor (n1156,n1153,n1154);
or (n1157,n1158,n1161);
and (n1158,n1159,n1160);
xor (n1159,n1077,n1078);
and (n1160,n213,n132);
and (n1161,n1162,n1163);
xor (n1162,n1159,n1160);
or (n1163,n1164,n1167);
and (n1164,n1165,n1166);
xor (n1165,n1083,n1084);
and (n1166,n53,n132);
and (n1167,n1168,n1169);
xor (n1168,n1165,n1166);
or (n1169,n1170,n1173);
and (n1170,n1171,n1172);
xor (n1171,n1088,n1089);
and (n1172,n62,n132);
and (n1173,n1174,n1175);
xor (n1174,n1171,n1172);
or (n1175,n1176,n1179);
and (n1176,n1177,n1178);
xor (n1177,n1093,n1094);
and (n1178,n89,n132);
and (n1179,n1180,n1181);
xor (n1180,n1177,n1178);
or (n1181,n1182,n1185);
and (n1182,n1183,n1184);
xor (n1183,n1099,n1100);
and (n1184,n83,n132);
and (n1185,n1186,n1187);
xor (n1186,n1183,n1184);
or (n1187,n1188,n1191);
and (n1188,n1189,n1190);
xor (n1189,n1104,n1105);
and (n1190,n167,n132);
and (n1191,n1192,n1193);
xor (n1192,n1189,n1190);
or (n1193,n1194,n1197);
and (n1194,n1195,n1196);
xor (n1195,n1110,n1111);
and (n1196,n152,n132);
and (n1197,n1198,n1199);
xor (n1198,n1195,n1196);
and (n1199,n1200,n949);
xor (n1200,n1116,n1117);
and (n1201,n141,n28);
or (n1202,n1203,n1205);
and (n1203,n1204,n299);
xor (n1204,n1126,n1127);
and (n1205,n1206,n1207);
xor (n1206,n1204,n299);
or (n1207,n1208,n1211);
and (n1208,n1209,n1210);
xor (n1209,n1132,n1133);
and (n1210,n18,n28);
and (n1211,n1212,n1213);
xor (n1212,n1209,n1210);
or (n1213,n1214,n1217);
and (n1214,n1215,n1216);
xor (n1215,n1138,n1139);
and (n1216,n175,n28);
and (n1217,n1218,n1219);
xor (n1218,n1215,n1216);
or (n1219,n1220,n1223);
and (n1220,n1221,n1222);
xor (n1221,n1144,n1145);
and (n1222,n188,n28);
and (n1223,n1224,n1225);
xor (n1224,n1221,n1222);
or (n1225,n1226,n1229);
and (n1226,n1227,n1228);
xor (n1227,n1150,n1151);
and (n1228,n220,n28);
and (n1229,n1230,n1231);
xor (n1230,n1227,n1228);
or (n1231,n1232,n1235);
and (n1232,n1233,n1234);
xor (n1233,n1156,n1157);
and (n1234,n213,n28);
and (n1235,n1236,n1237);
xor (n1236,n1233,n1234);
or (n1237,n1238,n1241);
and (n1238,n1239,n1240);
xor (n1239,n1162,n1163);
and (n1240,n53,n28);
and (n1241,n1242,n1243);
xor (n1242,n1239,n1240);
or (n1243,n1244,n1247);
and (n1244,n1245,n1246);
xor (n1245,n1168,n1169);
and (n1246,n62,n28);
and (n1247,n1248,n1249);
xor (n1248,n1245,n1246);
or (n1249,n1250,n1253);
and (n1250,n1251,n1252);
xor (n1251,n1174,n1175);
and (n1252,n89,n28);
and (n1253,n1254,n1255);
xor (n1254,n1251,n1252);
or (n1255,n1256,n1258);
and (n1256,n1257,n855);
xor (n1257,n1180,n1181);
and (n1258,n1259,n1260);
xor (n1259,n1257,n855);
or (n1260,n1261,n1263);
and (n1261,n1262,n899);
xor (n1262,n1186,n1187);
and (n1263,n1264,n1265);
xor (n1264,n1262,n899);
or (n1265,n1266,n1268);
and (n1266,n1267,n922);
xor (n1267,n1192,n1193);
and (n1268,n1269,n1270);
xor (n1269,n1267,n922);
and (n1270,n1271,n1272);
xor (n1271,n1198,n1199);
and (n1272,n101,n28);
and (n1273,n38,n26);
or (n1274,n1275,n1278);
and (n1275,n1276,n1277);
xor (n1276,n1206,n1207);
and (n1277,n18,n26);
and (n1278,n1279,n1280);
xor (n1279,n1276,n1277);
or (n1280,n1281,n1284);
and (n1281,n1282,n1283);
xor (n1282,n1212,n1213);
and (n1283,n175,n26);
and (n1284,n1285,n1286);
xor (n1285,n1282,n1283);
or (n1286,n1287,n1290);
and (n1287,n1288,n1289);
xor (n1288,n1218,n1219);
and (n1289,n188,n26);
and (n1290,n1291,n1292);
xor (n1291,n1288,n1289);
or (n1292,n1293,n1296);
and (n1293,n1294,n1295);
xor (n1294,n1224,n1225);
and (n1295,n220,n26);
and (n1296,n1297,n1298);
xor (n1297,n1294,n1295);
or (n1298,n1299,n1302);
and (n1299,n1300,n1301);
xor (n1300,n1230,n1231);
and (n1301,n213,n26);
and (n1302,n1303,n1304);
xor (n1303,n1300,n1301);
or (n1304,n1305,n1308);
and (n1305,n1306,n1307);
xor (n1306,n1236,n1237);
and (n1307,n53,n26);
and (n1308,n1309,n1310);
xor (n1309,n1306,n1307);
or (n1310,n1311,n1314);
and (n1311,n1312,n1313);
xor (n1312,n1242,n1243);
and (n1313,n62,n26);
and (n1314,n1315,n1316);
xor (n1315,n1312,n1313);
or (n1316,n1317,n1320);
and (n1317,n1318,n1319);
xor (n1318,n1248,n1249);
and (n1319,n89,n26);
and (n1320,n1321,n1322);
xor (n1321,n1318,n1319);
or (n1322,n1323,n1326);
and (n1323,n1324,n1325);
xor (n1324,n1254,n1255);
and (n1325,n83,n26);
and (n1326,n1327,n1328);
xor (n1327,n1324,n1325);
or (n1328,n1329,n1332);
and (n1329,n1330,n1331);
xor (n1330,n1259,n1260);
and (n1331,n167,n26);
and (n1332,n1333,n1334);
xor (n1333,n1330,n1331);
or (n1334,n1335,n1338);
and (n1335,n1336,n1337);
xor (n1336,n1264,n1265);
and (n1337,n152,n26);
and (n1338,n1339,n1340);
xor (n1339,n1336,n1337);
and (n1340,n1341,n873);
xor (n1341,n1269,n1270);
or (n1342,n1343,n1346);
and (n1343,n1344,n1345);
xor (n1344,n1279,n1280);
and (n1345,n175,n20);
and (n1346,n1347,n1348);
xor (n1347,n1344,n1345);
or (n1348,n1349,n1352);
and (n1349,n1350,n1351);
xor (n1350,n1285,n1286);
and (n1351,n188,n20);
and (n1352,n1353,n1354);
xor (n1353,n1350,n1351);
or (n1354,n1355,n1358);
and (n1355,n1356,n1357);
xor (n1356,n1291,n1292);
and (n1357,n220,n20);
and (n1358,n1359,n1360);
xor (n1359,n1356,n1357);
or (n1360,n1361,n1364);
and (n1361,n1362,n1363);
xor (n1362,n1297,n1298);
and (n1363,n213,n20);
and (n1364,n1365,n1366);
xor (n1365,n1362,n1363);
or (n1366,n1367,n1370);
and (n1367,n1368,n1369);
xor (n1368,n1303,n1304);
and (n1369,n53,n20);
and (n1370,n1371,n1372);
xor (n1371,n1368,n1369);
or (n1372,n1373,n1376);
and (n1373,n1374,n1375);
xor (n1374,n1309,n1310);
and (n1375,n62,n20);
and (n1376,n1377,n1378);
xor (n1377,n1374,n1375);
or (n1378,n1379,n1382);
and (n1379,n1380,n1381);
xor (n1380,n1315,n1316);
and (n1381,n89,n20);
and (n1382,n1383,n1384);
xor (n1383,n1380,n1381);
or (n1384,n1385,n1388);
and (n1385,n1386,n1387);
xor (n1386,n1321,n1322);
and (n1387,n83,n20);
and (n1388,n1389,n1390);
xor (n1389,n1386,n1387);
or (n1390,n1391,n1394);
and (n1391,n1392,n1393);
xor (n1392,n1327,n1328);
and (n1393,n167,n20);
and (n1394,n1395,n1396);
xor (n1395,n1392,n1393);
or (n1396,n1397,n1400);
and (n1397,n1398,n1399);
xor (n1398,n1333,n1334);
and (n1399,n152,n20);
and (n1400,n1401,n1402);
xor (n1401,n1398,n1399);
and (n1402,n1403,n1404);
xor (n1403,n1339,n1340);
and (n1404,n101,n20);
and (n1405,n175,n182);
or (n1406,n1407,n1410);
and (n1407,n1408,n1409);
xor (n1408,n1347,n1348);
and (n1409,n188,n182);
and (n1410,n1411,n1412);
xor (n1411,n1408,n1409);
or (n1412,n1413,n1416);
and (n1413,n1414,n1415);
xor (n1414,n1353,n1354);
and (n1415,n220,n182);
and (n1416,n1417,n1418);
xor (n1417,n1414,n1415);
or (n1418,n1419,n1422);
and (n1419,n1420,n1421);
xor (n1420,n1359,n1360);
and (n1421,n213,n182);
and (n1422,n1423,n1424);
xor (n1423,n1420,n1421);
or (n1424,n1425,n1428);
and (n1425,n1426,n1427);
xor (n1426,n1365,n1366);
and (n1427,n53,n182);
and (n1428,n1429,n1430);
xor (n1429,n1426,n1427);
or (n1430,n1431,n1434);
and (n1431,n1432,n1433);
xor (n1432,n1371,n1372);
and (n1433,n62,n182);
and (n1434,n1435,n1436);
xor (n1435,n1432,n1433);
or (n1436,n1437,n1440);
and (n1437,n1438,n1439);
xor (n1438,n1377,n1378);
and (n1439,n89,n182);
and (n1440,n1441,n1442);
xor (n1441,n1438,n1439);
or (n1442,n1443,n1446);
and (n1443,n1444,n1445);
xor (n1444,n1383,n1384);
and (n1445,n83,n182);
and (n1446,n1447,n1448);
xor (n1447,n1444,n1445);
or (n1448,n1449,n1452);
and (n1449,n1450,n1451);
xor (n1450,n1389,n1390);
and (n1451,n167,n182);
and (n1452,n1453,n1454);
xor (n1453,n1450,n1451);
or (n1454,n1455,n1458);
and (n1455,n1456,n1457);
xor (n1456,n1395,n1396);
and (n1457,n152,n182);
and (n1458,n1459,n1460);
xor (n1459,n1456,n1457);
and (n1460,n1461,n782);
xor (n1461,n1401,n1402);
and (n1462,n188,n177);
or (n1463,n1464,n1466);
and (n1464,n1465,n390);
xor (n1465,n1411,n1412);
and (n1466,n1467,n1468);
xor (n1467,n1465,n390);
or (n1468,n1469,n1471);
and (n1469,n1470,n319);
xor (n1470,n1417,n1418);
and (n1471,n1472,n1473);
xor (n1472,n1470,n319);
or (n1473,n1474,n1477);
and (n1474,n1475,n1476);
xor (n1475,n1423,n1424);
and (n1476,n53,n177);
and (n1477,n1478,n1479);
xor (n1478,n1475,n1476);
or (n1479,n1480,n1482);
and (n1480,n1481,n461);
xor (n1481,n1429,n1430);
and (n1482,n1483,n1484);
xor (n1483,n1481,n461);
or (n1484,n1485,n1488);
and (n1485,n1486,n1487);
xor (n1486,n1435,n1436);
and (n1487,n89,n177);
and (n1488,n1489,n1490);
xor (n1489,n1486,n1487);
or (n1490,n1491,n1494);
and (n1491,n1492,n1493);
xor (n1492,n1441,n1442);
and (n1493,n83,n177);
and (n1494,n1495,n1496);
xor (n1495,n1492,n1493);
or (n1496,n1497,n1500);
and (n1497,n1498,n1499);
xor (n1498,n1447,n1448);
and (n1499,n167,n177);
and (n1500,n1501,n1502);
xor (n1501,n1498,n1499);
or (n1502,n1503,n1506);
and (n1503,n1504,n1505);
xor (n1504,n1453,n1454);
and (n1505,n152,n177);
and (n1506,n1507,n1508);
xor (n1507,n1504,n1505);
and (n1508,n1509,n1510);
xor (n1509,n1459,n1460);
and (n1510,n101,n177);
and (n1511,n220,n202);
or (n1512,n1513,n1516);
and (n1513,n1514,n1515);
xor (n1514,n1467,n1468);
and (n1515,n213,n202);
and (n1516,n1517,n1518);
xor (n1517,n1514,n1515);
or (n1518,n1519,n1522);
and (n1519,n1520,n1521);
xor (n1520,n1472,n1473);
and (n1521,n53,n202);
and (n1522,n1523,n1524);
xor (n1523,n1520,n1521);
or (n1524,n1525,n1528);
and (n1525,n1526,n1527);
xor (n1526,n1478,n1479);
and (n1527,n62,n202);
and (n1528,n1529,n1530);
xor (n1529,n1526,n1527);
or (n1530,n1531,n1534);
and (n1531,n1532,n1533);
xor (n1532,n1483,n1484);
and (n1533,n89,n202);
and (n1534,n1535,n1536);
xor (n1535,n1532,n1533);
or (n1536,n1537,n1540);
and (n1537,n1538,n1539);
xor (n1538,n1489,n1490);
and (n1539,n83,n202);
and (n1540,n1541,n1542);
xor (n1541,n1538,n1539);
or (n1542,n1543,n1546);
and (n1543,n1544,n1545);
xor (n1544,n1495,n1496);
and (n1545,n167,n202);
and (n1546,n1547,n1548);
xor (n1547,n1544,n1545);
or (n1548,n1549,n1552);
and (n1549,n1550,n1551);
xor (n1550,n1501,n1502);
and (n1551,n152,n202);
and (n1552,n1553,n1554);
xor (n1553,n1550,n1551);
and (n1554,n1555,n665);
xor (n1555,n1507,n1508);
or (n1556,n1557,n1559);
and (n1557,n1558,n402);
xor (n1558,n1517,n1518);
and (n1559,n1560,n1561);
xor (n1560,n1558,n402);
or (n1561,n1562,n1565);
and (n1562,n1563,n1564);
xor (n1563,n1523,n1524);
and (n1564,n62,n47);
and (n1565,n1566,n1567);
xor (n1566,n1563,n1564);
or (n1567,n1568,n1571);
and (n1568,n1569,n1570);
xor (n1569,n1529,n1530);
and (n1570,n89,n47);
and (n1571,n1572,n1573);
xor (n1572,n1569,n1570);
or (n1573,n1574,n1577);
and (n1574,n1575,n1576);
xor (n1575,n1535,n1536);
and (n1576,n83,n47);
and (n1577,n1578,n1579);
xor (n1578,n1575,n1576);
or (n1579,n1580,n1583);
and (n1580,n1581,n1582);
xor (n1581,n1541,n1542);
and (n1582,n167,n47);
and (n1583,n1584,n1585);
xor (n1584,n1581,n1582);
or (n1585,n1586,n1589);
and (n1586,n1587,n1588);
xor (n1587,n1547,n1548);
and (n1588,n152,n47);
and (n1589,n1590,n1591);
xor (n1590,n1587,n1588);
and (n1591,n1592,n1593);
xor (n1592,n1553,n1554);
and (n1593,n101,n47);
and (n1594,n53,n46);
or (n1595,n1596,n1599);
and (n1596,n1597,n1598);
xor (n1597,n1560,n1561);
and (n1598,n62,n46);
and (n1599,n1600,n1601);
xor (n1600,n1597,n1598);
or (n1601,n1602,n1605);
and (n1602,n1603,n1604);
xor (n1603,n1566,n1567);
and (n1604,n89,n46);
and (n1605,n1606,n1607);
xor (n1606,n1603,n1604);
or (n1607,n1608,n1611);
and (n1608,n1609,n1610);
xor (n1609,n1572,n1573);
and (n1610,n83,n46);
and (n1611,n1612,n1613);
xor (n1612,n1609,n1610);
or (n1613,n1614,n1617);
and (n1614,n1615,n1616);
xor (n1615,n1578,n1579);
and (n1616,n167,n46);
and (n1617,n1618,n1619);
xor (n1618,n1615,n1616);
or (n1619,n1620,n1623);
and (n1620,n1621,n1622);
xor (n1621,n1584,n1585);
and (n1622,n152,n46);
and (n1623,n1624,n1625);
xor (n1624,n1621,n1622);
and (n1625,n1626,n534);
xor (n1626,n1590,n1591);
and (n1627,n62,n54);
or (n1628,n1629,n1632);
and (n1629,n1630,n1631);
xor (n1630,n1600,n1601);
and (n1631,n89,n54);
and (n1632,n1633,n1634);
xor (n1633,n1630,n1631);
or (n1634,n1635,n1638);
and (n1635,n1636,n1637);
xor (n1636,n1606,n1607);
and (n1637,n83,n54);
and (n1638,n1639,n1640);
xor (n1639,n1636,n1637);
or (n1640,n1641,n1644);
and (n1641,n1642,n1643);
xor (n1642,n1612,n1613);
and (n1643,n167,n54);
and (n1644,n1645,n1646);
xor (n1645,n1642,n1643);
or (n1646,n1647,n1650);
and (n1647,n1648,n1649);
xor (n1648,n1618,n1619);
and (n1649,n152,n54);
and (n1650,n1651,n1652);
xor (n1651,n1648,n1649);
and (n1652,n1653,n1654);
xor (n1653,n1624,n1625);
and (n1654,n101,n54);
and (n1655,n89,n74);
or (n1656,n1657,n1660);
and (n1657,n1658,n1659);
xor (n1658,n1633,n1634);
and (n1659,n83,n74);
and (n1660,n1661,n1662);
xor (n1661,n1658,n1659);
or (n1662,n1663,n1666);
and (n1663,n1664,n1665);
xor (n1664,n1639,n1640);
and (n1665,n167,n74);
and (n1666,n1667,n1668);
xor (n1667,n1664,n1665);
or (n1668,n1669,n1672);
and (n1669,n1670,n1671);
xor (n1670,n1645,n1646);
and (n1671,n152,n74);
and (n1672,n1673,n1674);
xor (n1673,n1670,n1671);
and (n1674,n1675,n1676);
xor (n1675,n1651,n1652);
not (n1676,n251);
and (n1677,n83,n79);
or (n1678,n1679,n1682);
and (n1679,n1680,n1681);
xor (n1680,n1661,n1662);
and (n1681,n167,n79);
and (n1682,n1683,n1684);
xor (n1683,n1680,n1681);
or (n1684,n1685,n1688);
and (n1685,n1686,n1687);
xor (n1686,n1667,n1668);
and (n1687,n152,n79);
and (n1688,n1689,n1690);
xor (n1689,n1686,n1687);
and (n1690,n1691,n1692);
xor (n1691,n1673,n1674);
and (n1692,n101,n79);
and (n1693,n167,n158);
or (n1694,n1695,n1698);
and (n1695,n1696,n1697);
xor (n1696,n1683,n1684);
and (n1697,n152,n158);
and (n1698,n1699,n1700);
xor (n1699,n1696,n1697);
and (n1700,n1701,n1702);
xor (n1701,n1689,n1690);
not (n1702,n274);
and (n1703,n1704,n1705);
xor (n1704,n1699,n1700);
and (n1705,n101,n98);
and (n1706,n101,n99);
endmodule
