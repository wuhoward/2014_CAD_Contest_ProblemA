module top (out,n20,n25,n26,n27,n29,n30,n41,n44,n47
        ,n50,n53,n56,n59,n62,n65,n68,n71,n74,n76
        ,n79,n96,n101,n104,n107,n110,n113,n116,n118,n120
        ,n129,n142,n147,n150,n153,n156,n169,n205,n210,n213
        ,n216,n219,n222,n225,n228,n231,n234,n250,n685,n698);
output out;
input n20;
input n25;
input n26;
input n27;
input n29;
input n30;
input n41;
input n44;
input n47;
input n50;
input n53;
input n56;
input n59;
input n62;
input n65;
input n68;
input n71;
input n74;
input n76;
input n79;
input n96;
input n101;
input n104;
input n107;
input n110;
input n113;
input n116;
input n118;
input n120;
input n129;
input n142;
input n147;
input n150;
input n153;
input n156;
input n169;
input n205;
input n210;
input n213;
input n216;
input n219;
input n222;
input n225;
input n228;
input n231;
input n234;
input n250;
input n685;
input n698;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n21;
wire n22;
wire n23;
wire n24;
wire n28;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n42;
wire n43;
wire n45;
wire n46;
wire n48;
wire n49;
wire n51;
wire n52;
wire n54;
wire n55;
wire n57;
wire n58;
wire n60;
wire n61;
wire n63;
wire n64;
wire n66;
wire n67;
wire n69;
wire n70;
wire n72;
wire n73;
wire n75;
wire n77;
wire n78;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n97;
wire n98;
wire n99;
wire n100;
wire n102;
wire n103;
wire n105;
wire n106;
wire n108;
wire n109;
wire n111;
wire n112;
wire n114;
wire n115;
wire n117;
wire n119;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n143;
wire n144;
wire n145;
wire n146;
wire n148;
wire n149;
wire n151;
wire n152;
wire n154;
wire n155;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n206;
wire n207;
wire n208;
wire n209;
wire n211;
wire n212;
wire n214;
wire n215;
wire n217;
wire n218;
wire n220;
wire n221;
wire n223;
wire n224;
wire n226;
wire n227;
wire n229;
wire n230;
wire n232;
wire n233;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
xor (out,n0,n1630);
nand (n0,n1,n1629);
or (n1,n2,n840);
not (n2,n3);
and (n3,n4,n839);
or (n4,n5,n755);
xor (n5,n6,n671);
xor (n6,n7,n537);
xor (n7,n8,n403);
xor (n8,n9,n256);
xor (n9,n10,n190);
xor (n10,n11,n135);
nand (n11,n12,n123);
or (n12,n13,n92);
or (n13,n14,n85);
nor (n14,n15,n83);
and (n15,n16,n80);
not (n16,n17);
wire s0n17,s1n17,notn17;
or (n17,s0n17,s1n17);
not(notn17,n77);
and (s0n17,notn17,n18);
and (s1n17,n77,n37);
wire s0n18,s1n18,notn18;
or (n18,s0n18,s1n18);
not(notn18,n21);
and (s0n18,notn18,1'b0);
and (s1n18,n21,n20);
or (n21,n22,n33);
or (n22,n23,n31);
nor (n23,n24,n26,n27,n28,n30);
not (n24,n25);
not (n28,n29);
nor (n31,n25,n32,n27,n28,n30);
not (n32,n26);
or (n33,n34,n36);
and (n34,n24,n26,n27,n28,n35);
not (n35,n30);
nor (n36,n24,n32,n27,n28,n30);
xor (n37,n38,n39);
not (n38,n20);
and (n39,n40,n42);
not (n40,n41);
and (n42,n43,n45);
not (n43,n44);
and (n45,n46,n48);
not (n46,n47);
and (n48,n49,n51);
not (n49,n50);
and (n51,n52,n54);
not (n52,n53);
and (n54,n55,n57);
not (n55,n56);
and (n57,n58,n60);
not (n58,n59);
and (n60,n61,n63);
not (n61,n62);
and (n63,n64,n66);
not (n64,n65);
and (n66,n67,n69);
not (n67,n68);
and (n69,n70,n72);
not (n70,n71);
and (n72,n73,n75);
not (n73,n74);
not (n75,n76);
and (n77,n78,n79);
or (n78,n23,n34);
wire s0n80,s1n80,notn80;
or (n80,s0n80,s1n80);
not(notn80,n77);
and (s0n80,notn80,n81);
and (s1n80,n77,n82);
wire s0n81,s1n81,notn81;
or (n81,s0n81,s1n81);
not(notn81,n21);
and (s0n81,notn81,1'b0);
and (s1n81,n21,n41);
xor (n82,n40,n42);
and (n83,n84,n17);
not (n84,n80);
nor (n85,n86,n90);
and (n86,n80,n87);
wire s0n87,s1n87,notn87;
or (n87,s0n87,s1n87);
not(notn87,n77);
and (s0n87,notn87,n88);
and (s1n87,n77,n89);
wire s0n88,s1n88,notn88;
or (n88,s0n88,s1n88);
not(notn88,n21);
and (s0n88,notn88,1'b0);
and (s1n88,n21,n44);
xor (n89,n43,n45);
and (n90,n84,n91);
not (n91,n87);
nor (n92,n93,n121);
and (n93,n16,n94);
wire s0n94,s1n94,notn94;
or (n94,s0n94,s1n94);
not(notn94,n119);
and (s0n94,notn94,n95);
and (s1n94,n119,n97);
wire s0n95,s1n95,notn95;
or (n95,s0n95,s1n95);
not(notn95,n21);
and (s0n95,notn95,1'b0);
and (s1n95,n21,n96);
xor (n97,n98,n99);
not (n98,n96);
and (n99,n100,n102);
not (n100,n101);
and (n102,n103,n105);
not (n103,n104);
and (n105,n106,n108);
not (n106,n107);
and (n108,n109,n111);
not (n109,n110);
and (n111,n112,n114);
not (n112,n113);
and (n114,n115,n117);
not (n115,n116);
not (n117,n118);
and (n119,n78,n120);
and (n121,n17,n122);
not (n122,n94);
or (n123,n124,n125);
not (n124,n85);
nor (n125,n126,n133);
and (n126,n16,n127);
wire s0n127,s1n127,notn127;
or (n127,s0n127,s1n127);
not(notn127,n119);
and (s0n127,notn127,n128);
and (s1n127,n119,n130);
wire s0n128,s1n128,notn128;
or (n128,s0n128,s1n128);
not(notn128,n21);
and (s0n128,notn128,1'b0);
and (s1n128,n21,n129);
xor (n130,n131,n132);
not (n131,n129);
and (n132,n98,n99);
and (n133,n17,n134);
not (n134,n127);
nand (n135,n136,n181);
or (n136,n137,n174);
or (n137,n138,n164);
nor (n138,n139,n161);
and (n139,n140,n158);
wire s0n140,s1n140,notn140;
or (n140,s0n140,s1n140);
not(notn140,n77);
and (s0n140,notn140,n141);
and (s1n140,n77,n143);
wire s0n141,s1n141,notn141;
or (n141,s0n141,s1n141);
not(notn141,n21);
and (s0n141,notn141,1'b0);
and (s1n141,n21,n142);
xor (n143,n144,n145);
not (n144,n142);
and (n145,n146,n148);
not (n146,n147);
and (n148,n149,n151);
not (n149,n150);
and (n151,n152,n154);
not (n152,n153);
and (n154,n155,n157);
not (n155,n156);
and (n157,n38,n39);
wire s0n158,s1n158,notn158;
or (n158,s0n158,s1n158);
not(notn158,n77);
and (s0n158,notn158,n159);
and (s1n158,n77,n160);
wire s0n159,s1n159,notn159;
or (n159,s0n159,s1n159);
not(notn159,n21);
and (s0n159,notn159,1'b0);
and (s1n159,n21,n147);
xor (n160,n146,n148);
and (n161,n162,n163);
not (n162,n140);
not (n163,n158);
nor (n164,n165,n173);
and (n165,n140,n166);
not (n166,n167);
wire s0n167,s1n167,notn167;
or (n167,s0n167,s1n167);
not(notn167,n77);
and (s0n167,notn167,n168);
and (s1n167,n77,n170);
wire s0n168,s1n168,notn168;
or (n168,s0n168,s1n168);
not(notn168,n21);
and (s0n168,notn168,1'b0);
and (s1n168,n21,n169);
xor (n170,n171,n172);
not (n171,n169);
and (n172,n144,n145);
and (n173,n162,n167);
nor (n174,n175,n179);
and (n175,n176,n166);
wire s0n176,s1n176,notn176;
or (n176,s0n176,s1n176);
not(notn176,n119);
and (s0n176,notn176,n177);
and (s1n176,n119,n178);
wire s0n177,s1n177,notn177;
or (n177,s0n177,s1n177);
not(notn177,n21);
and (s0n177,notn177,1'b0);
and (s1n177,n21,n116);
xor (n178,n115,n117);
and (n179,n180,n167);
not (n180,n176);
or (n181,n182,n183);
not (n182,n138);
nor (n183,n184,n188);
and (n184,n185,n166);
wire s0n185,s1n185,notn185;
or (n185,s0n185,s1n185);
not(notn185,n119);
and (s0n185,notn185,n186);
and (s1n185,n119,n187);
wire s0n186,s1n186,notn186;
or (n186,s0n186,s1n186);
not(notn186,n21);
and (s0n186,notn186,1'b0);
and (s1n186,n21,n113);
xor (n187,n112,n114);
and (n188,n189,n167);
not (n189,n185);
and (n190,n191,n199);
nor (n191,n192,n166);
nor (n192,n193,n197);
and (n193,n194,n163);
not (n194,n195);
and (n195,n196,n140);
wire s0n196,s1n196,notn196;
or (n196,s0n196,s1n196);
not(notn196,n21);
and (s0n196,notn196,1'b0);
and (s1n196,n21,n118);
and (n197,n162,n198);
not (n198,n196);
nand (n199,n200,n245);
or (n200,n201,n242);
nor (n201,n202,n240);
and (n202,n203,n236);
wire s0n203,s1n203,notn203;
or (n203,s0n203,s1n203);
not(notn203,n119);
and (s0n203,notn203,n204);
and (s1n203,n119,n206);
wire s0n204,s1n204,notn204;
or (n204,s0n204,s1n204);
not(notn204,n21);
and (s0n204,notn204,1'b0);
and (s1n204,n21,n205);
xor (n206,n207,n208);
not (n207,n205);
and (n208,n209,n211);
not (n209,n210);
and (n211,n212,n214);
not (n212,n213);
and (n214,n215,n217);
not (n215,n216);
and (n217,n218,n220);
not (n218,n219);
and (n220,n221,n223);
not (n221,n222);
and (n223,n224,n226);
not (n224,n225);
and (n226,n227,n229);
not (n227,n228);
and (n229,n230,n232);
not (n230,n231);
and (n232,n233,n235);
not (n233,n234);
and (n235,n131,n132);
not (n236,n237);
wire s0n237,s1n237,notn237;
or (n237,s0n237,s1n237);
not(notn237,n77);
and (s0n237,notn237,n238);
and (s1n237,n77,n239);
wire s0n238,s1n238,notn238;
or (n238,s0n238,s1n238);
not(notn238,n21);
and (s0n238,notn238,1'b0);
and (s1n238,n21,n74);
xor (n239,n73,n75);
and (n240,n241,n237);
not (n241,n203);
nand (n242,n237,n243);
not (n243,n244);
wire s0n244,s1n244,notn244;
or (n244,s0n244,s1n244);
not(notn244,n21);
and (s0n244,notn244,1'b0);
and (s1n244,n21,n76);
or (n245,n246,n243);
nor (n246,n247,n254);
and (n247,n248,n236);
wire s0n248,s1n248,notn248;
or (n248,s0n248,s1n248);
not(notn248,n119);
and (s0n248,notn248,n249);
and (s1n248,n119,n251);
wire s0n249,s1n249,notn249;
or (n249,s0n249,s1n249);
not(notn249,n21);
and (s0n249,notn249,1'b0);
and (s1n249,n21,n250);
xor (n251,n252,n253);
not (n252,n250);
and (n253,n207,n208);
and (n254,n255,n237);
not (n255,n248);
or (n256,n257,n402);
and (n257,n258,n311);
xor (n258,n259,n260);
xor (n259,n191,n199);
or (n260,n261,n310);
and (n261,n262,n274);
xor (n262,n263,n264);
nor (n263,n182,n198);
nand (n264,n265,n273);
or (n265,n266,n242);
nor (n266,n267,n271);
and (n267,n268,n236);
wire s0n268,s1n268,notn268;
or (n268,s0n268,s1n268);
not(notn268,n119);
and (s0n268,notn268,n269);
and (s1n268,n119,n270);
wire s0n269,s1n269,notn269;
or (n269,s0n269,s1n269);
not(notn269,n21);
and (s0n269,notn269,1'b0);
and (s1n269,n21,n210);
xor (n270,n209,n211);
and (n271,n272,n237);
not (n272,n268);
or (n273,n201,n243);
nand (n274,n275,n298);
or (n275,n276,n287);
nor (n276,n277,n285);
and (n277,n278,n281);
wire s0n278,s1n278,notn278;
or (n278,s0n278,s1n278);
not(notn278,n119);
and (s0n278,notn278,n279);
and (s1n278,n119,n280);
wire s0n279,s1n279,notn279;
or (n279,s0n279,s1n279);
not(notn279,n21);
and (s0n279,notn279,1'b0);
and (s1n279,n21,n225);
xor (n280,n224,n226);
not (n281,n282);
wire s0n282,s1n282,notn282;
or (n282,s0n282,s1n282);
not(notn282,n77);
and (s0n282,notn282,n283);
and (s1n282,n77,n284);
wire s0n283,s1n283,notn283;
or (n283,s0n283,s1n283);
not(notn283,n21);
and (s0n283,notn283,1'b0);
and (s1n283,n21,n56);
xor (n284,n55,n57);
and (n285,n286,n282);
not (n286,n278);
or (n287,n288,n295);
and (n288,n289,n292);
wire s0n289,s1n289,notn289;
or (n289,s0n289,s1n289);
not(notn289,n77);
and (s0n289,notn289,n290);
and (s1n289,n77,n291);
wire s0n290,s1n290,notn290;
or (n290,s0n290,s1n290);
not(notn290,n21);
and (s0n290,notn290,1'b0);
and (s1n290,n21,n62);
xor (n291,n61,n63);
wire s0n292,s1n292,notn292;
or (n292,s0n292,s1n292);
not(notn292,n77);
and (s0n292,notn292,n293);
and (s1n292,n77,n294);
wire s0n293,s1n293,notn293;
or (n293,s0n293,s1n293);
not(notn293,n21);
and (s0n293,notn293,1'b0);
and (s1n293,n21,n59);
xor (n294,n58,n60);
and (n295,n296,n297);
not (n296,n289);
not (n297,n292);
or (n298,n299,n303);
nand (n299,n287,n300);
nor (n300,n301,n302);
and (n301,n282,n292);
and (n302,n281,n297);
nor (n303,n304,n308);
and (n304,n305,n281);
wire s0n305,s1n305,notn305;
or (n305,s0n305,s1n305);
not(notn305,n119);
and (s0n305,notn305,n306);
and (s1n305,n119,n307);
wire s0n306,s1n306,notn306;
or (n306,s0n306,s1n306);
not(notn306,n21);
and (s0n306,notn306,1'b0);
and (s1n306,n21,n228);
xor (n307,n227,n229);
and (n308,n309,n282);
not (n309,n305);
and (n310,n263,n264);
or (n311,n312,n401);
and (n312,n313,n369);
xor (n313,n314,n348);
nand (n314,n315,n339);
or (n315,n316,n332);
not (n316,n317);
nor (n317,n318,n324);
nand (n318,n319,n323);
or (n319,n16,n320);
wire s0n320,s1n320,notn320;
or (n320,s0n320,s1n320);
not(notn320,n77);
and (s0n320,notn320,n321);
and (s1n320,n77,n322);
wire s0n321,s1n321,notn321;
or (n321,s0n321,s1n321);
not(notn321,n21);
and (s0n321,notn321,1'b0);
and (s1n321,n21,n156);
xor (n322,n155,n157);
nand (n323,n16,n320);
nor (n324,n325,n330);
and (n325,n326,n320);
not (n326,n327);
wire s0n327,s1n327,notn327;
or (n327,s0n327,s1n327);
not(notn327,n77);
and (s0n327,notn327,n328);
and (s1n327,n77,n329);
wire s0n328,s1n328,notn328;
or (n328,s0n328,s1n328);
not(notn328,n21);
and (s0n328,notn328,1'b0);
and (s1n328,n21,n153);
xor (n329,n152,n154);
and (n330,n331,n327);
not (n331,n320);
nor (n332,n333,n337);
and (n333,n334,n326);
wire s0n334,s1n334,notn334;
or (n334,s0n334,s1n334);
not(notn334,n119);
and (s0n334,notn334,n335);
and (s1n334,n119,n336);
wire s0n335,s1n335,notn335;
or (n335,s0n335,s1n335);
not(notn335,n21);
and (s0n335,notn335,1'b0);
and (s1n335,n21,n110);
xor (n336,n109,n111);
and (n337,n338,n327);
not (n338,n334);
or (n339,n340,n347);
nor (n340,n341,n345);
and (n341,n326,n342);
wire s0n342,s1n342,notn342;
or (n342,s0n342,s1n342);
not(notn342,n119);
and (s0n342,notn342,n343);
and (s1n342,n119,n344);
wire s0n343,s1n343,notn343;
or (n343,s0n343,s1n343);
not(notn343,n21);
and (s0n343,notn343,1'b0);
and (s1n343,n21,n107);
xor (n344,n106,n108);
and (n345,n346,n327);
not (n346,n342);
not (n347,n318);
nand (n348,n349,n365);
or (n349,n350,n362);
not (n350,n351);
and (n351,n352,n359);
nor (n352,n353,n358);
and (n353,n327,n354);
not (n354,n355);
wire s0n355,s1n355,notn355;
or (n355,s0n355,s1n355);
not(notn355,n77);
and (s0n355,notn355,n356);
and (s1n355,n77,n357);
wire s0n356,s1n356,notn356;
or (n356,s0n356,s1n356);
not(notn356,n21);
and (s0n356,notn356,1'b0);
and (s1n356,n21,n150);
xor (n357,n149,n151);
and (n358,n326,n355);
nand (n359,n360,n361);
or (n360,n354,n158);
or (n361,n163,n355);
nor (n362,n363,n364);
and (n363,n176,n163);
and (n364,n180,n158);
or (n365,n366,n352);
nor (n366,n367,n368);
and (n367,n185,n163);
and (n368,n189,n158);
nand (n369,n370,n393);
or (n370,n371,n386);
nand (n371,n372,n379);
nor (n372,n373,n377);
and (n373,n236,n374);
wire s0n374,s1n374,notn374;
or (n374,s0n374,s1n374);
not(notn374,n77);
and (s0n374,notn374,n375);
and (s1n374,n77,n376);
wire s0n375,s1n375,notn375;
or (n375,s0n375,s1n375);
not(notn375,n21);
and (s0n375,notn375,1'b0);
and (s1n375,n21,n71);
xor (n376,n70,n72);
and (n377,n237,n378);
not (n378,n374);
nand (n379,n380,n385);
or (n380,n381,n374);
not (n381,n382);
wire s0n382,s1n382,notn382;
or (n382,s0n382,s1n382);
not(notn382,n77);
and (s0n382,notn382,n383);
and (s1n382,n77,n384);
wire s0n383,s1n383,notn383;
or (n383,s0n383,s1n383);
not(notn383,n21);
and (s0n383,notn383,1'b0);
and (s1n383,n21,n68);
xor (n384,n67,n69);
nand (n385,n381,n374);
nor (n386,n387,n391);
and (n387,n381,n388);
wire s0n388,s1n388,notn388;
or (n388,s0n388,s1n388);
not(notn388,n119);
and (s0n388,notn388,n389);
and (s1n388,n119,n390);
wire s0n389,s1n389,notn389;
or (n389,s0n389,s1n389);
not(notn389,n21);
and (s0n389,notn389,1'b0);
and (s1n389,n21,n216);
xor (n390,n215,n217);
and (n391,n392,n382);
not (n392,n388);
or (n393,n372,n394);
nor (n394,n395,n399);
and (n395,n381,n396);
wire s0n396,s1n396,notn396;
or (n396,s0n396,s1n396);
not(notn396,n119);
and (s0n396,notn396,n397);
and (s1n396,n119,n398);
wire s0n397,s1n397,notn397;
or (n397,s0n397,s1n397);
not(notn397,n21);
and (s0n397,notn397,1'b0);
and (s1n397,n21,n213);
xor (n398,n212,n214);
and (n399,n400,n382);
not (n400,n396);
and (n401,n314,n348);
and (n402,n259,n260);
xor (n403,n404,n499);
xor (n404,n405,n435);
or (n405,n406,n434);
and (n406,n407,n428);
xor (n407,n408,n418);
nand (n408,n409,n410);
or (n409,n299,n276);
or (n410,n287,n411);
nor (n411,n412,n416);
and (n412,n413,n281);
wire s0n413,s1n413,notn413;
or (n413,s0n413,s1n413);
not(notn413,n119);
and (s0n413,notn413,n414);
and (s1n413,n119,n415);
wire s0n414,s1n414,notn414;
or (n414,s0n414,s1n414);
not(notn414,n21);
and (s0n414,notn414,1'b0);
and (s1n414,n21,n222);
xor (n415,n221,n223);
and (n416,n417,n282);
not (n417,n413);
nand (n418,n419,n420);
or (n419,n316,n340);
or (n420,n347,n421);
nor (n421,n422,n426);
and (n422,n423,n326);
wire s0n423,s1n423,notn423;
or (n423,s0n423,s1n423);
not(notn423,n119);
and (s0n423,notn423,n424);
and (s1n423,n119,n425);
wire s0n424,s1n424,notn424;
or (n424,s0n424,s1n424);
not(notn424,n21);
and (s0n424,notn424,1'b0);
and (s1n424,n21,n104);
xor (n425,n103,n105);
and (n426,n427,n327);
not (n427,n423);
nand (n428,n429,n430);
or (n429,n350,n366);
or (n430,n431,n352);
nor (n431,n432,n433);
and (n432,n334,n163);
and (n433,n338,n158);
and (n434,n408,n418);
or (n435,n436,n498);
and (n436,n437,n473);
xor (n437,n438,n444);
nand (n438,n439,n440);
or (n439,n371,n394);
or (n440,n441,n372);
nor (n441,n442,n443);
and (n442,n268,n381);
and (n443,n272,n382);
nand (n444,n445,n469);
or (n445,n446,n462);
nand (n446,n447,n458);
nor (n447,n448,n455);
and (n448,n449,n452);
wire s0n449,s1n449,notn449;
or (n449,s0n449,s1n449);
not(notn449,n77);
and (s0n449,notn449,n450);
and (s1n449,n77,n451);
wire s0n450,s1n450,notn450;
or (n450,s0n450,s1n450);
not(notn450,n21);
and (s0n450,notn450,1'b0);
and (s1n450,n21,n53);
xor (n451,n52,n54);
wire s0n452,s1n452,notn452;
or (n452,s0n452,s1n452);
not(notn452,n77);
and (s0n452,notn452,n453);
and (s1n452,n77,n454);
wire s0n453,s1n453,notn453;
or (n453,s0n453,s1n453);
not(notn453,n21);
and (s0n453,notn453,1'b0);
and (s1n453,n21,n50);
xor (n454,n49,n51);
and (n455,n456,n457);
not (n456,n449);
not (n457,n452);
not (n458,n459);
nor (n459,n460,n461);
and (n460,n282,n449);
and (n461,n281,n456);
nor (n462,n463,n467);
and (n463,n457,n464);
wire s0n464,s1n464,notn464;
or (n464,s0n464,s1n464);
not(notn464,n119);
and (s0n464,notn464,n465);
and (s1n464,n119,n466);
wire s0n465,s1n465,notn465;
or (n465,s0n465,s1n465);
not(notn465,n21);
and (s0n465,notn465,1'b0);
and (s1n465,n21,n231);
xor (n466,n230,n232);
and (n467,n452,n468);
not (n468,n464);
or (n469,n470,n458);
nor (n470,n471,n472);
and (n471,n457,n305);
and (n472,n452,n309);
nand (n473,n474,n494);
or (n474,n475,n487);
nand (n475,n476,n483);
not (n476,n477);
nand (n477,n478,n482);
or (n478,n381,n479);
wire s0n479,s1n479,notn479;
or (n479,s0n479,s1n479);
not(notn479,n77);
and (s0n479,notn479,n480);
and (s1n479,n77,n481);
wire s0n480,s1n480,notn480;
or (n480,s0n480,s1n480);
not(notn480,n21);
and (s0n480,notn480,1'b0);
and (s1n480,n21,n65);
xor (n481,n64,n66);
nand (n482,n479,n381);
nor (n483,n484,n486);
and (n484,n296,n485);
not (n485,n479);
and (n486,n289,n479);
nor (n487,n488,n492);
and (n488,n489,n296);
wire s0n489,s1n489,notn489;
or (n489,s0n489,s1n489);
not(notn489,n119);
and (s0n489,notn489,n490);
and (s1n489,n119,n491);
wire s0n490,s1n490,notn490;
or (n490,s0n490,s1n490);
not(notn490,n21);
and (s0n490,notn490,1'b0);
and (s1n490,n21,n219);
xor (n491,n218,n220);
and (n492,n493,n289);
not (n493,n489);
or (n494,n476,n495);
nor (n495,n496,n497);
and (n496,n388,n296);
and (n497,n392,n289);
and (n498,n438,n444);
xor (n499,n500,n513);
xor (n500,n501,n507);
nand (n501,n502,n503);
or (n502,n446,n470);
or (n503,n504,n458);
nor (n504,n505,n506);
and (n505,n457,n278);
and (n506,n452,n286);
nand (n507,n508,n509);
or (n508,n475,n495);
or (n509,n476,n510);
nor (n510,n511,n512);
and (n511,n396,n296);
and (n512,n400,n289);
nand (n513,n514,n533);
or (n514,n515,n526);
nand (n515,n516,n523);
or (n516,n517,n521);
and (n517,n518,n452);
wire s0n518,s1n518,notn518;
or (n518,s0n518,s1n518);
not(notn518,n77);
and (s0n518,notn518,n519);
and (s1n518,n77,n520);
wire s0n519,s1n519,notn519;
or (n519,s0n519,s1n519);
not(notn519,n21);
and (s0n519,notn519,1'b0);
and (s1n519,n21,n47);
xor (n520,n46,n48);
and (n521,n522,n457);
not (n522,n518);
nand (n523,n524,n525);
or (n524,n522,n87);
or (n525,n91,n518);
nor (n526,n527,n531);
and (n527,n91,n528);
wire s0n528,s1n528,notn528;
or (n528,s0n528,s1n528);
not(notn528,n119);
and (s0n528,notn528,n529);
and (s1n528,n119,n530);
wire s0n529,s1n529,notn529;
or (n529,s0n529,s1n529);
not(notn529,n21);
and (s0n529,notn529,1'b0);
and (s1n529,n21,n234);
xor (n530,n233,n235);
and (n531,n87,n532);
not (n532,n528);
or (n533,n516,n534);
nor (n534,n535,n536);
and (n535,n91,n464);
and (n536,n87,n468);
or (n537,n538,n670);
and (n538,n539,n597);
xor (n539,n540,n590);
or (n540,n541,n589);
and (n541,n542,n588);
xor (n542,n543,n571);
or (n543,n544,n570);
and (n544,n545,n561);
xor (n545,n546,n552);
nand (n546,n547,n551);
or (n547,n371,n548);
nor (n548,n549,n550);
and (n549,n381,n489);
and (n550,n493,n382);
or (n551,n372,n386);
nand (n552,n553,n557);
or (n553,n446,n554);
nor (n554,n555,n556);
and (n555,n457,n127);
and (n556,n452,n134);
or (n557,n558,n458);
nor (n558,n559,n560);
and (n559,n457,n528);
and (n560,n452,n532);
nand (n561,n562,n566);
or (n562,n563,n475);
nor (n563,n564,n565);
and (n564,n278,n296);
and (n565,n286,n289);
or (n566,n476,n567);
nor (n567,n568,n569);
and (n568,n413,n296);
and (n569,n417,n289);
and (n570,n546,n552);
xor (n571,n572,n579);
xor (n572,n573,n576);
nand (n573,n574,n575);
or (n574,n446,n558);
or (n575,n462,n458);
nand (n576,n577,n578);
or (n577,n475,n567);
or (n578,n476,n487);
nand (n579,n580,n584);
or (n580,n515,n581);
nor (n581,n582,n583);
and (n582,n91,n94);
and (n583,n87,n122);
or (n584,n516,n585);
nor (n585,n586,n587);
and (n586,n91,n127);
and (n587,n87,n134);
xor (n588,n262,n274);
and (n589,n543,n571);
xor (n590,n591,n596);
xor (n591,n592,n595);
or (n592,n593,n594);
and (n593,n572,n579);
and (n594,n573,n576);
xor (n595,n437,n473);
xor (n596,n407,n428);
or (n597,n598,n669);
and (n598,n599,n637);
xor (n599,n600,n601);
xor (n600,n313,n369);
or (n601,n602,n636);
and (n602,n603,n623);
xor (n603,n604,n614);
nand (n604,n605,n613);
or (n605,n515,n606);
nor (n606,n607,n611);
and (n607,n91,n608);
wire s0n608,s1n608,notn608;
or (n608,s0n608,s1n608);
not(notn608,n119);
and (s0n608,notn608,n609);
and (s1n608,n119,n610);
wire s0n609,s1n609,notn609;
or (n609,s0n609,s1n609);
not(notn609,n21);
and (s0n609,notn609,1'b0);
and (s1n609,n21,n101);
xor (n610,n100,n102);
and (n611,n87,n612);
not (n612,n608);
or (n613,n581,n516);
nand (n614,n615,n619);
or (n615,n13,n616);
nor (n616,n617,n618);
and (n617,n16,n342);
and (n618,n346,n17);
or (n619,n124,n620);
nor (n620,n621,n622);
and (n621,n16,n423);
and (n622,n17,n427);
xor (n623,n624,n630);
nor (n624,n625,n163);
nor (n625,n626,n629);
and (n626,n326,n627);
not (n627,n628);
and (n628,n196,n355);
and (n629,n354,n198);
nand (n630,n631,n635);
or (n631,n632,n242);
nor (n632,n633,n634);
and (n633,n396,n236);
and (n634,n400,n237);
or (n635,n266,n243);
and (n636,n604,n614);
xor (n637,n638,n646);
xor (n638,n639,n645);
nand (n639,n640,n641);
or (n640,n13,n620);
or (n641,n642,n124);
nor (n642,n643,n644);
and (n643,n16,n608);
and (n644,n17,n612);
and (n645,n624,n630);
or (n646,n647,n668);
and (n647,n648,n661);
xor (n648,n649,n655);
nand (n649,n650,n654);
or (n650,n299,n651);
nor (n651,n652,n653);
and (n652,n464,n281);
and (n653,n468,n282);
or (n654,n303,n287);
nand (n655,n656,n660);
or (n656,n316,n657);
nor (n657,n658,n659);
and (n658,n185,n326);
and (n659,n189,n327);
or (n660,n347,n332);
nand (n661,n662,n667);
or (n662,n663,n350);
not (n663,n664);
nand (n664,n665,n666);
or (n665,n163,n196);
or (n666,n158,n198);
or (n667,n362,n352);
and (n668,n649,n655);
and (n669,n600,n601);
and (n670,n540,n590);
xor (n671,n672,n746);
xor (n672,n673,n676);
or (n673,n674,n675);
and (n674,n591,n596);
and (n675,n592,n595);
xor (n676,n677,n730);
xor (n677,n678,n710);
xor (n678,n679,n704);
xor (n679,n680,n691);
nor (n680,n681,n198);
nor (n681,n682,n689);
and (n682,n166,n683);
wire s0n683,s1n683,notn683;
or (n683,s0n683,s1n683);
not(notn683,n77);
and (s0n683,notn683,n684);
and (s1n683,n77,n686);
wire s0n684,s1n684,notn684;
or (n684,s0n684,s1n684);
not(notn684,n21);
and (s0n684,notn684,1'b0);
and (s1n684,n21,n685);
xor (n686,n687,n688);
not (n687,n685);
and (n688,n171,n172);
and (n689,n167,n690);
not (n690,n683);
nand (n691,n692,n693);
or (n692,n246,n242);
or (n693,n694,n243);
nor (n694,n695,n702);
and (n695,n696,n236);
wire s0n696,s1n696,notn696;
or (n696,s0n696,s1n696);
not(notn696,n119);
and (s0n696,notn696,n697);
and (s1n696,n119,n699);
wire s0n697,s1n697,notn697;
or (n697,s0n697,s1n697);
not(notn697,n21);
and (s0n697,notn697,1'b0);
and (s1n697,n21,n698);
xor (n699,n700,n701);
not (n700,n698);
and (n701,n252,n253);
and (n702,n703,n237);
not (n703,n696);
nand (n704,n705,n706);
or (n705,n299,n411);
or (n706,n287,n707);
nor (n707,n708,n709);
and (n708,n489,n281);
and (n709,n493,n282);
xor (n710,n711,n724);
xor (n711,n712,n718);
nand (n712,n713,n714);
or (n713,n316,n421);
or (n714,n715,n347);
nor (n715,n716,n717);
and (n716,n326,n608);
and (n717,n327,n612);
nand (n718,n719,n720);
or (n719,n350,n431);
or (n720,n721,n352);
nor (n721,n722,n723);
and (n722,n163,n342);
and (n723,n158,n346);
nand (n724,n725,n726);
or (n725,n371,n441);
or (n726,n372,n727);
nor (n727,n728,n729);
and (n728,n203,n381);
and (n729,n241,n382);
or (n730,n731,n745);
and (n731,n732,n739);
xor (n732,n733,n736);
nand (n733,n734,n735);
or (n734,n515,n585);
or (n735,n516,n526);
nand (n736,n737,n738);
or (n737,n13,n642);
or (n738,n92,n124);
nand (n739,n740,n744);
or (n740,n137,n741);
nor (n741,n742,n743);
and (n742,n167,n198);
and (n743,n166,n196);
or (n744,n182,n174);
and (n745,n733,n736);
or (n746,n747,n754);
and (n747,n748,n753);
xor (n748,n749,n750);
xor (n749,n732,n739);
or (n750,n751,n752);
and (n751,n638,n646);
and (n752,n639,n645);
xor (n753,n258,n311);
and (n754,n749,n750);
or (n755,n756,n838);
and (n756,n757,n837);
xor (n757,n758,n759);
xor (n758,n748,n753);
or (n759,n760,n836);
and (n760,n761,n835);
xor (n761,n762,n828);
or (n762,n763,n827);
and (n763,n764,n805);
xor (n764,n765,n782);
or (n765,n766,n781);
and (n766,n767,n775);
xor (n767,n768,n769);
nor (n768,n352,n198);
nand (n769,n770,n774);
or (n770,n771,n242);
nor (n771,n772,n773);
and (n772,n388,n236);
and (n773,n392,n237);
or (n774,n632,n243);
nand (n775,n776,n780);
or (n776,n371,n777);
nor (n777,n778,n779);
and (n778,n381,n413);
and (n779,n417,n382);
or (n780,n372,n548);
and (n781,n768,n769);
or (n782,n783,n804);
and (n783,n784,n798);
xor (n784,n785,n791);
nand (n785,n786,n790);
or (n786,n475,n787);
nor (n787,n788,n789);
and (n788,n305,n296);
and (n789,n309,n289);
or (n790,n476,n563);
nand (n791,n792,n797);
or (n792,n793,n515);
not (n793,n794);
nand (n794,n795,n796);
or (n795,n427,n87);
or (n796,n91,n423);
or (n797,n606,n516);
nand (n798,n799,n803);
or (n799,n13,n800);
nor (n800,n801,n802);
and (n801,n334,n16);
and (n802,n338,n17);
or (n803,n616,n124);
and (n804,n785,n791);
or (n805,n806,n826);
and (n806,n807,n820);
xor (n807,n808,n814);
nand (n808,n809,n813);
or (n809,n316,n810);
nor (n810,n811,n812);
and (n811,n176,n326);
and (n812,n180,n327);
or (n813,n657,n347);
nand (n814,n815,n819);
or (n815,n299,n816);
nor (n816,n817,n818);
and (n817,n528,n281);
and (n818,n532,n282);
or (n819,n651,n287);
nand (n820,n821,n825);
or (n821,n446,n822);
nor (n822,n823,n824);
and (n823,n457,n94);
and (n824,n452,n122);
or (n825,n554,n458);
and (n826,n808,n814);
and (n827,n765,n782);
or (n828,n829,n834);
and (n829,n830,n833);
xor (n830,n831,n832);
xor (n831,n648,n661);
xor (n832,n545,n561);
xor (n833,n603,n623);
and (n834,n831,n832);
xor (n835,n542,n588);
and (n836,n762,n828);
xor (n837,n539,n597);
and (n838,n758,n759);
nand (n839,n5,n755);
not (n840,n841);
nor (n841,n842,n1618);
nor (n842,n843,n1601);
nand (n843,n844,n1550);
or (n844,n845,n1549);
and (n845,n846,n1139);
xor (n846,n847,n1078);
or (n847,n848,n1077);
and (n848,n849,n1026);
xor (n849,n850,n933);
xor (n850,n851,n902);
xor (n851,n852,n873);
xor (n852,n853,n864);
xor (n853,n854,n855);
nor (n854,n347,n198);
nand (n855,n856,n860);
or (n856,n857,n242);
nor (n857,n858,n859);
and (n858,n236,n413);
and (n859,n417,n237);
or (n860,n861,n243);
nor (n861,n862,n863);
and (n862,n489,n236);
and (n863,n493,n237);
nand (n864,n865,n869);
or (n865,n371,n866);
nor (n866,n867,n868);
and (n867,n381,n305);
and (n868,n309,n382);
or (n869,n372,n870);
nor (n870,n871,n872);
and (n871,n278,n381);
and (n872,n286,n382);
or (n873,n874,n901);
and (n874,n875,n891);
xor (n875,n876,n882);
nand (n876,n877,n881);
or (n877,n371,n878);
nor (n878,n879,n880);
and (n879,n381,n464);
and (n880,n468,n382);
or (n881,n372,n866);
nand (n882,n883,n887);
or (n883,n299,n884);
nor (n884,n885,n886);
and (n885,n608,n281);
and (n886,n612,n282);
or (n887,n287,n888);
nor (n888,n889,n890);
and (n889,n94,n281);
and (n890,n122,n282);
nand (n891,n892,n897);
or (n892,n893,n446);
not (n893,n894);
nand (n894,n895,n896);
or (n895,n452,n346);
or (n896,n457,n342);
or (n897,n898,n458);
nor (n898,n899,n900);
and (n899,n457,n423);
and (n900,n452,n427);
and (n901,n876,n882);
or (n902,n903,n932);
and (n903,n904,n923);
xor (n904,n905,n914);
nand (n905,n906,n910);
or (n906,n475,n907);
nor (n907,n908,n909);
and (n908,n127,n296);
and (n909,n134,n289);
or (n910,n911,n476);
nor (n911,n912,n913);
and (n912,n528,n296);
and (n913,n532,n289);
nand (n914,n915,n919);
or (n915,n515,n916);
nor (n916,n917,n918);
and (n917,n185,n91);
and (n918,n189,n87);
or (n919,n920,n516);
nor (n920,n921,n922);
and (n921,n334,n91);
and (n922,n338,n87);
nand (n923,n924,n928);
or (n924,n124,n925);
nor (n925,n926,n927);
and (n926,n176,n16);
and (n927,n180,n17);
or (n928,n13,n929);
nor (n929,n930,n931);
and (n930,n17,n198);
and (n931,n16,n196);
and (n932,n905,n914);
xor (n933,n934,n982);
xor (n934,n935,n962);
xor (n935,n936,n949);
xor (n936,n937,n943);
nand (n937,n938,n939);
or (n938,n515,n920);
or (n939,n940,n516);
nor (n940,n941,n942);
and (n941,n91,n342);
and (n942,n87,n346);
nand (n943,n944,n945);
or (n944,n13,n925);
or (n945,n946,n124);
nor (n946,n947,n948);
and (n947,n185,n16);
and (n948,n189,n17);
and (n949,n950,n956);
nand (n950,n951,n955);
or (n951,n952,n242);
nor (n952,n953,n954);
and (n953,n236,n278);
and (n954,n286,n237);
or (n955,n857,n243);
nor (n956,n957,n16);
nor (n957,n958,n961);
and (n958,n91,n959);
not (n959,n960);
and (n960,n196,n80);
and (n961,n84,n198);
xor (n962,n963,n976);
xor (n963,n964,n970);
nand (n964,n965,n966);
or (n965,n299,n888);
or (n966,n967,n287);
nor (n967,n968,n969);
and (n968,n127,n281);
and (n969,n134,n282);
nand (n970,n971,n972);
or (n971,n446,n898);
or (n972,n973,n458);
nor (n973,n974,n975);
and (n974,n457,n608);
and (n975,n452,n612);
nand (n976,n977,n981);
or (n977,n476,n978);
nor (n978,n979,n980);
and (n979,n464,n296);
and (n980,n468,n289);
or (n981,n475,n911);
or (n982,n983,n1025);
and (n983,n984,n1003);
xor (n984,n985,n986);
xor (n985,n950,n956);
or (n986,n987,n1002);
and (n987,n988,n996);
xor (n988,n989,n990);
nor (n989,n124,n198);
nand (n990,n991,n995);
or (n991,n992,n242);
nor (n992,n993,n994);
and (n993,n236,n305);
and (n994,n309,n237);
or (n995,n952,n243);
nand (n996,n997,n998);
or (n997,n372,n878);
or (n998,n371,n999);
nor (n999,n1000,n1001);
and (n1000,n528,n381);
and (n1001,n532,n382);
and (n1002,n989,n990);
or (n1003,n1004,n1024);
and (n1004,n1005,n1018);
xor (n1005,n1006,n1012);
nand (n1006,n1007,n1011);
or (n1007,n299,n1008);
nor (n1008,n1009,n1010);
and (n1009,n423,n281);
and (n1010,n427,n282);
or (n1011,n884,n287);
nand (n1012,n1013,n1014);
or (n1013,n458,n893);
or (n1014,n446,n1015);
nor (n1015,n1016,n1017);
and (n1016,n457,n334);
and (n1017,n452,n338);
nand (n1018,n1019,n1020);
or (n1019,n516,n916);
or (n1020,n515,n1021);
nor (n1021,n1022,n1023);
and (n1022,n176,n91);
and (n1023,n180,n87);
and (n1024,n1006,n1012);
and (n1025,n985,n986);
or (n1026,n1027,n1076);
and (n1027,n1028,n1031);
xor (n1028,n1029,n1030);
xor (n1029,n904,n923);
xor (n1030,n875,n891);
or (n1031,n1032,n1075);
and (n1032,n1033,n1053);
xor (n1033,n1034,n1040);
nand (n1034,n1035,n1039);
or (n1035,n475,n1036);
nor (n1036,n1037,n1038);
and (n1037,n94,n296);
and (n1038,n122,n289);
or (n1039,n476,n907);
and (n1040,n1041,n1047);
nand (n1041,n1042,n1046);
or (n1042,n1043,n242);
nor (n1043,n1044,n1045);
and (n1044,n464,n236);
and (n1045,n468,n237);
or (n1046,n992,n243);
nor (n1047,n1048,n91);
nor (n1048,n1049,n1052);
and (n1049,n457,n1050);
not (n1050,n1051);
and (n1051,n196,n518);
and (n1052,n522,n198);
or (n1053,n1054,n1074);
and (n1054,n1055,n1068);
xor (n1055,n1056,n1062);
nand (n1056,n1057,n1061);
or (n1057,n371,n1058);
nor (n1058,n1059,n1060);
and (n1059,n127,n381);
and (n1060,n134,n382);
or (n1061,n372,n999);
nand (n1062,n1063,n1067);
or (n1063,n299,n1064);
nor (n1064,n1065,n1066);
and (n1065,n342,n281);
and (n1066,n346,n282);
or (n1067,n1008,n287);
nand (n1068,n1069,n1073);
or (n1069,n446,n1070);
nor (n1070,n1071,n1072);
and (n1071,n185,n457);
and (n1072,n189,n452);
or (n1073,n1015,n458);
and (n1074,n1056,n1062);
and (n1075,n1034,n1040);
and (n1076,n1029,n1030);
and (n1077,n850,n933);
xor (n1078,n1079,n1102);
xor (n1079,n1080,n1099);
xor (n1080,n1081,n1088);
xor (n1081,n1082,n1085);
or (n1082,n1083,n1084);
and (n1083,n963,n976);
and (n1084,n964,n970);
or (n1085,n1086,n1087);
and (n1086,n936,n949);
and (n1087,n937,n943);
xor (n1088,n1089,n1096);
xor (n1089,n1090,n1093);
nand (n1090,n1091,n1092);
or (n1091,n446,n973);
or (n1092,n822,n458);
nand (n1093,n1094,n1095);
or (n1094,n475,n978);
or (n1095,n476,n787);
nand (n1096,n1097,n1098);
or (n1097,n516,n793);
or (n1098,n515,n940);
or (n1099,n1100,n1101);
and (n1100,n934,n982);
and (n1101,n935,n962);
xor (n1102,n1103,n1121);
xor (n1103,n1104,n1118);
xor (n1104,n1105,n1115);
xor (n1105,n1106,n1109);
nand (n1106,n1107,n1108);
or (n1107,n371,n870);
or (n1108,n372,n777);
nand (n1109,n1110,n1114);
or (n1110,n316,n1111);
nor (n1111,n1112,n1113);
and (n1112,n327,n198);
and (n1113,n326,n196);
or (n1114,n810,n347);
nand (n1115,n1116,n1117);
or (n1116,n816,n287);
or (n1117,n299,n967);
or (n1118,n1119,n1120);
and (n1119,n851,n902);
and (n1120,n852,n873);
xor (n1121,n1122,n1136);
xor (n1122,n1123,n1126);
nand (n1123,n1124,n1125);
or (n1124,n13,n946);
or (n1125,n800,n124);
xor (n1126,n1127,n1130);
nand (n1127,n1128,n1129);
or (n1128,n861,n242);
or (n1129,n771,n243);
nor (n1130,n1131,n326);
nor (n1131,n1132,n1135);
and (n1132,n16,n1133);
not (n1133,n1134);
and (n1134,n196,n320);
and (n1135,n331,n198);
or (n1136,n1137,n1138);
and (n1137,n853,n864);
and (n1138,n854,n855);
or (n1139,n1140,n1548);
and (n1140,n1141,n1172);
xor (n1141,n1142,n1171);
or (n1142,n1143,n1170);
and (n1143,n1144,n1169);
xor (n1144,n1145,n1168);
or (n1145,n1146,n1167);
and (n1146,n1147,n1150);
xor (n1147,n1148,n1149);
xor (n1148,n988,n996);
xor (n1149,n1005,n1018);
or (n1150,n1151,n1166);
and (n1151,n1152,n1165);
xor (n1152,n1153,n1159);
nand (n1153,n1154,n1158);
or (n1154,n515,n1155);
nor (n1155,n1156,n1157);
and (n1156,n87,n198);
and (n1157,n91,n196);
or (n1158,n1021,n516);
nand (n1159,n1160,n1164);
or (n1160,n475,n1161);
nor (n1161,n1162,n1163);
and (n1162,n608,n296);
and (n1163,n612,n289);
or (n1164,n1036,n476);
xor (n1165,n1041,n1047);
and (n1166,n1153,n1159);
and (n1167,n1148,n1149);
xor (n1168,n984,n1003);
xor (n1169,n1028,n1031);
and (n1170,n1145,n1168);
xor (n1171,n849,n1026);
nand (n1172,n1173,n1545,n1547);
or (n1173,n1174,n1540);
nand (n1174,n1175,n1529);
or (n1175,n1176,n1528);
and (n1176,n1177,n1298);
xor (n1177,n1178,n1283);
or (n1178,n1179,n1282);
and (n1179,n1180,n1248);
xor (n1180,n1181,n1203);
xor (n1181,n1182,n1197);
xor (n1182,n1183,n1190);
nand (n1183,n1184,n1189);
or (n1184,n299,n1185);
not (n1185,n1186);
nor (n1186,n1187,n1188);
and (n1187,n281,n338);
and (n1188,n334,n282);
or (n1189,n1064,n287);
nand (n1190,n1191,n1196);
or (n1191,n1192,n446);
not (n1192,n1193);
nand (n1193,n1194,n1195);
or (n1194,n180,n452);
or (n1195,n176,n457);
or (n1196,n1070,n458);
nand (n1197,n1198,n1202);
or (n1198,n475,n1199);
nor (n1199,n1200,n1201);
and (n1200,n423,n296);
and (n1201,n427,n289);
or (n1202,n476,n1161);
or (n1203,n1204,n1247);
and (n1204,n1205,n1227);
xor (n1205,n1206,n1212);
nand (n1206,n1207,n1211);
or (n1207,n475,n1208);
nor (n1208,n1209,n1210);
and (n1209,n342,n296);
and (n1210,n346,n289);
or (n1211,n1199,n476);
xor (n1212,n1213,n1219);
nor (n1213,n1214,n457);
nor (n1214,n1215,n1218);
and (n1215,n1216,n281);
not (n1216,n1217);
and (n1217,n196,n449);
and (n1218,n456,n198);
nand (n1219,n1220,n1223);
or (n1220,n242,n1221);
not (n1221,n1222);
xnor (n1222,n127,n236);
or (n1223,n1224,n243);
nor (n1224,n1225,n1226);
and (n1225,n236,n528);
and (n1226,n532,n237);
or (n1227,n1228,n1246);
and (n1228,n1229,n1237);
xor (n1229,n1230,n1231);
nor (n1230,n458,n198);
nand (n1231,n1232,n1233);
or (n1232,n243,n1221);
or (n1233,n1234,n242);
nor (n1234,n1235,n1236);
and (n1235,n236,n94);
and (n1236,n122,n237);
nand (n1237,n1238,n1242);
or (n1238,n299,n1239);
nor (n1239,n1240,n1241);
and (n1240,n176,n281);
and (n1241,n180,n282);
or (n1242,n1243,n287);
nor (n1243,n1244,n1245);
and (n1244,n185,n281);
and (n1245,n189,n282);
and (n1246,n1230,n1231);
and (n1247,n1206,n1212);
xor (n1248,n1249,n1263);
xor (n1249,n1250,n1251);
and (n1250,n1213,n1219);
xor (n1251,n1252,n1257);
xor (n1252,n1253,n1254);
nor (n1253,n516,n198);
nand (n1254,n1255,n1256);
or (n1255,n1224,n242);
or (n1256,n1043,n243);
nand (n1257,n1258,n1262);
or (n1258,n371,n1259);
nor (n1259,n1260,n1261);
and (n1260,n94,n381);
and (n1261,n122,n382);
or (n1262,n372,n1058);
or (n1263,n1264,n1281);
and (n1264,n1265,n1275);
xor (n1265,n1266,n1272);
nand (n1266,n1267,n1271);
or (n1267,n371,n1268);
nor (n1268,n1269,n1270);
and (n1269,n381,n608);
and (n1270,n612,n382);
or (n1271,n1259,n372);
nand (n1272,n1273,n1274);
or (n1273,n287,n1185);
or (n1274,n1243,n299);
nand (n1275,n1276,n1277);
or (n1276,n458,n1192);
or (n1277,n446,n1278);
nor (n1278,n1279,n1280);
and (n1279,n452,n198);
and (n1280,n457,n196);
and (n1281,n1266,n1272);
and (n1282,n1181,n1203);
xor (n1283,n1284,n1289);
xor (n1284,n1285,n1286);
xor (n1285,n1055,n1068);
or (n1286,n1287,n1288);
and (n1287,n1249,n1263);
and (n1288,n1250,n1251);
xor (n1289,n1290,n1297);
xor (n1290,n1291,n1294);
or (n1291,n1292,n1293);
and (n1292,n1252,n1257);
and (n1293,n1253,n1254);
or (n1294,n1295,n1296);
and (n1295,n1182,n1197);
and (n1296,n1183,n1190);
xor (n1297,n1152,n1165);
or (n1298,n1299,n1527);
and (n1299,n1300,n1337);
xor (n1300,n1301,n1336);
or (n1301,n1302,n1335);
and (n1302,n1303,n1334);
xor (n1303,n1304,n1333);
or (n1304,n1305,n1332);
and (n1305,n1306,n1319);
xor (n1306,n1307,n1313);
nand (n1307,n1308,n1312);
or (n1308,n371,n1309);
nor (n1309,n1310,n1311);
and (n1310,n423,n381);
and (n1311,n382,n427);
or (n1312,n1268,n372);
nand (n1313,n1314,n1318);
or (n1314,n475,n1315);
nor (n1315,n1316,n1317);
and (n1316,n334,n296);
and (n1317,n338,n289);
or (n1318,n1208,n476);
and (n1319,n1320,n1326);
nor (n1320,n1321,n281);
nor (n1321,n1322,n1325);
and (n1322,n1323,n296);
not (n1323,n1324);
and (n1324,n196,n292);
and (n1325,n297,n198);
nand (n1326,n1327,n1331);
or (n1327,n1328,n242);
nor (n1328,n1329,n1330);
and (n1329,n236,n608);
and (n1330,n612,n237);
or (n1331,n1234,n243);
and (n1332,n1307,n1313);
xor (n1333,n1265,n1275);
xor (n1334,n1205,n1227);
and (n1335,n1304,n1333);
xor (n1336,n1180,n1248);
nand (n1337,n1338,n1524,n1526);
or (n1338,n1339,n1397);
nand (n1339,n1340,n1392);
not (n1340,n1341);
nor (n1341,n1342,n1368);
xor (n1342,n1343,n1367);
xor (n1343,n1344,n1366);
or (n1344,n1345,n1365);
and (n1345,n1346,n1359);
xor (n1346,n1347,n1353);
nand (n1347,n1348,n1352);
or (n1348,n299,n1349);
nor (n1349,n1350,n1351);
and (n1350,n282,n198);
and (n1351,n281,n196);
or (n1352,n1239,n287);
nand (n1353,n1354,n1358);
or (n1354,n1355,n371);
nor (n1355,n1356,n1357);
and (n1356,n382,n346);
and (n1357,n381,n342);
or (n1358,n1309,n372);
nand (n1359,n1360,n1364);
or (n1360,n475,n1361);
nor (n1361,n1362,n1363);
and (n1362,n185,n296);
and (n1363,n189,n289);
or (n1364,n1315,n476);
and (n1365,n1347,n1353);
xor (n1366,n1229,n1237);
xor (n1367,n1306,n1319);
or (n1368,n1369,n1391);
and (n1369,n1370,n1390);
xor (n1370,n1371,n1372);
xor (n1371,n1320,n1326);
or (n1372,n1373,n1389);
and (n1373,n1374,n1383);
xor (n1374,n1375,n1376);
nor (n1375,n287,n198);
nand (n1376,n1377,n1382);
or (n1377,n1378,n242);
not (n1378,n1379);
nand (n1379,n1380,n1381);
or (n1380,n237,n427);
nand (n1381,n427,n237);
or (n1382,n1328,n243);
nand (n1383,n1384,n1388);
or (n1384,n371,n1385);
nor (n1385,n1386,n1387);
and (n1386,n381,n334);
and (n1387,n382,n338);
or (n1388,n1355,n372);
and (n1389,n1375,n1376);
xor (n1390,n1346,n1359);
and (n1391,n1371,n1372);
or (n1392,n1393,n1394);
xor (n1393,n1303,n1334);
or (n1394,n1395,n1396);
and (n1395,n1343,n1367);
and (n1396,n1344,n1366);
nor (n1397,n1398,n1523);
and (n1398,n1399,n1518);
or (n1399,n1400,n1517);
and (n1400,n1401,n1442);
xor (n1401,n1402,n1435);
or (n1402,n1403,n1434);
and (n1403,n1404,n1420);
xor (n1404,n1405,n1411);
nand (n1405,n1406,n1410);
or (n1406,n371,n1407);
nor (n1407,n1408,n1409);
and (n1408,n382,n189);
and (n1409,n381,n185);
or (n1410,n1385,n372);
or (n1411,n1412,n1416);
nor (n1412,n1413,n476);
nor (n1413,n1414,n1415);
and (n1414,n296,n176);
and (n1415,n289,n180);
nor (n1416,n475,n1417);
nor (n1417,n1418,n1419);
and (n1418,n289,n198);
and (n1419,n296,n196);
xor (n1420,n1421,n1427);
nor (n1421,n1422,n296);
nor (n1422,n1423,n1426);
and (n1423,n1424,n381);
not (n1424,n1425);
and (n1425,n196,n479);
and (n1426,n485,n198);
nand (n1427,n1428,n1433);
or (n1428,n242,n1429);
not (n1429,n1430);
nand (n1430,n1431,n1432);
or (n1431,n236,n342);
nand (n1432,n342,n236);
nand (n1433,n1379,n244);
and (n1434,n1405,n1411);
xor (n1435,n1436,n1441);
xor (n1436,n1437,n1440);
nand (n1437,n1438,n1439);
or (n1438,n475,n1413);
or (n1439,n1361,n476);
and (n1440,n1421,n1427);
xor (n1441,n1374,n1383);
or (n1442,n1443,n1516);
and (n1443,n1444,n1464);
xor (n1444,n1445,n1463);
or (n1445,n1446,n1462);
and (n1446,n1447,n1456);
xor (n1447,n1448,n1449);
and (n1448,n477,n196);
nand (n1449,n1450,n1455);
or (n1450,n242,n1451);
not (n1451,n1452);
nand (n1452,n1453,n1454);
or (n1453,n237,n338);
nand (n1454,n338,n237);
nand (n1455,n1430,n244);
nand (n1456,n1457,n1461);
or (n1457,n371,n1458);
nor (n1458,n1459,n1460);
and (n1459,n381,n176);
and (n1460,n382,n180);
or (n1461,n1407,n372);
and (n1462,n1448,n1449);
xor (n1463,n1404,n1420);
or (n1464,n1465,n1515);
and (n1465,n1466,n1483);
xor (n1466,n1467,n1482);
and (n1467,n1468,n1474);
and (n1468,n1469,n382);
nand (n1469,n1470,n1473);
nand (n1470,n1471,n236);
not (n1471,n1472);
and (n1472,n196,n374);
nand (n1473,n378,n198);
nand (n1474,n1475,n1476);
or (n1475,n243,n1451);
nand (n1476,n1477,n1481);
not (n1477,n1478);
nor (n1478,n1479,n1480);
and (n1479,n189,n237);
and (n1480,n185,n236);
not (n1481,n242);
xor (n1482,n1447,n1456);
or (n1483,n1484,n1514);
and (n1484,n1485,n1493);
xor (n1485,n1486,n1492);
nand (n1486,n1487,n1491);
or (n1487,n371,n1488);
nor (n1488,n1489,n1490);
and (n1489,n382,n198);
and (n1490,n381,n196);
or (n1491,n1458,n372);
xor (n1492,n1468,n1474);
or (n1493,n1494,n1513);
and (n1494,n1495,n1503);
xor (n1495,n1496,n1497);
nor (n1496,n372,n198);
nand (n1497,n1498,n1502);
or (n1498,n1499,n242);
or (n1499,n1500,n1501);
and (n1500,n236,n180);
and (n1501,n176,n237);
or (n1502,n1478,n243);
nor (n1503,n1504,n1511);
nor (n1504,n1505,n1507);
and (n1505,n1506,n244);
not (n1506,n1499);
and (n1507,n1508,n1481);
nand (n1508,n1509,n1510);
or (n1509,n236,n196);
or (n1510,n237,n198);
or (n1511,n236,n1512);
and (n1512,n196,n244);
and (n1513,n1496,n1497);
and (n1514,n1486,n1492);
and (n1515,n1467,n1482);
and (n1516,n1445,n1463);
and (n1517,n1402,n1435);
or (n1518,n1519,n1520);
xor (n1519,n1370,n1390);
or (n1520,n1521,n1522);
and (n1521,n1436,n1441);
and (n1522,n1437,n1440);
and (n1523,n1519,n1520);
nand (n1524,n1392,n1525);
and (n1525,n1342,n1368);
nand (n1526,n1393,n1394);
and (n1527,n1301,n1336);
and (n1528,n1178,n1283);
or (n1529,n1530,n1537);
xor (n1530,n1531,n1536);
xor (n1531,n1532,n1533);
xor (n1532,n1033,n1053);
or (n1533,n1534,n1535);
and (n1534,n1290,n1297);
and (n1535,n1291,n1294);
xor (n1536,n1147,n1150);
or (n1537,n1538,n1539);
and (n1538,n1284,n1289);
and (n1539,n1285,n1286);
nor (n1540,n1541,n1542);
xor (n1541,n1144,n1169);
or (n1542,n1543,n1544);
and (n1543,n1531,n1536);
and (n1544,n1532,n1533);
or (n1545,n1540,n1546);
nand (n1546,n1530,n1537);
nand (n1547,n1541,n1542);
and (n1548,n1142,n1171);
and (n1549,n847,n1078);
nor (n1550,n1551,n1596);
nor (n1551,n1552,n1587);
xor (n1552,n1553,n1572);
xor (n1553,n1554,n1555);
xor (n1554,n830,n833);
or (n1555,n1556,n1571);
and (n1556,n1557,n1564);
xor (n1557,n1558,n1561);
or (n1558,n1559,n1560);
and (n1559,n1122,n1136);
and (n1560,n1123,n1126);
or (n1561,n1562,n1563);
and (n1562,n1081,n1088);
and (n1563,n1082,n1085);
xor (n1564,n1565,n1568);
xor (n1565,n1566,n1567);
and (n1566,n1127,n1130);
xor (n1567,n767,n775);
or (n1568,n1569,n1570);
and (n1569,n1105,n1115);
and (n1570,n1106,n1109);
and (n1571,n1558,n1561);
xor (n1572,n1573,n1578);
xor (n1573,n1574,n1577);
or (n1574,n1575,n1576);
and (n1575,n1565,n1568);
and (n1576,n1566,n1567);
xor (n1577,n764,n805);
or (n1578,n1579,n1586);
and (n1579,n1580,n1585);
xor (n1580,n1581,n1584);
or (n1581,n1582,n1583);
and (n1582,n1089,n1096);
and (n1583,n1090,n1093);
xor (n1584,n784,n798);
xor (n1585,n807,n820);
and (n1586,n1581,n1584);
or (n1587,n1588,n1595);
and (n1588,n1589,n1594);
xor (n1589,n1590,n1591);
xor (n1590,n1580,n1585);
or (n1591,n1592,n1593);
and (n1592,n1103,n1121);
and (n1593,n1104,n1118);
xor (n1594,n1557,n1564);
and (n1595,n1590,n1591);
nor (n1596,n1597,n1598);
xor (n1597,n1589,n1594);
or (n1598,n1599,n1600);
and (n1599,n1079,n1102);
and (n1600,n1080,n1099);
or (n1601,n1602,n1613);
nor (n1602,n1603,n1604);
xor (n1603,n757,n837);
or (n1604,n1605,n1612);
and (n1605,n1606,n1611);
xor (n1606,n1607,n1608);
xor (n1607,n599,n637);
or (n1608,n1609,n1610);
and (n1609,n1573,n1578);
and (n1610,n1574,n1577);
xor (n1611,n761,n835);
and (n1612,n1607,n1608);
nor (n1613,n1614,n1617);
or (n1614,n1615,n1616);
and (n1615,n1553,n1572);
and (n1616,n1554,n1555);
xor (n1617,n1606,n1611);
nand (n1618,n1619,n1628);
or (n1619,n1620,n1602);
nor (n1620,n1621,n1627);
and (n1621,n1622,n1626);
nand (n1622,n1623,n1625);
or (n1623,n1551,n1624);
nand (n1624,n1597,n1598);
nand (n1625,n1552,n1587);
not (n1626,n1613);
and (n1627,n1614,n1617);
nand (n1628,n1603,n1604);
or (n1629,n841,n3);
xor (n1630,n1631,n2761);
xor (n1631,n1632,n2758);
xor (n1632,n1633,n2757);
xor (n1633,n1634,n2749);
xor (n1634,n1635,n2748);
xor (n1635,n1636,n2733);
xor (n1636,n1637,n2732);
xor (n1637,n1638,n2712);
xor (n1638,n1639,n2711);
xor (n1639,n1640,n2684);
xor (n1640,n1641,n2683);
xor (n1641,n1642,n2651);
xor (n1642,n1643,n2650);
xor (n1643,n1644,n2611);
xor (n1644,n1645,n2610);
xor (n1645,n1646,n2566);
xor (n1646,n1647,n2565);
xor (n1647,n1648,n2514);
xor (n1648,n1649,n2513);
xor (n1649,n1650,n2457);
xor (n1650,n1651,n2456);
xor (n1651,n1652,n2393);
xor (n1652,n1653,n2392);
xor (n1653,n1654,n2324);
xor (n1654,n1655,n2323);
xor (n1655,n1656,n2249);
xor (n1656,n1657,n2248);
xor (n1657,n1658,n2168);
xor (n1658,n1659,n2167);
xor (n1659,n1660,n2080);
xor (n1660,n1661,n2079);
xor (n1661,n1662,n1987);
xor (n1662,n1663,n1986);
xor (n1663,n1664,n1887);
xor (n1664,n1665,n1886);
xor (n1665,n1666,n1782);
xor (n1666,n1667,n1781);
xor (n1667,n1668,n1671);
xor (n1668,n1669,n1670);
and (n1669,n696,n244);
and (n1670,n248,n237);
or (n1671,n1672,n1675);
and (n1672,n1673,n1674);
and (n1673,n248,n244);
and (n1674,n203,n237);
and (n1675,n1676,n1677);
xor (n1676,n1673,n1674);
or (n1677,n1678,n1681);
and (n1678,n1679,n1680);
and (n1679,n203,n244);
and (n1680,n268,n237);
and (n1681,n1682,n1683);
xor (n1682,n1679,n1680);
or (n1683,n1684,n1687);
and (n1684,n1685,n1686);
and (n1685,n268,n244);
and (n1686,n396,n237);
and (n1687,n1688,n1689);
xor (n1688,n1685,n1686);
or (n1689,n1690,n1693);
and (n1690,n1691,n1692);
and (n1691,n396,n244);
and (n1692,n388,n237);
and (n1693,n1694,n1695);
xor (n1694,n1691,n1692);
or (n1695,n1696,n1699);
and (n1696,n1697,n1698);
and (n1697,n388,n244);
and (n1698,n489,n237);
and (n1699,n1700,n1701);
xor (n1700,n1697,n1698);
or (n1701,n1702,n1705);
and (n1702,n1703,n1704);
and (n1703,n489,n244);
and (n1704,n413,n237);
and (n1705,n1706,n1707);
xor (n1706,n1703,n1704);
or (n1707,n1708,n1711);
and (n1708,n1709,n1710);
and (n1709,n413,n244);
and (n1710,n278,n237);
and (n1711,n1712,n1713);
xor (n1712,n1709,n1710);
or (n1713,n1714,n1717);
and (n1714,n1715,n1716);
and (n1715,n278,n244);
and (n1716,n305,n237);
and (n1717,n1718,n1719);
xor (n1718,n1715,n1716);
or (n1719,n1720,n1723);
and (n1720,n1721,n1722);
and (n1721,n305,n244);
and (n1722,n464,n237);
and (n1723,n1724,n1725);
xor (n1724,n1721,n1722);
or (n1725,n1726,n1729);
and (n1726,n1727,n1728);
and (n1727,n464,n244);
and (n1728,n528,n237);
and (n1729,n1730,n1731);
xor (n1730,n1727,n1728);
or (n1731,n1732,n1735);
and (n1732,n1733,n1734);
and (n1733,n528,n244);
and (n1734,n127,n237);
and (n1735,n1736,n1737);
xor (n1736,n1733,n1734);
or (n1737,n1738,n1741);
and (n1738,n1739,n1740);
and (n1739,n127,n244);
and (n1740,n94,n237);
and (n1741,n1742,n1743);
xor (n1742,n1739,n1740);
or (n1743,n1744,n1747);
and (n1744,n1745,n1746);
and (n1745,n94,n244);
and (n1746,n608,n237);
and (n1747,n1748,n1749);
xor (n1748,n1745,n1746);
or (n1749,n1750,n1753);
and (n1750,n1751,n1752);
and (n1751,n608,n244);
and (n1752,n423,n237);
and (n1753,n1754,n1755);
xor (n1754,n1751,n1752);
or (n1755,n1756,n1759);
and (n1756,n1757,n1758);
and (n1757,n423,n244);
and (n1758,n342,n237);
and (n1759,n1760,n1761);
xor (n1760,n1757,n1758);
or (n1761,n1762,n1765);
and (n1762,n1763,n1764);
and (n1763,n342,n244);
and (n1764,n334,n237);
and (n1765,n1766,n1767);
xor (n1766,n1763,n1764);
or (n1767,n1768,n1771);
and (n1768,n1769,n1770);
and (n1769,n334,n244);
and (n1770,n185,n237);
and (n1771,n1772,n1773);
xor (n1772,n1769,n1770);
or (n1773,n1774,n1776);
and (n1774,n1775,n1501);
and (n1775,n185,n244);
and (n1776,n1777,n1778);
xor (n1777,n1775,n1501);
and (n1778,n1779,n1780);
and (n1779,n176,n244);
and (n1780,n196,n237);
and (n1781,n203,n374);
or (n1782,n1783,n1786);
and (n1783,n1784,n1785);
xor (n1784,n1676,n1677);
and (n1785,n268,n374);
and (n1786,n1787,n1788);
xor (n1787,n1784,n1785);
or (n1788,n1789,n1792);
and (n1789,n1790,n1791);
xor (n1790,n1682,n1683);
and (n1791,n396,n374);
and (n1792,n1793,n1794);
xor (n1793,n1790,n1791);
or (n1794,n1795,n1798);
and (n1795,n1796,n1797);
xor (n1796,n1688,n1689);
and (n1797,n388,n374);
and (n1798,n1799,n1800);
xor (n1799,n1796,n1797);
or (n1800,n1801,n1804);
and (n1801,n1802,n1803);
xor (n1802,n1694,n1695);
and (n1803,n489,n374);
and (n1804,n1805,n1806);
xor (n1805,n1802,n1803);
or (n1806,n1807,n1810);
and (n1807,n1808,n1809);
xor (n1808,n1700,n1701);
and (n1809,n413,n374);
and (n1810,n1811,n1812);
xor (n1811,n1808,n1809);
or (n1812,n1813,n1816);
and (n1813,n1814,n1815);
xor (n1814,n1706,n1707);
and (n1815,n278,n374);
and (n1816,n1817,n1818);
xor (n1817,n1814,n1815);
or (n1818,n1819,n1822);
and (n1819,n1820,n1821);
xor (n1820,n1712,n1713);
and (n1821,n305,n374);
and (n1822,n1823,n1824);
xor (n1823,n1820,n1821);
or (n1824,n1825,n1828);
and (n1825,n1826,n1827);
xor (n1826,n1718,n1719);
and (n1827,n464,n374);
and (n1828,n1829,n1830);
xor (n1829,n1826,n1827);
or (n1830,n1831,n1834);
and (n1831,n1832,n1833);
xor (n1832,n1724,n1725);
and (n1833,n528,n374);
and (n1834,n1835,n1836);
xor (n1835,n1832,n1833);
or (n1836,n1837,n1840);
and (n1837,n1838,n1839);
xor (n1838,n1730,n1731);
and (n1839,n127,n374);
and (n1840,n1841,n1842);
xor (n1841,n1838,n1839);
or (n1842,n1843,n1846);
and (n1843,n1844,n1845);
xor (n1844,n1736,n1737);
and (n1845,n94,n374);
and (n1846,n1847,n1848);
xor (n1847,n1844,n1845);
or (n1848,n1849,n1852);
and (n1849,n1850,n1851);
xor (n1850,n1742,n1743);
and (n1851,n608,n374);
and (n1852,n1853,n1854);
xor (n1853,n1850,n1851);
or (n1854,n1855,n1858);
and (n1855,n1856,n1857);
xor (n1856,n1748,n1749);
and (n1857,n423,n374);
and (n1858,n1859,n1860);
xor (n1859,n1856,n1857);
or (n1860,n1861,n1864);
and (n1861,n1862,n1863);
xor (n1862,n1754,n1755);
and (n1863,n342,n374);
and (n1864,n1865,n1866);
xor (n1865,n1862,n1863);
or (n1866,n1867,n1870);
and (n1867,n1868,n1869);
xor (n1868,n1760,n1761);
and (n1869,n334,n374);
and (n1870,n1871,n1872);
xor (n1871,n1868,n1869);
or (n1872,n1873,n1876);
and (n1873,n1874,n1875);
xor (n1874,n1766,n1767);
and (n1875,n185,n374);
and (n1876,n1877,n1878);
xor (n1877,n1874,n1875);
or (n1878,n1879,n1882);
and (n1879,n1880,n1881);
xor (n1880,n1772,n1773);
and (n1881,n176,n374);
and (n1882,n1883,n1884);
xor (n1883,n1880,n1881);
and (n1884,n1885,n1472);
xor (n1885,n1777,n1778);
and (n1886,n268,n382);
or (n1887,n1888,n1891);
and (n1888,n1889,n1890);
xor (n1889,n1787,n1788);
and (n1890,n396,n382);
and (n1891,n1892,n1893);
xor (n1892,n1889,n1890);
or (n1893,n1894,n1897);
and (n1894,n1895,n1896);
xor (n1895,n1793,n1794);
and (n1896,n388,n382);
and (n1897,n1898,n1899);
xor (n1898,n1895,n1896);
or (n1899,n1900,n1903);
and (n1900,n1901,n1902);
xor (n1901,n1799,n1800);
and (n1902,n489,n382);
and (n1903,n1904,n1905);
xor (n1904,n1901,n1902);
or (n1905,n1906,n1909);
and (n1906,n1907,n1908);
xor (n1907,n1805,n1806);
and (n1908,n413,n382);
and (n1909,n1910,n1911);
xor (n1910,n1907,n1908);
or (n1911,n1912,n1915);
and (n1912,n1913,n1914);
xor (n1913,n1811,n1812);
and (n1914,n278,n382);
and (n1915,n1916,n1917);
xor (n1916,n1913,n1914);
or (n1917,n1918,n1921);
and (n1918,n1919,n1920);
xor (n1919,n1817,n1818);
and (n1920,n305,n382);
and (n1921,n1922,n1923);
xor (n1922,n1919,n1920);
or (n1923,n1924,n1927);
and (n1924,n1925,n1926);
xor (n1925,n1823,n1824);
and (n1926,n464,n382);
and (n1927,n1928,n1929);
xor (n1928,n1925,n1926);
or (n1929,n1930,n1933);
and (n1930,n1931,n1932);
xor (n1931,n1829,n1830);
and (n1932,n528,n382);
and (n1933,n1934,n1935);
xor (n1934,n1931,n1932);
or (n1935,n1936,n1939);
and (n1936,n1937,n1938);
xor (n1937,n1835,n1836);
and (n1938,n127,n382);
and (n1939,n1940,n1941);
xor (n1940,n1937,n1938);
or (n1941,n1942,n1945);
and (n1942,n1943,n1944);
xor (n1943,n1841,n1842);
and (n1944,n94,n382);
and (n1945,n1946,n1947);
xor (n1946,n1943,n1944);
or (n1947,n1948,n1951);
and (n1948,n1949,n1950);
xor (n1949,n1847,n1848);
and (n1950,n608,n382);
and (n1951,n1952,n1953);
xor (n1952,n1949,n1950);
or (n1953,n1954,n1957);
and (n1954,n1955,n1956);
xor (n1955,n1853,n1854);
and (n1956,n423,n382);
and (n1957,n1958,n1959);
xor (n1958,n1955,n1956);
or (n1959,n1960,n1963);
and (n1960,n1961,n1962);
xor (n1961,n1859,n1860);
and (n1962,n342,n382);
and (n1963,n1964,n1965);
xor (n1964,n1961,n1962);
or (n1965,n1966,n1969);
and (n1966,n1967,n1968);
xor (n1967,n1865,n1866);
and (n1968,n334,n382);
and (n1969,n1970,n1971);
xor (n1970,n1967,n1968);
or (n1971,n1972,n1975);
and (n1972,n1973,n1974);
xor (n1973,n1871,n1872);
and (n1974,n185,n382);
and (n1975,n1976,n1977);
xor (n1976,n1973,n1974);
or (n1977,n1978,n1981);
and (n1978,n1979,n1980);
xor (n1979,n1877,n1878);
and (n1980,n176,n382);
and (n1981,n1982,n1983);
xor (n1982,n1979,n1980);
and (n1983,n1984,n1985);
xor (n1984,n1883,n1884);
and (n1985,n196,n382);
and (n1986,n396,n479);
or (n1987,n1988,n1991);
and (n1988,n1989,n1990);
xor (n1989,n1892,n1893);
and (n1990,n388,n479);
and (n1991,n1992,n1993);
xor (n1992,n1989,n1990);
or (n1993,n1994,n1997);
and (n1994,n1995,n1996);
xor (n1995,n1898,n1899);
and (n1996,n489,n479);
and (n1997,n1998,n1999);
xor (n1998,n1995,n1996);
or (n1999,n2000,n2003);
and (n2000,n2001,n2002);
xor (n2001,n1904,n1905);
and (n2002,n413,n479);
and (n2003,n2004,n2005);
xor (n2004,n2001,n2002);
or (n2005,n2006,n2009);
and (n2006,n2007,n2008);
xor (n2007,n1910,n1911);
and (n2008,n278,n479);
and (n2009,n2010,n2011);
xor (n2010,n2007,n2008);
or (n2011,n2012,n2015);
and (n2012,n2013,n2014);
xor (n2013,n1916,n1917);
and (n2014,n305,n479);
and (n2015,n2016,n2017);
xor (n2016,n2013,n2014);
or (n2017,n2018,n2021);
and (n2018,n2019,n2020);
xor (n2019,n1922,n1923);
and (n2020,n464,n479);
and (n2021,n2022,n2023);
xor (n2022,n2019,n2020);
or (n2023,n2024,n2027);
and (n2024,n2025,n2026);
xor (n2025,n1928,n1929);
and (n2026,n528,n479);
and (n2027,n2028,n2029);
xor (n2028,n2025,n2026);
or (n2029,n2030,n2033);
and (n2030,n2031,n2032);
xor (n2031,n1934,n1935);
and (n2032,n127,n479);
and (n2033,n2034,n2035);
xor (n2034,n2031,n2032);
or (n2035,n2036,n2039);
and (n2036,n2037,n2038);
xor (n2037,n1940,n1941);
and (n2038,n94,n479);
and (n2039,n2040,n2041);
xor (n2040,n2037,n2038);
or (n2041,n2042,n2045);
and (n2042,n2043,n2044);
xor (n2043,n1946,n1947);
and (n2044,n608,n479);
and (n2045,n2046,n2047);
xor (n2046,n2043,n2044);
or (n2047,n2048,n2051);
and (n2048,n2049,n2050);
xor (n2049,n1952,n1953);
and (n2050,n423,n479);
and (n2051,n2052,n2053);
xor (n2052,n2049,n2050);
or (n2053,n2054,n2057);
and (n2054,n2055,n2056);
xor (n2055,n1958,n1959);
and (n2056,n342,n479);
and (n2057,n2058,n2059);
xor (n2058,n2055,n2056);
or (n2059,n2060,n2063);
and (n2060,n2061,n2062);
xor (n2061,n1964,n1965);
and (n2062,n334,n479);
and (n2063,n2064,n2065);
xor (n2064,n2061,n2062);
or (n2065,n2066,n2069);
and (n2066,n2067,n2068);
xor (n2067,n1970,n1971);
and (n2068,n185,n479);
and (n2069,n2070,n2071);
xor (n2070,n2067,n2068);
or (n2071,n2072,n2075);
and (n2072,n2073,n2074);
xor (n2073,n1976,n1977);
and (n2074,n176,n479);
and (n2075,n2076,n2077);
xor (n2076,n2073,n2074);
and (n2077,n2078,n1425);
xor (n2078,n1982,n1983);
and (n2079,n388,n289);
or (n2080,n2081,n2084);
and (n2081,n2082,n2083);
xor (n2082,n1992,n1993);
and (n2083,n489,n289);
and (n2084,n2085,n2086);
xor (n2085,n2082,n2083);
or (n2086,n2087,n2090);
and (n2087,n2088,n2089);
xor (n2088,n1998,n1999);
and (n2089,n413,n289);
and (n2090,n2091,n2092);
xor (n2091,n2088,n2089);
or (n2092,n2093,n2096);
and (n2093,n2094,n2095);
xor (n2094,n2004,n2005);
and (n2095,n278,n289);
and (n2096,n2097,n2098);
xor (n2097,n2094,n2095);
or (n2098,n2099,n2102);
and (n2099,n2100,n2101);
xor (n2100,n2010,n2011);
and (n2101,n305,n289);
and (n2102,n2103,n2104);
xor (n2103,n2100,n2101);
or (n2104,n2105,n2108);
and (n2105,n2106,n2107);
xor (n2106,n2016,n2017);
and (n2107,n464,n289);
and (n2108,n2109,n2110);
xor (n2109,n2106,n2107);
or (n2110,n2111,n2114);
and (n2111,n2112,n2113);
xor (n2112,n2022,n2023);
and (n2113,n528,n289);
and (n2114,n2115,n2116);
xor (n2115,n2112,n2113);
or (n2116,n2117,n2120);
and (n2117,n2118,n2119);
xor (n2118,n2028,n2029);
and (n2119,n127,n289);
and (n2120,n2121,n2122);
xor (n2121,n2118,n2119);
or (n2122,n2123,n2126);
and (n2123,n2124,n2125);
xor (n2124,n2034,n2035);
and (n2125,n94,n289);
and (n2126,n2127,n2128);
xor (n2127,n2124,n2125);
or (n2128,n2129,n2132);
and (n2129,n2130,n2131);
xor (n2130,n2040,n2041);
and (n2131,n608,n289);
and (n2132,n2133,n2134);
xor (n2133,n2130,n2131);
or (n2134,n2135,n2138);
and (n2135,n2136,n2137);
xor (n2136,n2046,n2047);
and (n2137,n423,n289);
and (n2138,n2139,n2140);
xor (n2139,n2136,n2137);
or (n2140,n2141,n2144);
and (n2141,n2142,n2143);
xor (n2142,n2052,n2053);
and (n2143,n342,n289);
and (n2144,n2145,n2146);
xor (n2145,n2142,n2143);
or (n2146,n2147,n2150);
and (n2147,n2148,n2149);
xor (n2148,n2058,n2059);
and (n2149,n334,n289);
and (n2150,n2151,n2152);
xor (n2151,n2148,n2149);
or (n2152,n2153,n2156);
and (n2153,n2154,n2155);
xor (n2154,n2064,n2065);
and (n2155,n185,n289);
and (n2156,n2157,n2158);
xor (n2157,n2154,n2155);
or (n2158,n2159,n2162);
and (n2159,n2160,n2161);
xor (n2160,n2070,n2071);
and (n2161,n176,n289);
and (n2162,n2163,n2164);
xor (n2163,n2160,n2161);
and (n2164,n2165,n2166);
xor (n2165,n2076,n2077);
and (n2166,n196,n289);
and (n2167,n489,n292);
or (n2168,n2169,n2172);
and (n2169,n2170,n2171);
xor (n2170,n2085,n2086);
and (n2171,n413,n292);
and (n2172,n2173,n2174);
xor (n2173,n2170,n2171);
or (n2174,n2175,n2178);
and (n2175,n2176,n2177);
xor (n2176,n2091,n2092);
and (n2177,n278,n292);
and (n2178,n2179,n2180);
xor (n2179,n2176,n2177);
or (n2180,n2181,n2184);
and (n2181,n2182,n2183);
xor (n2182,n2097,n2098);
and (n2183,n305,n292);
and (n2184,n2185,n2186);
xor (n2185,n2182,n2183);
or (n2186,n2187,n2190);
and (n2187,n2188,n2189);
xor (n2188,n2103,n2104);
and (n2189,n464,n292);
and (n2190,n2191,n2192);
xor (n2191,n2188,n2189);
or (n2192,n2193,n2196);
and (n2193,n2194,n2195);
xor (n2194,n2109,n2110);
and (n2195,n528,n292);
and (n2196,n2197,n2198);
xor (n2197,n2194,n2195);
or (n2198,n2199,n2202);
and (n2199,n2200,n2201);
xor (n2200,n2115,n2116);
and (n2201,n127,n292);
and (n2202,n2203,n2204);
xor (n2203,n2200,n2201);
or (n2204,n2205,n2208);
and (n2205,n2206,n2207);
xor (n2206,n2121,n2122);
and (n2207,n94,n292);
and (n2208,n2209,n2210);
xor (n2209,n2206,n2207);
or (n2210,n2211,n2214);
and (n2211,n2212,n2213);
xor (n2212,n2127,n2128);
and (n2213,n608,n292);
and (n2214,n2215,n2216);
xor (n2215,n2212,n2213);
or (n2216,n2217,n2220);
and (n2217,n2218,n2219);
xor (n2218,n2133,n2134);
and (n2219,n423,n292);
and (n2220,n2221,n2222);
xor (n2221,n2218,n2219);
or (n2222,n2223,n2226);
and (n2223,n2224,n2225);
xor (n2224,n2139,n2140);
and (n2225,n342,n292);
and (n2226,n2227,n2228);
xor (n2227,n2224,n2225);
or (n2228,n2229,n2232);
and (n2229,n2230,n2231);
xor (n2230,n2145,n2146);
and (n2231,n334,n292);
and (n2232,n2233,n2234);
xor (n2233,n2230,n2231);
or (n2234,n2235,n2238);
and (n2235,n2236,n2237);
xor (n2236,n2151,n2152);
and (n2237,n185,n292);
and (n2238,n2239,n2240);
xor (n2239,n2236,n2237);
or (n2240,n2241,n2244);
and (n2241,n2242,n2243);
xor (n2242,n2157,n2158);
and (n2243,n176,n292);
and (n2244,n2245,n2246);
xor (n2245,n2242,n2243);
and (n2246,n2247,n1324);
xor (n2247,n2163,n2164);
and (n2248,n413,n282);
or (n2249,n2250,n2253);
and (n2250,n2251,n2252);
xor (n2251,n2173,n2174);
and (n2252,n278,n282);
and (n2253,n2254,n2255);
xor (n2254,n2251,n2252);
or (n2255,n2256,n2259);
and (n2256,n2257,n2258);
xor (n2257,n2179,n2180);
and (n2258,n305,n282);
and (n2259,n2260,n2261);
xor (n2260,n2257,n2258);
or (n2261,n2262,n2265);
and (n2262,n2263,n2264);
xor (n2263,n2185,n2186);
and (n2264,n464,n282);
and (n2265,n2266,n2267);
xor (n2266,n2263,n2264);
or (n2267,n2268,n2271);
and (n2268,n2269,n2270);
xor (n2269,n2191,n2192);
and (n2270,n528,n282);
and (n2271,n2272,n2273);
xor (n2272,n2269,n2270);
or (n2273,n2274,n2277);
and (n2274,n2275,n2276);
xor (n2275,n2197,n2198);
and (n2276,n127,n282);
and (n2277,n2278,n2279);
xor (n2278,n2275,n2276);
or (n2279,n2280,n2283);
and (n2280,n2281,n2282);
xor (n2281,n2203,n2204);
and (n2282,n94,n282);
and (n2283,n2284,n2285);
xor (n2284,n2281,n2282);
or (n2285,n2286,n2289);
and (n2286,n2287,n2288);
xor (n2287,n2209,n2210);
and (n2288,n608,n282);
and (n2289,n2290,n2291);
xor (n2290,n2287,n2288);
or (n2291,n2292,n2295);
and (n2292,n2293,n2294);
xor (n2293,n2215,n2216);
and (n2294,n423,n282);
and (n2295,n2296,n2297);
xor (n2296,n2293,n2294);
or (n2297,n2298,n2301);
and (n2298,n2299,n2300);
xor (n2299,n2221,n2222);
and (n2300,n342,n282);
and (n2301,n2302,n2303);
xor (n2302,n2299,n2300);
or (n2303,n2304,n2306);
and (n2304,n2305,n1188);
xor (n2305,n2227,n2228);
and (n2306,n2307,n2308);
xor (n2307,n2305,n1188);
or (n2308,n2309,n2312);
and (n2309,n2310,n2311);
xor (n2310,n2233,n2234);
and (n2311,n185,n282);
and (n2312,n2313,n2314);
xor (n2313,n2310,n2311);
or (n2314,n2315,n2318);
and (n2315,n2316,n2317);
xor (n2316,n2239,n2240);
and (n2317,n176,n282);
and (n2318,n2319,n2320);
xor (n2319,n2316,n2317);
and (n2320,n2321,n2322);
xor (n2321,n2245,n2246);
and (n2322,n196,n282);
and (n2323,n278,n449);
or (n2324,n2325,n2328);
and (n2325,n2326,n2327);
xor (n2326,n2254,n2255);
and (n2327,n305,n449);
and (n2328,n2329,n2330);
xor (n2329,n2326,n2327);
or (n2330,n2331,n2334);
and (n2331,n2332,n2333);
xor (n2332,n2260,n2261);
and (n2333,n464,n449);
and (n2334,n2335,n2336);
xor (n2335,n2332,n2333);
or (n2336,n2337,n2340);
and (n2337,n2338,n2339);
xor (n2338,n2266,n2267);
and (n2339,n528,n449);
and (n2340,n2341,n2342);
xor (n2341,n2338,n2339);
or (n2342,n2343,n2346);
and (n2343,n2344,n2345);
xor (n2344,n2272,n2273);
and (n2345,n127,n449);
and (n2346,n2347,n2348);
xor (n2347,n2344,n2345);
or (n2348,n2349,n2352);
and (n2349,n2350,n2351);
xor (n2350,n2278,n2279);
and (n2351,n94,n449);
and (n2352,n2353,n2354);
xor (n2353,n2350,n2351);
or (n2354,n2355,n2358);
and (n2355,n2356,n2357);
xor (n2356,n2284,n2285);
and (n2357,n608,n449);
and (n2358,n2359,n2360);
xor (n2359,n2356,n2357);
or (n2360,n2361,n2364);
and (n2361,n2362,n2363);
xor (n2362,n2290,n2291);
and (n2363,n423,n449);
and (n2364,n2365,n2366);
xor (n2365,n2362,n2363);
or (n2366,n2367,n2370);
and (n2367,n2368,n2369);
xor (n2368,n2296,n2297);
and (n2369,n342,n449);
and (n2370,n2371,n2372);
xor (n2371,n2368,n2369);
or (n2372,n2373,n2376);
and (n2373,n2374,n2375);
xor (n2374,n2302,n2303);
and (n2375,n334,n449);
and (n2376,n2377,n2378);
xor (n2377,n2374,n2375);
or (n2378,n2379,n2382);
and (n2379,n2380,n2381);
xor (n2380,n2307,n2308);
and (n2381,n185,n449);
and (n2382,n2383,n2384);
xor (n2383,n2380,n2381);
or (n2384,n2385,n2388);
and (n2385,n2386,n2387);
xor (n2386,n2313,n2314);
and (n2387,n176,n449);
and (n2388,n2389,n2390);
xor (n2389,n2386,n2387);
and (n2390,n2391,n1217);
xor (n2391,n2319,n2320);
and (n2392,n305,n452);
or (n2393,n2394,n2397);
and (n2394,n2395,n2396);
xor (n2395,n2329,n2330);
and (n2396,n464,n452);
and (n2397,n2398,n2399);
xor (n2398,n2395,n2396);
or (n2399,n2400,n2403);
and (n2400,n2401,n2402);
xor (n2401,n2335,n2336);
and (n2402,n528,n452);
and (n2403,n2404,n2405);
xor (n2404,n2401,n2402);
or (n2405,n2406,n2409);
and (n2406,n2407,n2408);
xor (n2407,n2341,n2342);
and (n2408,n127,n452);
and (n2409,n2410,n2411);
xor (n2410,n2407,n2408);
or (n2411,n2412,n2415);
and (n2412,n2413,n2414);
xor (n2413,n2347,n2348);
and (n2414,n94,n452);
and (n2415,n2416,n2417);
xor (n2416,n2413,n2414);
or (n2417,n2418,n2421);
and (n2418,n2419,n2420);
xor (n2419,n2353,n2354);
and (n2420,n608,n452);
and (n2421,n2422,n2423);
xor (n2422,n2419,n2420);
or (n2423,n2424,n2427);
and (n2424,n2425,n2426);
xor (n2425,n2359,n2360);
and (n2426,n423,n452);
and (n2427,n2428,n2429);
xor (n2428,n2425,n2426);
or (n2429,n2430,n2433);
and (n2430,n2431,n2432);
xor (n2431,n2365,n2366);
and (n2432,n342,n452);
and (n2433,n2434,n2435);
xor (n2434,n2431,n2432);
or (n2435,n2436,n2439);
and (n2436,n2437,n2438);
xor (n2437,n2371,n2372);
and (n2438,n334,n452);
and (n2439,n2440,n2441);
xor (n2440,n2437,n2438);
or (n2441,n2442,n2445);
and (n2442,n2443,n2444);
xor (n2443,n2377,n2378);
and (n2444,n185,n452);
and (n2445,n2446,n2447);
xor (n2446,n2443,n2444);
or (n2447,n2448,n2451);
and (n2448,n2449,n2450);
xor (n2449,n2383,n2384);
and (n2450,n176,n452);
and (n2451,n2452,n2453);
xor (n2452,n2449,n2450);
and (n2453,n2454,n2455);
xor (n2454,n2389,n2390);
and (n2455,n196,n452);
and (n2456,n464,n518);
or (n2457,n2458,n2461);
and (n2458,n2459,n2460);
xor (n2459,n2398,n2399);
and (n2460,n528,n518);
and (n2461,n2462,n2463);
xor (n2462,n2459,n2460);
or (n2463,n2464,n2467);
and (n2464,n2465,n2466);
xor (n2465,n2404,n2405);
and (n2466,n127,n518);
and (n2467,n2468,n2469);
xor (n2468,n2465,n2466);
or (n2469,n2470,n2473);
and (n2470,n2471,n2472);
xor (n2471,n2410,n2411);
and (n2472,n94,n518);
and (n2473,n2474,n2475);
xor (n2474,n2471,n2472);
or (n2475,n2476,n2479);
and (n2476,n2477,n2478);
xor (n2477,n2416,n2417);
and (n2478,n608,n518);
and (n2479,n2480,n2481);
xor (n2480,n2477,n2478);
or (n2481,n2482,n2485);
and (n2482,n2483,n2484);
xor (n2483,n2422,n2423);
and (n2484,n423,n518);
and (n2485,n2486,n2487);
xor (n2486,n2483,n2484);
or (n2487,n2488,n2491);
and (n2488,n2489,n2490);
xor (n2489,n2428,n2429);
and (n2490,n342,n518);
and (n2491,n2492,n2493);
xor (n2492,n2489,n2490);
or (n2493,n2494,n2497);
and (n2494,n2495,n2496);
xor (n2495,n2434,n2435);
and (n2496,n334,n518);
and (n2497,n2498,n2499);
xor (n2498,n2495,n2496);
or (n2499,n2500,n2503);
and (n2500,n2501,n2502);
xor (n2501,n2440,n2441);
and (n2502,n185,n518);
and (n2503,n2504,n2505);
xor (n2504,n2501,n2502);
or (n2505,n2506,n2509);
and (n2506,n2507,n2508);
xor (n2507,n2446,n2447);
and (n2508,n176,n518);
and (n2509,n2510,n2511);
xor (n2510,n2507,n2508);
and (n2511,n2512,n1051);
xor (n2512,n2452,n2453);
and (n2513,n528,n87);
or (n2514,n2515,n2518);
and (n2515,n2516,n2517);
xor (n2516,n2462,n2463);
and (n2517,n127,n87);
and (n2518,n2519,n2520);
xor (n2519,n2516,n2517);
or (n2520,n2521,n2524);
and (n2521,n2522,n2523);
xor (n2522,n2468,n2469);
and (n2523,n94,n87);
and (n2524,n2525,n2526);
xor (n2525,n2522,n2523);
or (n2526,n2527,n2530);
and (n2527,n2528,n2529);
xor (n2528,n2474,n2475);
and (n2529,n608,n87);
and (n2530,n2531,n2532);
xor (n2531,n2528,n2529);
or (n2532,n2533,n2536);
and (n2533,n2534,n2535);
xor (n2534,n2480,n2481);
and (n2535,n423,n87);
and (n2536,n2537,n2538);
xor (n2537,n2534,n2535);
or (n2538,n2539,n2542);
and (n2539,n2540,n2541);
xor (n2540,n2486,n2487);
and (n2541,n342,n87);
and (n2542,n2543,n2544);
xor (n2543,n2540,n2541);
or (n2544,n2545,n2548);
and (n2545,n2546,n2547);
xor (n2546,n2492,n2493);
and (n2547,n334,n87);
and (n2548,n2549,n2550);
xor (n2549,n2546,n2547);
or (n2550,n2551,n2554);
and (n2551,n2552,n2553);
xor (n2552,n2498,n2499);
and (n2553,n185,n87);
and (n2554,n2555,n2556);
xor (n2555,n2552,n2553);
or (n2556,n2557,n2560);
and (n2557,n2558,n2559);
xor (n2558,n2504,n2505);
and (n2559,n176,n87);
and (n2560,n2561,n2562);
xor (n2561,n2558,n2559);
and (n2562,n2563,n2564);
xor (n2563,n2510,n2511);
and (n2564,n196,n87);
and (n2565,n127,n80);
or (n2566,n2567,n2570);
and (n2567,n2568,n2569);
xor (n2568,n2519,n2520);
and (n2569,n94,n80);
and (n2570,n2571,n2572);
xor (n2571,n2568,n2569);
or (n2572,n2573,n2576);
and (n2573,n2574,n2575);
xor (n2574,n2525,n2526);
and (n2575,n608,n80);
and (n2576,n2577,n2578);
xor (n2577,n2574,n2575);
or (n2578,n2579,n2582);
and (n2579,n2580,n2581);
xor (n2580,n2531,n2532);
and (n2581,n423,n80);
and (n2582,n2583,n2584);
xor (n2583,n2580,n2581);
or (n2584,n2585,n2588);
and (n2585,n2586,n2587);
xor (n2586,n2537,n2538);
and (n2587,n342,n80);
and (n2588,n2589,n2590);
xor (n2589,n2586,n2587);
or (n2590,n2591,n2594);
and (n2591,n2592,n2593);
xor (n2592,n2543,n2544);
and (n2593,n334,n80);
and (n2594,n2595,n2596);
xor (n2595,n2592,n2593);
or (n2596,n2597,n2600);
and (n2597,n2598,n2599);
xor (n2598,n2549,n2550);
and (n2599,n185,n80);
and (n2600,n2601,n2602);
xor (n2601,n2598,n2599);
or (n2602,n2603,n2606);
and (n2603,n2604,n2605);
xor (n2604,n2555,n2556);
and (n2605,n176,n80);
and (n2606,n2607,n2608);
xor (n2607,n2604,n2605);
and (n2608,n2609,n960);
xor (n2609,n2561,n2562);
and (n2610,n94,n17);
or (n2611,n2612,n2615);
and (n2612,n2613,n2614);
xor (n2613,n2571,n2572);
and (n2614,n608,n17);
and (n2615,n2616,n2617);
xor (n2616,n2613,n2614);
or (n2617,n2618,n2621);
and (n2618,n2619,n2620);
xor (n2619,n2577,n2578);
and (n2620,n423,n17);
and (n2621,n2622,n2623);
xor (n2622,n2619,n2620);
or (n2623,n2624,n2627);
and (n2624,n2625,n2626);
xor (n2625,n2583,n2584);
and (n2626,n342,n17);
and (n2627,n2628,n2629);
xor (n2628,n2625,n2626);
or (n2629,n2630,n2633);
and (n2630,n2631,n2632);
xor (n2631,n2589,n2590);
and (n2632,n334,n17);
and (n2633,n2634,n2635);
xor (n2634,n2631,n2632);
or (n2635,n2636,n2639);
and (n2636,n2637,n2638);
xor (n2637,n2595,n2596);
and (n2638,n185,n17);
and (n2639,n2640,n2641);
xor (n2640,n2637,n2638);
or (n2641,n2642,n2645);
and (n2642,n2643,n2644);
xor (n2643,n2601,n2602);
and (n2644,n176,n17);
and (n2645,n2646,n2647);
xor (n2646,n2643,n2644);
and (n2647,n2648,n2649);
xor (n2648,n2607,n2608);
and (n2649,n196,n17);
and (n2650,n608,n320);
or (n2651,n2652,n2655);
and (n2652,n2653,n2654);
xor (n2653,n2616,n2617);
and (n2654,n423,n320);
and (n2655,n2656,n2657);
xor (n2656,n2653,n2654);
or (n2657,n2658,n2661);
and (n2658,n2659,n2660);
xor (n2659,n2622,n2623);
and (n2660,n342,n320);
and (n2661,n2662,n2663);
xor (n2662,n2659,n2660);
or (n2663,n2664,n2667);
and (n2664,n2665,n2666);
xor (n2665,n2628,n2629);
and (n2666,n334,n320);
and (n2667,n2668,n2669);
xor (n2668,n2665,n2666);
or (n2669,n2670,n2673);
and (n2670,n2671,n2672);
xor (n2671,n2634,n2635);
and (n2672,n185,n320);
and (n2673,n2674,n2675);
xor (n2674,n2671,n2672);
or (n2675,n2676,n2679);
and (n2676,n2677,n2678);
xor (n2677,n2640,n2641);
and (n2678,n176,n320);
and (n2679,n2680,n2681);
xor (n2680,n2677,n2678);
and (n2681,n2682,n1134);
xor (n2682,n2646,n2647);
and (n2683,n423,n327);
or (n2684,n2685,n2688);
and (n2685,n2686,n2687);
xor (n2686,n2656,n2657);
and (n2687,n342,n327);
and (n2688,n2689,n2690);
xor (n2689,n2686,n2687);
or (n2690,n2691,n2694);
and (n2691,n2692,n2693);
xor (n2692,n2662,n2663);
and (n2693,n334,n327);
and (n2694,n2695,n2696);
xor (n2695,n2692,n2693);
or (n2696,n2697,n2700);
and (n2697,n2698,n2699);
xor (n2698,n2668,n2669);
and (n2699,n185,n327);
and (n2700,n2701,n2702);
xor (n2701,n2698,n2699);
or (n2702,n2703,n2706);
and (n2703,n2704,n2705);
xor (n2704,n2674,n2675);
and (n2705,n176,n327);
and (n2706,n2707,n2708);
xor (n2707,n2704,n2705);
and (n2708,n2709,n2710);
xor (n2709,n2680,n2681);
and (n2710,n196,n327);
and (n2711,n342,n355);
or (n2712,n2713,n2716);
and (n2713,n2714,n2715);
xor (n2714,n2689,n2690);
and (n2715,n334,n355);
and (n2716,n2717,n2718);
xor (n2717,n2714,n2715);
or (n2718,n2719,n2722);
and (n2719,n2720,n2721);
xor (n2720,n2695,n2696);
and (n2721,n185,n355);
and (n2722,n2723,n2724);
xor (n2723,n2720,n2721);
or (n2724,n2725,n2728);
and (n2725,n2726,n2727);
xor (n2726,n2701,n2702);
and (n2727,n176,n355);
and (n2728,n2729,n2730);
xor (n2729,n2726,n2727);
and (n2730,n2731,n628);
xor (n2731,n2707,n2708);
and (n2732,n334,n158);
or (n2733,n2734,n2737);
and (n2734,n2735,n2736);
xor (n2735,n2717,n2718);
and (n2736,n185,n158);
and (n2737,n2738,n2739);
xor (n2738,n2735,n2736);
or (n2739,n2740,n2743);
and (n2740,n2741,n2742);
xor (n2741,n2723,n2724);
and (n2742,n176,n158);
and (n2743,n2744,n2745);
xor (n2744,n2741,n2742);
and (n2745,n2746,n2747);
xor (n2746,n2729,n2730);
and (n2747,n196,n158);
and (n2748,n185,n140);
or (n2749,n2750,n2753);
and (n2750,n2751,n2752);
xor (n2751,n2738,n2739);
and (n2752,n176,n140);
and (n2753,n2754,n2755);
xor (n2754,n2751,n2752);
and (n2755,n2756,n195);
xor (n2756,n2744,n2745);
and (n2757,n176,n167);
and (n2758,n2759,n2760);
xor (n2759,n2754,n2755);
and (n2760,n196,n167);
and (n2761,n196,n683);
endmodule
