module top (out,n3,n4,n5,n22,n24,n31,n32,n39,n51
        ,n53,n58,n63,n70,n90,n97,n98,n107,n129,n131
        ,n136,n146,n163,n173,n183,n187,n194,n222);
output out;
input n3;
input n4;
input n5;
input n22;
input n24;
input n31;
input n32;
input n39;
input n51;
input n53;
input n58;
input n63;
input n70;
input n90;
input n97;
input n98;
input n107;
input n129;
input n131;
input n136;
input n146;
input n163;
input n173;
input n183;
input n187;
input n194;
input n222;
wire n0;
wire n1;
wire n2;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n23;
wire n25;
wire n26;
wire n27;
wire n28;
wire n29;
wire n30;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n52;
wire n54;
wire n55;
wire n56;
wire n57;
wire n59;
wire n60;
wire n61;
wire n62;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n130;
wire n132;
wire n133;
wire n134;
wire n135;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n184;
wire n185;
wire n186;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
xnor (out,n0,n556);
nor (n0,n1,n6);
and (n1,n2,n5);
nor (n2,n3,n4);
and (n6,n7,n553);
nand (n7,n8,n552);
or (n8,n9,n305);
not (n9,n10);
nand (n10,n11,n304);
nand (n11,n12,n269);
not (n12,n13);
xor (n13,n14,n224);
xor (n14,n15,n110);
xor (n15,n16,n73);
xor (n16,n17,n45);
nand (n17,n18,n34);
or (n18,n19,n27);
not (n19,n20);
nand (n20,n21,n25);
or (n21,n22,n23);
not (n23,n24);
or (n25,n26,n24);
not (n26,n22);
not (n27,n28);
nand (n28,n29,n33);
or (n29,n30,n32);
not (n30,n31);
nand (n33,n32,n30);
nand (n34,n35,n41);
not (n35,n36);
nor (n36,n37,n40);
and (n37,n38,n22);
not (n38,n39);
and (n40,n26,n39);
and (n41,n27,n42);
nand (n42,n43,n44);
nand (n43,n22,n30);
nand (n44,n31,n26);
nand (n45,n46,n66);
or (n46,n47,n61);
not (n47,n48);
nor (n48,n49,n55);
nand (n49,n50,n54);
or (n50,n51,n52);
not (n52,n53);
nand (n54,n51,n52);
nor (n55,n56,n59);
and (n56,n57,n58);
not (n57,n51);
and (n59,n51,n60);
not (n60,n58);
nor (n61,n62,n64);
and (n62,n60,n63);
and (n64,n58,n65);
not (n65,n63);
or (n66,n67,n68);
not (n67,n49);
nor (n68,n69,n71);
and (n69,n60,n70);
and (n71,n58,n72);
not (n72,n70);
nand (n73,n74,n109);
or (n74,n75,n83);
not (n75,n76);
nand (n76,n77,n22);
nand (n77,n78,n79);
or (n78,n39,n31);
nand (n79,n80,n82);
not (n80,n81);
and (n81,n39,n31);
not (n82,n32);
not (n83,n84);
nand (n84,n85,n103);
or (n85,n86,n92);
not (n86,n87);
nand (n87,n88,n91);
or (n88,n53,n89);
not (n89,n90);
or (n91,n52,n90);
nand (n92,n93,n100);
not (n93,n94);
nand (n94,n95,n99);
or (n95,n96,n98);
not (n96,n97);
nand (n99,n98,n96);
nand (n100,n101,n102);
or (n101,n96,n53);
nand (n102,n96,n53);
nand (n103,n94,n104);
nor (n104,n105,n108);
and (n105,n106,n52);
not (n106,n107);
and (n108,n107,n53);
or (n109,n84,n76);
xor (n110,n111,n199);
xor (n111,n112,n150);
or (n112,n113,n149);
and (n113,n114,n123);
xor (n114,n115,n116);
and (n115,n28,n39);
nand (n116,n117,n122);
or (n117,n118,n92);
not (n118,n119);
nand (n119,n120,n121);
or (n120,n53,n72);
or (n121,n52,n70);
nand (n122,n94,n87);
nand (n123,n124,n142);
or (n124,n125,n133);
not (n125,n126);
nor (n126,n127,n132);
and (n127,n128,n130);
not (n128,n129);
not (n130,n131);
and (n132,n129,n131);
nand (n133,n134,n138);
nand (n134,n135,n137);
or (n135,n136,n130);
nand (n137,n130,n136);
not (n138,n139);
nand (n139,n140,n141);
or (n140,n60,n136);
nand (n141,n136,n60);
nand (n142,n143,n139);
not (n143,n144);
nor (n144,n145,n147);
and (n145,n130,n146);
and (n147,n131,n148);
not (n148,n146);
and (n149,n115,n116);
or (n150,n151,n198);
and (n151,n152,n190);
xor (n152,n153,n175);
nand (n153,n154,n169);
or (n154,n155,n159);
not (n155,n156);
nor (n156,n157,n158);
and (n157,n23,n82);
and (n158,n24,n32);
not (n159,n160);
nor (n160,n161,n165);
nand (n161,n162,n164);
or (n162,n130,n163);
nand (n164,n130,n163);
nor (n165,n166,n167);
and (n166,n82,n163);
and (n167,n32,n168);
not (n168,n163);
nand (n169,n161,n170);
nand (n170,n171,n174);
or (n171,n32,n172);
not (n172,n173);
or (n174,n82,n173);
nand (n175,n176,n184);
or (n176,n177,n181);
nor (n177,n178,n180);
and (n178,n179,n107);
not (n179,n98);
and (n180,n98,n106);
nand (n181,n182,n98);
not (n182,n183);
or (n184,n185,n182);
nor (n185,n186,n188);
and (n186,n179,n187);
and (n188,n98,n189);
not (n189,n187);
nand (n190,n191,n197);
or (n191,n47,n192);
nor (n192,n193,n195);
and (n193,n60,n194);
and (n195,n58,n196);
not (n196,n194);
or (n197,n61,n67);
and (n198,n153,n175);
xor (n199,n200,n215);
xor (n200,n201,n207);
nand (n201,n202,n203);
or (n202,n133,n144);
or (n203,n204,n138);
nor (n204,n205,n206);
and (n205,n130,n194);
and (n206,n131,n196);
nand (n207,n208,n214);
or (n208,n209,n213);
not (n209,n210);
nand (n210,n211,n212);
or (n211,n128,n32);
or (n212,n82,n129);
not (n213,n161);
nand (n214,n160,n170);
nand (n215,n216,n217);
or (n216,n185,n181);
or (n217,n218,n182);
not (n218,n219);
nor (n219,n220,n223);
and (n220,n221,n179);
not (n221,n222);
and (n223,n222,n98);
or (n224,n225,n268);
and (n225,n226,n267);
xor (n226,n227,n242);
and (n227,n228,n234);
and (n228,n229,n32);
nand (n229,n230,n231);
or (n230,n39,n163);
nand (n231,n232,n130);
not (n232,n233);
and (n233,n39,n163);
nand (n234,n235,n236);
or (n235,n118,n93);
nand (n236,n237,n241);
not (n237,n238);
nor (n238,n239,n240);
and (n239,n52,n63);
and (n240,n53,n65);
not (n241,n92);
or (n242,n243,n266);
and (n243,n244,n259);
xor (n244,n245,n252);
nand (n245,n246,n251);
or (n246,n247,n133);
not (n247,n248);
nor (n248,n249,n250);
and (n249,n173,n131);
and (n250,n172,n130);
nand (n251,n139,n126);
nand (n252,n253,n258);
or (n253,n254,n159);
not (n254,n255);
nand (n255,n256,n257);
or (n256,n82,n39);
or (n257,n38,n32);
nand (n258,n161,n156);
nand (n259,n260,n265);
or (n260,n181,n261);
not (n261,n262);
nor (n262,n263,n264);
and (n263,n89,n179);
and (n264,n90,n98);
or (n265,n177,n182);
and (n266,n245,n252);
xor (n267,n114,n123);
and (n268,n227,n242);
not (n269,n270);
or (n270,n271,n303);
and (n271,n272,n302);
xor (n272,n273,n274);
xor (n273,n152,n190);
or (n274,n275,n301);
and (n275,n276,n284);
xor (n276,n277,n283);
nand (n277,n278,n282);
or (n278,n47,n279);
nor (n279,n280,n281);
and (n280,n60,n146);
and (n281,n58,n148);
or (n282,n67,n192);
xor (n283,n228,n234);
or (n284,n285,n300);
and (n285,n286,n294);
xor (n286,n287,n288);
and (n287,n161,n39);
nand (n288,n289,n290);
or (n289,n182,n261);
or (n290,n291,n181);
nor (n291,n292,n293);
and (n292,n179,n70);
and (n293,n98,n72);
nand (n294,n295,n299);
or (n295,n133,n296);
nor (n296,n297,n298);
and (n297,n130,n24);
and (n298,n131,n23);
or (n299,n138,n247);
and (n300,n287,n288);
and (n301,n277,n283);
xor (n302,n226,n267);
and (n303,n273,n274);
nand (n304,n13,n270);
not (n305,n306);
nand (n306,n307,n551);
or (n307,n308,n545);
nor (n308,n309,n541);
and (n309,n310,n407);
not (n310,n311);
nand (n311,n312,n395);
not (n312,n313);
nor (n313,n314,n370);
xor (n314,n315,n347);
xor (n315,n316,n346);
or (n316,n317,n345);
and (n317,n318,n336);
xor (n318,n319,n327);
nand (n319,n320,n325);
or (n320,n321,n133);
not (n321,n322);
nand (n322,n323,n324);
or (n323,n130,n39);
or (n324,n131,n38);
nand (n325,n326,n139);
not (n326,n296);
nand (n327,n328,n332);
or (n328,n92,n329);
nor (n329,n330,n331);
and (n330,n52,n146);
and (n331,n53,n148);
or (n332,n333,n93);
nor (n333,n334,n335);
and (n334,n52,n194);
and (n335,n53,n196);
nand (n336,n337,n341);
or (n337,n47,n338);
nor (n338,n339,n340);
and (n339,n60,n173);
and (n340,n58,n172);
or (n341,n342,n67);
nor (n342,n343,n344);
and (n343,n60,n129);
and (n344,n58,n128);
and (n345,n319,n327);
xor (n346,n286,n294);
xor (n347,n348,n355);
xor (n348,n349,n352);
nand (n349,n350,n351);
or (n350,n92,n333);
or (n351,n93,n238);
nand (n352,n353,n354);
or (n353,n47,n342);
or (n354,n279,n67);
and (n355,n356,n363);
nor (n356,n357,n130);
nor (n357,n358,n361);
and (n358,n359,n60);
not (n359,n360);
and (n360,n39,n136);
and (n361,n38,n362);
not (n362,n136);
nand (n363,n364,n369);
or (n364,n365,n181);
not (n365,n366);
nor (n366,n367,n368);
and (n367,n65,n179);
and (n368,n63,n98);
or (n369,n291,n182);
or (n370,n371,n394);
and (n371,n372,n393);
xor (n372,n373,n374);
xor (n373,n356,n363);
or (n374,n375,n392);
and (n375,n376,n385);
xor (n376,n377,n378);
and (n377,n139,n39);
nand (n378,n379,n384);
or (n379,n181,n380);
not (n380,n381);
nor (n381,n382,n383);
and (n382,n194,n98);
and (n383,n196,n179);
nand (n384,n366,n183);
nand (n385,n386,n391);
or (n386,n92,n387);
not (n387,n388);
nor (n388,n389,n390);
and (n389,n128,n52);
and (n390,n129,n53);
or (n391,n93,n329);
and (n392,n377,n378);
xor (n393,n318,n336);
and (n394,n373,n374);
not (n395,n396);
nor (n396,n397,n404);
xor (n397,n398,n403);
xor (n398,n399,n400);
xor (n399,n244,n259);
or (n400,n401,n402);
and (n401,n348,n355);
and (n402,n349,n352);
xor (n403,n276,n284);
or (n404,n405,n406);
and (n405,n315,n347);
and (n406,n316,n346);
or (n407,n408,n540);
and (n408,n409,n437);
xor (n409,n410,n436);
or (n410,n411,n435);
and (n411,n412,n434);
xor (n412,n413,n420);
nand (n413,n414,n419);
or (n414,n47,n415);
not (n415,n416);
nor (n416,n417,n418);
and (n417,n24,n58);
and (n418,n23,n60);
or (n419,n338,n67);
and (n420,n421,n427);
nor (n421,n422,n60);
nor (n422,n423,n426);
and (n423,n424,n52);
not (n424,n425);
and (n425,n39,n51);
and (n426,n38,n57);
nand (n427,n428,n429);
or (n428,n182,n380);
nand (n429,n430,n433);
nand (n430,n431,n432);
or (n431,n146,n179);
nand (n432,n179,n146);
not (n433,n181);
xor (n434,n376,n385);
and (n435,n413,n420);
xor (n436,n372,n393);
or (n437,n438,n539);
and (n438,n439,n458);
xor (n439,n440,n457);
or (n440,n441,n456);
and (n441,n442,n455);
xor (n442,n443,n448);
nand (n443,n444,n447);
or (n444,n445,n92);
not (n445,n446);
xor (n446,n172,n52);
nand (n447,n94,n388);
nand (n448,n449,n454);
or (n449,n450,n47);
not (n450,n451);
nand (n451,n452,n453);
or (n452,n60,n39);
or (n453,n38,n58);
nand (n454,n416,n49);
xor (n455,n421,n427);
and (n456,n443,n448);
xor (n457,n412,n434);
or (n458,n459,n538);
and (n459,n460,n482);
xor (n460,n461,n481);
or (n461,n462,n480);
and (n462,n463,n472);
xor (n463,n464,n465);
and (n464,n49,n39);
nand (n465,n466,n471);
or (n466,n467,n92);
not (n467,n468);
nor (n468,n469,n470);
and (n469,n23,n52);
and (n470,n24,n53);
nand (n471,n94,n446);
nand (n472,n473,n478);
or (n473,n181,n474);
not (n474,n475);
nand (n475,n476,n477);
or (n476,n129,n179);
nand (n477,n179,n129);
or (n478,n479,n182);
not (n479,n430);
and (n480,n464,n465);
xor (n481,n442,n455);
nand (n482,n483,n537);
or (n483,n484,n499);
nor (n484,n485,n486);
xor (n485,n463,n472);
nor (n486,n487,n494);
not (n487,n488);
nand (n488,n489,n493);
or (n489,n181,n490);
nor (n490,n491,n492);
and (n491,n172,n98);
and (n492,n173,n179);
nand (n493,n475,n183);
nand (n494,n495,n53);
nand (n495,n496,n498);
or (n496,n497,n98);
and (n497,n39,n97);
or (n498,n39,n97);
nor (n499,n500,n536);
and (n500,n501,n512);
nand (n501,n502,n506);
nor (n502,n503,n504);
and (n503,n494,n488);
and (n504,n505,n487);
not (n505,n494);
nor (n506,n507,n511);
and (n507,n241,n508);
nand (n508,n509,n510);
or (n509,n52,n39);
or (n510,n38,n53);
and (n511,n94,n468);
nand (n512,n513,n535);
or (n513,n514,n529);
not (n514,n515);
nor (n515,n516,n527);
not (n516,n517);
nand (n517,n518,n523);
or (n518,n182,n519);
not (n519,n520);
nor (n520,n521,n522);
and (n521,n23,n179);
and (n522,n24,n98);
nand (n523,n524,n433);
nor (n524,n525,n526);
and (n525,n38,n179);
and (n526,n39,n98);
nand (n527,n528,n98);
nand (n528,n39,n183);
not (n529,n530);
nand (n530,n531,n534);
nor (n531,n532,n533);
nor (n532,n519,n181);
nor (n533,n490,n182);
nand (n534,n39,n94);
or (n535,n531,n534);
nor (n536,n506,n502);
nand (n537,n485,n486);
and (n538,n461,n481);
and (n539,n440,n457);
and (n540,n410,n436);
nand (n541,n542,n544);
or (n542,n396,n543);
nand (n543,n314,n370);
nand (n544,n397,n404);
not (n545,n546);
or (n546,n547,n548);
xor (n547,n272,n302);
or (n548,n549,n550);
and (n549,n398,n403);
and (n550,n399,n400);
nand (n551,n547,n548);
or (n552,n306,n10);
not (n553,n554);
nand (n554,n555,n3);
not (n555,n4);
wire s0n556,s1n556,notn556;
or (n556,s0n556,s1n556);
not(notn556,n4);
and (s0n556,notn556,n557);
and (s1n556,n4,1'b0);
wire s0n557,s1n557,notn557;
or (n557,s0n557,s1n557);
not(notn557,n3);
and (s0n557,notn557,n5);
and (s1n557,n3,n558);
xor (n558,n559,n874);
xor (n559,n560,n872);
xor (n560,n561,n871);
xor (n561,n562,n863);
xor (n562,n563,n862);
xor (n563,n564,n848);
xor (n564,n565,n847);
xor (n565,n566,n828);
xor (n566,n567,n827);
xor (n567,n568,n801);
xor (n568,n569,n800);
xor (n569,n570,n768);
xor (n570,n571,n767);
xor (n571,n572,n729);
xor (n572,n573,n728);
xor (n573,n574,n685);
xor (n574,n575,n684);
xor (n575,n576,n634);
xor (n576,n577,n633);
xor (n577,n578,n581);
xor (n578,n579,n580);
and (n579,n222,n183);
and (n580,n187,n98);
or (n581,n582,n585);
and (n582,n583,n584);
and (n583,n187,n183);
and (n584,n107,n98);
and (n585,n586,n587);
xor (n586,n583,n584);
or (n587,n588,n590);
and (n588,n589,n264);
and (n589,n107,n183);
and (n590,n591,n592);
xor (n591,n589,n264);
or (n592,n593,n596);
and (n593,n594,n595);
and (n594,n90,n183);
and (n595,n70,n98);
and (n596,n597,n598);
xor (n597,n594,n595);
or (n598,n599,n601);
and (n599,n600,n368);
and (n600,n70,n183);
and (n601,n602,n603);
xor (n602,n600,n368);
or (n603,n604,n606);
and (n604,n605,n382);
and (n605,n63,n183);
and (n606,n607,n608);
xor (n607,n605,n382);
or (n608,n609,n612);
and (n609,n610,n611);
and (n610,n194,n183);
and (n611,n146,n98);
and (n612,n613,n614);
xor (n613,n610,n611);
or (n614,n615,n618);
and (n615,n616,n617);
and (n616,n146,n183);
and (n617,n129,n98);
and (n618,n619,n620);
xor (n619,n616,n617);
or (n620,n621,n624);
and (n621,n622,n623);
and (n622,n129,n183);
and (n623,n173,n98);
and (n624,n625,n626);
xor (n625,n622,n623);
or (n626,n627,n629);
and (n627,n628,n522);
and (n628,n173,n183);
and (n629,n630,n631);
xor (n630,n628,n522);
and (n631,n632,n526);
and (n632,n24,n183);
and (n633,n107,n97);
or (n634,n635,n638);
and (n635,n636,n637);
xor (n636,n586,n587);
and (n637,n90,n97);
and (n638,n639,n640);
xor (n639,n636,n637);
or (n640,n641,n644);
and (n641,n642,n643);
xor (n642,n591,n592);
and (n643,n70,n97);
and (n644,n645,n646);
xor (n645,n642,n643);
or (n646,n647,n650);
and (n647,n648,n649);
xor (n648,n597,n598);
and (n649,n63,n97);
and (n650,n651,n652);
xor (n651,n648,n649);
or (n652,n653,n656);
and (n653,n654,n655);
xor (n654,n602,n603);
and (n655,n194,n97);
and (n656,n657,n658);
xor (n657,n654,n655);
or (n658,n659,n662);
and (n659,n660,n661);
xor (n660,n607,n608);
and (n661,n146,n97);
and (n662,n663,n664);
xor (n663,n660,n661);
or (n664,n665,n668);
and (n665,n666,n667);
xor (n666,n613,n614);
and (n667,n129,n97);
and (n668,n669,n670);
xor (n669,n666,n667);
or (n670,n671,n674);
and (n671,n672,n673);
xor (n672,n619,n620);
and (n673,n173,n97);
and (n674,n675,n676);
xor (n675,n672,n673);
or (n676,n677,n680);
and (n677,n678,n679);
xor (n678,n625,n626);
and (n679,n24,n97);
and (n680,n681,n682);
xor (n681,n678,n679);
and (n682,n683,n497);
xor (n683,n630,n631);
and (n684,n90,n53);
or (n685,n686,n689);
and (n686,n687,n688);
xor (n687,n639,n640);
and (n688,n70,n53);
and (n689,n690,n691);
xor (n690,n687,n688);
or (n691,n692,n695);
and (n692,n693,n694);
xor (n693,n645,n646);
and (n694,n63,n53);
and (n695,n696,n697);
xor (n696,n693,n694);
or (n697,n698,n701);
and (n698,n699,n700);
xor (n699,n651,n652);
and (n700,n194,n53);
and (n701,n702,n703);
xor (n702,n699,n700);
or (n703,n704,n707);
and (n704,n705,n706);
xor (n705,n657,n658);
and (n706,n146,n53);
and (n707,n708,n709);
xor (n708,n705,n706);
or (n709,n710,n712);
and (n710,n711,n390);
xor (n711,n663,n664);
and (n712,n713,n714);
xor (n713,n711,n390);
or (n714,n715,n718);
and (n715,n716,n717);
xor (n716,n669,n670);
and (n717,n173,n53);
and (n718,n719,n720);
xor (n719,n716,n717);
or (n720,n721,n723);
and (n721,n722,n470);
xor (n722,n675,n676);
and (n723,n724,n725);
xor (n724,n722,n470);
and (n725,n726,n727);
xor (n726,n681,n682);
and (n727,n39,n53);
and (n728,n70,n51);
or (n729,n730,n733);
and (n730,n731,n732);
xor (n731,n690,n691);
and (n732,n63,n51);
and (n733,n734,n735);
xor (n734,n731,n732);
or (n735,n736,n739);
and (n736,n737,n738);
xor (n737,n696,n697);
and (n738,n194,n51);
and (n739,n740,n741);
xor (n740,n737,n738);
or (n741,n742,n745);
and (n742,n743,n744);
xor (n743,n702,n703);
and (n744,n146,n51);
and (n745,n746,n747);
xor (n746,n743,n744);
or (n747,n748,n751);
and (n748,n749,n750);
xor (n749,n708,n709);
and (n750,n129,n51);
and (n751,n752,n753);
xor (n752,n749,n750);
or (n753,n754,n757);
and (n754,n755,n756);
xor (n755,n713,n714);
and (n756,n173,n51);
and (n757,n758,n759);
xor (n758,n755,n756);
or (n759,n760,n763);
and (n760,n761,n762);
xor (n761,n719,n720);
and (n762,n24,n51);
and (n763,n764,n765);
xor (n764,n761,n762);
and (n765,n766,n425);
xor (n766,n724,n725);
and (n767,n63,n58);
or (n768,n769,n772);
and (n769,n770,n771);
xor (n770,n734,n735);
and (n771,n194,n58);
and (n772,n773,n774);
xor (n773,n770,n771);
or (n774,n775,n778);
and (n775,n776,n777);
xor (n776,n740,n741);
and (n777,n146,n58);
and (n778,n779,n780);
xor (n779,n776,n777);
or (n780,n781,n784);
and (n781,n782,n783);
xor (n782,n746,n747);
and (n783,n129,n58);
and (n784,n785,n786);
xor (n785,n782,n783);
or (n786,n787,n790);
and (n787,n788,n789);
xor (n788,n752,n753);
and (n789,n173,n58);
and (n790,n791,n792);
xor (n791,n788,n789);
or (n792,n793,n795);
and (n793,n794,n417);
xor (n794,n758,n759);
and (n795,n796,n797);
xor (n796,n794,n417);
and (n797,n798,n799);
xor (n798,n764,n765);
and (n799,n39,n58);
and (n800,n194,n136);
or (n801,n802,n805);
and (n802,n803,n804);
xor (n803,n773,n774);
and (n804,n146,n136);
and (n805,n806,n807);
xor (n806,n803,n804);
or (n807,n808,n811);
and (n808,n809,n810);
xor (n809,n779,n780);
and (n810,n129,n136);
and (n811,n812,n813);
xor (n812,n809,n810);
or (n813,n814,n817);
and (n814,n815,n816);
xor (n815,n785,n786);
and (n816,n173,n136);
and (n817,n818,n819);
xor (n818,n815,n816);
or (n819,n820,n823);
and (n820,n821,n822);
xor (n821,n791,n792);
and (n822,n24,n136);
and (n823,n824,n825);
xor (n824,n821,n822);
and (n825,n826,n360);
xor (n826,n796,n797);
and (n827,n146,n131);
or (n828,n829,n831);
and (n829,n830,n132);
xor (n830,n806,n807);
and (n831,n832,n833);
xor (n832,n830,n132);
or (n833,n834,n836);
and (n834,n835,n249);
xor (n835,n812,n813);
and (n836,n837,n838);
xor (n837,n835,n249);
or (n838,n839,n842);
and (n839,n840,n841);
xor (n840,n818,n819);
and (n841,n24,n131);
and (n842,n843,n844);
xor (n843,n840,n841);
and (n844,n845,n846);
xor (n845,n824,n825);
and (n846,n39,n131);
and (n847,n129,n163);
or (n848,n849,n852);
and (n849,n850,n851);
xor (n850,n832,n833);
and (n851,n173,n163);
and (n852,n853,n854);
xor (n853,n850,n851);
or (n854,n855,n858);
and (n855,n856,n857);
xor (n856,n837,n838);
and (n857,n24,n163);
and (n858,n859,n860);
xor (n859,n856,n857);
and (n860,n861,n233);
xor (n861,n843,n844);
and (n862,n173,n32);
or (n863,n864,n866);
and (n864,n865,n158);
xor (n865,n853,n854);
and (n866,n867,n868);
xor (n867,n865,n158);
and (n868,n869,n870);
xor (n869,n859,n860);
and (n870,n39,n32);
and (n871,n24,n31);
and (n872,n873,n81);
xor (n873,n867,n868);
and (n874,n39,n22);
endmodule
