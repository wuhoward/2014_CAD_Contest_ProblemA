module top (out,n6,n23,n24,n27,n28,n35,n36,n38,n39
        ,n56,n74,n75,n77,n78,n97,n137,n143,n152,n161
        ,n162,n168,n169,n174,n181,n187,n200,n201,n205,n210
        ,n228,n271,n352,n402,n601,n1022);
output out;
input n6;
input n23;
input n24;
input n27;
input n28;
input n35;
input n36;
input n38;
input n39;
input n56;
input n74;
input n75;
input n77;
input n78;
input n97;
input n137;
input n143;
input n152;
input n161;
input n162;
input n168;
input n169;
input n174;
input n181;
input n187;
input n200;
input n201;
input n205;
input n210;
input n228;
input n271;
input n352;
input n402;
input n601;
input n1022;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n25;
wire n26;
wire n29;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n37;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n55;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n76;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n170;
wire n171;
wire n172;
wire n173;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n202;
wire n203;
wire n204;
wire n206;
wire n207;
wire n208;
wire n209;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
xor (out,n0,n1024);
nor (n0,n1,n1023);
not (n1,n2);
nand (n2,n3,n1022);
nand (n3,n4,n1020);
or (n4,n5,n7);
not (n5,n6);
not (n7,n8);
nand (n8,n9,n1019);
or (n9,n10,n114);
not (n10,n11);
nor (n11,n12,n113);
and (n12,n13,n101);
not (n13,n14);
or (n14,n15,n100);
and (n15,n16,n62);
xor (n16,n17,n51);
nand (n17,n18,n42);
or (n18,n19,n31);
not (n19,n20);
nand (n20,n21,n29);
or (n21,n22,n25);
wire s0n22,s1n22,notn22;
or (n22,s0n22,s1n22);
not(notn22,n6);
and (s0n22,notn22,n23);
and (s1n22,n6,n24);
not (n25,n26);
and (n26,n27,n28);
or (n29,n30,n26);
not (n30,n22);
nor (n31,n32,n40);
and (n32,n33,n37);
not (n33,n34);
wire s0n34,s1n34,notn34;
or (n34,s0n34,s1n34);
not(notn34,n6);
and (s0n34,notn34,n35);
and (s1n34,n6,n36);
wire s0n37,s1n37,notn37;
or (n37,s0n37,s1n37);
not(notn37,n6);
and (s0n37,notn37,n38);
and (s1n37,n6,n39);
and (n40,n34,n41);
not (n41,n37);
or (n42,n43,n47);
nand (n43,n31,n44);
nand (n44,n45,n46);
or (n45,n33,n22);
nand (n46,n22,n33);
nor (n47,n48,n49);
and (n48,n30,n28);
and (n49,n22,n50);
not (n50,n28);
nand (n51,n52,n57,n59);
or (n52,n53,n56);
wire s0n53,s1n53,notn53;
or (n53,s0n53,s1n53);
not(notn53,n6);
and (s0n53,notn53,1'b0);
and (s1n53,n6,n55);
and (n55,n27,n24);
not (n57,n58);
and (n58,n56,n53);
not (n59,n60);
nand (n60,n22,n61);
not (n61,n53);
or (n62,n63,n99);
and (n63,n64,n93);
xor (n64,n65,n86);
nand (n65,n66,n83);
or (n66,n67,n70);
not (n67,n68);
nand (n68,n69,n80);
not (n69,n70);
nand (n70,n71,n79);
or (n71,n72,n76);
not (n72,n73);
wire s0n73,s1n73,notn73;
or (n73,s0n73,s1n73);
not(notn73,n6);
and (s0n73,notn73,n74);
and (s1n73,n6,n75);
wire s0n76,s1n76,notn76;
or (n76,s0n76,s1n76);
not(notn76,n6);
and (s0n76,notn76,n77);
and (s1n76,n6,n78);
nand (n79,n76,n72);
nand (n80,n81,n82);
or (n81,n72,n37);
nand (n82,n37,n72);
nand (n83,n84,n85);
or (n84,n37,n25);
or (n85,n41,n26);
nand (n86,n87,n92);
or (n87,n43,n88);
nor (n88,n89,n90);
and (n89,n30,n56);
and (n90,n22,n91);
not (n91,n56);
or (n92,n31,n47);
nor (n93,n60,n94);
nor (n94,n95,n98);
and (n95,n53,n96);
not (n96,n97);
and (n98,n61,n97);
and (n99,n65,n86);
and (n100,n17,n51);
not (n101,n102);
xor (n102,n103,n112);
xor (n103,n104,n108);
nand (n104,n105,n20);
or (n105,n106,n107);
not (n106,n43);
not (n107,n31);
nor (n108,n60,n109);
nor (n109,n110,n111);
and (n110,n53,n50);
and (n111,n61,n28);
not (n112,n51);
and (n113,n14,n102);
nand (n114,n115,n995,n1018);
nand (n115,n116,n772);
nand (n116,n117,n761,n771);
nand (n117,n118,n564);
nand (n118,n119,n420,n563);
nand (n119,n120,n371);
nand (n120,n121,n370);
or (n121,n122,n323);
nor (n122,n123,n322);
and (n123,n124,n294);
not (n124,n125);
nor (n125,n126,n252);
or (n126,n127,n251);
and (n127,n128,n220);
xor (n128,n129,n191);
or (n129,n130,n190);
and (n130,n131,n177);
xor (n131,n132,n146);
nand (n132,n133,n140);
or (n133,n134,n43);
not (n134,n135);
nand (n135,n136,n138);
or (n136,n30,n137);
or (n138,n22,n139);
not (n139,n137);
or (n140,n31,n141);
nor (n141,n142,n144);
and (n142,n143,n30);
and (n144,n145,n22);
not (n145,n143);
nand (n146,n147,n171);
or (n147,n148,n155);
not (n148,n149);
nand (n149,n150,n153);
or (n150,n76,n151);
not (n151,n152);
or (n153,n154,n152);
not (n154,n76);
not (n155,n156);
and (n156,n157,n164);
nand (n157,n158,n163);
or (n158,n159,n76);
not (n159,n160);
wire s0n160,s1n160,notn160;
or (n160,s0n160,s1n160);
not(notn160,n6);
and (s0n160,notn160,n161);
and (s1n160,n6,n162);
nand (n163,n76,n159);
not (n164,n165);
nand (n165,n166,n170);
or (n166,n159,n167);
wire s0n167,s1n167,notn167;
or (n167,s0n167,s1n167);
not(notn167,n6);
and (s0n167,notn167,n168);
and (s1n167,n6,n169);
nand (n170,n167,n159);
nand (n171,n165,n172);
nor (n172,n173,n175);
and (n173,n174,n76);
and (n175,n176,n154);
not (n176,n174);
nand (n177,n178,n184);
or (n178,n68,n179);
nor (n179,n180,n182);
and (n180,n41,n181);
and (n182,n37,n183);
not (n183,n181);
or (n184,n69,n185);
nor (n185,n186,n188);
and (n186,n41,n187);
and (n188,n37,n189);
not (n189,n187);
and (n190,n132,n146);
xor (n191,n192,n214);
xor (n192,n193,n194);
and (n193,n59,n137);
nand (n194,n195,n207);
or (n195,n196,n202);
not (n196,n197);
nor (n197,n198,n199);
not (n198,n167);
wire s0n199,s1n199,notn199;
or (n199,s0n199,s1n199);
not(notn199,n6);
and (s0n199,notn199,n200);
and (s1n199,n6,n201);
nor (n202,n203,n206);
and (n203,n204,n167);
not (n204,n205);
and (n206,n205,n198);
or (n207,n208,n213);
nor (n208,n209,n211);
and (n209,n198,n210);
and (n211,n167,n212);
not (n212,n210);
not (n213,n199);
nand (n214,n215,n216);
or (n215,n43,n141);
or (n216,n31,n217);
nor (n217,n218,n219);
and (n218,n181,n30);
and (n219,n183,n22);
xor (n220,n221,n237);
xor (n221,n222,n231);
nand (n222,n223,n225);
or (n223,n155,n224);
not (n224,n172);
or (n225,n164,n226);
nor (n226,n227,n229);
and (n227,n154,n228);
and (n229,n76,n230);
not (n230,n228);
nand (n231,n232,n233);
or (n232,n68,n185);
or (n233,n69,n234);
nor (n234,n235,n236);
and (n235,n41,n152);
and (n236,n37,n151);
and (n237,n238,n243);
nor (n238,n239,n30);
nor (n239,n240,n242);
and (n240,n41,n241);
nand (n241,n34,n137);
and (n242,n33,n139);
nand (n243,n244,n249);
or (n244,n245,n196);
not (n245,n246);
nor (n246,n247,n248);
and (n247,n228,n167);
and (n248,n230,n198);
nand (n249,n250,n199);
not (n250,n202);
and (n251,n129,n191);
xor (n252,n253,n277);
xor (n253,n254,n274);
xor (n254,n255,n266);
xor (n255,n256,n262);
nand (n256,n257,n258);
or (n257,n217,n43);
nand (n258,n259,n107);
nor (n259,n260,n261);
and (n260,n187,n22);
and (n261,n189,n30);
nor (n262,n60,n263);
nor (n263,n264,n265);
and (n264,n53,n145);
and (n265,n61,n143);
nand (n266,n267,n268);
or (n267,n196,n208);
or (n268,n269,n213);
nor (n269,n270,n272);
and (n270,n198,n271);
and (n272,n167,n273);
not (n273,n271);
or (n274,n275,n276);
and (n275,n221,n237);
and (n276,n222,n231);
xor (n277,n278,n291);
xor (n278,n279,n285);
nand (n279,n280,n281);
or (n280,n68,n234);
or (n281,n69,n282);
nor (n282,n283,n284);
and (n283,n41,n174);
and (n284,n37,n176);
nand (n285,n286,n287);
or (n286,n155,n226);
or (n287,n288,n164);
nor (n288,n289,n290);
and (n289,n154,n205);
and (n290,n76,n204);
or (n291,n292,n293);
and (n292,n192,n214);
and (n293,n193,n194);
not (n294,n295);
nand (n295,n296,n297);
xor (n296,n128,n220);
or (n297,n298,n321);
and (n298,n299,n320);
xor (n299,n300,n301);
xor (n300,n238,n243);
or (n301,n302,n319);
and (n302,n303,n312);
xor (n303,n304,n305);
and (n304,n107,n137);
nand (n305,n306,n307);
or (n306,n213,n245);
nand (n307,n308,n197);
not (n308,n309);
nor (n309,n310,n311);
and (n310,n174,n198);
and (n311,n176,n167);
nand (n312,n313,n318);
or (n313,n314,n155);
not (n314,n315);
nor (n315,n316,n317);
and (n316,n187,n76);
and (n317,n154,n189);
nand (n318,n165,n149);
and (n319,n304,n305);
xor (n320,n131,n177);
and (n321,n300,n301);
and (n322,n126,n252);
nor (n323,n324,n367);
xor (n324,n325,n364);
xor (n325,n326,n345);
xor (n326,n327,n339);
xor (n327,n328,n335);
nand (n328,n329,n331);
or (n329,n330,n43);
not (n330,n259);
nand (n331,n107,n332);
nor (n332,n333,n334);
and (n333,n152,n22);
and (n334,n151,n30);
nor (n335,n60,n336);
nor (n336,n337,n338);
and (n337,n53,n183);
and (n338,n61,n181);
nand (n339,n340,n341);
or (n340,n68,n282);
or (n341,n69,n342);
nor (n342,n343,n344);
and (n343,n41,n228);
and (n344,n37,n230);
xor (n345,n346,n361);
xor (n346,n347,n355);
nand (n347,n348,n349);
or (n348,n196,n269);
or (n349,n350,n213);
nor (n350,n351,n353);
and (n351,n198,n352);
and (n353,n167,n354);
not (n354,n352);
nand (n355,n356,n357);
or (n356,n155,n288);
or (n357,n358,n164);
nor (n358,n359,n360);
and (n359,n154,n210);
and (n360,n76,n212);
or (n361,n362,n363);
and (n362,n255,n266);
and (n363,n256,n262);
or (n364,n365,n366);
and (n365,n278,n291);
and (n366,n279,n285);
or (n367,n368,n369);
and (n368,n253,n277);
and (n369,n254,n274);
nand (n370,n324,n367);
nand (n371,n372,n416);
not (n372,n373);
xor (n373,n374,n415);
xor (n374,n375,n394);
xor (n375,n376,n388);
xor (n376,n377,n384);
nand (n377,n378,n380);
or (n378,n379,n43);
not (n379,n332);
nand (n380,n107,n381);
nor (n381,n382,n383);
and (n382,n174,n22);
and (n383,n176,n30);
nor (n384,n60,n385);
nor (n385,n386,n387);
and (n386,n53,n189);
and (n387,n61,n187);
nand (n388,n389,n390);
or (n389,n68,n342);
or (n390,n69,n391);
nor (n391,n392,n393);
and (n392,n41,n205);
and (n393,n37,n204);
xor (n394,n395,n412);
xor (n395,n396,n411);
xor (n396,n397,n405);
nand (n397,n398,n399);
or (n398,n196,n350);
or (n399,n400,n213);
nor (n400,n401,n403);
and (n401,n198,n402);
and (n403,n167,n404);
not (n404,n402);
nand (n405,n406,n407);
or (n406,n155,n358);
or (n407,n164,n408);
nor (n408,n409,n410);
and (n409,n154,n271);
and (n410,n76,n273);
and (n411,n347,n355);
or (n412,n413,n414);
and (n413,n327,n339);
and (n414,n328,n335);
and (n415,n346,n361);
not (n416,n417);
or (n417,n418,n419);
and (n418,n325,n364);
and (n419,n326,n345);
nand (n420,n371,n421,n562);
nor (n421,n422,n559);
nor (n422,n423,n557);
and (n423,n424,n552);
or (n424,n425,n551);
and (n425,n426,n467);
xor (n426,n427,n460);
or (n427,n428,n459);
and (n428,n429,n447);
xor (n429,n430,n437);
nand (n430,n431,n436);
or (n431,n432,n155);
not (n432,n433);
nor (n433,n434,n435);
and (n434,n183,n154);
and (n435,n181,n76);
nand (n436,n165,n315);
nand (n437,n438,n443);
or (n438,n439,n69);
not (n439,n440);
nor (n440,n441,n442);
and (n441,n143,n37);
and (n442,n145,n41);
nand (n443,n67,n444);
nand (n444,n445,n446);
or (n445,n41,n137);
or (n446,n37,n139);
xor (n447,n448,n453);
and (n448,n449,n37);
nand (n449,n450,n452);
or (n450,n76,n451);
and (n451,n137,n73);
or (n452,n73,n137);
nand (n453,n454,n458);
or (n454,n196,n455);
nor (n455,n456,n457);
and (n456,n198,n152);
and (n457,n167,n151);
or (n458,n309,n213);
and (n459,n430,n437);
xor (n460,n461,n466);
xor (n461,n462,n465);
nand (n462,n463,n464);
or (n463,n439,n68);
or (n464,n69,n179);
and (n465,n448,n453);
xor (n466,n303,n312);
or (n467,n468,n550);
and (n468,n469,n490);
xor (n469,n470,n489);
or (n470,n471,n488);
and (n471,n472,n481);
xor (n472,n473,n474);
and (n473,n70,n137);
nand (n474,n475,n480);
or (n475,n476,n155);
not (n476,n477);
nor (n477,n478,n479);
and (n478,n143,n76);
and (n479,n145,n154);
nand (n480,n433,n165);
nand (n481,n482,n487);
or (n482,n196,n483);
not (n483,n484);
nor (n484,n485,n486);
and (n485,n189,n198);
and (n486,n187,n167);
or (n487,n455,n213);
and (n488,n473,n474);
xor (n489,n429,n447);
or (n490,n491,n549);
and (n491,n492,n548);
xor (n492,n493,n507);
nor (n493,n494,n502);
not (n494,n495);
nand (n495,n496,n501);
or (n496,n497,n196);
not (n497,n498);
nand (n498,n499,n500);
or (n499,n183,n167);
nand (n500,n167,n183);
nand (n501,n484,n199);
nand (n502,n503,n76);
nand (n503,n504,n506);
or (n504,n167,n505);
and (n505,n137,n160);
or (n506,n160,n137);
nand (n507,n508,n546);
or (n508,n509,n532);
not (n509,n510);
nand (n510,n511,n531);
or (n511,n512,n521);
nor (n512,n513,n520);
nand (n513,n514,n519);
or (n514,n515,n196);
not (n515,n516);
nand (n516,n517,n518);
or (n517,n145,n167);
nand (n518,n167,n145);
nand (n519,n498,n199);
nor (n520,n164,n139);
nand (n521,n522,n529);
nand (n522,n523,n528);
or (n523,n524,n196);
not (n524,n525);
nand (n525,n526,n527);
or (n526,n198,n137);
or (n527,n167,n139);
nand (n528,n516,n199);
nor (n529,n530,n198);
and (n530,n137,n199);
nand (n531,n513,n520);
not (n532,n533);
nand (n533,n534,n542);
not (n534,n535);
nand (n535,n536,n541);
or (n536,n537,n155);
not (n537,n538);
nand (n538,n539,n540);
or (n539,n154,n137);
or (n540,n76,n139);
nand (n541,n165,n477);
nor (n542,n543,n545);
and (n543,n494,n544);
not (n544,n502);
and (n545,n495,n502);
nand (n546,n547,n535);
not (n547,n542);
xor (n548,n472,n481);
and (n549,n493,n507);
and (n550,n470,n489);
and (n551,n427,n460);
or (n552,n553,n554);
xor (n553,n299,n320);
or (n554,n555,n556);
and (n555,n461,n466);
and (n556,n462,n465);
not (n557,n558);
nand (n558,n553,n554);
nand (n559,n560,n124);
not (n560,n561);
nor (n561,n296,n297);
not (n562,n323);
nand (n563,n373,n417);
nor (n564,n565,n665);
nand (n565,n566,n658);
not (n566,n567);
nor (n567,n568,n649);
xor (n568,n569,n640);
xor (n569,n570,n594);
xor (n570,n571,n585);
xor (n571,n572,n581);
nand (n572,n573,n577);
or (n573,n43,n574);
nor (n574,n575,n576);
and (n575,n30,n228);
and (n576,n22,n230);
or (n577,n31,n578);
nor (n578,n579,n580);
and (n579,n205,n30);
and (n580,n204,n22);
nor (n581,n60,n582);
nor (n582,n583,n584);
and (n583,n53,n176);
and (n584,n61,n174);
nand (n585,n586,n590);
or (n586,n587,n69);
nor (n587,n588,n589);
and (n588,n41,n271);
and (n589,n37,n273);
or (n590,n68,n591);
nor (n591,n592,n593);
and (n592,n41,n210);
and (n593,n37,n212);
xor (n594,n595,n624);
xor (n595,n596,n617);
xor (n596,n597,n608);
nand (n597,n598,n604);
or (n598,n196,n599);
nor (n599,n600,n602);
and (n600,n198,n601);
and (n602,n167,n603);
not (n603,n601);
or (n604,n605,n213);
nor (n605,n606,n607);
and (n606,n198,n97);
and (n607,n167,n96);
nand (n608,n609,n613);
or (n609,n155,n610);
nor (n610,n611,n612);
and (n611,n154,n352);
and (n612,n76,n354);
or (n613,n614,n164);
nor (n614,n615,n616);
and (n615,n154,n402);
and (n616,n76,n404);
and (n617,n618,n621);
nand (n618,n619,n620);
or (n619,n196,n400);
or (n620,n599,n213);
nand (n621,n622,n623);
or (n622,n155,n408);
or (n623,n610,n164);
or (n624,n625,n639);
and (n625,n626,n636);
xor (n626,n627,n632);
nand (n627,n628,n630);
or (n628,n629,n43);
not (n629,n381);
nand (n630,n631,n107);
not (n631,n574);
nor (n632,n60,n633);
nor (n633,n634,n635);
and (n634,n53,n151);
and (n635,n61,n152);
nand (n636,n637,n638);
or (n637,n68,n391);
or (n638,n69,n591);
and (n639,n627,n632);
or (n640,n641,n648);
and (n641,n642,n645);
xor (n642,n643,n644);
xor (n643,n618,n621);
and (n644,n397,n405);
or (n645,n646,n647);
and (n646,n376,n388);
and (n647,n377,n384);
and (n648,n643,n644);
or (n649,n650,n657);
and (n650,n651,n654);
xor (n651,n652,n653);
xor (n652,n626,n636);
xor (n653,n642,n645);
or (n654,n655,n656);
and (n655,n395,n412);
and (n656,n396,n411);
and (n657,n652,n653);
nand (n658,n659,n661);
not (n659,n660);
xor (n660,n651,n654);
not (n661,n662);
or (n662,n663,n664);
and (n663,n374,n415);
and (n664,n375,n394);
nand (n665,n666,n714);
nand (n666,n667,n710);
not (n667,n668);
xor (n668,n669,n707);
xor (n669,n670,n688);
xor (n670,n671,n682);
xor (n671,n672,n678);
nand (n672,n673,n674);
or (n673,n578,n43);
nand (n674,n107,n675);
nor (n675,n676,n677);
and (n676,n210,n22);
and (n677,n212,n30);
nor (n678,n60,n679);
nor (n679,n680,n681);
and (n680,n53,n230);
and (n681,n61,n228);
nand (n682,n683,n684);
or (n683,n68,n587);
or (n684,n69,n685);
nor (n685,n686,n687);
and (n686,n41,n352);
and (n687,n37,n354);
xor (n688,n689,n704);
xor (n689,n690,n703);
xor (n690,n691,n697);
nand (n691,n692,n693);
or (n692,n196,n605);
or (n693,n694,n213);
nor (n694,n695,n696);
and (n695,n198,n56);
and (n696,n167,n91);
nand (n697,n698,n699);
or (n698,n155,n614);
or (n699,n164,n700);
nor (n700,n701,n702);
and (n701,n154,n601);
and (n702,n76,n603);
and (n703,n597,n608);
or (n704,n705,n706);
and (n705,n571,n585);
and (n706,n572,n581);
or (n707,n708,n709);
and (n708,n595,n624);
and (n709,n596,n617);
not (n710,n711);
or (n711,n712,n713);
and (n712,n569,n640);
and (n713,n570,n594);
nand (n714,n715,n757);
not (n715,n716);
xor (n716,n717,n754);
xor (n717,n718,n737);
xor (n718,n719,n731);
xor (n719,n720,n727);
nand (n720,n721,n723);
or (n721,n722,n43);
not (n722,n675);
nand (n723,n107,n724);
nor (n724,n725,n726);
and (n725,n271,n22);
and (n726,n273,n30);
nor (n727,n60,n728);
nor (n728,n729,n730);
and (n729,n53,n204);
and (n730,n61,n205);
nand (n731,n732,n733);
or (n732,n68,n685);
or (n733,n69,n734);
nor (n734,n735,n736);
and (n735,n41,n402);
and (n736,n37,n404);
xor (n737,n738,n751);
xor (n738,n739,n750);
xor (n739,n740,n746);
nand (n740,n741,n742);
or (n741,n196,n694);
or (n742,n743,n213);
nor (n743,n744,n745);
and (n744,n198,n28);
and (n745,n167,n50);
nand (n746,n747,n748);
or (n747,n155,n700);
or (n748,n749,n164);
xor (n749,n97,n154);
and (n750,n691,n697);
or (n751,n752,n753);
and (n752,n671,n682);
and (n753,n672,n678);
or (n754,n755,n756);
and (n755,n689,n704);
and (n756,n690,n703);
not (n757,n758);
or (n758,n759,n760);
and (n759,n669,n707);
and (n760,n670,n688);
nand (n761,n762,n714);
nand (n762,n763,n770);
or (n763,n764,n765);
not (n764,n666);
not (n765,n766);
nand (n766,n767,n769);
or (n767,n567,n768);
nand (n768,n660,n662);
nand (n769,n568,n649);
nand (n770,n668,n711);
nand (n771,n758,n716);
and (n772,n773,n951,n990);
and (n773,n774,n873,n945);
nor (n774,n775,n822);
nor (n775,n776,n779);
or (n776,n777,n778);
and (n777,n717,n754);
and (n778,n718,n737);
xor (n779,n780,n819);
xor (n780,n781,n800);
xor (n781,n782,n794);
xor (n782,n783,n790);
nand (n783,n784,n786);
or (n784,n785,n43);
not (n785,n724);
or (n786,n31,n787);
nor (n787,n788,n789);
and (n788,n30,n352);
and (n789,n22,n354);
nor (n790,n60,n791);
nor (n791,n792,n793);
and (n792,n53,n212);
and (n793,n61,n210);
nand (n794,n795,n796);
or (n795,n68,n734);
or (n796,n69,n797);
nor (n797,n798,n799);
and (n798,n41,n601);
and (n799,n37,n603);
xor (n800,n801,n816);
xor (n801,n802,n815);
xor (n802,n803,n809);
nand (n803,n804,n805);
or (n804,n196,n743);
or (n805,n806,n213);
nor (n806,n807,n808);
and (n807,n198,n26);
and (n808,n167,n25);
nand (n809,n810,n811);
or (n810,n749,n155);
nand (n811,n165,n812);
nand (n812,n813,n814);
or (n813,n76,n91);
or (n814,n154,n56);
and (n815,n740,n746);
or (n816,n817,n818);
and (n817,n719,n731);
and (n818,n720,n727);
or (n819,n820,n821);
and (n820,n738,n751);
and (n821,n739,n750);
not (n822,n823);
nand (n823,n824,n869);
not (n824,n825);
xor (n825,n826,n845);
xor (n826,n827,n842);
xor (n827,n828,n836);
xor (n828,n829,n833);
nor (n829,n60,n830);
nor (n830,n831,n832);
and (n831,n53,n273);
and (n832,n61,n271);
nand (n833,n834,n835);
or (n834,n199,n197);
not (n835,n806);
nand (n836,n837,n841);
or (n837,n838,n69);
nor (n838,n839,n840);
and (n839,n97,n41);
and (n840,n96,n37);
or (n841,n68,n797);
or (n842,n843,n844);
and (n843,n801,n816);
and (n844,n802,n815);
xor (n845,n846,n851);
xor (n846,n847,n848);
and (n847,n803,n809);
or (n848,n849,n850);
and (n849,n782,n794);
and (n850,n783,n790);
nand (n851,n852,n868);
or (n852,n853,n861);
not (n853,n854);
nand (n854,n855,n857);
or (n855,n155,n856);
not (n856,n812);
or (n857,n164,n858);
nor (n858,n859,n860);
and (n859,n154,n28);
and (n860,n76,n50);
not (n861,n862);
nand (n862,n863,n864);
or (n863,n43,n787);
or (n864,n31,n865);
nor (n865,n866,n867);
and (n866,n30,n402);
and (n867,n22,n404);
or (n868,n862,n854);
not (n869,n870);
or (n870,n871,n872);
and (n871,n780,n819);
and (n872,n781,n800);
nand (n873,n874,n935);
not (n874,n875);
xor (n875,n876,n927);
xor (n876,n877,n897);
xor (n877,n878,n893);
xor (n878,n879,n884);
nand (n879,n880,n881);
or (n880,n156,n165);
nand (n881,n882,n883);
or (n882,n76,n25);
or (n883,n154,n26);
nand (n884,n885,n889);
or (n885,n68,n886);
nor (n886,n887,n888);
and (n887,n41,n56);
and (n888,n37,n91);
or (n889,n69,n890);
nor (n890,n891,n892);
and (n891,n41,n28);
and (n892,n37,n50);
nor (n893,n60,n894);
nor (n894,n895,n896);
and (n895,n53,n404);
and (n896,n61,n402);
xor (n897,n898,n913);
xor (n898,n899,n908);
nand (n899,n900,n904);
or (n900,n43,n901);
nor (n901,n902,n903);
and (n902,n30,n601);
and (n903,n22,n603);
or (n904,n31,n905);
nor (n905,n906,n907);
and (n906,n30,n97);
and (n907,n22,n96);
nand (n908,n909,n911);
or (n909,n910,n164);
not (n910,n881);
nand (n911,n912,n156);
not (n912,n858);
or (n913,n914,n926);
and (n914,n915,n923);
xor (n915,n916,n920);
nor (n916,n60,n917);
nor (n917,n918,n919);
and (n918,n53,n354);
and (n919,n61,n352);
nand (n920,n921,n922);
or (n921,n68,n838);
or (n922,n69,n886);
nand (n923,n924,n925);
or (n924,n43,n865);
or (n925,n31,n901);
and (n926,n916,n920);
or (n927,n928,n934);
and (n928,n929,n931);
xor (n929,n930,n868);
not (n930,n908);
or (n931,n932,n933);
and (n932,n828,n836);
and (n933,n829,n833);
and (n934,n930,n868);
not (n935,n936);
or (n936,n937,n944);
and (n937,n938,n941);
xor (n938,n939,n940);
xor (n939,n915,n923);
xor (n940,n929,n931);
or (n941,n942,n943);
and (n942,n846,n851);
and (n943,n847,n848);
and (n944,n939,n940);
not (n945,n946);
nor (n946,n947,n948);
xor (n947,n938,n941);
or (n948,n949,n950);
and (n949,n826,n845);
and (n950,n827,n842);
nor (n951,n952,n977);
nor (n952,n953,n956);
or (n953,n954,n955);
and (n954,n876,n927);
and (n955,n877,n897);
xor (n956,n957,n974);
xor (n957,n958,n961);
or (n958,n959,n960);
and (n959,n878,n893);
and (n960,n879,n884);
xor (n961,n962,n970);
xor (n962,n963,n966);
nand (n963,n964,n965);
or (n964,n43,n905);
or (n965,n31,n88);
nor (n966,n60,n967);
nor (n967,n968,n969);
and (n968,n53,n603);
and (n969,n61,n601);
nor (n970,n971,n973);
and (n971,n67,n972);
not (n972,n890);
and (n973,n70,n83);
or (n974,n975,n976);
and (n975,n898,n913);
and (n976,n899,n908);
and (n977,n978,n982);
not (n978,n979);
or (n979,n980,n981);
and (n980,n957,n974);
and (n981,n958,n961);
not (n982,n983);
xor (n983,n984,n987);
xor (n984,n985,n986);
not (n985,n970);
xor (n986,n64,n93);
or (n987,n988,n989);
and (n988,n962,n970);
and (n989,n963,n966);
or (n990,n991,n994);
or (n991,n992,n993);
and (n992,n984,n987);
and (n993,n985,n986);
xor (n994,n16,n62);
nand (n995,n996,n990);
nand (n996,n997,n1012);
or (n997,n998,n999);
not (n998,n951);
not (n999,n1000);
nand (n1000,n1001,n1011);
or (n1001,n1002,n1003);
not (n1002,n873);
not (n1003,n1004);
nand (n1004,n1005,n1010);
or (n1005,n1006,n946);
nor (n1006,n1007,n1009);
and (n1007,n1008,n823);
and (n1008,n776,n779);
nor (n1009,n824,n869);
nand (n1010,n947,n948);
or (n1011,n874,n935);
nor (n1012,n1013,n1017);
and (n1013,n1014,n1016);
not (n1014,n1015);
nand (n1015,n953,n956);
not (n1016,n977);
nor (n1017,n978,n982);
nand (n1018,n991,n994);
nand (n1019,n10,n114);
not (n1020,n1021);
and (n1021,n8,n5,n27);
nor (n1023,n3,n1022);
xor (n1024,n1022,n1025);
wire s0n1025,s1n1025,notn1025;
or (n1025,s0n1025,s1n1025);
not(notn1025,n6);
and (s0n1025,notn1025,n1026);
and (s1n1025,n6,n1027);
and (n1026,n27,n1027);
xor (n1027,n1028,n1842);
xor (n1028,n1029,n2324);
xor (n1029,n1030,n1837);
xor (n1030,n1031,n2317);
xor (n1031,n1032,n1831);
xor (n1032,n1033,n2305);
xor (n1033,n1034,n1825);
xor (n1034,n1035,n2288);
xor (n1035,n1036,n1819);
xor (n1036,n1037,n2266);
xor (n1037,n1038,n1813);
xor (n1038,n1039,n2239);
xor (n1039,n1040,n1807);
xor (n1040,n1041,n2207);
xor (n1041,n1042,n1801);
xor (n1042,n1043,n2170);
xor (n1043,n1044,n1795);
xor (n1044,n1045,n2128);
xor (n1045,n1046,n1789);
xor (n1046,n1047,n2081);
xor (n1047,n1048,n1783);
xor (n1048,n1049,n2029);
xor (n1049,n1050,n1777);
xor (n1050,n1051,n1972);
xor (n1051,n1052,n1771);
xor (n1052,n1053,n1910);
xor (n1053,n1054,n1765);
xor (n1054,n1055,n1843);
xor (n1055,n1056,n58);
xor (n1056,n1057,n1757);
xor (n1057,n1058,n1756);
xor (n1058,n1059,n1668);
xor (n1059,n1060,n1667);
xor (n1060,n1061,n1569);
xor (n1061,n1062,n1568);
xor (n1062,n1063,n1466);
xor (n1063,n1064,n1465);
xor (n1064,n1065,n1358);
xor (n1065,n1066,n1357);
xor (n1066,n1067,n1078);
xor (n1067,n1068,n1077);
xor (n1068,n1069,n1076);
xor (n1069,n1070,n1075);
xor (n1070,n1071,n1074);
xor (n1071,n1072,n1073);
and (n1072,n26,n199);
and (n1073,n26,n167);
and (n1074,n1072,n1073);
and (n1075,n26,n160);
and (n1076,n1070,n1075);
and (n1077,n26,n76);
or (n1078,n1079,n1080);
and (n1079,n1068,n1077);
and (n1080,n1067,n1081);
or (n1081,n1079,n1082);
and (n1082,n1067,n1083);
or (n1083,n1079,n1084);
and (n1084,n1067,n1085);
or (n1085,n1079,n1086);
and (n1086,n1067,n1087);
or (n1087,n1088,n1272);
and (n1088,n1089,n1271);
xor (n1089,n1069,n1090);
or (n1090,n1091,n1183);
and (n1091,n1092,n1182);
xor (n1092,n1071,n1093);
or (n1093,n1074,n1094);
and (n1094,n1095,n1097);
xor (n1095,n1072,n1096);
and (n1096,n28,n167);
or (n1097,n1098,n1101);
and (n1098,n1099,n1100);
and (n1099,n28,n199);
and (n1100,n56,n167);
and (n1101,n1102,n1103);
xor (n1102,n1099,n1100);
or (n1103,n1104,n1107);
and (n1104,n1105,n1106);
and (n1105,n56,n199);
and (n1106,n97,n167);
and (n1107,n1108,n1109);
xor (n1108,n1105,n1106);
or (n1109,n1110,n1113);
and (n1110,n1111,n1112);
and (n1111,n97,n199);
and (n1112,n601,n167);
and (n1113,n1114,n1115);
xor (n1114,n1111,n1112);
or (n1115,n1116,n1119);
and (n1116,n1117,n1118);
and (n1117,n601,n199);
and (n1118,n402,n167);
and (n1119,n1120,n1121);
xor (n1120,n1117,n1118);
or (n1121,n1122,n1125);
and (n1122,n1123,n1124);
and (n1123,n402,n199);
and (n1124,n352,n167);
and (n1125,n1126,n1127);
xor (n1126,n1123,n1124);
or (n1127,n1128,n1131);
and (n1128,n1129,n1130);
and (n1129,n352,n199);
and (n1130,n271,n167);
and (n1131,n1132,n1133);
xor (n1132,n1129,n1130);
or (n1133,n1134,n1137);
and (n1134,n1135,n1136);
and (n1135,n271,n199);
and (n1136,n210,n167);
and (n1137,n1138,n1139);
xor (n1138,n1135,n1136);
or (n1139,n1140,n1143);
and (n1140,n1141,n1142);
and (n1141,n210,n199);
and (n1142,n205,n167);
and (n1143,n1144,n1145);
xor (n1144,n1141,n1142);
or (n1145,n1146,n1148);
and (n1146,n1147,n247);
and (n1147,n205,n199);
and (n1148,n1149,n1150);
xor (n1149,n1147,n247);
or (n1150,n1151,n1154);
and (n1151,n1152,n1153);
and (n1152,n228,n199);
and (n1153,n174,n167);
and (n1154,n1155,n1156);
xor (n1155,n1152,n1153);
or (n1156,n1157,n1160);
and (n1157,n1158,n1159);
and (n1158,n174,n199);
and (n1159,n152,n167);
and (n1160,n1161,n1162);
xor (n1161,n1158,n1159);
or (n1162,n1163,n1165);
and (n1163,n1164,n486);
and (n1164,n152,n199);
and (n1165,n1166,n1167);
xor (n1166,n1164,n486);
or (n1167,n1168,n1171);
and (n1168,n1169,n1170);
and (n1169,n187,n199);
and (n1170,n181,n167);
and (n1171,n1172,n1173);
xor (n1172,n1169,n1170);
or (n1173,n1174,n1177);
and (n1174,n1175,n1176);
and (n1175,n181,n199);
and (n1176,n143,n167);
and (n1177,n1178,n1179);
xor (n1178,n1175,n1176);
and (n1179,n1180,n1181);
and (n1180,n143,n199);
and (n1181,n137,n167);
and (n1182,n28,n160);
and (n1183,n1184,n1185);
xor (n1184,n1092,n1182);
or (n1185,n1186,n1189);
and (n1186,n1187,n1188);
xor (n1187,n1095,n1097);
and (n1188,n56,n160);
and (n1189,n1190,n1191);
xor (n1190,n1187,n1188);
or (n1191,n1192,n1195);
and (n1192,n1193,n1194);
xor (n1193,n1102,n1103);
and (n1194,n97,n160);
and (n1195,n1196,n1197);
xor (n1196,n1193,n1194);
or (n1197,n1198,n1201);
and (n1198,n1199,n1200);
xor (n1199,n1108,n1109);
and (n1200,n601,n160);
and (n1201,n1202,n1203);
xor (n1202,n1199,n1200);
or (n1203,n1204,n1207);
and (n1204,n1205,n1206);
xor (n1205,n1114,n1115);
and (n1206,n402,n160);
and (n1207,n1208,n1209);
xor (n1208,n1205,n1206);
or (n1209,n1210,n1213);
and (n1210,n1211,n1212);
xor (n1211,n1120,n1121);
and (n1212,n352,n160);
and (n1213,n1214,n1215);
xor (n1214,n1211,n1212);
or (n1215,n1216,n1219);
and (n1216,n1217,n1218);
xor (n1217,n1126,n1127);
and (n1218,n271,n160);
and (n1219,n1220,n1221);
xor (n1220,n1217,n1218);
or (n1221,n1222,n1225);
and (n1222,n1223,n1224);
xor (n1223,n1132,n1133);
and (n1224,n210,n160);
and (n1225,n1226,n1227);
xor (n1226,n1223,n1224);
or (n1227,n1228,n1231);
and (n1228,n1229,n1230);
xor (n1229,n1138,n1139);
and (n1230,n205,n160);
and (n1231,n1232,n1233);
xor (n1232,n1229,n1230);
or (n1233,n1234,n1237);
and (n1234,n1235,n1236);
xor (n1235,n1144,n1145);
and (n1236,n228,n160);
and (n1237,n1238,n1239);
xor (n1238,n1235,n1236);
or (n1239,n1240,n1243);
and (n1240,n1241,n1242);
xor (n1241,n1149,n1150);
and (n1242,n174,n160);
and (n1243,n1244,n1245);
xor (n1244,n1241,n1242);
or (n1245,n1246,n1249);
and (n1246,n1247,n1248);
xor (n1247,n1155,n1156);
and (n1248,n152,n160);
and (n1249,n1250,n1251);
xor (n1250,n1247,n1248);
or (n1251,n1252,n1255);
and (n1252,n1253,n1254);
xor (n1253,n1161,n1162);
and (n1254,n187,n160);
and (n1255,n1256,n1257);
xor (n1256,n1253,n1254);
or (n1257,n1258,n1261);
and (n1258,n1259,n1260);
xor (n1259,n1166,n1167);
and (n1260,n181,n160);
and (n1261,n1262,n1263);
xor (n1262,n1259,n1260);
or (n1263,n1264,n1267);
and (n1264,n1265,n1266);
xor (n1265,n1172,n1173);
and (n1266,n143,n160);
and (n1267,n1268,n1269);
xor (n1268,n1265,n1266);
and (n1269,n1270,n505);
xor (n1270,n1178,n1179);
and (n1271,n28,n76);
and (n1272,n1273,n1274);
xor (n1273,n1089,n1271);
or (n1274,n1275,n1278);
and (n1275,n1276,n1277);
xor (n1276,n1184,n1185);
and (n1277,n56,n76);
and (n1278,n1279,n1280);
xor (n1279,n1276,n1277);
or (n1280,n1281,n1284);
and (n1281,n1282,n1283);
xor (n1282,n1190,n1191);
and (n1283,n97,n76);
and (n1284,n1285,n1286);
xor (n1285,n1282,n1283);
or (n1286,n1287,n1290);
and (n1287,n1288,n1289);
xor (n1288,n1196,n1197);
and (n1289,n601,n76);
and (n1290,n1291,n1292);
xor (n1291,n1288,n1289);
or (n1292,n1293,n1296);
and (n1293,n1294,n1295);
xor (n1294,n1202,n1203);
and (n1295,n402,n76);
and (n1296,n1297,n1298);
xor (n1297,n1294,n1295);
or (n1298,n1299,n1302);
and (n1299,n1300,n1301);
xor (n1300,n1208,n1209);
and (n1301,n352,n76);
and (n1302,n1303,n1304);
xor (n1303,n1300,n1301);
or (n1304,n1305,n1308);
and (n1305,n1306,n1307);
xor (n1306,n1214,n1215);
and (n1307,n271,n76);
and (n1308,n1309,n1310);
xor (n1309,n1306,n1307);
or (n1310,n1311,n1314);
and (n1311,n1312,n1313);
xor (n1312,n1220,n1221);
and (n1313,n210,n76);
and (n1314,n1315,n1316);
xor (n1315,n1312,n1313);
or (n1316,n1317,n1320);
and (n1317,n1318,n1319);
xor (n1318,n1226,n1227);
and (n1319,n205,n76);
and (n1320,n1321,n1322);
xor (n1321,n1318,n1319);
or (n1322,n1323,n1326);
and (n1323,n1324,n1325);
xor (n1324,n1232,n1233);
and (n1325,n228,n76);
and (n1326,n1327,n1328);
xor (n1327,n1324,n1325);
or (n1328,n1329,n1331);
and (n1329,n1330,n173);
xor (n1330,n1238,n1239);
and (n1331,n1332,n1333);
xor (n1332,n1330,n173);
or (n1333,n1334,n1337);
and (n1334,n1335,n1336);
xor (n1335,n1244,n1245);
and (n1336,n152,n76);
and (n1337,n1338,n1339);
xor (n1338,n1335,n1336);
or (n1339,n1340,n1342);
and (n1340,n1341,n316);
xor (n1341,n1250,n1251);
and (n1342,n1343,n1344);
xor (n1343,n1341,n316);
or (n1344,n1345,n1347);
and (n1345,n1346,n435);
xor (n1346,n1256,n1257);
and (n1347,n1348,n1349);
xor (n1348,n1346,n435);
or (n1349,n1350,n1352);
and (n1350,n1351,n478);
xor (n1351,n1262,n1263);
and (n1352,n1353,n1354);
xor (n1353,n1351,n478);
and (n1354,n1355,n1356);
xor (n1355,n1268,n1269);
and (n1356,n137,n76);
and (n1357,n26,n73);
or (n1358,n1359,n1361);
and (n1359,n1360,n1357);
xor (n1360,n1067,n1081);
and (n1361,n1362,n1363);
xor (n1362,n1360,n1357);
or (n1363,n1364,n1366);
and (n1364,n1365,n1357);
xor (n1365,n1067,n1083);
and (n1366,n1367,n1368);
xor (n1367,n1365,n1357);
or (n1368,n1369,n1371);
and (n1369,n1370,n1357);
xor (n1370,n1067,n1085);
and (n1371,n1372,n1373);
xor (n1372,n1370,n1357);
or (n1373,n1374,n1377);
and (n1374,n1375,n1376);
xor (n1375,n1067,n1087);
and (n1376,n28,n73);
and (n1377,n1378,n1379);
xor (n1378,n1375,n1376);
or (n1379,n1380,n1383);
and (n1380,n1381,n1382);
xor (n1381,n1273,n1274);
and (n1382,n56,n73);
and (n1383,n1384,n1385);
xor (n1384,n1381,n1382);
or (n1385,n1386,n1389);
and (n1386,n1387,n1388);
xor (n1387,n1279,n1280);
and (n1388,n97,n73);
and (n1389,n1390,n1391);
xor (n1390,n1387,n1388);
or (n1391,n1392,n1395);
and (n1392,n1393,n1394);
xor (n1393,n1285,n1286);
and (n1394,n601,n73);
and (n1395,n1396,n1397);
xor (n1396,n1393,n1394);
or (n1397,n1398,n1401);
and (n1398,n1399,n1400);
xor (n1399,n1291,n1292);
and (n1400,n402,n73);
and (n1401,n1402,n1403);
xor (n1402,n1399,n1400);
or (n1403,n1404,n1407);
and (n1404,n1405,n1406);
xor (n1405,n1297,n1298);
and (n1406,n352,n73);
and (n1407,n1408,n1409);
xor (n1408,n1405,n1406);
or (n1409,n1410,n1413);
and (n1410,n1411,n1412);
xor (n1411,n1303,n1304);
and (n1412,n271,n73);
and (n1413,n1414,n1415);
xor (n1414,n1411,n1412);
or (n1415,n1416,n1419);
and (n1416,n1417,n1418);
xor (n1417,n1309,n1310);
and (n1418,n210,n73);
and (n1419,n1420,n1421);
xor (n1420,n1417,n1418);
or (n1421,n1422,n1425);
and (n1422,n1423,n1424);
xor (n1423,n1315,n1316);
and (n1424,n205,n73);
and (n1425,n1426,n1427);
xor (n1426,n1423,n1424);
or (n1427,n1428,n1431);
and (n1428,n1429,n1430);
xor (n1429,n1321,n1322);
and (n1430,n228,n73);
and (n1431,n1432,n1433);
xor (n1432,n1429,n1430);
or (n1433,n1434,n1437);
and (n1434,n1435,n1436);
xor (n1435,n1327,n1328);
and (n1436,n174,n73);
and (n1437,n1438,n1439);
xor (n1438,n1435,n1436);
or (n1439,n1440,n1443);
and (n1440,n1441,n1442);
xor (n1441,n1332,n1333);
and (n1442,n152,n73);
and (n1443,n1444,n1445);
xor (n1444,n1441,n1442);
or (n1445,n1446,n1449);
and (n1446,n1447,n1448);
xor (n1447,n1338,n1339);
and (n1448,n187,n73);
and (n1449,n1450,n1451);
xor (n1450,n1447,n1448);
or (n1451,n1452,n1455);
and (n1452,n1453,n1454);
xor (n1453,n1343,n1344);
and (n1454,n181,n73);
and (n1455,n1456,n1457);
xor (n1456,n1453,n1454);
or (n1457,n1458,n1461);
and (n1458,n1459,n1460);
xor (n1459,n1348,n1349);
and (n1460,n143,n73);
and (n1461,n1462,n1463);
xor (n1462,n1459,n1460);
and (n1463,n1464,n451);
xor (n1464,n1353,n1354);
and (n1465,n26,n37);
or (n1466,n1467,n1469);
and (n1467,n1468,n1465);
xor (n1468,n1362,n1363);
and (n1469,n1470,n1471);
xor (n1470,n1468,n1465);
or (n1471,n1472,n1474);
and (n1472,n1473,n1465);
xor (n1473,n1367,n1368);
and (n1474,n1475,n1476);
xor (n1475,n1473,n1465);
or (n1476,n1477,n1480);
and (n1477,n1478,n1479);
xor (n1478,n1372,n1373);
and (n1479,n28,n37);
and (n1480,n1481,n1482);
xor (n1481,n1478,n1479);
or (n1482,n1483,n1486);
and (n1483,n1484,n1485);
xor (n1484,n1378,n1379);
and (n1485,n56,n37);
and (n1486,n1487,n1488);
xor (n1487,n1484,n1485);
or (n1488,n1489,n1492);
and (n1489,n1490,n1491);
xor (n1490,n1384,n1385);
and (n1491,n97,n37);
and (n1492,n1493,n1494);
xor (n1493,n1490,n1491);
or (n1494,n1495,n1498);
and (n1495,n1496,n1497);
xor (n1496,n1390,n1391);
and (n1497,n601,n37);
and (n1498,n1499,n1500);
xor (n1499,n1496,n1497);
or (n1500,n1501,n1504);
and (n1501,n1502,n1503);
xor (n1502,n1396,n1397);
and (n1503,n402,n37);
and (n1504,n1505,n1506);
xor (n1505,n1502,n1503);
or (n1506,n1507,n1510);
and (n1507,n1508,n1509);
xor (n1508,n1402,n1403);
and (n1509,n352,n37);
and (n1510,n1511,n1512);
xor (n1511,n1508,n1509);
or (n1512,n1513,n1516);
and (n1513,n1514,n1515);
xor (n1514,n1408,n1409);
and (n1515,n271,n37);
and (n1516,n1517,n1518);
xor (n1517,n1514,n1515);
or (n1518,n1519,n1522);
and (n1519,n1520,n1521);
xor (n1520,n1414,n1415);
and (n1521,n210,n37);
and (n1522,n1523,n1524);
xor (n1523,n1520,n1521);
or (n1524,n1525,n1528);
and (n1525,n1526,n1527);
xor (n1526,n1420,n1421);
and (n1527,n205,n37);
and (n1528,n1529,n1530);
xor (n1529,n1526,n1527);
or (n1530,n1531,n1534);
and (n1531,n1532,n1533);
xor (n1532,n1426,n1427);
and (n1533,n228,n37);
and (n1534,n1535,n1536);
xor (n1535,n1532,n1533);
or (n1536,n1537,n1540);
and (n1537,n1538,n1539);
xor (n1538,n1432,n1433);
and (n1539,n174,n37);
and (n1540,n1541,n1542);
xor (n1541,n1538,n1539);
or (n1542,n1543,n1546);
and (n1543,n1544,n1545);
xor (n1544,n1438,n1439);
and (n1545,n152,n37);
and (n1546,n1547,n1548);
xor (n1547,n1544,n1545);
or (n1548,n1549,n1552);
and (n1549,n1550,n1551);
xor (n1550,n1444,n1445);
and (n1551,n187,n37);
and (n1552,n1553,n1554);
xor (n1553,n1550,n1551);
or (n1554,n1555,n1558);
and (n1555,n1556,n1557);
xor (n1556,n1450,n1451);
and (n1557,n181,n37);
and (n1558,n1559,n1560);
xor (n1559,n1556,n1557);
or (n1560,n1561,n1563);
and (n1561,n1562,n441);
xor (n1562,n1456,n1457);
and (n1563,n1564,n1565);
xor (n1564,n1562,n441);
and (n1565,n1566,n1567);
xor (n1566,n1462,n1463);
and (n1567,n137,n37);
and (n1568,n26,n34);
or (n1569,n1570,n1572);
and (n1570,n1571,n1568);
xor (n1571,n1470,n1471);
and (n1572,n1573,n1574);
xor (n1573,n1571,n1568);
or (n1574,n1575,n1578);
and (n1575,n1576,n1577);
xor (n1576,n1475,n1476);
and (n1577,n28,n34);
and (n1578,n1579,n1580);
xor (n1579,n1576,n1577);
or (n1580,n1581,n1584);
and (n1581,n1582,n1583);
xor (n1582,n1481,n1482);
and (n1583,n56,n34);
and (n1584,n1585,n1586);
xor (n1585,n1582,n1583);
or (n1586,n1587,n1590);
and (n1587,n1588,n1589);
xor (n1588,n1487,n1488);
and (n1589,n97,n34);
and (n1590,n1591,n1592);
xor (n1591,n1588,n1589);
or (n1592,n1593,n1596);
and (n1593,n1594,n1595);
xor (n1594,n1493,n1494);
and (n1595,n601,n34);
and (n1596,n1597,n1598);
xor (n1597,n1594,n1595);
or (n1598,n1599,n1602);
and (n1599,n1600,n1601);
xor (n1600,n1499,n1500);
and (n1601,n402,n34);
and (n1602,n1603,n1604);
xor (n1603,n1600,n1601);
or (n1604,n1605,n1608);
and (n1605,n1606,n1607);
xor (n1606,n1505,n1506);
and (n1607,n352,n34);
and (n1608,n1609,n1610);
xor (n1609,n1606,n1607);
or (n1610,n1611,n1614);
and (n1611,n1612,n1613);
xor (n1612,n1511,n1512);
and (n1613,n271,n34);
and (n1614,n1615,n1616);
xor (n1615,n1612,n1613);
or (n1616,n1617,n1620);
and (n1617,n1618,n1619);
xor (n1618,n1517,n1518);
and (n1619,n210,n34);
and (n1620,n1621,n1622);
xor (n1621,n1618,n1619);
or (n1622,n1623,n1626);
and (n1623,n1624,n1625);
xor (n1624,n1523,n1524);
and (n1625,n205,n34);
and (n1626,n1627,n1628);
xor (n1627,n1624,n1625);
or (n1628,n1629,n1632);
and (n1629,n1630,n1631);
xor (n1630,n1529,n1530);
and (n1631,n228,n34);
and (n1632,n1633,n1634);
xor (n1633,n1630,n1631);
or (n1634,n1635,n1638);
and (n1635,n1636,n1637);
xor (n1636,n1535,n1536);
and (n1637,n174,n34);
and (n1638,n1639,n1640);
xor (n1639,n1636,n1637);
or (n1640,n1641,n1644);
and (n1641,n1642,n1643);
xor (n1642,n1541,n1542);
and (n1643,n152,n34);
and (n1644,n1645,n1646);
xor (n1645,n1642,n1643);
or (n1646,n1647,n1650);
and (n1647,n1648,n1649);
xor (n1648,n1547,n1548);
and (n1649,n187,n34);
and (n1650,n1651,n1652);
xor (n1651,n1648,n1649);
or (n1652,n1653,n1656);
and (n1653,n1654,n1655);
xor (n1654,n1553,n1554);
and (n1655,n181,n34);
and (n1656,n1657,n1658);
xor (n1657,n1654,n1655);
or (n1658,n1659,n1662);
and (n1659,n1660,n1661);
xor (n1660,n1559,n1560);
and (n1661,n143,n34);
and (n1662,n1663,n1664);
xor (n1663,n1660,n1661);
and (n1664,n1665,n1666);
xor (n1665,n1564,n1565);
not (n1666,n241);
and (n1667,n26,n22);
or (n1668,n1669,n1672);
and (n1669,n1670,n1671);
xor (n1670,n1573,n1574);
and (n1671,n28,n22);
and (n1672,n1673,n1674);
xor (n1673,n1670,n1671);
or (n1674,n1675,n1678);
and (n1675,n1676,n1677);
xor (n1676,n1579,n1580);
and (n1677,n56,n22);
and (n1678,n1679,n1680);
xor (n1679,n1676,n1677);
or (n1680,n1681,n1684);
and (n1681,n1682,n1683);
xor (n1682,n1585,n1586);
and (n1683,n97,n22);
and (n1684,n1685,n1686);
xor (n1685,n1682,n1683);
or (n1686,n1687,n1690);
and (n1687,n1688,n1689);
xor (n1688,n1591,n1592);
and (n1689,n601,n22);
and (n1690,n1691,n1692);
xor (n1691,n1688,n1689);
or (n1692,n1693,n1696);
and (n1693,n1694,n1695);
xor (n1694,n1597,n1598);
and (n1695,n402,n22);
and (n1696,n1697,n1698);
xor (n1697,n1694,n1695);
or (n1698,n1699,n1702);
and (n1699,n1700,n1701);
xor (n1700,n1603,n1604);
and (n1701,n352,n22);
and (n1702,n1703,n1704);
xor (n1703,n1700,n1701);
or (n1704,n1705,n1707);
and (n1705,n1706,n725);
xor (n1706,n1609,n1610);
and (n1707,n1708,n1709);
xor (n1708,n1706,n725);
or (n1709,n1710,n1712);
and (n1710,n1711,n676);
xor (n1711,n1615,n1616);
and (n1712,n1713,n1714);
xor (n1713,n1711,n676);
or (n1714,n1715,n1718);
and (n1715,n1716,n1717);
xor (n1716,n1621,n1622);
and (n1717,n205,n22);
and (n1718,n1719,n1720);
xor (n1719,n1716,n1717);
or (n1720,n1721,n1724);
and (n1721,n1722,n1723);
xor (n1722,n1627,n1628);
and (n1723,n228,n22);
and (n1724,n1725,n1726);
xor (n1725,n1722,n1723);
or (n1726,n1727,n1729);
and (n1727,n1728,n382);
xor (n1728,n1633,n1634);
and (n1729,n1730,n1731);
xor (n1730,n1728,n382);
or (n1731,n1732,n1734);
and (n1732,n1733,n333);
xor (n1733,n1639,n1640);
and (n1734,n1735,n1736);
xor (n1735,n1733,n333);
or (n1736,n1737,n1739);
and (n1737,n1738,n260);
xor (n1738,n1645,n1646);
and (n1739,n1740,n1741);
xor (n1740,n1738,n260);
or (n1741,n1742,n1745);
and (n1742,n1743,n1744);
xor (n1743,n1651,n1652);
and (n1744,n181,n22);
and (n1745,n1746,n1747);
xor (n1746,n1743,n1744);
or (n1747,n1748,n1751);
and (n1748,n1749,n1750);
xor (n1749,n1657,n1658);
and (n1750,n143,n22);
and (n1751,n1752,n1753);
xor (n1752,n1749,n1750);
and (n1753,n1754,n1755);
xor (n1754,n1663,n1664);
and (n1755,n137,n22);
and (n1756,n28,n53);
or (n1757,n1758,n1760);
and (n1758,n1759,n58);
xor (n1759,n1673,n1674);
and (n1760,n1761,n1762);
xor (n1761,n1759,n58);
or (n1762,n1763,n1766);
and (n1763,n1764,n1765);
xor (n1764,n1679,n1680);
and (n1765,n97,n53);
and (n1766,n1767,n1768);
xor (n1767,n1764,n1765);
or (n1768,n1769,n1772);
and (n1769,n1770,n1771);
xor (n1770,n1685,n1686);
and (n1771,n601,n53);
and (n1772,n1773,n1774);
xor (n1773,n1770,n1771);
or (n1774,n1775,n1778);
and (n1775,n1776,n1777);
xor (n1776,n1691,n1692);
and (n1777,n402,n53);
and (n1778,n1779,n1780);
xor (n1779,n1776,n1777);
or (n1780,n1781,n1784);
and (n1781,n1782,n1783);
xor (n1782,n1697,n1698);
and (n1783,n352,n53);
and (n1784,n1785,n1786);
xor (n1785,n1782,n1783);
or (n1786,n1787,n1790);
and (n1787,n1788,n1789);
xor (n1788,n1703,n1704);
and (n1789,n271,n53);
and (n1790,n1791,n1792);
xor (n1791,n1788,n1789);
or (n1792,n1793,n1796);
and (n1793,n1794,n1795);
xor (n1794,n1708,n1709);
and (n1795,n210,n53);
and (n1796,n1797,n1798);
xor (n1797,n1794,n1795);
or (n1798,n1799,n1802);
and (n1799,n1800,n1801);
xor (n1800,n1713,n1714);
and (n1801,n205,n53);
and (n1802,n1803,n1804);
xor (n1803,n1800,n1801);
or (n1804,n1805,n1808);
and (n1805,n1806,n1807);
xor (n1806,n1719,n1720);
and (n1807,n228,n53);
and (n1808,n1809,n1810);
xor (n1809,n1806,n1807);
or (n1810,n1811,n1814);
and (n1811,n1812,n1813);
xor (n1812,n1725,n1726);
and (n1813,n174,n53);
and (n1814,n1815,n1816);
xor (n1815,n1812,n1813);
or (n1816,n1817,n1820);
and (n1817,n1818,n1819);
xor (n1818,n1730,n1731);
and (n1819,n152,n53);
and (n1820,n1821,n1822);
xor (n1821,n1818,n1819);
or (n1822,n1823,n1826);
and (n1823,n1824,n1825);
xor (n1824,n1735,n1736);
and (n1825,n187,n53);
and (n1826,n1827,n1828);
xor (n1827,n1824,n1825);
or (n1828,n1829,n1832);
and (n1829,n1830,n1831);
xor (n1830,n1740,n1741);
and (n1831,n181,n53);
and (n1832,n1833,n1834);
xor (n1833,n1830,n1831);
or (n1834,n1835,n1838);
and (n1835,n1836,n1837);
xor (n1836,n1746,n1747);
and (n1837,n143,n53);
and (n1838,n1839,n1840);
xor (n1839,n1836,n1837);
and (n1840,n1841,n1842);
xor (n1841,n1752,n1753);
and (n1842,n137,n53);
or (n1843,n1844,n1846);
and (n1844,n1845,n1765);
xor (n1845,n1761,n1762);
and (n1846,n1847,n1848);
xor (n1847,n1845,n1765);
or (n1848,n1849,n1851);
and (n1849,n1850,n1771);
xor (n1850,n1767,n1768);
and (n1851,n1852,n1853);
xor (n1852,n1850,n1771);
or (n1853,n1854,n1856);
and (n1854,n1855,n1777);
xor (n1855,n1773,n1774);
and (n1856,n1857,n1858);
xor (n1857,n1855,n1777);
or (n1858,n1859,n1861);
and (n1859,n1860,n1783);
xor (n1860,n1779,n1780);
and (n1861,n1862,n1863);
xor (n1862,n1860,n1783);
or (n1863,n1864,n1866);
and (n1864,n1865,n1789);
xor (n1865,n1785,n1786);
and (n1866,n1867,n1868);
xor (n1867,n1865,n1789);
or (n1868,n1869,n1871);
and (n1869,n1870,n1795);
xor (n1870,n1791,n1792);
and (n1871,n1872,n1873);
xor (n1872,n1870,n1795);
or (n1873,n1874,n1876);
and (n1874,n1875,n1801);
xor (n1875,n1797,n1798);
and (n1876,n1877,n1878);
xor (n1877,n1875,n1801);
or (n1878,n1879,n1881);
and (n1879,n1880,n1807);
xor (n1880,n1803,n1804);
and (n1881,n1882,n1883);
xor (n1882,n1880,n1807);
or (n1883,n1884,n1886);
and (n1884,n1885,n1813);
xor (n1885,n1809,n1810);
and (n1886,n1887,n1888);
xor (n1887,n1885,n1813);
or (n1888,n1889,n1891);
and (n1889,n1890,n1819);
xor (n1890,n1815,n1816);
and (n1891,n1892,n1893);
xor (n1892,n1890,n1819);
or (n1893,n1894,n1896);
and (n1894,n1895,n1825);
xor (n1895,n1821,n1822);
and (n1896,n1897,n1898);
xor (n1897,n1895,n1825);
or (n1898,n1899,n1901);
and (n1899,n1900,n1831);
xor (n1900,n1827,n1828);
and (n1901,n1902,n1903);
xor (n1902,n1900,n1831);
or (n1903,n1904,n1906);
and (n1904,n1905,n1837);
xor (n1905,n1833,n1834);
and (n1906,n1907,n1908);
xor (n1907,n1905,n1837);
and (n1908,n1909,n1842);
xor (n1909,n1839,n1840);
or (n1910,n1911,n1913);
and (n1911,n1912,n1771);
xor (n1912,n1847,n1848);
and (n1913,n1914,n1915);
xor (n1914,n1912,n1771);
or (n1915,n1916,n1918);
and (n1916,n1917,n1777);
xor (n1917,n1852,n1853);
and (n1918,n1919,n1920);
xor (n1919,n1917,n1777);
or (n1920,n1921,n1923);
and (n1921,n1922,n1783);
xor (n1922,n1857,n1858);
and (n1923,n1924,n1925);
xor (n1924,n1922,n1783);
or (n1925,n1926,n1928);
and (n1926,n1927,n1789);
xor (n1927,n1862,n1863);
and (n1928,n1929,n1930);
xor (n1929,n1927,n1789);
or (n1930,n1931,n1933);
and (n1931,n1932,n1795);
xor (n1932,n1867,n1868);
and (n1933,n1934,n1935);
xor (n1934,n1932,n1795);
or (n1935,n1936,n1938);
and (n1936,n1937,n1801);
xor (n1937,n1872,n1873);
and (n1938,n1939,n1940);
xor (n1939,n1937,n1801);
or (n1940,n1941,n1943);
and (n1941,n1942,n1807);
xor (n1942,n1877,n1878);
and (n1943,n1944,n1945);
xor (n1944,n1942,n1807);
or (n1945,n1946,n1948);
and (n1946,n1947,n1813);
xor (n1947,n1882,n1883);
and (n1948,n1949,n1950);
xor (n1949,n1947,n1813);
or (n1950,n1951,n1953);
and (n1951,n1952,n1819);
xor (n1952,n1887,n1888);
and (n1953,n1954,n1955);
xor (n1954,n1952,n1819);
or (n1955,n1956,n1958);
and (n1956,n1957,n1825);
xor (n1957,n1892,n1893);
and (n1958,n1959,n1960);
xor (n1959,n1957,n1825);
or (n1960,n1961,n1963);
and (n1961,n1962,n1831);
xor (n1962,n1897,n1898);
and (n1963,n1964,n1965);
xor (n1964,n1962,n1831);
or (n1965,n1966,n1968);
and (n1966,n1967,n1837);
xor (n1967,n1902,n1903);
and (n1968,n1969,n1970);
xor (n1969,n1967,n1837);
and (n1970,n1971,n1842);
xor (n1971,n1907,n1908);
or (n1972,n1973,n1975);
and (n1973,n1974,n1777);
xor (n1974,n1914,n1915);
and (n1975,n1976,n1977);
xor (n1976,n1974,n1777);
or (n1977,n1978,n1980);
and (n1978,n1979,n1783);
xor (n1979,n1919,n1920);
and (n1980,n1981,n1982);
xor (n1981,n1979,n1783);
or (n1982,n1983,n1985);
and (n1983,n1984,n1789);
xor (n1984,n1924,n1925);
and (n1985,n1986,n1987);
xor (n1986,n1984,n1789);
or (n1987,n1988,n1990);
and (n1988,n1989,n1795);
xor (n1989,n1929,n1930);
and (n1990,n1991,n1992);
xor (n1991,n1989,n1795);
or (n1992,n1993,n1995);
and (n1993,n1994,n1801);
xor (n1994,n1934,n1935);
and (n1995,n1996,n1997);
xor (n1996,n1994,n1801);
or (n1997,n1998,n2000);
and (n1998,n1999,n1807);
xor (n1999,n1939,n1940);
and (n2000,n2001,n2002);
xor (n2001,n1999,n1807);
or (n2002,n2003,n2005);
and (n2003,n2004,n1813);
xor (n2004,n1944,n1945);
and (n2005,n2006,n2007);
xor (n2006,n2004,n1813);
or (n2007,n2008,n2010);
and (n2008,n2009,n1819);
xor (n2009,n1949,n1950);
and (n2010,n2011,n2012);
xor (n2011,n2009,n1819);
or (n2012,n2013,n2015);
and (n2013,n2014,n1825);
xor (n2014,n1954,n1955);
and (n2015,n2016,n2017);
xor (n2016,n2014,n1825);
or (n2017,n2018,n2020);
and (n2018,n2019,n1831);
xor (n2019,n1959,n1960);
and (n2020,n2021,n2022);
xor (n2021,n2019,n1831);
or (n2022,n2023,n2025);
and (n2023,n2024,n1837);
xor (n2024,n1964,n1965);
and (n2025,n2026,n2027);
xor (n2026,n2024,n1837);
and (n2027,n2028,n1842);
xor (n2028,n1969,n1970);
or (n2029,n2030,n2032);
and (n2030,n2031,n1783);
xor (n2031,n1976,n1977);
and (n2032,n2033,n2034);
xor (n2033,n2031,n1783);
or (n2034,n2035,n2037);
and (n2035,n2036,n1789);
xor (n2036,n1981,n1982);
and (n2037,n2038,n2039);
xor (n2038,n2036,n1789);
or (n2039,n2040,n2042);
and (n2040,n2041,n1795);
xor (n2041,n1986,n1987);
and (n2042,n2043,n2044);
xor (n2043,n2041,n1795);
or (n2044,n2045,n2047);
and (n2045,n2046,n1801);
xor (n2046,n1991,n1992);
and (n2047,n2048,n2049);
xor (n2048,n2046,n1801);
or (n2049,n2050,n2052);
and (n2050,n2051,n1807);
xor (n2051,n1996,n1997);
and (n2052,n2053,n2054);
xor (n2053,n2051,n1807);
or (n2054,n2055,n2057);
and (n2055,n2056,n1813);
xor (n2056,n2001,n2002);
and (n2057,n2058,n2059);
xor (n2058,n2056,n1813);
or (n2059,n2060,n2062);
and (n2060,n2061,n1819);
xor (n2061,n2006,n2007);
and (n2062,n2063,n2064);
xor (n2063,n2061,n1819);
or (n2064,n2065,n2067);
and (n2065,n2066,n1825);
xor (n2066,n2011,n2012);
and (n2067,n2068,n2069);
xor (n2068,n2066,n1825);
or (n2069,n2070,n2072);
and (n2070,n2071,n1831);
xor (n2071,n2016,n2017);
and (n2072,n2073,n2074);
xor (n2073,n2071,n1831);
or (n2074,n2075,n2077);
and (n2075,n2076,n1837);
xor (n2076,n2021,n2022);
and (n2077,n2078,n2079);
xor (n2078,n2076,n1837);
and (n2079,n2080,n1842);
xor (n2080,n2026,n2027);
or (n2081,n2082,n2084);
and (n2082,n2083,n1789);
xor (n2083,n2033,n2034);
and (n2084,n2085,n2086);
xor (n2085,n2083,n1789);
or (n2086,n2087,n2089);
and (n2087,n2088,n1795);
xor (n2088,n2038,n2039);
and (n2089,n2090,n2091);
xor (n2090,n2088,n1795);
or (n2091,n2092,n2094);
and (n2092,n2093,n1801);
xor (n2093,n2043,n2044);
and (n2094,n2095,n2096);
xor (n2095,n2093,n1801);
or (n2096,n2097,n2099);
and (n2097,n2098,n1807);
xor (n2098,n2048,n2049);
and (n2099,n2100,n2101);
xor (n2100,n2098,n1807);
or (n2101,n2102,n2104);
and (n2102,n2103,n1813);
xor (n2103,n2053,n2054);
and (n2104,n2105,n2106);
xor (n2105,n2103,n1813);
or (n2106,n2107,n2109);
and (n2107,n2108,n1819);
xor (n2108,n2058,n2059);
and (n2109,n2110,n2111);
xor (n2110,n2108,n1819);
or (n2111,n2112,n2114);
and (n2112,n2113,n1825);
xor (n2113,n2063,n2064);
and (n2114,n2115,n2116);
xor (n2115,n2113,n1825);
or (n2116,n2117,n2119);
and (n2117,n2118,n1831);
xor (n2118,n2068,n2069);
and (n2119,n2120,n2121);
xor (n2120,n2118,n1831);
or (n2121,n2122,n2124);
and (n2122,n2123,n1837);
xor (n2123,n2073,n2074);
and (n2124,n2125,n2126);
xor (n2125,n2123,n1837);
and (n2126,n2127,n1842);
xor (n2127,n2078,n2079);
or (n2128,n2129,n2131);
and (n2129,n2130,n1795);
xor (n2130,n2085,n2086);
and (n2131,n2132,n2133);
xor (n2132,n2130,n1795);
or (n2133,n2134,n2136);
and (n2134,n2135,n1801);
xor (n2135,n2090,n2091);
and (n2136,n2137,n2138);
xor (n2137,n2135,n1801);
or (n2138,n2139,n2141);
and (n2139,n2140,n1807);
xor (n2140,n2095,n2096);
and (n2141,n2142,n2143);
xor (n2142,n2140,n1807);
or (n2143,n2144,n2146);
and (n2144,n2145,n1813);
xor (n2145,n2100,n2101);
and (n2146,n2147,n2148);
xor (n2147,n2145,n1813);
or (n2148,n2149,n2151);
and (n2149,n2150,n1819);
xor (n2150,n2105,n2106);
and (n2151,n2152,n2153);
xor (n2152,n2150,n1819);
or (n2153,n2154,n2156);
and (n2154,n2155,n1825);
xor (n2155,n2110,n2111);
and (n2156,n2157,n2158);
xor (n2157,n2155,n1825);
or (n2158,n2159,n2161);
and (n2159,n2160,n1831);
xor (n2160,n2115,n2116);
and (n2161,n2162,n2163);
xor (n2162,n2160,n1831);
or (n2163,n2164,n2166);
and (n2164,n2165,n1837);
xor (n2165,n2120,n2121);
and (n2166,n2167,n2168);
xor (n2167,n2165,n1837);
and (n2168,n2169,n1842);
xor (n2169,n2125,n2126);
or (n2170,n2171,n2173);
and (n2171,n2172,n1801);
xor (n2172,n2132,n2133);
and (n2173,n2174,n2175);
xor (n2174,n2172,n1801);
or (n2175,n2176,n2178);
and (n2176,n2177,n1807);
xor (n2177,n2137,n2138);
and (n2178,n2179,n2180);
xor (n2179,n2177,n1807);
or (n2180,n2181,n2183);
and (n2181,n2182,n1813);
xor (n2182,n2142,n2143);
and (n2183,n2184,n2185);
xor (n2184,n2182,n1813);
or (n2185,n2186,n2188);
and (n2186,n2187,n1819);
xor (n2187,n2147,n2148);
and (n2188,n2189,n2190);
xor (n2189,n2187,n1819);
or (n2190,n2191,n2193);
and (n2191,n2192,n1825);
xor (n2192,n2152,n2153);
and (n2193,n2194,n2195);
xor (n2194,n2192,n1825);
or (n2195,n2196,n2198);
and (n2196,n2197,n1831);
xor (n2197,n2157,n2158);
and (n2198,n2199,n2200);
xor (n2199,n2197,n1831);
or (n2200,n2201,n2203);
and (n2201,n2202,n1837);
xor (n2202,n2162,n2163);
and (n2203,n2204,n2205);
xor (n2204,n2202,n1837);
and (n2205,n2206,n1842);
xor (n2206,n2167,n2168);
or (n2207,n2208,n2210);
and (n2208,n2209,n1807);
xor (n2209,n2174,n2175);
and (n2210,n2211,n2212);
xor (n2211,n2209,n1807);
or (n2212,n2213,n2215);
and (n2213,n2214,n1813);
xor (n2214,n2179,n2180);
and (n2215,n2216,n2217);
xor (n2216,n2214,n1813);
or (n2217,n2218,n2220);
and (n2218,n2219,n1819);
xor (n2219,n2184,n2185);
and (n2220,n2221,n2222);
xor (n2221,n2219,n1819);
or (n2222,n2223,n2225);
and (n2223,n2224,n1825);
xor (n2224,n2189,n2190);
and (n2225,n2226,n2227);
xor (n2226,n2224,n1825);
or (n2227,n2228,n2230);
and (n2228,n2229,n1831);
xor (n2229,n2194,n2195);
and (n2230,n2231,n2232);
xor (n2231,n2229,n1831);
or (n2232,n2233,n2235);
and (n2233,n2234,n1837);
xor (n2234,n2199,n2200);
and (n2235,n2236,n2237);
xor (n2236,n2234,n1837);
and (n2237,n2238,n1842);
xor (n2238,n2204,n2205);
or (n2239,n2240,n2242);
and (n2240,n2241,n1813);
xor (n2241,n2211,n2212);
and (n2242,n2243,n2244);
xor (n2243,n2241,n1813);
or (n2244,n2245,n2247);
and (n2245,n2246,n1819);
xor (n2246,n2216,n2217);
and (n2247,n2248,n2249);
xor (n2248,n2246,n1819);
or (n2249,n2250,n2252);
and (n2250,n2251,n1825);
xor (n2251,n2221,n2222);
and (n2252,n2253,n2254);
xor (n2253,n2251,n1825);
or (n2254,n2255,n2257);
and (n2255,n2256,n1831);
xor (n2256,n2226,n2227);
and (n2257,n2258,n2259);
xor (n2258,n2256,n1831);
or (n2259,n2260,n2262);
and (n2260,n2261,n1837);
xor (n2261,n2231,n2232);
and (n2262,n2263,n2264);
xor (n2263,n2261,n1837);
and (n2264,n2265,n1842);
xor (n2265,n2236,n2237);
or (n2266,n2267,n2269);
and (n2267,n2268,n1819);
xor (n2268,n2243,n2244);
and (n2269,n2270,n2271);
xor (n2270,n2268,n1819);
or (n2271,n2272,n2274);
and (n2272,n2273,n1825);
xor (n2273,n2248,n2249);
and (n2274,n2275,n2276);
xor (n2275,n2273,n1825);
or (n2276,n2277,n2279);
and (n2277,n2278,n1831);
xor (n2278,n2253,n2254);
and (n2279,n2280,n2281);
xor (n2280,n2278,n1831);
or (n2281,n2282,n2284);
and (n2282,n2283,n1837);
xor (n2283,n2258,n2259);
and (n2284,n2285,n2286);
xor (n2285,n2283,n1837);
and (n2286,n2287,n1842);
xor (n2287,n2263,n2264);
or (n2288,n2289,n2291);
and (n2289,n2290,n1825);
xor (n2290,n2270,n2271);
and (n2291,n2292,n2293);
xor (n2292,n2290,n1825);
or (n2293,n2294,n2296);
and (n2294,n2295,n1831);
xor (n2295,n2275,n2276);
and (n2296,n2297,n2298);
xor (n2297,n2295,n1831);
or (n2298,n2299,n2301);
and (n2299,n2300,n1837);
xor (n2300,n2280,n2281);
and (n2301,n2302,n2303);
xor (n2302,n2300,n1837);
and (n2303,n2304,n1842);
xor (n2304,n2285,n2286);
or (n2305,n2306,n2308);
and (n2306,n2307,n1831);
xor (n2307,n2292,n2293);
and (n2308,n2309,n2310);
xor (n2309,n2307,n1831);
or (n2310,n2311,n2313);
and (n2311,n2312,n1837);
xor (n2312,n2297,n2298);
and (n2313,n2314,n2315);
xor (n2314,n2312,n1837);
and (n2315,n2316,n1842);
xor (n2316,n2302,n2303);
or (n2317,n2318,n2320);
and (n2318,n2319,n1837);
xor (n2319,n2309,n2310);
and (n2320,n2321,n2322);
xor (n2321,n2319,n1837);
and (n2322,n2323,n1842);
xor (n2323,n2314,n2315);
and (n2324,n2325,n1842);
xor (n2325,n2321,n2322);
endmodule
