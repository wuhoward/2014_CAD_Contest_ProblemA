module top (out,n4,n5,n23,n24,n28,n32,n39,n47,n49
        ,n56,n57,n66,n74,n80,n86,n91,n104,n111,n117
        ,n125,n131,n135,n141,n150,n151,n160,n165,n174,n182
        ,n186,n190,n199,n402,n444,n892);
output out;
input n4;
input n5;
input n23;
input n24;
input n28;
input n32;
input n39;
input n47;
input n49;
input n56;
input n57;
input n66;
input n74;
input n80;
input n86;
input n91;
input n104;
input n111;
input n117;
input n125;
input n131;
input n135;
input n141;
input n150;
input n151;
input n160;
input n165;
input n174;
input n182;
input n186;
input n190;
input n199;
input n402;
input n444;
input n892;
wire n0;
wire n1;
wire n2;
wire n3;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n25;
wire n26;
wire n27;
wire n29;
wire n30;
wire n31;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n48;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n87;
wire n88;
wire n89;
wire n90;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n132;
wire n133;
wire n134;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n161;
wire n162;
wire n163;
wire n164;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n183;
wire n184;
wire n185;
wire n187;
wire n188;
wire n189;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
xor (out,n0,n894);
or (n0,n1,n891);
and (n1,n2,n6);
nor (n2,n3,n5);
not (n3,n4);
xor (n6,n7,n453);
xor (n7,n8,n360);
or (n8,n9,n359);
and (n9,n10,n303);
xor (n10,n11,n202);
xor (n11,n12,n169);
xor (n12,n13,n95);
or (n13,n14,n94);
and (n14,n15,n69);
xor (n15,n16,n42);
nand (n16,n17,n36);
or (n17,n18,n30);
nand (n18,n19,n26);
not (n19,n20);
nand (n20,n21,n25);
or (n21,n22,n24);
not (n22,n23);
nand (n25,n22,n24);
nand (n26,n27,n29);
or (n27,n22,n28);
nand (n29,n28,n22);
nor (n30,n31,n34);
and (n31,n32,n33);
not (n33,n28);
and (n34,n35,n28);
not (n35,n32);
or (n36,n19,n37);
nor (n37,n38,n40);
and (n38,n33,n39);
and (n40,n28,n41);
not (n41,n39);
nand (n42,n43,n63);
or (n43,n44,n52);
not (n44,n45);
nand (n45,n46,n50);
or (n46,n47,n48);
not (n48,n49);
or (n50,n51,n49);
not (n51,n47);
nand (n52,n53,n60);
nor (n53,n54,n58);
and (n54,n55,n57);
not (n55,n56);
and (n58,n56,n59);
not (n59,n57);
nand (n60,n61,n62);
or (n61,n57,n51);
nand (n62,n51,n57);
or (n63,n64,n53);
nor (n64,n65,n67);
and (n65,n66,n51);
and (n67,n47,n68);
not (n68,n66);
nand (n69,n70,n88);
or (n70,n71,n82);
nand (n71,n72,n77);
nor (n72,n73,n75);
and (n73,n51,n74);
and (n75,n47,n76);
not (n76,n74);
nand (n77,n78,n81);
or (n78,n79,n74);
not (n79,n80);
nand (n81,n79,n74);
not (n82,n83);
nor (n83,n84,n87);
and (n84,n85,n79);
not (n85,n86);
and (n87,n86,n80);
or (n88,n89,n72);
nor (n89,n90,n92);
and (n90,n79,n91);
and (n92,n80,n93);
not (n93,n91);
and (n94,n16,n42);
or (n95,n96,n168);
and (n96,n97,n144);
xor (n97,n98,n120);
nand (n98,n99,n114);
or (n99,n100,n109);
nand (n100,n101,n106);
nor (n101,n102,n105);
and (n102,n103,n28);
not (n103,n104);
and (n105,n104,n33);
nand (n106,n107,n108);
or (n107,n104,n55);
nand (n108,n55,n104);
nor (n109,n110,n112);
and (n110,n55,n111);
and (n112,n56,n113);
not (n113,n111);
or (n114,n101,n115);
nor (n115,n116,n118);
and (n116,n55,n117);
and (n118,n56,n119);
not (n119,n117);
nand (n120,n121,n138);
or (n121,n122,n133);
nand (n122,n123,n128);
nor (n123,n124,n126);
and (n124,n79,n125);
and (n126,n80,n127);
not (n127,n125);
nand (n128,n129,n132);
nand (n129,n130,n125);
not (n130,n131);
nand (n132,n131,n127);
nor (n133,n134,n136);
and (n134,n135,n130);
and (n136,n131,n137);
not (n137,n135);
or (n138,n139,n123);
nor (n139,n140,n142);
and (n140,n141,n130);
and (n142,n131,n143);
not (n143,n141);
nand (n144,n145,n162);
or (n145,n146,n157);
nand (n146,n147,n154);
or (n147,n148,n152);
and (n148,n149,n151);
not (n149,n150);
and (n152,n150,n153);
not (n153,n151);
nor (n154,n155,n156);
and (n155,n131,n149);
and (n156,n130,n150);
nor (n157,n158,n161);
and (n158,n159,n151);
not (n159,n160);
and (n161,n160,n153);
or (n162,n163,n154);
nor (n163,n164,n166);
and (n164,n153,n165);
and (n166,n167,n151);
not (n167,n165);
and (n168,n98,n120);
xor (n169,n170,n194);
xor (n170,n171,n177);
nor (n171,n172,n159);
nor (n172,n173,n175);
and (n173,n153,n174);
and (n175,n151,n176);
not (n176,n174);
nand (n177,n178,n187);
or (n178,n179,n184);
nor (n179,n180,n183);
and (n180,n24,n181);
not (n181,n182);
nor (n183,n24,n181);
nand (n184,n185,n24);
not (n185,n186);
or (n187,n188,n185);
nor (n188,n189,n192);
and (n189,n190,n191);
not (n191,n24);
and (n192,n193,n24);
not (n193,n190);
nand (n194,n195,n196);
or (n195,n18,n37);
or (n196,n19,n197);
nor (n197,n198,n200);
and (n198,n33,n199);
and (n200,n28,n201);
not (n201,n199);
xor (n202,n203,n253);
xor (n203,n204,n224);
xor (n204,n205,n218);
xor (n205,n206,n212);
nand (n206,n207,n208);
or (n207,n52,n64);
or (n208,n209,n53);
nor (n209,n210,n211);
and (n210,n51,n111);
and (n211,n47,n113);
nand (n212,n213,n214);
or (n213,n71,n89);
or (n214,n215,n72);
nor (n215,n216,n217);
and (n216,n79,n49);
and (n217,n80,n48);
nand (n218,n219,n220);
or (n219,n100,n115);
or (n220,n101,n221);
nor (n221,n222,n223);
and (n222,n55,n32);
and (n223,n56,n35);
xor (n224,n225,n241);
xor (n225,n226,n232);
nand (n226,n227,n228);
or (n227,n122,n139);
or (n228,n123,n229);
nor (n229,n230,n231);
and (n230,n130,n86);
and (n231,n131,n85);
nand (n232,n233,n238);
or (n233,n154,n234);
not (n234,n235);
nand (n235,n236,n237);
or (n236,n137,n151);
or (n237,n153,n135);
nand (n238,n239,n240);
not (n239,n163);
not (n240,n146);
and (n241,n242,n247);
nor (n242,n243,n153);
nor (n243,n244,n246);
and (n244,n245,n130);
nand (n245,n150,n160);
and (n246,n159,n149);
nand (n247,n248,n252);
or (n248,n249,n184);
nor (n249,n250,n251);
and (n250,n191,n199);
and (n251,n24,n201);
or (n252,n179,n185);
or (n253,n254,n302);
and (n254,n255,n278);
xor (n255,n256,n257);
xor (n256,n242,n247);
or (n257,n258,n277);
and (n258,n259,n270);
xor (n259,n260,n262);
and (n260,n261,n160);
not (n261,n154);
nand (n262,n263,n268);
or (n263,n264,n18);
not (n264,n265);
nand (n265,n266,n267);
or (n266,n28,n119);
or (n267,n33,n117);
nand (n268,n269,n20);
not (n269,n30);
nand (n270,n271,n276);
or (n271,n52,n272);
not (n272,n273);
nand (n273,n274,n275);
or (n274,n47,n93);
or (n275,n51,n91);
or (n276,n53,n44);
and (n277,n260,n262);
or (n278,n279,n301);
and (n279,n280,n295);
xor (n280,n281,n289);
nand (n281,n282,n287);
or (n282,n283,n71);
not (n283,n284);
nand (n284,n285,n286);
or (n285,n80,n143);
or (n286,n79,n141);
nand (n287,n83,n288);
not (n288,n72);
nand (n289,n290,n291);
or (n290,n185,n249);
or (n291,n292,n184);
nor (n292,n293,n294);
and (n293,n191,n39);
and (n294,n24,n41);
nand (n295,n296,n300);
or (n296,n297,n122);
nor (n297,n298,n299);
and (n298,n165,n130);
and (n299,n131,n167);
or (n300,n133,n123);
and (n301,n281,n289);
and (n302,n256,n257);
or (n303,n304,n358);
and (n304,n305,n308);
xor (n305,n306,n307);
xor (n306,n97,n144);
xor (n307,n15,n69);
or (n308,n309,n357);
and (n309,n310,n331);
xor (n310,n311,n317);
nand (n311,n312,n316);
or (n312,n100,n313);
nor (n313,n314,n315);
and (n314,n55,n66);
and (n315,n56,n68);
or (n316,n101,n109);
nor (n317,n318,n325);
not (n318,n319);
nand (n319,n320,n324);
or (n320,n321,n18);
nor (n321,n322,n323);
and (n322,n111,n33);
and (n323,n113,n28);
nand (n324,n20,n265);
nand (n325,n326,n131);
nand (n326,n327,n328);
or (n327,n160,n125);
nand (n328,n329,n79);
not (n329,n330);
and (n330,n160,n125);
or (n331,n332,n356);
and (n332,n333,n349);
xor (n333,n334,n342);
nand (n334,n335,n336);
or (n335,n53,n272);
nand (n336,n337,n341);
not (n337,n338);
nor (n338,n339,n340);
and (n339,n85,n47);
and (n340,n86,n51);
not (n341,n52);
nand (n342,n343,n348);
or (n343,n344,n71);
not (n344,n345);
nor (n345,n346,n347);
and (n346,n79,n137);
and (n347,n80,n135);
nand (n348,n288,n284);
nand (n349,n350,n355);
or (n350,n351,n184);
not (n351,n352);
or (n352,n353,n354);
and (n353,n35,n24);
and (n354,n32,n191);
or (n355,n292,n185);
and (n356,n334,n342);
and (n357,n311,n317);
and (n358,n306,n307);
and (n359,n11,n202);
xor (n360,n361,n420);
xor (n361,n362,n417);
xor (n362,n363,n388);
xor (n363,n364,n367);
or (n364,n365,n366);
and (n365,n205,n218);
and (n366,n206,n212);
xor (n367,n368,n382);
xor (n368,n369,n376);
nand (n369,n370,n375);
or (n370,n72,n371);
not (n371,n372);
nor (n372,n373,n374);
and (n373,n68,n79);
and (n374,n66,n80);
or (n375,n71,n215);
nand (n376,n377,n378);
or (n377,n100,n221);
or (n378,n101,n379);
nor (n379,n380,n381);
and (n380,n39,n55);
and (n381,n41,n56);
nand (n382,n383,n384);
or (n383,n122,n229);
or (n384,n123,n385);
nor (n385,n386,n387);
and (n386,n91,n130);
and (n387,n131,n93);
xor (n388,n389,n411);
xor (n389,n390,n396);
nand (n390,n391,n392);
or (n391,n18,n197);
or (n392,n19,n393);
nor (n393,n394,n395);
and (n394,n33,n182);
and (n395,n28,n181);
nand (n396,n397,n407);
or (n397,n398,n404);
nand (n398,n172,n399);
nand (n399,n400,n403);
or (n400,n401,n174);
not (n401,n402);
nand (n403,n401,n174);
nor (n404,n405,n406);
and (n405,n159,n402);
and (n406,n160,n401);
or (n407,n408,n172);
nor (n408,n409,n410);
and (n409,n165,n401);
and (n410,n167,n402);
nand (n411,n412,n413);
or (n412,n52,n209);
or (n413,n53,n414);
nor (n414,n415,n416);
and (n415,n51,n117);
and (n416,n47,n119);
or (n417,n418,n419);
and (n418,n203,n253);
and (n419,n204,n224);
xor (n420,n421,n450);
xor (n421,n422,n425);
or (n422,n423,n424);
and (n423,n225,n241);
and (n424,n226,n232);
xor (n425,n426,n447);
xor (n426,n427,n433);
nand (n427,n428,n429);
or (n428,n146,n234);
or (n429,n430,n154);
nor (n430,n431,n432);
and (n431,n141,n153);
and (n432,n151,n143);
xor (n433,n434,n439);
nor (n434,n435,n401);
nor (n435,n436,n438);
and (n436,n437,n153);
nand (n437,n160,n174);
and (n438,n159,n176);
nand (n439,n440,n441);
or (n440,n188,n184);
or (n441,n442,n185);
nor (n442,n443,n445);
and (n443,n191,n444);
and (n445,n24,n446);
not (n446,n444);
or (n447,n448,n449);
and (n448,n170,n194);
and (n449,n171,n177);
or (n450,n451,n452);
and (n451,n12,n169);
and (n452,n13,n95);
or (n453,n454,n890);
and (n454,n455,n489);
xor (n455,n456,n488);
or (n456,n457,n487);
and (n457,n458,n486);
xor (n458,n459,n460);
xor (n459,n255,n278);
or (n460,n461,n485);
and (n461,n462,n465);
xor (n462,n463,n464);
xor (n463,n280,n295);
xor (n464,n259,n270);
or (n465,n466,n484);
and (n466,n467,n480);
xor (n467,n468,n474);
nand (n468,n469,n473);
or (n469,n122,n470);
nor (n470,n471,n472);
and (n471,n159,n131);
and (n472,n160,n130);
or (n473,n297,n123);
nand (n474,n475,n479);
or (n475,n100,n476);
nor (n476,n477,n478);
and (n477,n55,n49);
and (n478,n56,n48);
or (n479,n101,n313);
nand (n480,n481,n483);
or (n481,n482,n318);
not (n482,n325);
or (n483,n319,n325);
and (n484,n468,n474);
and (n485,n463,n464);
xor (n486,n305,n308);
and (n487,n459,n460);
xor (n488,n10,n303);
nand (n489,n490,n886);
or (n490,n491,n864);
nor (n491,n492,n863);
and (n492,n493,n844);
or (n493,n494,n843);
and (n494,n495,n638);
xor (n495,n496,n607);
or (n496,n497,n606);
and (n497,n498,n568);
xor (n498,n499,n529);
xor (n499,n500,n519);
xor (n500,n501,n510);
nand (n501,n502,n506);
or (n502,n52,n503);
nor (n503,n504,n505);
and (n504,n135,n51);
and (n505,n137,n47);
or (n506,n507,n53);
nor (n507,n508,n509);
and (n508,n51,n141);
and (n509,n47,n143);
nand (n510,n511,n515);
or (n511,n71,n512);
nor (n512,n513,n514);
and (n513,n159,n80);
and (n514,n160,n79);
or (n515,n516,n72);
nor (n516,n517,n518);
and (n517,n165,n79);
and (n518,n167,n80);
nand (n519,n520,n525);
or (n520,n184,n521);
not (n521,n522);
nor (n522,n523,n524);
and (n523,n111,n24);
and (n524,n113,n191);
or (n525,n526,n185);
nor (n526,n527,n528);
and (n527,n117,n191);
and (n528,n119,n24);
or (n529,n530,n567);
and (n530,n531,n550);
xor (n531,n532,n541);
nand (n532,n533,n537);
or (n533,n18,n534);
nor (n534,n535,n536);
and (n535,n33,n91);
and (n536,n28,n93);
or (n537,n19,n538);
nor (n538,n539,n540);
and (n539,n48,n28);
and (n540,n49,n33);
nand (n541,n542,n546);
or (n542,n100,n543);
nor (n543,n544,n545);
and (n544,n141,n55);
and (n545,n56,n143);
or (n546,n101,n547);
nor (n547,n548,n549);
and (n548,n55,n86);
and (n549,n56,n85);
and (n550,n551,n557);
nor (n551,n552,n51);
nor (n552,n553,n556);
and (n553,n554,n55);
not (n554,n555);
and (n555,n160,n57);
and (n556,n159,n59);
nand (n557,n558,n563);
or (n558,n559,n184);
not (n559,n560);
nor (n560,n561,n562);
and (n561,n48,n191);
and (n562,n49,n24);
or (n563,n564,n185);
nor (n564,n565,n566);
and (n565,n66,n191);
and (n566,n68,n24);
and (n567,n532,n541);
xor (n568,n569,n591);
xor (n569,n570,n576);
nand (n570,n571,n572);
or (n571,n100,n547);
or (n572,n101,n573);
nor (n573,n574,n575);
and (n574,n55,n91);
and (n575,n56,n93);
xor (n576,n577,n582);
nor (n577,n578,n79);
nor (n578,n579,n581);
and (n579,n580,n51);
nand (n580,n160,n74);
and (n581,n159,n76);
nand (n582,n583,n588);
or (n583,n19,n584);
not (n584,n585);
nand (n585,n586,n587);
or (n586,n28,n68);
or (n587,n33,n66);
nand (n588,n589,n590);
not (n589,n538);
not (n590,n18);
or (n591,n592,n605);
and (n592,n593,n598);
xor (n593,n594,n595);
nor (n594,n72,n159);
nand (n595,n596,n597);
or (n596,n185,n521);
or (n597,n564,n184);
nand (n598,n599,n600);
or (n599,n53,n503);
nand (n600,n601,n341);
not (n601,n602);
or (n602,n603,n604);
and (n603,n167,n51);
and (n604,n165,n47);
and (n605,n594,n595);
and (n606,n499,n529);
xor (n607,n608,n623);
xor (n608,n609,n620);
xor (n609,n610,n617);
xor (n610,n611,n614);
nand (n611,n612,n613);
or (n612,n72,n344);
or (n613,n71,n516);
nand (n614,n615,n616);
or (n615,n526,n184);
nand (n616,n352,n186);
nand (n617,n618,n619);
or (n618,n100,n573);
or (n619,n101,n476);
or (n620,n621,n622);
and (n621,n569,n591);
and (n622,n570,n576);
xor (n623,n624,n629);
xor (n624,n625,n626);
and (n625,n577,n582);
or (n626,n627,n628);
and (n627,n500,n519);
and (n628,n501,n510);
xor (n629,n630,n635);
xor (n630,n631,n632);
nor (n631,n123,n159);
nand (n632,n633,n634);
or (n633,n584,n18);
or (n634,n19,n321);
nand (n635,n636,n637);
or (n636,n52,n507);
or (n637,n53,n338);
nand (n638,n639,n839,n842);
nand (n639,n640,n695,n832);
not (n640,n641);
nor (n641,n642,n669);
xor (n642,n643,n668);
xor (n643,n644,n667);
or (n644,n645,n666);
and (n645,n646,n660);
xor (n646,n647,n653);
nand (n647,n648,n652);
or (n648,n52,n649);
nor (n649,n650,n651);
and (n650,n159,n47);
and (n651,n160,n51);
or (n652,n602,n53);
nand (n653,n654,n659);
or (n654,n655,n18);
not (n655,n656);
nor (n656,n657,n658);
and (n657,n86,n28);
and (n658,n85,n33);
or (n659,n19,n534);
nand (n660,n661,n665);
or (n661,n100,n662);
nor (n662,n663,n664);
and (n663,n135,n55);
and (n664,n56,n137);
or (n665,n101,n543);
and (n666,n647,n653);
xor (n667,n593,n598);
xor (n668,n531,n550);
or (n669,n670,n694);
and (n670,n671,n693);
xor (n671,n672,n673);
xor (n672,n551,n557);
or (n673,n674,n692);
and (n674,n675,n685);
xor (n675,n676,n678);
and (n676,n677,n160);
not (n677,n53);
nand (n678,n679,n684);
or (n679,n184,n680);
not (n680,n681);
nor (n681,n682,n683);
and (n682,n93,n191);
and (n683,n91,n24);
nand (n684,n560,n186);
nand (n685,n686,n691);
or (n686,n687,n18);
not (n687,n688);
nor (n688,n689,n690);
and (n689,n143,n33);
and (n690,n141,n28);
nand (n691,n656,n20);
and (n692,n676,n678);
xor (n693,n646,n660);
and (n694,n672,n673);
or (n695,n696,n831);
and (n696,n697,n723);
xor (n697,n698,n722);
or (n698,n699,n721);
and (n699,n700,n720);
xor (n700,n701,n707);
nand (n701,n702,n706);
or (n702,n100,n703);
nor (n703,n704,n705);
and (n704,n55,n165);
and (n705,n56,n167);
or (n706,n662,n101);
and (n707,n708,n714);
and (n708,n709,n56);
nand (n709,n710,n711);
or (n710,n160,n104);
nand (n711,n712,n33);
not (n712,n713);
and (n713,n160,n104);
nand (n714,n715,n716);
or (n715,n185,n680);
or (n716,n717,n184);
nor (n717,n718,n719);
and (n718,n191,n86);
and (n719,n24,n85);
xor (n720,n675,n685);
and (n721,n701,n707);
xor (n722,n671,n693);
nand (n723,n724,n830);
or (n724,n725,n825);
nor (n725,n726,n824);
and (n726,n727,n803);
nand (n727,n728,n801);
or (n728,n729,n784);
not (n729,n730);
or (n730,n731,n783);
and (n731,n732,n761);
xor (n732,n733,n742);
nand (n733,n734,n738);
or (n734,n18,n735);
nor (n735,n736,n737);
and (n736,n28,n159);
and (n737,n160,n33);
or (n738,n19,n739);
nor (n739,n740,n741);
and (n740,n167,n28);
and (n741,n165,n33);
nand (n742,n743,n760);
or (n743,n744,n750);
not (n744,n745);
nand (n745,n746,n28);
nand (n746,n747,n749);
or (n747,n748,n24);
and (n748,n160,n23);
nand (n749,n159,n22);
not (n750,n751);
nand (n751,n752,n756);
or (n752,n753,n184);
or (n753,n754,n755);
and (n754,n135,n24);
and (n755,n137,n191);
or (n756,n757,n185);
nor (n757,n758,n759);
and (n758,n143,n24);
and (n759,n141,n191);
or (n760,n751,n745);
or (n761,n762,n782);
and (n762,n763,n771);
xor (n763,n764,n765);
nor (n764,n19,n159);
nand (n765,n766,n770);
or (n766,n767,n184);
nor (n767,n768,n769);
and (n768,n167,n24);
and (n769,n165,n191);
or (n770,n753,n185);
nor (n771,n772,n780);
nor (n772,n773,n775);
and (n773,n774,n186);
not (n774,n767);
and (n775,n776,n779);
nand (n776,n777,n778);
or (n777,n159,n24);
nand (n778,n24,n159);
not (n779,n184);
or (n780,n781,n191);
and (n781,n160,n186);
and (n782,n764,n765);
and (n783,n733,n742);
not (n784,n785);
nand (n785,n786,n800);
not (n786,n787);
xor (n787,n788,n797);
xor (n788,n789,n791);
and (n789,n790,n160);
not (n790,n101);
nand (n791,n792,n793);
or (n792,n739,n18);
nand (n793,n794,n20);
nor (n794,n795,n796);
and (n795,n137,n33);
and (n796,n135,n28);
nand (n797,n798,n799);
or (n798,n757,n184);
or (n799,n717,n185);
nand (n800,n744,n751);
nand (n801,n802,n787);
not (n802,n800);
nand (n803,n804,n820);
not (n804,n805);
xor (n805,n806,n819);
xor (n806,n807,n811);
nand (n807,n808,n810);
or (n808,n809,n18);
not (n809,n794);
nand (n810,n688,n20);
nand (n811,n812,n817);
or (n812,n813,n100);
not (n813,n814);
nand (n814,n815,n816);
or (n815,n160,n55);
or (n816,n159,n56);
nand (n817,n818,n790);
not (n818,n703);
xor (n819,n708,n714);
not (n820,n821);
or (n821,n822,n823);
and (n822,n788,n797);
and (n823,n789,n791);
nor (n824,n804,n820);
nor (n825,n826,n827);
xor (n826,n700,n720);
or (n827,n828,n829);
and (n828,n806,n819);
and (n829,n807,n811);
nand (n830,n826,n827);
and (n831,n698,n722);
nand (n832,n833,n837);
not (n833,n834);
or (n834,n835,n836);
and (n835,n643,n668);
and (n836,n644,n667);
not (n837,n838);
xor (n838,n498,n568);
nand (n839,n840,n832);
not (n840,n841);
nand (n841,n642,n669);
nand (n842,n838,n834);
and (n843,n496,n607);
or (n844,n845,n860);
xor (n845,n846,n857);
xor (n846,n847,n848);
xor (n847,n467,n480);
xor (n848,n849,n856);
xor (n849,n850,n853);
or (n850,n851,n852);
and (n851,n630,n635);
and (n852,n631,n632);
or (n853,n854,n855);
and (n854,n610,n617);
and (n855,n611,n614);
xor (n856,n333,n349);
or (n857,n858,n859);
and (n858,n624,n629);
and (n859,n625,n626);
or (n860,n861,n862);
and (n861,n608,n623);
and (n862,n609,n620);
and (n863,n845,n860);
nand (n864,n865,n879);
not (n865,n866);
and (n866,n867,n875);
not (n867,n868);
xor (n868,n869,n874);
xor (n869,n870,n871);
xor (n870,n310,n331);
or (n871,n872,n873);
and (n872,n849,n856);
and (n873,n850,n853);
xor (n874,n462,n465);
not (n875,n876);
or (n876,n877,n878);
and (n877,n846,n857);
and (n878,n847,n848);
nand (n879,n880,n882);
not (n880,n881);
xor (n881,n458,n486);
not (n882,n883);
or (n883,n884,n885);
and (n884,n869,n874);
and (n885,n870,n871);
nor (n886,n887,n889);
and (n887,n879,n888);
nor (n888,n867,n875);
nor (n889,n880,n882);
and (n890,n456,n488);
and (n891,n892,n893);
not (n893,n2);
or (n894,n895,n891);
and (n895,n896,n2);
xor (n896,n897,n1514);
xor (n897,n898,n1511);
xor (n898,n899,n1510);
xor (n899,n900,n1501);
xor (n900,n901,n1500);
xor (n901,n902,n1485);
xor (n902,n903,n1484);
xor (n903,n904,n1463);
xor (n904,n905,n1462);
xor (n905,n906,n1436);
xor (n906,n907,n1435);
xor (n907,n908,n1404);
xor (n908,n909,n1403);
xor (n909,n910,n1364);
xor (n910,n911,n1363);
xor (n911,n912,n1319);
xor (n912,n913,n1318);
xor (n913,n914,n1268);
xor (n914,n915,n1267);
xor (n915,n916,n1210);
xor (n916,n917,n1209);
xor (n917,n918,n1147);
xor (n918,n919,n1146);
xor (n919,n920,n1080);
xor (n920,n921,n1079);
xor (n921,n922,n1005);
xor (n922,n923,n1004);
xor (n923,n924,n927);
xor (n924,n925,n926);
and (n925,n444,n186);
and (n926,n190,n24);
or (n927,n928,n931);
and (n928,n929,n930);
and (n929,n190,n186);
and (n930,n182,n24);
and (n931,n932,n933);
xor (n932,n929,n930);
or (n933,n934,n937);
and (n934,n935,n936);
and (n935,n182,n186);
and (n936,n199,n24);
and (n937,n938,n939);
xor (n938,n935,n936);
or (n939,n940,n943);
and (n940,n941,n942);
and (n941,n199,n186);
and (n942,n39,n24);
and (n943,n944,n945);
xor (n944,n941,n942);
or (n945,n946,n949);
and (n946,n947,n948);
and (n947,n39,n186);
and (n948,n32,n24);
and (n949,n950,n951);
xor (n950,n947,n948);
or (n951,n952,n955);
and (n952,n953,n954);
and (n953,n32,n186);
and (n954,n117,n24);
and (n955,n956,n957);
xor (n956,n953,n954);
or (n957,n958,n960);
and (n958,n959,n523);
and (n959,n117,n186);
and (n960,n961,n962);
xor (n961,n959,n523);
or (n962,n963,n966);
and (n963,n964,n965);
and (n964,n111,n186);
and (n965,n66,n24);
and (n966,n967,n968);
xor (n967,n964,n965);
or (n968,n969,n971);
and (n969,n970,n562);
and (n970,n66,n186);
and (n971,n972,n973);
xor (n972,n970,n562);
or (n973,n974,n976);
and (n974,n975,n683);
and (n975,n49,n186);
and (n976,n977,n978);
xor (n977,n975,n683);
or (n978,n979,n982);
and (n979,n980,n981);
and (n980,n91,n186);
and (n981,n86,n24);
and (n982,n983,n984);
xor (n983,n980,n981);
or (n984,n985,n988);
and (n985,n986,n987);
and (n986,n86,n186);
and (n987,n141,n24);
and (n988,n989,n990);
xor (n989,n986,n987);
or (n990,n991,n993);
and (n991,n992,n754);
and (n992,n141,n186);
and (n993,n994,n995);
xor (n994,n992,n754);
or (n995,n996,n999);
and (n996,n997,n998);
and (n997,n135,n186);
and (n998,n165,n24);
and (n999,n1000,n1001);
xor (n1000,n997,n998);
and (n1001,n1002,n1003);
and (n1002,n165,n186);
and (n1003,n160,n24);
and (n1004,n182,n23);
or (n1005,n1006,n1009);
and (n1006,n1007,n1008);
xor (n1007,n932,n933);
and (n1008,n199,n23);
and (n1009,n1010,n1011);
xor (n1010,n1007,n1008);
or (n1011,n1012,n1015);
and (n1012,n1013,n1014);
xor (n1013,n938,n939);
and (n1014,n39,n23);
and (n1015,n1016,n1017);
xor (n1016,n1013,n1014);
or (n1017,n1018,n1021);
and (n1018,n1019,n1020);
xor (n1019,n944,n945);
and (n1020,n32,n23);
and (n1021,n1022,n1023);
xor (n1022,n1019,n1020);
or (n1023,n1024,n1027);
and (n1024,n1025,n1026);
xor (n1025,n950,n951);
and (n1026,n117,n23);
and (n1027,n1028,n1029);
xor (n1028,n1025,n1026);
or (n1029,n1030,n1033);
and (n1030,n1031,n1032);
xor (n1031,n956,n957);
and (n1032,n111,n23);
and (n1033,n1034,n1035);
xor (n1034,n1031,n1032);
or (n1035,n1036,n1039);
and (n1036,n1037,n1038);
xor (n1037,n961,n962);
and (n1038,n66,n23);
and (n1039,n1040,n1041);
xor (n1040,n1037,n1038);
or (n1041,n1042,n1045);
and (n1042,n1043,n1044);
xor (n1043,n967,n968);
and (n1044,n49,n23);
and (n1045,n1046,n1047);
xor (n1046,n1043,n1044);
or (n1047,n1048,n1051);
and (n1048,n1049,n1050);
xor (n1049,n972,n973);
and (n1050,n91,n23);
and (n1051,n1052,n1053);
xor (n1052,n1049,n1050);
or (n1053,n1054,n1057);
and (n1054,n1055,n1056);
xor (n1055,n977,n978);
and (n1056,n86,n23);
and (n1057,n1058,n1059);
xor (n1058,n1055,n1056);
or (n1059,n1060,n1063);
and (n1060,n1061,n1062);
xor (n1061,n983,n984);
and (n1062,n141,n23);
and (n1063,n1064,n1065);
xor (n1064,n1061,n1062);
or (n1065,n1066,n1069);
and (n1066,n1067,n1068);
xor (n1067,n989,n990);
and (n1068,n135,n23);
and (n1069,n1070,n1071);
xor (n1070,n1067,n1068);
or (n1071,n1072,n1075);
and (n1072,n1073,n1074);
xor (n1073,n994,n995);
and (n1074,n165,n23);
and (n1075,n1076,n1077);
xor (n1076,n1073,n1074);
and (n1077,n1078,n748);
xor (n1078,n1000,n1001);
and (n1079,n199,n28);
or (n1080,n1081,n1084);
and (n1081,n1082,n1083);
xor (n1082,n1010,n1011);
and (n1083,n39,n28);
and (n1084,n1085,n1086);
xor (n1085,n1082,n1083);
or (n1086,n1087,n1090);
and (n1087,n1088,n1089);
xor (n1088,n1016,n1017);
and (n1089,n32,n28);
and (n1090,n1091,n1092);
xor (n1091,n1088,n1089);
or (n1092,n1093,n1096);
and (n1093,n1094,n1095);
xor (n1094,n1022,n1023);
and (n1095,n117,n28);
and (n1096,n1097,n1098);
xor (n1097,n1094,n1095);
or (n1098,n1099,n1102);
and (n1099,n1100,n1101);
xor (n1100,n1028,n1029);
and (n1101,n111,n28);
and (n1102,n1103,n1104);
xor (n1103,n1100,n1101);
or (n1104,n1105,n1108);
and (n1105,n1106,n1107);
xor (n1106,n1034,n1035);
and (n1107,n66,n28);
and (n1108,n1109,n1110);
xor (n1109,n1106,n1107);
or (n1110,n1111,n1114);
and (n1111,n1112,n1113);
xor (n1112,n1040,n1041);
and (n1113,n49,n28);
and (n1114,n1115,n1116);
xor (n1115,n1112,n1113);
or (n1116,n1117,n1120);
and (n1117,n1118,n1119);
xor (n1118,n1046,n1047);
and (n1119,n91,n28);
and (n1120,n1121,n1122);
xor (n1121,n1118,n1119);
or (n1122,n1123,n1125);
and (n1123,n1124,n657);
xor (n1124,n1052,n1053);
and (n1125,n1126,n1127);
xor (n1126,n1124,n657);
or (n1127,n1128,n1130);
and (n1128,n1129,n690);
xor (n1129,n1058,n1059);
and (n1130,n1131,n1132);
xor (n1131,n1129,n690);
or (n1132,n1133,n1135);
and (n1133,n1134,n796);
xor (n1134,n1064,n1065);
and (n1135,n1136,n1137);
xor (n1136,n1134,n796);
or (n1137,n1138,n1141);
and (n1138,n1139,n1140);
xor (n1139,n1070,n1071);
and (n1140,n165,n28);
and (n1141,n1142,n1143);
xor (n1142,n1139,n1140);
and (n1143,n1144,n1145);
xor (n1144,n1076,n1077);
and (n1145,n160,n28);
and (n1146,n39,n104);
or (n1147,n1148,n1151);
and (n1148,n1149,n1150);
xor (n1149,n1085,n1086);
and (n1150,n32,n104);
and (n1151,n1152,n1153);
xor (n1152,n1149,n1150);
or (n1153,n1154,n1157);
and (n1154,n1155,n1156);
xor (n1155,n1091,n1092);
and (n1156,n117,n104);
and (n1157,n1158,n1159);
xor (n1158,n1155,n1156);
or (n1159,n1160,n1163);
and (n1160,n1161,n1162);
xor (n1161,n1097,n1098);
and (n1162,n111,n104);
and (n1163,n1164,n1165);
xor (n1164,n1161,n1162);
or (n1165,n1166,n1169);
and (n1166,n1167,n1168);
xor (n1167,n1103,n1104);
and (n1168,n66,n104);
and (n1169,n1170,n1171);
xor (n1170,n1167,n1168);
or (n1171,n1172,n1175);
and (n1172,n1173,n1174);
xor (n1173,n1109,n1110);
and (n1174,n49,n104);
and (n1175,n1176,n1177);
xor (n1176,n1173,n1174);
or (n1177,n1178,n1181);
and (n1178,n1179,n1180);
xor (n1179,n1115,n1116);
and (n1180,n91,n104);
and (n1181,n1182,n1183);
xor (n1182,n1179,n1180);
or (n1183,n1184,n1187);
and (n1184,n1185,n1186);
xor (n1185,n1121,n1122);
and (n1186,n86,n104);
and (n1187,n1188,n1189);
xor (n1188,n1185,n1186);
or (n1189,n1190,n1193);
and (n1190,n1191,n1192);
xor (n1191,n1126,n1127);
and (n1192,n141,n104);
and (n1193,n1194,n1195);
xor (n1194,n1191,n1192);
or (n1195,n1196,n1199);
and (n1196,n1197,n1198);
xor (n1197,n1131,n1132);
and (n1198,n135,n104);
and (n1199,n1200,n1201);
xor (n1200,n1197,n1198);
or (n1201,n1202,n1205);
and (n1202,n1203,n1204);
xor (n1203,n1136,n1137);
and (n1204,n165,n104);
and (n1205,n1206,n1207);
xor (n1206,n1203,n1204);
and (n1207,n1208,n713);
xor (n1208,n1142,n1143);
and (n1209,n32,n56);
or (n1210,n1211,n1214);
and (n1211,n1212,n1213);
xor (n1212,n1152,n1153);
and (n1213,n117,n56);
and (n1214,n1215,n1216);
xor (n1215,n1212,n1213);
or (n1216,n1217,n1220);
and (n1217,n1218,n1219);
xor (n1218,n1158,n1159);
and (n1219,n111,n56);
and (n1220,n1221,n1222);
xor (n1221,n1218,n1219);
or (n1222,n1223,n1226);
and (n1223,n1224,n1225);
xor (n1224,n1164,n1165);
and (n1225,n66,n56);
and (n1226,n1227,n1228);
xor (n1227,n1224,n1225);
or (n1228,n1229,n1232);
and (n1229,n1230,n1231);
xor (n1230,n1170,n1171);
and (n1231,n49,n56);
and (n1232,n1233,n1234);
xor (n1233,n1230,n1231);
or (n1234,n1235,n1238);
and (n1235,n1236,n1237);
xor (n1236,n1176,n1177);
and (n1237,n91,n56);
and (n1238,n1239,n1240);
xor (n1239,n1236,n1237);
or (n1240,n1241,n1244);
and (n1241,n1242,n1243);
xor (n1242,n1182,n1183);
and (n1243,n86,n56);
and (n1244,n1245,n1246);
xor (n1245,n1242,n1243);
or (n1246,n1247,n1250);
and (n1247,n1248,n1249);
xor (n1248,n1188,n1189);
and (n1249,n141,n56);
and (n1250,n1251,n1252);
xor (n1251,n1248,n1249);
or (n1252,n1253,n1256);
and (n1253,n1254,n1255);
xor (n1254,n1194,n1195);
and (n1255,n135,n56);
and (n1256,n1257,n1258);
xor (n1257,n1254,n1255);
or (n1258,n1259,n1262);
and (n1259,n1260,n1261);
xor (n1260,n1200,n1201);
and (n1261,n165,n56);
and (n1262,n1263,n1264);
xor (n1263,n1260,n1261);
and (n1264,n1265,n1266);
xor (n1265,n1206,n1207);
and (n1266,n160,n56);
and (n1267,n117,n57);
or (n1268,n1269,n1272);
and (n1269,n1270,n1271);
xor (n1270,n1215,n1216);
and (n1271,n111,n57);
and (n1272,n1273,n1274);
xor (n1273,n1270,n1271);
or (n1274,n1275,n1278);
and (n1275,n1276,n1277);
xor (n1276,n1221,n1222);
and (n1277,n66,n57);
and (n1278,n1279,n1280);
xor (n1279,n1276,n1277);
or (n1280,n1281,n1284);
and (n1281,n1282,n1283);
xor (n1282,n1227,n1228);
and (n1283,n49,n57);
and (n1284,n1285,n1286);
xor (n1285,n1282,n1283);
or (n1286,n1287,n1290);
and (n1287,n1288,n1289);
xor (n1288,n1233,n1234);
and (n1289,n91,n57);
and (n1290,n1291,n1292);
xor (n1291,n1288,n1289);
or (n1292,n1293,n1296);
and (n1293,n1294,n1295);
xor (n1294,n1239,n1240);
and (n1295,n86,n57);
and (n1296,n1297,n1298);
xor (n1297,n1294,n1295);
or (n1298,n1299,n1302);
and (n1299,n1300,n1301);
xor (n1300,n1245,n1246);
and (n1301,n141,n57);
and (n1302,n1303,n1304);
xor (n1303,n1300,n1301);
or (n1304,n1305,n1308);
and (n1305,n1306,n1307);
xor (n1306,n1251,n1252);
and (n1307,n135,n57);
and (n1308,n1309,n1310);
xor (n1309,n1306,n1307);
or (n1310,n1311,n1314);
and (n1311,n1312,n1313);
xor (n1312,n1257,n1258);
and (n1313,n165,n57);
and (n1314,n1315,n1316);
xor (n1315,n1312,n1313);
and (n1316,n1317,n555);
xor (n1317,n1263,n1264);
and (n1318,n111,n47);
or (n1319,n1320,n1323);
and (n1320,n1321,n1322);
xor (n1321,n1273,n1274);
and (n1322,n66,n47);
and (n1323,n1324,n1325);
xor (n1324,n1321,n1322);
or (n1325,n1326,n1329);
and (n1326,n1327,n1328);
xor (n1327,n1279,n1280);
and (n1328,n49,n47);
and (n1329,n1330,n1331);
xor (n1330,n1327,n1328);
or (n1331,n1332,n1335);
and (n1332,n1333,n1334);
xor (n1333,n1285,n1286);
and (n1334,n91,n47);
and (n1335,n1336,n1337);
xor (n1336,n1333,n1334);
or (n1337,n1338,n1341);
and (n1338,n1339,n1340);
xor (n1339,n1291,n1292);
and (n1340,n86,n47);
and (n1341,n1342,n1343);
xor (n1342,n1339,n1340);
or (n1343,n1344,n1347);
and (n1344,n1345,n1346);
xor (n1345,n1297,n1298);
and (n1346,n141,n47);
and (n1347,n1348,n1349);
xor (n1348,n1345,n1346);
or (n1349,n1350,n1353);
and (n1350,n1351,n1352);
xor (n1351,n1303,n1304);
and (n1352,n135,n47);
and (n1353,n1354,n1355);
xor (n1354,n1351,n1352);
or (n1355,n1356,n1358);
and (n1356,n1357,n604);
xor (n1357,n1309,n1310);
and (n1358,n1359,n1360);
xor (n1359,n1357,n604);
and (n1360,n1361,n1362);
xor (n1361,n1315,n1316);
and (n1362,n160,n47);
and (n1363,n66,n74);
or (n1364,n1365,n1368);
and (n1365,n1366,n1367);
xor (n1366,n1324,n1325);
and (n1367,n49,n74);
and (n1368,n1369,n1370);
xor (n1369,n1366,n1367);
or (n1370,n1371,n1374);
and (n1371,n1372,n1373);
xor (n1372,n1330,n1331);
and (n1373,n91,n74);
and (n1374,n1375,n1376);
xor (n1375,n1372,n1373);
or (n1376,n1377,n1380);
and (n1377,n1378,n1379);
xor (n1378,n1336,n1337);
and (n1379,n86,n74);
and (n1380,n1381,n1382);
xor (n1381,n1378,n1379);
or (n1382,n1383,n1386);
and (n1383,n1384,n1385);
xor (n1384,n1342,n1343);
and (n1385,n141,n74);
and (n1386,n1387,n1388);
xor (n1387,n1384,n1385);
or (n1388,n1389,n1392);
and (n1389,n1390,n1391);
xor (n1390,n1348,n1349);
and (n1391,n135,n74);
and (n1392,n1393,n1394);
xor (n1393,n1390,n1391);
or (n1394,n1395,n1398);
and (n1395,n1396,n1397);
xor (n1396,n1354,n1355);
and (n1397,n165,n74);
and (n1398,n1399,n1400);
xor (n1399,n1396,n1397);
and (n1400,n1401,n1402);
xor (n1401,n1359,n1360);
not (n1402,n580);
and (n1403,n49,n80);
or (n1404,n1405,n1408);
and (n1405,n1406,n1407);
xor (n1406,n1369,n1370);
and (n1407,n91,n80);
and (n1408,n1409,n1410);
xor (n1409,n1406,n1407);
or (n1410,n1411,n1413);
and (n1411,n1412,n87);
xor (n1412,n1375,n1376);
and (n1413,n1414,n1415);
xor (n1414,n1412,n87);
or (n1415,n1416,n1419);
and (n1416,n1417,n1418);
xor (n1417,n1381,n1382);
and (n1418,n141,n80);
and (n1419,n1420,n1421);
xor (n1420,n1417,n1418);
or (n1421,n1422,n1424);
and (n1422,n1423,n347);
xor (n1423,n1387,n1388);
and (n1424,n1425,n1426);
xor (n1425,n1423,n347);
or (n1426,n1427,n1430);
and (n1427,n1428,n1429);
xor (n1428,n1393,n1394);
and (n1429,n165,n80);
and (n1430,n1431,n1432);
xor (n1431,n1428,n1429);
and (n1432,n1433,n1434);
xor (n1433,n1399,n1400);
and (n1434,n160,n80);
and (n1435,n91,n125);
or (n1436,n1437,n1440);
and (n1437,n1438,n1439);
xor (n1438,n1409,n1410);
and (n1439,n86,n125);
and (n1440,n1441,n1442);
xor (n1441,n1438,n1439);
or (n1442,n1443,n1446);
and (n1443,n1444,n1445);
xor (n1444,n1414,n1415);
and (n1445,n141,n125);
and (n1446,n1447,n1448);
xor (n1447,n1444,n1445);
or (n1448,n1449,n1452);
and (n1449,n1450,n1451);
xor (n1450,n1420,n1421);
and (n1451,n135,n125);
and (n1452,n1453,n1454);
xor (n1453,n1450,n1451);
or (n1454,n1455,n1458);
and (n1455,n1456,n1457);
xor (n1456,n1425,n1426);
and (n1457,n165,n125);
and (n1458,n1459,n1460);
xor (n1459,n1456,n1457);
and (n1460,n1461,n330);
xor (n1461,n1431,n1432);
and (n1462,n86,n131);
or (n1463,n1464,n1467);
and (n1464,n1465,n1466);
xor (n1465,n1441,n1442);
and (n1466,n141,n131);
and (n1467,n1468,n1469);
xor (n1468,n1465,n1466);
or (n1469,n1470,n1473);
and (n1470,n1471,n1472);
xor (n1471,n1447,n1448);
and (n1472,n135,n131);
and (n1473,n1474,n1475);
xor (n1474,n1471,n1472);
or (n1475,n1476,n1479);
and (n1476,n1477,n1478);
xor (n1477,n1453,n1454);
and (n1478,n165,n131);
and (n1479,n1480,n1481);
xor (n1480,n1477,n1478);
and (n1481,n1482,n1483);
xor (n1482,n1459,n1460);
and (n1483,n160,n131);
and (n1484,n141,n150);
or (n1485,n1486,n1489);
and (n1486,n1487,n1488);
xor (n1487,n1468,n1469);
and (n1488,n135,n150);
and (n1489,n1490,n1491);
xor (n1490,n1487,n1488);
or (n1491,n1492,n1495);
and (n1492,n1493,n1494);
xor (n1493,n1474,n1475);
and (n1494,n165,n150);
and (n1495,n1496,n1497);
xor (n1496,n1493,n1494);
and (n1497,n1498,n1499);
xor (n1498,n1480,n1481);
not (n1499,n245);
and (n1500,n135,n151);
or (n1501,n1502,n1505);
and (n1502,n1503,n1504);
xor (n1503,n1490,n1491);
and (n1504,n165,n151);
and (n1505,n1506,n1507);
xor (n1506,n1503,n1504);
and (n1507,n1508,n1509);
xor (n1508,n1496,n1497);
and (n1509,n160,n151);
and (n1510,n165,n174);
and (n1511,n1512,n1513);
xor (n1512,n1506,n1507);
not (n1513,n437);
and (n1514,n160,n402);
endmodule
