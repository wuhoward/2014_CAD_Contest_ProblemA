module top (out,n23,n24,n28,n30,n37,n44,n51,n58,n65
        ,n72,n79,n86,n93,n99,n101,n168,n235,n302,n369
        ,n436,n503,n570,n637,n702,n782,n783,n787,n789,n796
        ,n803,n810,n817,n824,n831,n838,n845,n852,n858,n860
        ,n927,n994,n1061,n1128,n1195,n1262,n1329,n1396,n1461,n1519);
output out;
input n23;
input n24;
input n28;
input n30;
input n37;
input n44;
input n51;
input n58;
input n65;
input n72;
input n79;
input n86;
input n93;
input n99;
input n101;
input n168;
input n235;
input n302;
input n369;
input n436;
input n503;
input n570;
input n637;
input n702;
input n782;
input n783;
input n787;
input n789;
input n796;
input n803;
input n810;
input n817;
input n824;
input n831;
input n838;
input n845;
input n852;
input n858;
input n860;
input n927;
input n994;
input n1061;
input n1128;
input n1195;
input n1262;
input n1329;
input n1396;
input n1461;
input n1519;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n25;
wire n26;
wire n27;
wire n29;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n100;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n784;
wire n785;
wire n786;
wire n788;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n859;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
xor (out,n0,n1520);
wire s0n0,s1n0,notn0;
or (n0,s0n0,s1n0);
not(notn0,n1519);
and (s0n0,notn0,n1);
and (s1n0,n1519,n760);
xor (n1,n2,n703);
xor (n2,n3,n701);
xor (n3,n4,n638);
xor (n4,n5,n636);
or (n5,n6,n571);
and (n6,n7,n569);
or (n7,n8,n504);
and (n8,n9,n502);
or (n9,n10,n437);
and (n10,n11,n435);
or (n11,n12,n370);
and (n12,n13,n368);
or (n13,n14,n303);
and (n14,n15,n301);
or (n15,n16,n236);
and (n16,n17,n234);
or (n17,n18,n169);
and (n18,n19,n167);
or (n19,n20,n102);
and (n20,n21,n100);
and (n21,n22,n25);
and (n22,n23,n24);
or (n25,n26,n31);
and (n26,n27,n29);
and (n27,n23,n28);
and (n29,n30,n24);
and (n31,n32,n33);
xor (n32,n27,n29);
or (n33,n34,n38);
and (n34,n35,n36);
and (n35,n30,n28);
and (n36,n37,n24);
and (n38,n39,n40);
xor (n39,n35,n36);
or (n40,n41,n45);
and (n41,n42,n43);
and (n42,n37,n28);
and (n43,n44,n24);
and (n45,n46,n47);
xor (n46,n42,n43);
or (n47,n48,n52);
and (n48,n49,n50);
and (n49,n44,n28);
and (n50,n51,n24);
and (n52,n53,n54);
xor (n53,n49,n50);
or (n54,n55,n59);
and (n55,n56,n57);
and (n56,n51,n28);
and (n57,n58,n24);
and (n59,n60,n61);
xor (n60,n56,n57);
or (n61,n62,n66);
and (n62,n63,n64);
and (n63,n58,n28);
and (n64,n65,n24);
and (n66,n67,n68);
xor (n67,n63,n64);
or (n68,n69,n73);
and (n69,n70,n71);
and (n70,n65,n28);
and (n71,n72,n24);
and (n73,n74,n75);
xor (n74,n70,n71);
or (n75,n76,n80);
and (n76,n77,n78);
and (n77,n72,n28);
and (n78,n79,n24);
and (n80,n81,n82);
xor (n81,n77,n78);
or (n82,n83,n87);
and (n83,n84,n85);
and (n84,n79,n28);
and (n85,n86,n24);
and (n87,n88,n89);
xor (n88,n84,n85);
or (n89,n90,n94);
and (n90,n91,n92);
and (n91,n86,n28);
and (n92,n93,n24);
and (n94,n95,n96);
xor (n95,n91,n92);
and (n96,n97,n98);
and (n97,n93,n28);
and (n98,n99,n24);
and (n100,n23,n101);
and (n102,n103,n104);
xor (n103,n21,n100);
or (n104,n105,n108);
and (n105,n106,n107);
xor (n106,n22,n25);
and (n107,n30,n101);
and (n108,n109,n110);
xor (n109,n106,n107);
or (n110,n111,n114);
and (n111,n112,n113);
xor (n112,n32,n33);
and (n113,n37,n101);
and (n114,n115,n116);
xor (n115,n112,n113);
or (n116,n117,n120);
and (n117,n118,n119);
xor (n118,n39,n40);
and (n119,n44,n101);
and (n120,n121,n122);
xor (n121,n118,n119);
or (n122,n123,n126);
and (n123,n124,n125);
xor (n124,n46,n47);
and (n125,n51,n101);
and (n126,n127,n128);
xor (n127,n124,n125);
or (n128,n129,n132);
and (n129,n130,n131);
xor (n130,n53,n54);
and (n131,n58,n101);
and (n132,n133,n134);
xor (n133,n130,n131);
or (n134,n135,n138);
and (n135,n136,n137);
xor (n136,n60,n61);
and (n137,n65,n101);
and (n138,n139,n140);
xor (n139,n136,n137);
or (n140,n141,n144);
and (n141,n142,n143);
xor (n142,n67,n68);
and (n143,n72,n101);
and (n144,n145,n146);
xor (n145,n142,n143);
or (n146,n147,n150);
and (n147,n148,n149);
xor (n148,n74,n75);
and (n149,n79,n101);
and (n150,n151,n152);
xor (n151,n148,n149);
or (n152,n153,n156);
and (n153,n154,n155);
xor (n154,n81,n82);
and (n155,n86,n101);
and (n156,n157,n158);
xor (n157,n154,n155);
or (n158,n159,n162);
and (n159,n160,n161);
xor (n160,n88,n89);
and (n161,n93,n101);
and (n162,n163,n164);
xor (n163,n160,n161);
and (n164,n165,n166);
xor (n165,n95,n96);
and (n166,n99,n101);
and (n167,n23,n168);
and (n169,n170,n171);
xor (n170,n19,n167);
or (n171,n172,n175);
and (n172,n173,n174);
xor (n173,n103,n104);
and (n174,n30,n168);
and (n175,n176,n177);
xor (n176,n173,n174);
or (n177,n178,n181);
and (n178,n179,n180);
xor (n179,n109,n110);
and (n180,n37,n168);
and (n181,n182,n183);
xor (n182,n179,n180);
or (n183,n184,n187);
and (n184,n185,n186);
xor (n185,n115,n116);
and (n186,n44,n168);
and (n187,n188,n189);
xor (n188,n185,n186);
or (n189,n190,n193);
and (n190,n191,n192);
xor (n191,n121,n122);
and (n192,n51,n168);
and (n193,n194,n195);
xor (n194,n191,n192);
or (n195,n196,n199);
and (n196,n197,n198);
xor (n197,n127,n128);
and (n198,n58,n168);
and (n199,n200,n201);
xor (n200,n197,n198);
or (n201,n202,n205);
and (n202,n203,n204);
xor (n203,n133,n134);
and (n204,n65,n168);
and (n205,n206,n207);
xor (n206,n203,n204);
or (n207,n208,n211);
and (n208,n209,n210);
xor (n209,n139,n140);
and (n210,n72,n168);
and (n211,n212,n213);
xor (n212,n209,n210);
or (n213,n214,n217);
and (n214,n215,n216);
xor (n215,n145,n146);
and (n216,n79,n168);
and (n217,n218,n219);
xor (n218,n215,n216);
or (n219,n220,n223);
and (n220,n221,n222);
xor (n221,n151,n152);
and (n222,n86,n168);
and (n223,n224,n225);
xor (n224,n221,n222);
or (n225,n226,n229);
and (n226,n227,n228);
xor (n227,n157,n158);
and (n228,n93,n168);
and (n229,n230,n231);
xor (n230,n227,n228);
and (n231,n232,n233);
xor (n232,n163,n164);
and (n233,n99,n168);
and (n234,n23,n235);
and (n236,n237,n238);
xor (n237,n17,n234);
or (n238,n239,n242);
and (n239,n240,n241);
xor (n240,n170,n171);
and (n241,n30,n235);
and (n242,n243,n244);
xor (n243,n240,n241);
or (n244,n245,n248);
and (n245,n246,n247);
xor (n246,n176,n177);
and (n247,n37,n235);
and (n248,n249,n250);
xor (n249,n246,n247);
or (n250,n251,n254);
and (n251,n252,n253);
xor (n252,n182,n183);
and (n253,n44,n235);
and (n254,n255,n256);
xor (n255,n252,n253);
or (n256,n257,n260);
and (n257,n258,n259);
xor (n258,n188,n189);
and (n259,n51,n235);
and (n260,n261,n262);
xor (n261,n258,n259);
or (n262,n263,n266);
and (n263,n264,n265);
xor (n264,n194,n195);
and (n265,n58,n235);
and (n266,n267,n268);
xor (n267,n264,n265);
or (n268,n269,n272);
and (n269,n270,n271);
xor (n270,n200,n201);
and (n271,n65,n235);
and (n272,n273,n274);
xor (n273,n270,n271);
or (n274,n275,n278);
and (n275,n276,n277);
xor (n276,n206,n207);
and (n277,n72,n235);
and (n278,n279,n280);
xor (n279,n276,n277);
or (n280,n281,n284);
and (n281,n282,n283);
xor (n282,n212,n213);
and (n283,n79,n235);
and (n284,n285,n286);
xor (n285,n282,n283);
or (n286,n287,n290);
and (n287,n288,n289);
xor (n288,n218,n219);
and (n289,n86,n235);
and (n290,n291,n292);
xor (n291,n288,n289);
or (n292,n293,n296);
and (n293,n294,n295);
xor (n294,n224,n225);
and (n295,n93,n235);
and (n296,n297,n298);
xor (n297,n294,n295);
and (n298,n299,n300);
xor (n299,n230,n231);
and (n300,n99,n235);
and (n301,n23,n302);
and (n303,n304,n305);
xor (n304,n15,n301);
or (n305,n306,n309);
and (n306,n307,n308);
xor (n307,n237,n238);
and (n308,n30,n302);
and (n309,n310,n311);
xor (n310,n307,n308);
or (n311,n312,n315);
and (n312,n313,n314);
xor (n313,n243,n244);
and (n314,n37,n302);
and (n315,n316,n317);
xor (n316,n313,n314);
or (n317,n318,n321);
and (n318,n319,n320);
xor (n319,n249,n250);
and (n320,n44,n302);
and (n321,n322,n323);
xor (n322,n319,n320);
or (n323,n324,n327);
and (n324,n325,n326);
xor (n325,n255,n256);
and (n326,n51,n302);
and (n327,n328,n329);
xor (n328,n325,n326);
or (n329,n330,n333);
and (n330,n331,n332);
xor (n331,n261,n262);
and (n332,n58,n302);
and (n333,n334,n335);
xor (n334,n331,n332);
or (n335,n336,n339);
and (n336,n337,n338);
xor (n337,n267,n268);
and (n338,n65,n302);
and (n339,n340,n341);
xor (n340,n337,n338);
or (n341,n342,n345);
and (n342,n343,n344);
xor (n343,n273,n274);
and (n344,n72,n302);
and (n345,n346,n347);
xor (n346,n343,n344);
or (n347,n348,n351);
and (n348,n349,n350);
xor (n349,n279,n280);
and (n350,n79,n302);
and (n351,n352,n353);
xor (n352,n349,n350);
or (n353,n354,n357);
and (n354,n355,n356);
xor (n355,n285,n286);
and (n356,n86,n302);
and (n357,n358,n359);
xor (n358,n355,n356);
or (n359,n360,n363);
and (n360,n361,n362);
xor (n361,n291,n292);
and (n362,n93,n302);
and (n363,n364,n365);
xor (n364,n361,n362);
and (n365,n366,n367);
xor (n366,n297,n298);
and (n367,n99,n302);
and (n368,n23,n369);
and (n370,n371,n372);
xor (n371,n13,n368);
or (n372,n373,n376);
and (n373,n374,n375);
xor (n374,n304,n305);
and (n375,n30,n369);
and (n376,n377,n378);
xor (n377,n374,n375);
or (n378,n379,n382);
and (n379,n380,n381);
xor (n380,n310,n311);
and (n381,n37,n369);
and (n382,n383,n384);
xor (n383,n380,n381);
or (n384,n385,n388);
and (n385,n386,n387);
xor (n386,n316,n317);
and (n387,n44,n369);
and (n388,n389,n390);
xor (n389,n386,n387);
or (n390,n391,n394);
and (n391,n392,n393);
xor (n392,n322,n323);
and (n393,n51,n369);
and (n394,n395,n396);
xor (n395,n392,n393);
or (n396,n397,n400);
and (n397,n398,n399);
xor (n398,n328,n329);
and (n399,n58,n369);
and (n400,n401,n402);
xor (n401,n398,n399);
or (n402,n403,n406);
and (n403,n404,n405);
xor (n404,n334,n335);
and (n405,n65,n369);
and (n406,n407,n408);
xor (n407,n404,n405);
or (n408,n409,n412);
and (n409,n410,n411);
xor (n410,n340,n341);
and (n411,n72,n369);
and (n412,n413,n414);
xor (n413,n410,n411);
or (n414,n415,n418);
and (n415,n416,n417);
xor (n416,n346,n347);
and (n417,n79,n369);
and (n418,n419,n420);
xor (n419,n416,n417);
or (n420,n421,n424);
and (n421,n422,n423);
xor (n422,n352,n353);
and (n423,n86,n369);
and (n424,n425,n426);
xor (n425,n422,n423);
or (n426,n427,n430);
and (n427,n428,n429);
xor (n428,n358,n359);
and (n429,n93,n369);
and (n430,n431,n432);
xor (n431,n428,n429);
and (n432,n433,n434);
xor (n433,n364,n365);
and (n434,n99,n369);
and (n435,n23,n436);
and (n437,n438,n439);
xor (n438,n11,n435);
or (n439,n440,n443);
and (n440,n441,n442);
xor (n441,n371,n372);
and (n442,n30,n436);
and (n443,n444,n445);
xor (n444,n441,n442);
or (n445,n446,n449);
and (n446,n447,n448);
xor (n447,n377,n378);
and (n448,n37,n436);
and (n449,n450,n451);
xor (n450,n447,n448);
or (n451,n452,n455);
and (n452,n453,n454);
xor (n453,n383,n384);
and (n454,n44,n436);
and (n455,n456,n457);
xor (n456,n453,n454);
or (n457,n458,n461);
and (n458,n459,n460);
xor (n459,n389,n390);
and (n460,n51,n436);
and (n461,n462,n463);
xor (n462,n459,n460);
or (n463,n464,n467);
and (n464,n465,n466);
xor (n465,n395,n396);
and (n466,n58,n436);
and (n467,n468,n469);
xor (n468,n465,n466);
or (n469,n470,n473);
and (n470,n471,n472);
xor (n471,n401,n402);
and (n472,n65,n436);
and (n473,n474,n475);
xor (n474,n471,n472);
or (n475,n476,n479);
and (n476,n477,n478);
xor (n477,n407,n408);
and (n478,n72,n436);
and (n479,n480,n481);
xor (n480,n477,n478);
or (n481,n482,n485);
and (n482,n483,n484);
xor (n483,n413,n414);
and (n484,n79,n436);
and (n485,n486,n487);
xor (n486,n483,n484);
or (n487,n488,n491);
and (n488,n489,n490);
xor (n489,n419,n420);
and (n490,n86,n436);
and (n491,n492,n493);
xor (n492,n489,n490);
or (n493,n494,n497);
and (n494,n495,n496);
xor (n495,n425,n426);
and (n496,n93,n436);
and (n497,n498,n499);
xor (n498,n495,n496);
and (n499,n500,n501);
xor (n500,n431,n432);
and (n501,n99,n436);
and (n502,n23,n503);
and (n504,n505,n506);
xor (n505,n9,n502);
or (n506,n507,n510);
and (n507,n508,n509);
xor (n508,n438,n439);
and (n509,n30,n503);
and (n510,n511,n512);
xor (n511,n508,n509);
or (n512,n513,n516);
and (n513,n514,n515);
xor (n514,n444,n445);
and (n515,n37,n503);
and (n516,n517,n518);
xor (n517,n514,n515);
or (n518,n519,n522);
and (n519,n520,n521);
xor (n520,n450,n451);
and (n521,n44,n503);
and (n522,n523,n524);
xor (n523,n520,n521);
or (n524,n525,n528);
and (n525,n526,n527);
xor (n526,n456,n457);
and (n527,n51,n503);
and (n528,n529,n530);
xor (n529,n526,n527);
or (n530,n531,n534);
and (n531,n532,n533);
xor (n532,n462,n463);
and (n533,n58,n503);
and (n534,n535,n536);
xor (n535,n532,n533);
or (n536,n537,n540);
and (n537,n538,n539);
xor (n538,n468,n469);
and (n539,n65,n503);
and (n540,n541,n542);
xor (n541,n538,n539);
or (n542,n543,n546);
and (n543,n544,n545);
xor (n544,n474,n475);
and (n545,n72,n503);
and (n546,n547,n548);
xor (n547,n544,n545);
or (n548,n549,n552);
and (n549,n550,n551);
xor (n550,n480,n481);
and (n551,n79,n503);
and (n552,n553,n554);
xor (n553,n550,n551);
or (n554,n555,n558);
and (n555,n556,n557);
xor (n556,n486,n487);
and (n557,n86,n503);
and (n558,n559,n560);
xor (n559,n556,n557);
or (n560,n561,n564);
and (n561,n562,n563);
xor (n562,n492,n493);
and (n563,n93,n503);
and (n564,n565,n566);
xor (n565,n562,n563);
and (n566,n567,n568);
xor (n567,n498,n499);
and (n568,n99,n503);
and (n569,n23,n570);
and (n571,n572,n573);
xor (n572,n7,n569);
or (n573,n574,n577);
and (n574,n575,n576);
xor (n575,n505,n506);
and (n576,n30,n570);
and (n577,n578,n579);
xor (n578,n575,n576);
or (n579,n580,n583);
and (n580,n581,n582);
xor (n581,n511,n512);
and (n582,n37,n570);
and (n583,n584,n585);
xor (n584,n581,n582);
or (n585,n586,n589);
and (n586,n587,n588);
xor (n587,n517,n518);
and (n588,n44,n570);
and (n589,n590,n591);
xor (n590,n587,n588);
or (n591,n592,n595);
and (n592,n593,n594);
xor (n593,n523,n524);
and (n594,n51,n570);
and (n595,n596,n597);
xor (n596,n593,n594);
or (n597,n598,n601);
and (n598,n599,n600);
xor (n599,n529,n530);
and (n600,n58,n570);
and (n601,n602,n603);
xor (n602,n599,n600);
or (n603,n604,n607);
and (n604,n605,n606);
xor (n605,n535,n536);
and (n606,n65,n570);
and (n607,n608,n609);
xor (n608,n605,n606);
or (n609,n610,n613);
and (n610,n611,n612);
xor (n611,n541,n542);
and (n612,n72,n570);
and (n613,n614,n615);
xor (n614,n611,n612);
or (n615,n616,n619);
and (n616,n617,n618);
xor (n617,n547,n548);
and (n618,n79,n570);
and (n619,n620,n621);
xor (n620,n617,n618);
or (n621,n622,n625);
and (n622,n623,n624);
xor (n623,n553,n554);
and (n624,n86,n570);
and (n625,n626,n627);
xor (n626,n623,n624);
or (n627,n628,n631);
and (n628,n629,n630);
xor (n629,n559,n560);
and (n630,n93,n570);
and (n631,n632,n633);
xor (n632,n629,n630);
and (n633,n634,n635);
xor (n634,n565,n566);
and (n635,n99,n570);
and (n636,n23,n637);
or (n638,n639,n642);
and (n639,n640,n641);
xor (n640,n572,n573);
and (n641,n30,n637);
and (n642,n643,n644);
xor (n643,n640,n641);
or (n644,n645,n648);
and (n645,n646,n647);
xor (n646,n578,n579);
and (n647,n37,n637);
and (n648,n649,n650);
xor (n649,n646,n647);
or (n650,n651,n654);
and (n651,n652,n653);
xor (n652,n584,n585);
and (n653,n44,n637);
and (n654,n655,n656);
xor (n655,n652,n653);
or (n656,n657,n660);
and (n657,n658,n659);
xor (n658,n590,n591);
and (n659,n51,n637);
and (n660,n661,n662);
xor (n661,n658,n659);
or (n662,n663,n666);
and (n663,n664,n665);
xor (n664,n596,n597);
and (n665,n58,n637);
and (n666,n667,n668);
xor (n667,n664,n665);
or (n668,n669,n672);
and (n669,n670,n671);
xor (n670,n602,n603);
and (n671,n65,n637);
and (n672,n673,n674);
xor (n673,n670,n671);
or (n674,n675,n678);
and (n675,n676,n677);
xor (n676,n608,n609);
and (n677,n72,n637);
and (n678,n679,n680);
xor (n679,n676,n677);
or (n680,n681,n684);
and (n681,n682,n683);
xor (n682,n614,n615);
and (n683,n79,n637);
and (n684,n685,n686);
xor (n685,n682,n683);
or (n686,n687,n690);
and (n687,n688,n689);
xor (n688,n620,n621);
and (n689,n86,n637);
and (n690,n691,n692);
xor (n691,n688,n689);
or (n692,n693,n696);
and (n693,n694,n695);
xor (n694,n626,n627);
and (n695,n93,n637);
and (n696,n697,n698);
xor (n697,n694,n695);
and (n698,n699,n700);
xor (n699,n632,n633);
and (n700,n99,n637);
and (n701,n30,n702);
or (n703,n704,n707);
and (n704,n705,n706);
xor (n705,n643,n644);
and (n706,n37,n702);
and (n707,n708,n709);
xor (n708,n705,n706);
or (n709,n710,n713);
and (n710,n711,n712);
xor (n711,n649,n650);
and (n712,n44,n702);
and (n713,n714,n715);
xor (n714,n711,n712);
or (n715,n716,n719);
and (n716,n717,n718);
xor (n717,n655,n656);
and (n718,n51,n702);
and (n719,n720,n721);
xor (n720,n717,n718);
or (n721,n722,n725);
and (n722,n723,n724);
xor (n723,n661,n662);
and (n724,n58,n702);
and (n725,n726,n727);
xor (n726,n723,n724);
or (n727,n728,n731);
and (n728,n729,n730);
xor (n729,n667,n668);
and (n730,n65,n702);
and (n731,n732,n733);
xor (n732,n729,n730);
or (n733,n734,n737);
and (n734,n735,n736);
xor (n735,n673,n674);
and (n736,n72,n702);
and (n737,n738,n739);
xor (n738,n735,n736);
or (n739,n740,n743);
and (n740,n741,n742);
xor (n741,n679,n680);
and (n742,n79,n702);
and (n743,n744,n745);
xor (n744,n741,n742);
or (n745,n746,n749);
and (n746,n747,n748);
xor (n747,n685,n686);
and (n748,n86,n702);
and (n749,n750,n751);
xor (n750,n747,n748);
or (n751,n752,n755);
and (n752,n753,n754);
xor (n753,n691,n692);
and (n754,n93,n702);
and (n755,n756,n757);
xor (n756,n753,n754);
and (n757,n758,n759);
xor (n758,n697,n698);
and (n759,n99,n702);
xor (n760,n761,n1462);
xor (n761,n762,n1460);
xor (n762,n763,n1397);
xor (n763,n764,n1395);
or (n764,n765,n1330);
and (n765,n766,n1328);
or (n766,n767,n1263);
and (n767,n768,n1261);
or (n768,n769,n1196);
and (n769,n770,n1194);
or (n770,n771,n1129);
and (n771,n772,n1127);
or (n772,n773,n1062);
and (n773,n774,n1060);
or (n774,n775,n995);
and (n775,n776,n993);
or (n776,n777,n928);
and (n777,n778,n926);
or (n778,n779,n861);
and (n779,n780,n859);
and (n780,n781,n784);
and (n781,n782,n783);
or (n784,n785,n790);
and (n785,n786,n788);
and (n786,n782,n787);
and (n788,n789,n783);
and (n790,n791,n792);
xor (n791,n786,n788);
or (n792,n793,n797);
and (n793,n794,n795);
and (n794,n789,n787);
and (n795,n796,n783);
and (n797,n798,n799);
xor (n798,n794,n795);
or (n799,n800,n804);
and (n800,n801,n802);
and (n801,n796,n787);
and (n802,n803,n783);
and (n804,n805,n806);
xor (n805,n801,n802);
or (n806,n807,n811);
and (n807,n808,n809);
and (n808,n803,n787);
and (n809,n810,n783);
and (n811,n812,n813);
xor (n812,n808,n809);
or (n813,n814,n818);
and (n814,n815,n816);
and (n815,n810,n787);
and (n816,n817,n783);
and (n818,n819,n820);
xor (n819,n815,n816);
or (n820,n821,n825);
and (n821,n822,n823);
and (n822,n817,n787);
and (n823,n824,n783);
and (n825,n826,n827);
xor (n826,n822,n823);
or (n827,n828,n832);
and (n828,n829,n830);
and (n829,n824,n787);
and (n830,n831,n783);
and (n832,n833,n834);
xor (n833,n829,n830);
or (n834,n835,n839);
and (n835,n836,n837);
and (n836,n831,n787);
and (n837,n838,n783);
and (n839,n840,n841);
xor (n840,n836,n837);
or (n841,n842,n846);
and (n842,n843,n844);
and (n843,n838,n787);
and (n844,n845,n783);
and (n846,n847,n848);
xor (n847,n843,n844);
or (n848,n849,n853);
and (n849,n850,n851);
and (n850,n845,n787);
and (n851,n852,n783);
and (n853,n854,n855);
xor (n854,n850,n851);
and (n855,n856,n857);
and (n856,n852,n787);
and (n857,n858,n783);
and (n859,n782,n860);
and (n861,n862,n863);
xor (n862,n780,n859);
or (n863,n864,n867);
and (n864,n865,n866);
xor (n865,n781,n784);
and (n866,n789,n860);
and (n867,n868,n869);
xor (n868,n865,n866);
or (n869,n870,n873);
and (n870,n871,n872);
xor (n871,n791,n792);
and (n872,n796,n860);
and (n873,n874,n875);
xor (n874,n871,n872);
or (n875,n876,n879);
and (n876,n877,n878);
xor (n877,n798,n799);
and (n878,n803,n860);
and (n879,n880,n881);
xor (n880,n877,n878);
or (n881,n882,n885);
and (n882,n883,n884);
xor (n883,n805,n806);
and (n884,n810,n860);
and (n885,n886,n887);
xor (n886,n883,n884);
or (n887,n888,n891);
and (n888,n889,n890);
xor (n889,n812,n813);
and (n890,n817,n860);
and (n891,n892,n893);
xor (n892,n889,n890);
or (n893,n894,n897);
and (n894,n895,n896);
xor (n895,n819,n820);
and (n896,n824,n860);
and (n897,n898,n899);
xor (n898,n895,n896);
or (n899,n900,n903);
and (n900,n901,n902);
xor (n901,n826,n827);
and (n902,n831,n860);
and (n903,n904,n905);
xor (n904,n901,n902);
or (n905,n906,n909);
and (n906,n907,n908);
xor (n907,n833,n834);
and (n908,n838,n860);
and (n909,n910,n911);
xor (n910,n907,n908);
or (n911,n912,n915);
and (n912,n913,n914);
xor (n913,n840,n841);
and (n914,n845,n860);
and (n915,n916,n917);
xor (n916,n913,n914);
or (n917,n918,n921);
and (n918,n919,n920);
xor (n919,n847,n848);
and (n920,n852,n860);
and (n921,n922,n923);
xor (n922,n919,n920);
and (n923,n924,n925);
xor (n924,n854,n855);
and (n925,n858,n860);
and (n926,n782,n927);
and (n928,n929,n930);
xor (n929,n778,n926);
or (n930,n931,n934);
and (n931,n932,n933);
xor (n932,n862,n863);
and (n933,n789,n927);
and (n934,n935,n936);
xor (n935,n932,n933);
or (n936,n937,n940);
and (n937,n938,n939);
xor (n938,n868,n869);
and (n939,n796,n927);
and (n940,n941,n942);
xor (n941,n938,n939);
or (n942,n943,n946);
and (n943,n944,n945);
xor (n944,n874,n875);
and (n945,n803,n927);
and (n946,n947,n948);
xor (n947,n944,n945);
or (n948,n949,n952);
and (n949,n950,n951);
xor (n950,n880,n881);
and (n951,n810,n927);
and (n952,n953,n954);
xor (n953,n950,n951);
or (n954,n955,n958);
and (n955,n956,n957);
xor (n956,n886,n887);
and (n957,n817,n927);
and (n958,n959,n960);
xor (n959,n956,n957);
or (n960,n961,n964);
and (n961,n962,n963);
xor (n962,n892,n893);
and (n963,n824,n927);
and (n964,n965,n966);
xor (n965,n962,n963);
or (n966,n967,n970);
and (n967,n968,n969);
xor (n968,n898,n899);
and (n969,n831,n927);
and (n970,n971,n972);
xor (n971,n968,n969);
or (n972,n973,n976);
and (n973,n974,n975);
xor (n974,n904,n905);
and (n975,n838,n927);
and (n976,n977,n978);
xor (n977,n974,n975);
or (n978,n979,n982);
and (n979,n980,n981);
xor (n980,n910,n911);
and (n981,n845,n927);
and (n982,n983,n984);
xor (n983,n980,n981);
or (n984,n985,n988);
and (n985,n986,n987);
xor (n986,n916,n917);
and (n987,n852,n927);
and (n988,n989,n990);
xor (n989,n986,n987);
and (n990,n991,n992);
xor (n991,n922,n923);
and (n992,n858,n927);
and (n993,n782,n994);
and (n995,n996,n997);
xor (n996,n776,n993);
or (n997,n998,n1001);
and (n998,n999,n1000);
xor (n999,n929,n930);
and (n1000,n789,n994);
and (n1001,n1002,n1003);
xor (n1002,n999,n1000);
or (n1003,n1004,n1007);
and (n1004,n1005,n1006);
xor (n1005,n935,n936);
and (n1006,n796,n994);
and (n1007,n1008,n1009);
xor (n1008,n1005,n1006);
or (n1009,n1010,n1013);
and (n1010,n1011,n1012);
xor (n1011,n941,n942);
and (n1012,n803,n994);
and (n1013,n1014,n1015);
xor (n1014,n1011,n1012);
or (n1015,n1016,n1019);
and (n1016,n1017,n1018);
xor (n1017,n947,n948);
and (n1018,n810,n994);
and (n1019,n1020,n1021);
xor (n1020,n1017,n1018);
or (n1021,n1022,n1025);
and (n1022,n1023,n1024);
xor (n1023,n953,n954);
and (n1024,n817,n994);
and (n1025,n1026,n1027);
xor (n1026,n1023,n1024);
or (n1027,n1028,n1031);
and (n1028,n1029,n1030);
xor (n1029,n959,n960);
and (n1030,n824,n994);
and (n1031,n1032,n1033);
xor (n1032,n1029,n1030);
or (n1033,n1034,n1037);
and (n1034,n1035,n1036);
xor (n1035,n965,n966);
and (n1036,n831,n994);
and (n1037,n1038,n1039);
xor (n1038,n1035,n1036);
or (n1039,n1040,n1043);
and (n1040,n1041,n1042);
xor (n1041,n971,n972);
and (n1042,n838,n994);
and (n1043,n1044,n1045);
xor (n1044,n1041,n1042);
or (n1045,n1046,n1049);
and (n1046,n1047,n1048);
xor (n1047,n977,n978);
and (n1048,n845,n994);
and (n1049,n1050,n1051);
xor (n1050,n1047,n1048);
or (n1051,n1052,n1055);
and (n1052,n1053,n1054);
xor (n1053,n983,n984);
and (n1054,n852,n994);
and (n1055,n1056,n1057);
xor (n1056,n1053,n1054);
and (n1057,n1058,n1059);
xor (n1058,n989,n990);
and (n1059,n858,n994);
and (n1060,n782,n1061);
and (n1062,n1063,n1064);
xor (n1063,n774,n1060);
or (n1064,n1065,n1068);
and (n1065,n1066,n1067);
xor (n1066,n996,n997);
and (n1067,n789,n1061);
and (n1068,n1069,n1070);
xor (n1069,n1066,n1067);
or (n1070,n1071,n1074);
and (n1071,n1072,n1073);
xor (n1072,n1002,n1003);
and (n1073,n796,n1061);
and (n1074,n1075,n1076);
xor (n1075,n1072,n1073);
or (n1076,n1077,n1080);
and (n1077,n1078,n1079);
xor (n1078,n1008,n1009);
and (n1079,n803,n1061);
and (n1080,n1081,n1082);
xor (n1081,n1078,n1079);
or (n1082,n1083,n1086);
and (n1083,n1084,n1085);
xor (n1084,n1014,n1015);
and (n1085,n810,n1061);
and (n1086,n1087,n1088);
xor (n1087,n1084,n1085);
or (n1088,n1089,n1092);
and (n1089,n1090,n1091);
xor (n1090,n1020,n1021);
and (n1091,n817,n1061);
and (n1092,n1093,n1094);
xor (n1093,n1090,n1091);
or (n1094,n1095,n1098);
and (n1095,n1096,n1097);
xor (n1096,n1026,n1027);
and (n1097,n824,n1061);
and (n1098,n1099,n1100);
xor (n1099,n1096,n1097);
or (n1100,n1101,n1104);
and (n1101,n1102,n1103);
xor (n1102,n1032,n1033);
and (n1103,n831,n1061);
and (n1104,n1105,n1106);
xor (n1105,n1102,n1103);
or (n1106,n1107,n1110);
and (n1107,n1108,n1109);
xor (n1108,n1038,n1039);
and (n1109,n838,n1061);
and (n1110,n1111,n1112);
xor (n1111,n1108,n1109);
or (n1112,n1113,n1116);
and (n1113,n1114,n1115);
xor (n1114,n1044,n1045);
and (n1115,n845,n1061);
and (n1116,n1117,n1118);
xor (n1117,n1114,n1115);
or (n1118,n1119,n1122);
and (n1119,n1120,n1121);
xor (n1120,n1050,n1051);
and (n1121,n852,n1061);
and (n1122,n1123,n1124);
xor (n1123,n1120,n1121);
and (n1124,n1125,n1126);
xor (n1125,n1056,n1057);
and (n1126,n858,n1061);
and (n1127,n782,n1128);
and (n1129,n1130,n1131);
xor (n1130,n772,n1127);
or (n1131,n1132,n1135);
and (n1132,n1133,n1134);
xor (n1133,n1063,n1064);
and (n1134,n789,n1128);
and (n1135,n1136,n1137);
xor (n1136,n1133,n1134);
or (n1137,n1138,n1141);
and (n1138,n1139,n1140);
xor (n1139,n1069,n1070);
and (n1140,n796,n1128);
and (n1141,n1142,n1143);
xor (n1142,n1139,n1140);
or (n1143,n1144,n1147);
and (n1144,n1145,n1146);
xor (n1145,n1075,n1076);
and (n1146,n803,n1128);
and (n1147,n1148,n1149);
xor (n1148,n1145,n1146);
or (n1149,n1150,n1153);
and (n1150,n1151,n1152);
xor (n1151,n1081,n1082);
and (n1152,n810,n1128);
and (n1153,n1154,n1155);
xor (n1154,n1151,n1152);
or (n1155,n1156,n1159);
and (n1156,n1157,n1158);
xor (n1157,n1087,n1088);
and (n1158,n817,n1128);
and (n1159,n1160,n1161);
xor (n1160,n1157,n1158);
or (n1161,n1162,n1165);
and (n1162,n1163,n1164);
xor (n1163,n1093,n1094);
and (n1164,n824,n1128);
and (n1165,n1166,n1167);
xor (n1166,n1163,n1164);
or (n1167,n1168,n1171);
and (n1168,n1169,n1170);
xor (n1169,n1099,n1100);
and (n1170,n831,n1128);
and (n1171,n1172,n1173);
xor (n1172,n1169,n1170);
or (n1173,n1174,n1177);
and (n1174,n1175,n1176);
xor (n1175,n1105,n1106);
and (n1176,n838,n1128);
and (n1177,n1178,n1179);
xor (n1178,n1175,n1176);
or (n1179,n1180,n1183);
and (n1180,n1181,n1182);
xor (n1181,n1111,n1112);
and (n1182,n845,n1128);
and (n1183,n1184,n1185);
xor (n1184,n1181,n1182);
or (n1185,n1186,n1189);
and (n1186,n1187,n1188);
xor (n1187,n1117,n1118);
and (n1188,n852,n1128);
and (n1189,n1190,n1191);
xor (n1190,n1187,n1188);
and (n1191,n1192,n1193);
xor (n1192,n1123,n1124);
and (n1193,n858,n1128);
and (n1194,n782,n1195);
and (n1196,n1197,n1198);
xor (n1197,n770,n1194);
or (n1198,n1199,n1202);
and (n1199,n1200,n1201);
xor (n1200,n1130,n1131);
and (n1201,n789,n1195);
and (n1202,n1203,n1204);
xor (n1203,n1200,n1201);
or (n1204,n1205,n1208);
and (n1205,n1206,n1207);
xor (n1206,n1136,n1137);
and (n1207,n796,n1195);
and (n1208,n1209,n1210);
xor (n1209,n1206,n1207);
or (n1210,n1211,n1214);
and (n1211,n1212,n1213);
xor (n1212,n1142,n1143);
and (n1213,n803,n1195);
and (n1214,n1215,n1216);
xor (n1215,n1212,n1213);
or (n1216,n1217,n1220);
and (n1217,n1218,n1219);
xor (n1218,n1148,n1149);
and (n1219,n810,n1195);
and (n1220,n1221,n1222);
xor (n1221,n1218,n1219);
or (n1222,n1223,n1226);
and (n1223,n1224,n1225);
xor (n1224,n1154,n1155);
and (n1225,n817,n1195);
and (n1226,n1227,n1228);
xor (n1227,n1224,n1225);
or (n1228,n1229,n1232);
and (n1229,n1230,n1231);
xor (n1230,n1160,n1161);
and (n1231,n824,n1195);
and (n1232,n1233,n1234);
xor (n1233,n1230,n1231);
or (n1234,n1235,n1238);
and (n1235,n1236,n1237);
xor (n1236,n1166,n1167);
and (n1237,n831,n1195);
and (n1238,n1239,n1240);
xor (n1239,n1236,n1237);
or (n1240,n1241,n1244);
and (n1241,n1242,n1243);
xor (n1242,n1172,n1173);
and (n1243,n838,n1195);
and (n1244,n1245,n1246);
xor (n1245,n1242,n1243);
or (n1246,n1247,n1250);
and (n1247,n1248,n1249);
xor (n1248,n1178,n1179);
and (n1249,n845,n1195);
and (n1250,n1251,n1252);
xor (n1251,n1248,n1249);
or (n1252,n1253,n1256);
and (n1253,n1254,n1255);
xor (n1254,n1184,n1185);
and (n1255,n852,n1195);
and (n1256,n1257,n1258);
xor (n1257,n1254,n1255);
and (n1258,n1259,n1260);
xor (n1259,n1190,n1191);
and (n1260,n858,n1195);
and (n1261,n782,n1262);
and (n1263,n1264,n1265);
xor (n1264,n768,n1261);
or (n1265,n1266,n1269);
and (n1266,n1267,n1268);
xor (n1267,n1197,n1198);
and (n1268,n789,n1262);
and (n1269,n1270,n1271);
xor (n1270,n1267,n1268);
or (n1271,n1272,n1275);
and (n1272,n1273,n1274);
xor (n1273,n1203,n1204);
and (n1274,n796,n1262);
and (n1275,n1276,n1277);
xor (n1276,n1273,n1274);
or (n1277,n1278,n1281);
and (n1278,n1279,n1280);
xor (n1279,n1209,n1210);
and (n1280,n803,n1262);
and (n1281,n1282,n1283);
xor (n1282,n1279,n1280);
or (n1283,n1284,n1287);
and (n1284,n1285,n1286);
xor (n1285,n1215,n1216);
and (n1286,n810,n1262);
and (n1287,n1288,n1289);
xor (n1288,n1285,n1286);
or (n1289,n1290,n1293);
and (n1290,n1291,n1292);
xor (n1291,n1221,n1222);
and (n1292,n817,n1262);
and (n1293,n1294,n1295);
xor (n1294,n1291,n1292);
or (n1295,n1296,n1299);
and (n1296,n1297,n1298);
xor (n1297,n1227,n1228);
and (n1298,n824,n1262);
and (n1299,n1300,n1301);
xor (n1300,n1297,n1298);
or (n1301,n1302,n1305);
and (n1302,n1303,n1304);
xor (n1303,n1233,n1234);
and (n1304,n831,n1262);
and (n1305,n1306,n1307);
xor (n1306,n1303,n1304);
or (n1307,n1308,n1311);
and (n1308,n1309,n1310);
xor (n1309,n1239,n1240);
and (n1310,n838,n1262);
and (n1311,n1312,n1313);
xor (n1312,n1309,n1310);
or (n1313,n1314,n1317);
and (n1314,n1315,n1316);
xor (n1315,n1245,n1246);
and (n1316,n845,n1262);
and (n1317,n1318,n1319);
xor (n1318,n1315,n1316);
or (n1319,n1320,n1323);
and (n1320,n1321,n1322);
xor (n1321,n1251,n1252);
and (n1322,n852,n1262);
and (n1323,n1324,n1325);
xor (n1324,n1321,n1322);
and (n1325,n1326,n1327);
xor (n1326,n1257,n1258);
and (n1327,n858,n1262);
and (n1328,n782,n1329);
and (n1330,n1331,n1332);
xor (n1331,n766,n1328);
or (n1332,n1333,n1336);
and (n1333,n1334,n1335);
xor (n1334,n1264,n1265);
and (n1335,n789,n1329);
and (n1336,n1337,n1338);
xor (n1337,n1334,n1335);
or (n1338,n1339,n1342);
and (n1339,n1340,n1341);
xor (n1340,n1270,n1271);
and (n1341,n796,n1329);
and (n1342,n1343,n1344);
xor (n1343,n1340,n1341);
or (n1344,n1345,n1348);
and (n1345,n1346,n1347);
xor (n1346,n1276,n1277);
and (n1347,n803,n1329);
and (n1348,n1349,n1350);
xor (n1349,n1346,n1347);
or (n1350,n1351,n1354);
and (n1351,n1352,n1353);
xor (n1352,n1282,n1283);
and (n1353,n810,n1329);
and (n1354,n1355,n1356);
xor (n1355,n1352,n1353);
or (n1356,n1357,n1360);
and (n1357,n1358,n1359);
xor (n1358,n1288,n1289);
and (n1359,n817,n1329);
and (n1360,n1361,n1362);
xor (n1361,n1358,n1359);
or (n1362,n1363,n1366);
and (n1363,n1364,n1365);
xor (n1364,n1294,n1295);
and (n1365,n824,n1329);
and (n1366,n1367,n1368);
xor (n1367,n1364,n1365);
or (n1368,n1369,n1372);
and (n1369,n1370,n1371);
xor (n1370,n1300,n1301);
and (n1371,n831,n1329);
and (n1372,n1373,n1374);
xor (n1373,n1370,n1371);
or (n1374,n1375,n1378);
and (n1375,n1376,n1377);
xor (n1376,n1306,n1307);
and (n1377,n838,n1329);
and (n1378,n1379,n1380);
xor (n1379,n1376,n1377);
or (n1380,n1381,n1384);
and (n1381,n1382,n1383);
xor (n1382,n1312,n1313);
and (n1383,n845,n1329);
and (n1384,n1385,n1386);
xor (n1385,n1382,n1383);
or (n1386,n1387,n1390);
and (n1387,n1388,n1389);
xor (n1388,n1318,n1319);
and (n1389,n852,n1329);
and (n1390,n1391,n1392);
xor (n1391,n1388,n1389);
and (n1392,n1393,n1394);
xor (n1393,n1324,n1325);
and (n1394,n858,n1329);
and (n1395,n782,n1396);
or (n1397,n1398,n1401);
and (n1398,n1399,n1400);
xor (n1399,n1331,n1332);
and (n1400,n789,n1396);
and (n1401,n1402,n1403);
xor (n1402,n1399,n1400);
or (n1403,n1404,n1407);
and (n1404,n1405,n1406);
xor (n1405,n1337,n1338);
and (n1406,n796,n1396);
and (n1407,n1408,n1409);
xor (n1408,n1405,n1406);
or (n1409,n1410,n1413);
and (n1410,n1411,n1412);
xor (n1411,n1343,n1344);
and (n1412,n803,n1396);
and (n1413,n1414,n1415);
xor (n1414,n1411,n1412);
or (n1415,n1416,n1419);
and (n1416,n1417,n1418);
xor (n1417,n1349,n1350);
and (n1418,n810,n1396);
and (n1419,n1420,n1421);
xor (n1420,n1417,n1418);
or (n1421,n1422,n1425);
and (n1422,n1423,n1424);
xor (n1423,n1355,n1356);
and (n1424,n817,n1396);
and (n1425,n1426,n1427);
xor (n1426,n1423,n1424);
or (n1427,n1428,n1431);
and (n1428,n1429,n1430);
xor (n1429,n1361,n1362);
and (n1430,n824,n1396);
and (n1431,n1432,n1433);
xor (n1432,n1429,n1430);
or (n1433,n1434,n1437);
and (n1434,n1435,n1436);
xor (n1435,n1367,n1368);
and (n1436,n831,n1396);
and (n1437,n1438,n1439);
xor (n1438,n1435,n1436);
or (n1439,n1440,n1443);
and (n1440,n1441,n1442);
xor (n1441,n1373,n1374);
and (n1442,n838,n1396);
and (n1443,n1444,n1445);
xor (n1444,n1441,n1442);
or (n1445,n1446,n1449);
and (n1446,n1447,n1448);
xor (n1447,n1379,n1380);
and (n1448,n845,n1396);
and (n1449,n1450,n1451);
xor (n1450,n1447,n1448);
or (n1451,n1452,n1455);
and (n1452,n1453,n1454);
xor (n1453,n1385,n1386);
and (n1454,n852,n1396);
and (n1455,n1456,n1457);
xor (n1456,n1453,n1454);
and (n1457,n1458,n1459);
xor (n1458,n1391,n1392);
and (n1459,n858,n1396);
and (n1460,n789,n1461);
or (n1462,n1463,n1466);
and (n1463,n1464,n1465);
xor (n1464,n1402,n1403);
and (n1465,n796,n1461);
and (n1466,n1467,n1468);
xor (n1467,n1464,n1465);
or (n1468,n1469,n1472);
and (n1469,n1470,n1471);
xor (n1470,n1408,n1409);
and (n1471,n803,n1461);
and (n1472,n1473,n1474);
xor (n1473,n1470,n1471);
or (n1474,n1475,n1478);
and (n1475,n1476,n1477);
xor (n1476,n1414,n1415);
and (n1477,n810,n1461);
and (n1478,n1479,n1480);
xor (n1479,n1476,n1477);
or (n1480,n1481,n1484);
and (n1481,n1482,n1483);
xor (n1482,n1420,n1421);
and (n1483,n817,n1461);
and (n1484,n1485,n1486);
xor (n1485,n1482,n1483);
or (n1486,n1487,n1490);
and (n1487,n1488,n1489);
xor (n1488,n1426,n1427);
and (n1489,n824,n1461);
and (n1490,n1491,n1492);
xor (n1491,n1488,n1489);
or (n1492,n1493,n1496);
and (n1493,n1494,n1495);
xor (n1494,n1432,n1433);
and (n1495,n831,n1461);
and (n1496,n1497,n1498);
xor (n1497,n1494,n1495);
or (n1498,n1499,n1502);
and (n1499,n1500,n1501);
xor (n1500,n1438,n1439);
and (n1501,n838,n1461);
and (n1502,n1503,n1504);
xor (n1503,n1500,n1501);
or (n1504,n1505,n1508);
and (n1505,n1506,n1507);
xor (n1506,n1444,n1445);
and (n1507,n845,n1461);
and (n1508,n1509,n1510);
xor (n1509,n1506,n1507);
or (n1510,n1511,n1514);
and (n1511,n1512,n1513);
xor (n1512,n1450,n1451);
and (n1513,n852,n1461);
and (n1514,n1515,n1516);
xor (n1515,n1512,n1513);
and (n1516,n1517,n1518);
xor (n1517,n1456,n1457);
and (n1518,n858,n1461);
xor (n1520,n1521,n2222);
xor (n1521,n1522,n2220);
xor (n1522,n1523,n2157);
xor (n1523,n1524,n2155);
or (n1524,n1525,n2090);
and (n1525,n1526,n2088);
or (n1526,n1527,n2023);
and (n1527,n1528,n2021);
or (n1528,n1529,n1956);
and (n1529,n1530,n1954);
or (n1530,n1531,n1889);
and (n1531,n1532,n1887);
or (n1532,n1533,n1822);
and (n1533,n1534,n1820);
or (n1534,n1535,n1755);
and (n1535,n1536,n1753);
or (n1536,n1537,n1688);
and (n1537,n1538,n1686);
or (n1538,n1539,n1621);
and (n1539,n1540,n1619);
and (n1540,n1541,n1544);
and (n1541,n1542,n1543);
wire s0n1542,s1n1542,notn1542;
or (n1542,s0n1542,s1n1542);
not(notn1542,n1519);
and (s0n1542,notn1542,n23);
and (s1n1542,n1519,n782);
wire s0n1543,s1n1543,notn1543;
or (n1543,s0n1543,s1n1543);
not(notn1543,n1519);
and (s0n1543,notn1543,n24);
and (s1n1543,n1519,n783);
or (n1544,n1545,n1550);
and (n1545,n1546,n1548);
and (n1546,n1542,n1547);
wire s0n1547,s1n1547,notn1547;
or (n1547,s0n1547,s1n1547);
not(notn1547,n1519);
and (s0n1547,notn1547,n28);
and (s1n1547,n1519,n787);
and (n1548,n1549,n1543);
wire s0n1549,s1n1549,notn1549;
or (n1549,s0n1549,s1n1549);
not(notn1549,n1519);
and (s0n1549,notn1549,n30);
and (s1n1549,n1519,n789);
and (n1550,n1551,n1552);
xor (n1551,n1546,n1548);
or (n1552,n1553,n1557);
and (n1553,n1554,n1555);
and (n1554,n1549,n1547);
and (n1555,n1556,n1543);
wire s0n1556,s1n1556,notn1556;
or (n1556,s0n1556,s1n1556);
not(notn1556,n1519);
and (s0n1556,notn1556,n37);
and (s1n1556,n1519,n796);
and (n1557,n1558,n1559);
xor (n1558,n1554,n1555);
or (n1559,n1560,n1564);
and (n1560,n1561,n1562);
and (n1561,n1556,n1547);
and (n1562,n1563,n1543);
wire s0n1563,s1n1563,notn1563;
or (n1563,s0n1563,s1n1563);
not(notn1563,n1519);
and (s0n1563,notn1563,n44);
and (s1n1563,n1519,n803);
and (n1564,n1565,n1566);
xor (n1565,n1561,n1562);
or (n1566,n1567,n1571);
and (n1567,n1568,n1569);
and (n1568,n1563,n1547);
and (n1569,n1570,n1543);
wire s0n1570,s1n1570,notn1570;
or (n1570,s0n1570,s1n1570);
not(notn1570,n1519);
and (s0n1570,notn1570,n51);
and (s1n1570,n1519,n810);
and (n1571,n1572,n1573);
xor (n1572,n1568,n1569);
or (n1573,n1574,n1578);
and (n1574,n1575,n1576);
and (n1575,n1570,n1547);
and (n1576,n1577,n1543);
wire s0n1577,s1n1577,notn1577;
or (n1577,s0n1577,s1n1577);
not(notn1577,n1519);
and (s0n1577,notn1577,n58);
and (s1n1577,n1519,n817);
and (n1578,n1579,n1580);
xor (n1579,n1575,n1576);
or (n1580,n1581,n1585);
and (n1581,n1582,n1583);
and (n1582,n1577,n1547);
and (n1583,n1584,n1543);
wire s0n1584,s1n1584,notn1584;
or (n1584,s0n1584,s1n1584);
not(notn1584,n1519);
and (s0n1584,notn1584,n65);
and (s1n1584,n1519,n824);
and (n1585,n1586,n1587);
xor (n1586,n1582,n1583);
or (n1587,n1588,n1592);
and (n1588,n1589,n1590);
and (n1589,n1584,n1547);
and (n1590,n1591,n1543);
wire s0n1591,s1n1591,notn1591;
or (n1591,s0n1591,s1n1591);
not(notn1591,n1519);
and (s0n1591,notn1591,n72);
and (s1n1591,n1519,n831);
and (n1592,n1593,n1594);
xor (n1593,n1589,n1590);
or (n1594,n1595,n1599);
and (n1595,n1596,n1597);
and (n1596,n1591,n1547);
and (n1597,n1598,n1543);
wire s0n1598,s1n1598,notn1598;
or (n1598,s0n1598,s1n1598);
not(notn1598,n1519);
and (s0n1598,notn1598,n79);
and (s1n1598,n1519,n838);
and (n1599,n1600,n1601);
xor (n1600,n1596,n1597);
or (n1601,n1602,n1606);
and (n1602,n1603,n1604);
and (n1603,n1598,n1547);
and (n1604,n1605,n1543);
wire s0n1605,s1n1605,notn1605;
or (n1605,s0n1605,s1n1605);
not(notn1605,n1519);
and (s0n1605,notn1605,n86);
and (s1n1605,n1519,n845);
and (n1606,n1607,n1608);
xor (n1607,n1603,n1604);
or (n1608,n1609,n1613);
and (n1609,n1610,n1611);
and (n1610,n1605,n1547);
and (n1611,n1612,n1543);
wire s0n1612,s1n1612,notn1612;
or (n1612,s0n1612,s1n1612);
not(notn1612,n1519);
and (s0n1612,notn1612,n93);
and (s1n1612,n1519,n852);
and (n1613,n1614,n1615);
xor (n1614,n1610,n1611);
and (n1615,n1616,n1617);
and (n1616,n1612,n1547);
and (n1617,n1618,n1543);
wire s0n1618,s1n1618,notn1618;
or (n1618,s0n1618,s1n1618);
not(notn1618,n1519);
and (s0n1618,notn1618,n99);
and (s1n1618,n1519,n858);
and (n1619,n1542,n1620);
wire s0n1620,s1n1620,notn1620;
or (n1620,s0n1620,s1n1620);
not(notn1620,n1519);
and (s0n1620,notn1620,n101);
and (s1n1620,n1519,n860);
and (n1621,n1622,n1623);
xor (n1622,n1540,n1619);
or (n1623,n1624,n1627);
and (n1624,n1625,n1626);
xor (n1625,n1541,n1544);
and (n1626,n1549,n1620);
and (n1627,n1628,n1629);
xor (n1628,n1625,n1626);
or (n1629,n1630,n1633);
and (n1630,n1631,n1632);
xor (n1631,n1551,n1552);
and (n1632,n1556,n1620);
and (n1633,n1634,n1635);
xor (n1634,n1631,n1632);
or (n1635,n1636,n1639);
and (n1636,n1637,n1638);
xor (n1637,n1558,n1559);
and (n1638,n1563,n1620);
and (n1639,n1640,n1641);
xor (n1640,n1637,n1638);
or (n1641,n1642,n1645);
and (n1642,n1643,n1644);
xor (n1643,n1565,n1566);
and (n1644,n1570,n1620);
and (n1645,n1646,n1647);
xor (n1646,n1643,n1644);
or (n1647,n1648,n1651);
and (n1648,n1649,n1650);
xor (n1649,n1572,n1573);
and (n1650,n1577,n1620);
and (n1651,n1652,n1653);
xor (n1652,n1649,n1650);
or (n1653,n1654,n1657);
and (n1654,n1655,n1656);
xor (n1655,n1579,n1580);
and (n1656,n1584,n1620);
and (n1657,n1658,n1659);
xor (n1658,n1655,n1656);
or (n1659,n1660,n1663);
and (n1660,n1661,n1662);
xor (n1661,n1586,n1587);
and (n1662,n1591,n1620);
and (n1663,n1664,n1665);
xor (n1664,n1661,n1662);
or (n1665,n1666,n1669);
and (n1666,n1667,n1668);
xor (n1667,n1593,n1594);
and (n1668,n1598,n1620);
and (n1669,n1670,n1671);
xor (n1670,n1667,n1668);
or (n1671,n1672,n1675);
and (n1672,n1673,n1674);
xor (n1673,n1600,n1601);
and (n1674,n1605,n1620);
and (n1675,n1676,n1677);
xor (n1676,n1673,n1674);
or (n1677,n1678,n1681);
and (n1678,n1679,n1680);
xor (n1679,n1607,n1608);
and (n1680,n1612,n1620);
and (n1681,n1682,n1683);
xor (n1682,n1679,n1680);
and (n1683,n1684,n1685);
xor (n1684,n1614,n1615);
and (n1685,n1618,n1620);
and (n1686,n1542,n1687);
wire s0n1687,s1n1687,notn1687;
or (n1687,s0n1687,s1n1687);
not(notn1687,n1519);
and (s0n1687,notn1687,n168);
and (s1n1687,n1519,n927);
and (n1688,n1689,n1690);
xor (n1689,n1538,n1686);
or (n1690,n1691,n1694);
and (n1691,n1692,n1693);
xor (n1692,n1622,n1623);
and (n1693,n1549,n1687);
and (n1694,n1695,n1696);
xor (n1695,n1692,n1693);
or (n1696,n1697,n1700);
and (n1697,n1698,n1699);
xor (n1698,n1628,n1629);
and (n1699,n1556,n1687);
and (n1700,n1701,n1702);
xor (n1701,n1698,n1699);
or (n1702,n1703,n1706);
and (n1703,n1704,n1705);
xor (n1704,n1634,n1635);
and (n1705,n1563,n1687);
and (n1706,n1707,n1708);
xor (n1707,n1704,n1705);
or (n1708,n1709,n1712);
and (n1709,n1710,n1711);
xor (n1710,n1640,n1641);
and (n1711,n1570,n1687);
and (n1712,n1713,n1714);
xor (n1713,n1710,n1711);
or (n1714,n1715,n1718);
and (n1715,n1716,n1717);
xor (n1716,n1646,n1647);
and (n1717,n1577,n1687);
and (n1718,n1719,n1720);
xor (n1719,n1716,n1717);
or (n1720,n1721,n1724);
and (n1721,n1722,n1723);
xor (n1722,n1652,n1653);
and (n1723,n1584,n1687);
and (n1724,n1725,n1726);
xor (n1725,n1722,n1723);
or (n1726,n1727,n1730);
and (n1727,n1728,n1729);
xor (n1728,n1658,n1659);
and (n1729,n1591,n1687);
and (n1730,n1731,n1732);
xor (n1731,n1728,n1729);
or (n1732,n1733,n1736);
and (n1733,n1734,n1735);
xor (n1734,n1664,n1665);
and (n1735,n1598,n1687);
and (n1736,n1737,n1738);
xor (n1737,n1734,n1735);
or (n1738,n1739,n1742);
and (n1739,n1740,n1741);
xor (n1740,n1670,n1671);
and (n1741,n1605,n1687);
and (n1742,n1743,n1744);
xor (n1743,n1740,n1741);
or (n1744,n1745,n1748);
and (n1745,n1746,n1747);
xor (n1746,n1676,n1677);
and (n1747,n1612,n1687);
and (n1748,n1749,n1750);
xor (n1749,n1746,n1747);
and (n1750,n1751,n1752);
xor (n1751,n1682,n1683);
and (n1752,n1618,n1687);
and (n1753,n1542,n1754);
wire s0n1754,s1n1754,notn1754;
or (n1754,s0n1754,s1n1754);
not(notn1754,n1519);
and (s0n1754,notn1754,n235);
and (s1n1754,n1519,n994);
and (n1755,n1756,n1757);
xor (n1756,n1536,n1753);
or (n1757,n1758,n1761);
and (n1758,n1759,n1760);
xor (n1759,n1689,n1690);
and (n1760,n1549,n1754);
and (n1761,n1762,n1763);
xor (n1762,n1759,n1760);
or (n1763,n1764,n1767);
and (n1764,n1765,n1766);
xor (n1765,n1695,n1696);
and (n1766,n1556,n1754);
and (n1767,n1768,n1769);
xor (n1768,n1765,n1766);
or (n1769,n1770,n1773);
and (n1770,n1771,n1772);
xor (n1771,n1701,n1702);
and (n1772,n1563,n1754);
and (n1773,n1774,n1775);
xor (n1774,n1771,n1772);
or (n1775,n1776,n1779);
and (n1776,n1777,n1778);
xor (n1777,n1707,n1708);
and (n1778,n1570,n1754);
and (n1779,n1780,n1781);
xor (n1780,n1777,n1778);
or (n1781,n1782,n1785);
and (n1782,n1783,n1784);
xor (n1783,n1713,n1714);
and (n1784,n1577,n1754);
and (n1785,n1786,n1787);
xor (n1786,n1783,n1784);
or (n1787,n1788,n1791);
and (n1788,n1789,n1790);
xor (n1789,n1719,n1720);
and (n1790,n1584,n1754);
and (n1791,n1792,n1793);
xor (n1792,n1789,n1790);
or (n1793,n1794,n1797);
and (n1794,n1795,n1796);
xor (n1795,n1725,n1726);
and (n1796,n1591,n1754);
and (n1797,n1798,n1799);
xor (n1798,n1795,n1796);
or (n1799,n1800,n1803);
and (n1800,n1801,n1802);
xor (n1801,n1731,n1732);
and (n1802,n1598,n1754);
and (n1803,n1804,n1805);
xor (n1804,n1801,n1802);
or (n1805,n1806,n1809);
and (n1806,n1807,n1808);
xor (n1807,n1737,n1738);
and (n1808,n1605,n1754);
and (n1809,n1810,n1811);
xor (n1810,n1807,n1808);
or (n1811,n1812,n1815);
and (n1812,n1813,n1814);
xor (n1813,n1743,n1744);
and (n1814,n1612,n1754);
and (n1815,n1816,n1817);
xor (n1816,n1813,n1814);
and (n1817,n1818,n1819);
xor (n1818,n1749,n1750);
and (n1819,n1618,n1754);
and (n1820,n1542,n1821);
wire s0n1821,s1n1821,notn1821;
or (n1821,s0n1821,s1n1821);
not(notn1821,n1519);
and (s0n1821,notn1821,n302);
and (s1n1821,n1519,n1061);
and (n1822,n1823,n1824);
xor (n1823,n1534,n1820);
or (n1824,n1825,n1828);
and (n1825,n1826,n1827);
xor (n1826,n1756,n1757);
and (n1827,n1549,n1821);
and (n1828,n1829,n1830);
xor (n1829,n1826,n1827);
or (n1830,n1831,n1834);
and (n1831,n1832,n1833);
xor (n1832,n1762,n1763);
and (n1833,n1556,n1821);
and (n1834,n1835,n1836);
xor (n1835,n1832,n1833);
or (n1836,n1837,n1840);
and (n1837,n1838,n1839);
xor (n1838,n1768,n1769);
and (n1839,n1563,n1821);
and (n1840,n1841,n1842);
xor (n1841,n1838,n1839);
or (n1842,n1843,n1846);
and (n1843,n1844,n1845);
xor (n1844,n1774,n1775);
and (n1845,n1570,n1821);
and (n1846,n1847,n1848);
xor (n1847,n1844,n1845);
or (n1848,n1849,n1852);
and (n1849,n1850,n1851);
xor (n1850,n1780,n1781);
and (n1851,n1577,n1821);
and (n1852,n1853,n1854);
xor (n1853,n1850,n1851);
or (n1854,n1855,n1858);
and (n1855,n1856,n1857);
xor (n1856,n1786,n1787);
and (n1857,n1584,n1821);
and (n1858,n1859,n1860);
xor (n1859,n1856,n1857);
or (n1860,n1861,n1864);
and (n1861,n1862,n1863);
xor (n1862,n1792,n1793);
and (n1863,n1591,n1821);
and (n1864,n1865,n1866);
xor (n1865,n1862,n1863);
or (n1866,n1867,n1870);
and (n1867,n1868,n1869);
xor (n1868,n1798,n1799);
and (n1869,n1598,n1821);
and (n1870,n1871,n1872);
xor (n1871,n1868,n1869);
or (n1872,n1873,n1876);
and (n1873,n1874,n1875);
xor (n1874,n1804,n1805);
and (n1875,n1605,n1821);
and (n1876,n1877,n1878);
xor (n1877,n1874,n1875);
or (n1878,n1879,n1882);
and (n1879,n1880,n1881);
xor (n1880,n1810,n1811);
and (n1881,n1612,n1821);
and (n1882,n1883,n1884);
xor (n1883,n1880,n1881);
and (n1884,n1885,n1886);
xor (n1885,n1816,n1817);
and (n1886,n1618,n1821);
and (n1887,n1542,n1888);
wire s0n1888,s1n1888,notn1888;
or (n1888,s0n1888,s1n1888);
not(notn1888,n1519);
and (s0n1888,notn1888,n369);
and (s1n1888,n1519,n1128);
and (n1889,n1890,n1891);
xor (n1890,n1532,n1887);
or (n1891,n1892,n1895);
and (n1892,n1893,n1894);
xor (n1893,n1823,n1824);
and (n1894,n1549,n1888);
and (n1895,n1896,n1897);
xor (n1896,n1893,n1894);
or (n1897,n1898,n1901);
and (n1898,n1899,n1900);
xor (n1899,n1829,n1830);
and (n1900,n1556,n1888);
and (n1901,n1902,n1903);
xor (n1902,n1899,n1900);
or (n1903,n1904,n1907);
and (n1904,n1905,n1906);
xor (n1905,n1835,n1836);
and (n1906,n1563,n1888);
and (n1907,n1908,n1909);
xor (n1908,n1905,n1906);
or (n1909,n1910,n1913);
and (n1910,n1911,n1912);
xor (n1911,n1841,n1842);
and (n1912,n1570,n1888);
and (n1913,n1914,n1915);
xor (n1914,n1911,n1912);
or (n1915,n1916,n1919);
and (n1916,n1917,n1918);
xor (n1917,n1847,n1848);
and (n1918,n1577,n1888);
and (n1919,n1920,n1921);
xor (n1920,n1917,n1918);
or (n1921,n1922,n1925);
and (n1922,n1923,n1924);
xor (n1923,n1853,n1854);
and (n1924,n1584,n1888);
and (n1925,n1926,n1927);
xor (n1926,n1923,n1924);
or (n1927,n1928,n1931);
and (n1928,n1929,n1930);
xor (n1929,n1859,n1860);
and (n1930,n1591,n1888);
and (n1931,n1932,n1933);
xor (n1932,n1929,n1930);
or (n1933,n1934,n1937);
and (n1934,n1935,n1936);
xor (n1935,n1865,n1866);
and (n1936,n1598,n1888);
and (n1937,n1938,n1939);
xor (n1938,n1935,n1936);
or (n1939,n1940,n1943);
and (n1940,n1941,n1942);
xor (n1941,n1871,n1872);
and (n1942,n1605,n1888);
and (n1943,n1944,n1945);
xor (n1944,n1941,n1942);
or (n1945,n1946,n1949);
and (n1946,n1947,n1948);
xor (n1947,n1877,n1878);
and (n1948,n1612,n1888);
and (n1949,n1950,n1951);
xor (n1950,n1947,n1948);
and (n1951,n1952,n1953);
xor (n1952,n1883,n1884);
and (n1953,n1618,n1888);
and (n1954,n1542,n1955);
wire s0n1955,s1n1955,notn1955;
or (n1955,s0n1955,s1n1955);
not(notn1955,n1519);
and (s0n1955,notn1955,n436);
and (s1n1955,n1519,n1195);
and (n1956,n1957,n1958);
xor (n1957,n1530,n1954);
or (n1958,n1959,n1962);
and (n1959,n1960,n1961);
xor (n1960,n1890,n1891);
and (n1961,n1549,n1955);
and (n1962,n1963,n1964);
xor (n1963,n1960,n1961);
or (n1964,n1965,n1968);
and (n1965,n1966,n1967);
xor (n1966,n1896,n1897);
and (n1967,n1556,n1955);
and (n1968,n1969,n1970);
xor (n1969,n1966,n1967);
or (n1970,n1971,n1974);
and (n1971,n1972,n1973);
xor (n1972,n1902,n1903);
and (n1973,n1563,n1955);
and (n1974,n1975,n1976);
xor (n1975,n1972,n1973);
or (n1976,n1977,n1980);
and (n1977,n1978,n1979);
xor (n1978,n1908,n1909);
and (n1979,n1570,n1955);
and (n1980,n1981,n1982);
xor (n1981,n1978,n1979);
or (n1982,n1983,n1986);
and (n1983,n1984,n1985);
xor (n1984,n1914,n1915);
and (n1985,n1577,n1955);
and (n1986,n1987,n1988);
xor (n1987,n1984,n1985);
or (n1988,n1989,n1992);
and (n1989,n1990,n1991);
xor (n1990,n1920,n1921);
and (n1991,n1584,n1955);
and (n1992,n1993,n1994);
xor (n1993,n1990,n1991);
or (n1994,n1995,n1998);
and (n1995,n1996,n1997);
xor (n1996,n1926,n1927);
and (n1997,n1591,n1955);
and (n1998,n1999,n2000);
xor (n1999,n1996,n1997);
or (n2000,n2001,n2004);
and (n2001,n2002,n2003);
xor (n2002,n1932,n1933);
and (n2003,n1598,n1955);
and (n2004,n2005,n2006);
xor (n2005,n2002,n2003);
or (n2006,n2007,n2010);
and (n2007,n2008,n2009);
xor (n2008,n1938,n1939);
and (n2009,n1605,n1955);
and (n2010,n2011,n2012);
xor (n2011,n2008,n2009);
or (n2012,n2013,n2016);
and (n2013,n2014,n2015);
xor (n2014,n1944,n1945);
and (n2015,n1612,n1955);
and (n2016,n2017,n2018);
xor (n2017,n2014,n2015);
and (n2018,n2019,n2020);
xor (n2019,n1950,n1951);
and (n2020,n1618,n1955);
and (n2021,n1542,n2022);
wire s0n2022,s1n2022,notn2022;
or (n2022,s0n2022,s1n2022);
not(notn2022,n1519);
and (s0n2022,notn2022,n503);
and (s1n2022,n1519,n1262);
and (n2023,n2024,n2025);
xor (n2024,n1528,n2021);
or (n2025,n2026,n2029);
and (n2026,n2027,n2028);
xor (n2027,n1957,n1958);
and (n2028,n1549,n2022);
and (n2029,n2030,n2031);
xor (n2030,n2027,n2028);
or (n2031,n2032,n2035);
and (n2032,n2033,n2034);
xor (n2033,n1963,n1964);
and (n2034,n1556,n2022);
and (n2035,n2036,n2037);
xor (n2036,n2033,n2034);
or (n2037,n2038,n2041);
and (n2038,n2039,n2040);
xor (n2039,n1969,n1970);
and (n2040,n1563,n2022);
and (n2041,n2042,n2043);
xor (n2042,n2039,n2040);
or (n2043,n2044,n2047);
and (n2044,n2045,n2046);
xor (n2045,n1975,n1976);
and (n2046,n1570,n2022);
and (n2047,n2048,n2049);
xor (n2048,n2045,n2046);
or (n2049,n2050,n2053);
and (n2050,n2051,n2052);
xor (n2051,n1981,n1982);
and (n2052,n1577,n2022);
and (n2053,n2054,n2055);
xor (n2054,n2051,n2052);
or (n2055,n2056,n2059);
and (n2056,n2057,n2058);
xor (n2057,n1987,n1988);
and (n2058,n1584,n2022);
and (n2059,n2060,n2061);
xor (n2060,n2057,n2058);
or (n2061,n2062,n2065);
and (n2062,n2063,n2064);
xor (n2063,n1993,n1994);
and (n2064,n1591,n2022);
and (n2065,n2066,n2067);
xor (n2066,n2063,n2064);
or (n2067,n2068,n2071);
and (n2068,n2069,n2070);
xor (n2069,n1999,n2000);
and (n2070,n1598,n2022);
and (n2071,n2072,n2073);
xor (n2072,n2069,n2070);
or (n2073,n2074,n2077);
and (n2074,n2075,n2076);
xor (n2075,n2005,n2006);
and (n2076,n1605,n2022);
and (n2077,n2078,n2079);
xor (n2078,n2075,n2076);
or (n2079,n2080,n2083);
and (n2080,n2081,n2082);
xor (n2081,n2011,n2012);
and (n2082,n1612,n2022);
and (n2083,n2084,n2085);
xor (n2084,n2081,n2082);
and (n2085,n2086,n2087);
xor (n2086,n2017,n2018);
and (n2087,n1618,n2022);
and (n2088,n1542,n2089);
wire s0n2089,s1n2089,notn2089;
or (n2089,s0n2089,s1n2089);
not(notn2089,n1519);
and (s0n2089,notn2089,n570);
and (s1n2089,n1519,n1329);
and (n2090,n2091,n2092);
xor (n2091,n1526,n2088);
or (n2092,n2093,n2096);
and (n2093,n2094,n2095);
xor (n2094,n2024,n2025);
and (n2095,n1549,n2089);
and (n2096,n2097,n2098);
xor (n2097,n2094,n2095);
or (n2098,n2099,n2102);
and (n2099,n2100,n2101);
xor (n2100,n2030,n2031);
and (n2101,n1556,n2089);
and (n2102,n2103,n2104);
xor (n2103,n2100,n2101);
or (n2104,n2105,n2108);
and (n2105,n2106,n2107);
xor (n2106,n2036,n2037);
and (n2107,n1563,n2089);
and (n2108,n2109,n2110);
xor (n2109,n2106,n2107);
or (n2110,n2111,n2114);
and (n2111,n2112,n2113);
xor (n2112,n2042,n2043);
and (n2113,n1570,n2089);
and (n2114,n2115,n2116);
xor (n2115,n2112,n2113);
or (n2116,n2117,n2120);
and (n2117,n2118,n2119);
xor (n2118,n2048,n2049);
and (n2119,n1577,n2089);
and (n2120,n2121,n2122);
xor (n2121,n2118,n2119);
or (n2122,n2123,n2126);
and (n2123,n2124,n2125);
xor (n2124,n2054,n2055);
and (n2125,n1584,n2089);
and (n2126,n2127,n2128);
xor (n2127,n2124,n2125);
or (n2128,n2129,n2132);
and (n2129,n2130,n2131);
xor (n2130,n2060,n2061);
and (n2131,n1591,n2089);
and (n2132,n2133,n2134);
xor (n2133,n2130,n2131);
or (n2134,n2135,n2138);
and (n2135,n2136,n2137);
xor (n2136,n2066,n2067);
and (n2137,n1598,n2089);
and (n2138,n2139,n2140);
xor (n2139,n2136,n2137);
or (n2140,n2141,n2144);
and (n2141,n2142,n2143);
xor (n2142,n2072,n2073);
and (n2143,n1605,n2089);
and (n2144,n2145,n2146);
xor (n2145,n2142,n2143);
or (n2146,n2147,n2150);
and (n2147,n2148,n2149);
xor (n2148,n2078,n2079);
and (n2149,n1612,n2089);
and (n2150,n2151,n2152);
xor (n2151,n2148,n2149);
and (n2152,n2153,n2154);
xor (n2153,n2084,n2085);
and (n2154,n1618,n2089);
and (n2155,n1542,n2156);
wire s0n2156,s1n2156,notn2156;
or (n2156,s0n2156,s1n2156);
not(notn2156,n1519);
and (s0n2156,notn2156,n637);
and (s1n2156,n1519,n1396);
or (n2157,n2158,n2161);
and (n2158,n2159,n2160);
xor (n2159,n2091,n2092);
and (n2160,n1549,n2156);
and (n2161,n2162,n2163);
xor (n2162,n2159,n2160);
or (n2163,n2164,n2167);
and (n2164,n2165,n2166);
xor (n2165,n2097,n2098);
and (n2166,n1556,n2156);
and (n2167,n2168,n2169);
xor (n2168,n2165,n2166);
or (n2169,n2170,n2173);
and (n2170,n2171,n2172);
xor (n2171,n2103,n2104);
and (n2172,n1563,n2156);
and (n2173,n2174,n2175);
xor (n2174,n2171,n2172);
or (n2175,n2176,n2179);
and (n2176,n2177,n2178);
xor (n2177,n2109,n2110);
and (n2178,n1570,n2156);
and (n2179,n2180,n2181);
xor (n2180,n2177,n2178);
or (n2181,n2182,n2185);
and (n2182,n2183,n2184);
xor (n2183,n2115,n2116);
and (n2184,n1577,n2156);
and (n2185,n2186,n2187);
xor (n2186,n2183,n2184);
or (n2187,n2188,n2191);
and (n2188,n2189,n2190);
xor (n2189,n2121,n2122);
and (n2190,n1584,n2156);
and (n2191,n2192,n2193);
xor (n2192,n2189,n2190);
or (n2193,n2194,n2197);
and (n2194,n2195,n2196);
xor (n2195,n2127,n2128);
and (n2196,n1591,n2156);
and (n2197,n2198,n2199);
xor (n2198,n2195,n2196);
or (n2199,n2200,n2203);
and (n2200,n2201,n2202);
xor (n2201,n2133,n2134);
and (n2202,n1598,n2156);
and (n2203,n2204,n2205);
xor (n2204,n2201,n2202);
or (n2205,n2206,n2209);
and (n2206,n2207,n2208);
xor (n2207,n2139,n2140);
and (n2208,n1605,n2156);
and (n2209,n2210,n2211);
xor (n2210,n2207,n2208);
or (n2211,n2212,n2215);
and (n2212,n2213,n2214);
xor (n2213,n2145,n2146);
and (n2214,n1612,n2156);
and (n2215,n2216,n2217);
xor (n2216,n2213,n2214);
and (n2217,n2218,n2219);
xor (n2218,n2151,n2152);
and (n2219,n1618,n2156);
and (n2220,n1549,n2221);
wire s0n2221,s1n2221,notn2221;
or (n2221,s0n2221,s1n2221);
not(notn2221,n1519);
and (s0n2221,notn2221,n702);
and (s1n2221,n1519,n1461);
or (n2222,n2223,n2226);
and (n2223,n2224,n2225);
xor (n2224,n2162,n2163);
and (n2225,n1556,n2221);
and (n2226,n2227,n2228);
xor (n2227,n2224,n2225);
or (n2228,n2229,n2232);
and (n2229,n2230,n2231);
xor (n2230,n2168,n2169);
and (n2231,n1563,n2221);
and (n2232,n2233,n2234);
xor (n2233,n2230,n2231);
or (n2234,n2235,n2238);
and (n2235,n2236,n2237);
xor (n2236,n2174,n2175);
and (n2237,n1570,n2221);
and (n2238,n2239,n2240);
xor (n2239,n2236,n2237);
or (n2240,n2241,n2244);
and (n2241,n2242,n2243);
xor (n2242,n2180,n2181);
and (n2243,n1577,n2221);
and (n2244,n2245,n2246);
xor (n2245,n2242,n2243);
or (n2246,n2247,n2250);
and (n2247,n2248,n2249);
xor (n2248,n2186,n2187);
and (n2249,n1584,n2221);
and (n2250,n2251,n2252);
xor (n2251,n2248,n2249);
or (n2252,n2253,n2256);
and (n2253,n2254,n2255);
xor (n2254,n2192,n2193);
and (n2255,n1591,n2221);
and (n2256,n2257,n2258);
xor (n2257,n2254,n2255);
or (n2258,n2259,n2262);
and (n2259,n2260,n2261);
xor (n2260,n2198,n2199);
and (n2261,n1598,n2221);
and (n2262,n2263,n2264);
xor (n2263,n2260,n2261);
or (n2264,n2265,n2268);
and (n2265,n2266,n2267);
xor (n2266,n2204,n2205);
and (n2267,n1605,n2221);
and (n2268,n2269,n2270);
xor (n2269,n2266,n2267);
or (n2270,n2271,n2274);
and (n2271,n2272,n2273);
xor (n2272,n2210,n2211);
and (n2273,n1612,n2221);
and (n2274,n2275,n2276);
xor (n2275,n2272,n2273);
and (n2276,n2277,n2278);
xor (n2277,n2216,n2217);
and (n2278,n1618,n2221);
endmodule
