module top (out,n14,n16,n17,n19,n22,n23,n29,n31,n32
        ,n34,n37,n41,n43,n44,n46,n49,n54,n56,n58
        ,n70,n79,n81,n83,n86,n98,n105,n107,n109,n112
        ,n120,n121,n133,n145,n183,n187,n189,n191,n219,n220
        ,n327,n344,n345,n578,n582,n584,n595,n607,n621);
output out;
input n14;
input n16;
input n17;
input n19;
input n22;
input n23;
input n29;
input n31;
input n32;
input n34;
input n37;
input n41;
input n43;
input n44;
input n46;
input n49;
input n54;
input n56;
input n58;
input n70;
input n79;
input n81;
input n83;
input n86;
input n98;
input n105;
input n107;
input n109;
input n112;
input n120;
input n121;
input n133;
input n145;
input n183;
input n187;
input n189;
input n191;
input n219;
input n220;
input n327;
input n344;
input n345;
input n578;
input n582;
input n584;
input n595;
input n607;
input n621;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n15;
wire n18;
wire n20;
wire n21;
wire n24;
wire n25;
wire n26;
wire n27;
wire n28;
wire n30;
wire n33;
wire n35;
wire n36;
wire n38;
wire n39;
wire n40;
wire n42;
wire n45;
wire n47;
wire n48;
wire n50;
wire n51;
wire n52;
wire n53;
wire n55;
wire n57;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n80;
wire n82;
wire n84;
wire n85;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n106;
wire n108;
wire n110;
wire n111;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n184;
wire n185;
wire n186;
wire n188;
wire n190;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n579;
wire n580;
wire n581;
wire n583;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2988;
wire n2989;
wire n2990;
wire n2991;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2996;
wire n2997;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3003;
wire n3004;
wire n3005;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3010;
wire n3011;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3038;
wire n3039;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
wire n3056;
xor (out,n0,n2593);
xnor (n0,n1,n2517);
nand (n1,n2,n557);
nor (n2,n3,n555);
nor (n3,n4,n478);
nand (n4,n5,n398);
nand (n5,n6,n314,n397);
nand (n6,n7,n173);
xor (n7,n8,n137);
xor (n8,n9,n62);
xor (n9,n10,n24);
xor (n10,n11,n23);
xor (n11,n12,n22);
or (n12,n13,n18);
and (n13,n14,n15);
xor (n15,n16,n17);
and (n18,n19,n20);
nor (n20,n15,n21);
xnor (n21,n22,n16);
nand (n24,n25,n50,n61);
nand (n25,n26,n38);
xor (n26,n27,n37);
or (n27,n28,n33);
and (n28,n29,n30);
xor (n30,n31,n32);
and (n33,n34,n35);
nor (n35,n30,n36);
xnor (n36,n37,n31);
xor (n38,n39,n49);
or (n39,n40,n45);
and (n40,n41,n42);
xor (n42,n43,n44);
and (n45,n46,n47);
nor (n47,n42,n48);
xnor (n48,n49,n43);
nand (n50,n51,n38);
xor (n51,n52,n32);
or (n52,n53,n57);
and (n53,n54,n55);
xor (n55,n56,n49);
and (n57,n58,n59);
nor (n59,n55,n60);
xnor (n60,n32,n56);
nand (n61,n26,n51);
nand (n62,n63,n113,n136);
nand (n63,n64,n88);
nand (n64,n65,n75,n87);
nand (n65,n66,n71);
xor (n66,n67,n37);
or (n67,n68,n69);
and (n68,n34,n30);
and (n69,n70,n35);
xor (n71,n72,n49);
or (n72,n73,n74);
and (n73,n46,n42);
and (n74,n54,n47);
nand (n75,n76,n71);
xor (n76,n77,n86);
or (n77,n78,n82);
and (n78,n79,n80);
xor (n80,n81,n37);
and (n82,n83,n84);
nor (n84,n80,n85);
xnor (n85,n86,n81);
nand (n87,n66,n76);
xor (n88,n89,n102);
xor (n89,n90,n94);
xor (n90,n91,n86);
or (n91,n92,n93);
and (n92,n70,n80);
and (n93,n79,n84);
xor (n94,n95,n17);
or (n95,n96,n99);
and (n96,n83,n97);
xor (n97,n98,n86);
and (n99,n14,n100);
nor (n100,n97,n101);
xnor (n101,n17,n98);
xor (n102,n103,n112);
or (n103,n104,n108);
and (n104,n105,n106);
xor (n106,n107,n22);
and (n108,n109,n110);
nor (n110,n106,n111);
xnor (n111,n112,n107);
nand (n113,n114,n88);
nand (n114,n115,n129,n135);
nand (n115,n116,n125);
xor (n116,n117,n44);
or (n117,n118,n122);
and (n118,n41,n119);
xor (n119,n120,n121);
and (n122,n46,n123);
nor (n123,n119,n124);
xnor (n124,n44,n120);
xor (n125,n126,n17);
or (n126,n127,n128);
and (n127,n14,n97);
and (n128,n19,n100);
nand (n129,n130,n125);
xor (n130,n131,n22);
or (n131,n132,n134);
and (n132,n133,n15);
and (n134,n105,n20);
nand (n135,n116,n130);
nand (n136,n64,n114);
xor (n137,n138,n169);
xor (n138,n139,n155);
xor (n139,n140,n151);
xor (n140,n141,n147);
not (n141,n142);
xor (n142,n143,n44);
or (n143,n144,n146);
and (n144,n145,n119);
and (n146,n145,n123);
xor (n147,n148,n49);
or (n148,n149,n150);
and (n149,n145,n42);
and (n150,n41,n47);
xor (n151,n152,n37);
or (n152,n153,n154);
and (n153,n58,n30);
and (n154,n29,n35);
xor (n155,n156,n165);
xor (n156,n157,n161);
xor (n157,n158,n32);
or (n158,n159,n160);
and (n159,n46,n55);
and (n160,n54,n59);
xor (n161,n162,n86);
or (n162,n163,n164);
and (n163,n34,n80);
and (n164,n70,n84);
xor (n165,n166,n17);
or (n166,n167,n168);
and (n167,n79,n97);
and (n168,n83,n100);
nand (n169,n170,n171,n172);
nand (n170,n90,n94);
nand (n171,n102,n94);
nand (n172,n90,n102);
xor (n173,n174,n253);
xor (n174,n175,n233);
nand (n175,n176,n206,n232);
nand (n176,n177,n196);
nand (n177,n178,n194,n195);
nand (n178,n179,n184);
xor (n179,n180,n112);
or (n180,n181,n182);
and (n181,n109,n106);
and (n182,n183,n110);
xor (n184,n185,n23);
or (n185,n186,n190);
and (n186,n187,n188);
xor (n188,n189,n112);
and (n190,n191,n192);
nor (n192,n188,n193);
xnor (n193,n23,n189);
nand (n194,n23,n184);
nand (n195,n179,n23);
xor (n196,n197,n202);
xor (n197,n198,n141);
xor (n198,n199,n23);
or (n199,n200,n201);
and (n200,n183,n188);
and (n201,n187,n192);
xor (n202,n203,n22);
or (n203,n204,n205);
and (n204,n19,n15);
and (n205,n133,n20);
nand (n206,n207,n196);
xor (n207,n208,n230);
xor (n208,n23,n209);
nand (n209,n210,n224,n229);
nand (n210,n211,n214);
xor (n211,n212,n44);
or (n212,n144,n213);
and (n213,n41,n123);
not (n214,n215);
xor (n215,n216,n121);
or (n216,n217,n221);
and (n217,n145,n218);
xor (n218,n219,n220);
and (n221,n145,n222);
nor (n222,n218,n223);
xnor (n223,n121,n219);
nand (n224,n225,n214);
xor (n225,n226,n32);
or (n226,n227,n228);
and (n227,n58,n55);
and (n228,n29,n59);
nand (n229,n211,n225);
xor (n230,n231,n51);
xor (n231,n26,n38);
nand (n232,n177,n207);
xor (n233,n234,n249);
xor (n234,n235,n239);
nand (n235,n236,n237,n238);
nand (n236,n198,n141);
nand (n237,n202,n141);
nand (n238,n198,n202);
xor (n239,n240,n142);
xor (n240,n241,n245);
xor (n241,n242,n112);
or (n242,n243,n244);
and (n243,n133,n106);
and (n244,n105,n110);
xor (n245,n246,n23);
or (n246,n247,n248);
and (n247,n109,n188);
and (n248,n183,n192);
nand (n249,n250,n251,n252);
nand (n250,n23,n209);
nand (n251,n230,n209);
nand (n252,n23,n230);
nand (n253,n254,n310,n313);
nand (n254,n255,n275);
nand (n255,n256,n271,n274);
nand (n256,n257,n269);
nand (n257,n258,n263,n268);
nand (n258,n215,n259);
xor (n259,n260,n32);
or (n260,n261,n262);
and (n261,n29,n55);
and (n262,n34,n59);
nand (n263,n264,n259);
xor (n264,n265,n37);
or (n265,n266,n267);
and (n266,n70,n30);
and (n267,n79,n35);
nand (n268,n215,n264);
xor (n269,n270,n76);
xor (n270,n66,n71);
nand (n271,n272,n269);
xor (n272,n273,n225);
xor (n273,n211,n214);
nand (n274,n257,n272);
nand (n275,n276,n306,n309);
nand (n276,n277,n290);
nand (n277,n278,n284,n289);
nand (n278,n279,n283);
xor (n279,n280,n49);
or (n280,n281,n282);
and (n281,n54,n42);
and (n282,n58,n47);
not (n283,n116);
nand (n284,n285,n283);
xor (n285,n286,n86);
or (n286,n287,n288);
and (n287,n83,n80);
and (n288,n14,n84);
nand (n289,n279,n285);
nand (n290,n291,n300,n305);
nand (n291,n292,n296);
xor (n292,n293,n17);
or (n293,n294,n295);
and (n294,n19,n97);
and (n295,n133,n100);
xor (n296,n297,n22);
or (n297,n298,n299);
and (n298,n105,n15);
and (n299,n109,n20);
nand (n300,n301,n296);
xor (n301,n302,n112);
or (n302,n303,n304);
and (n303,n183,n106);
and (n304,n187,n110);
nand (n305,n292,n301);
nand (n306,n307,n290);
xor (n307,n308,n130);
xor (n308,n116,n125);
nand (n309,n277,n307);
nand (n310,n311,n275);
xor (n311,n312,n114);
xor (n312,n64,n88);
nand (n313,n255,n311);
nand (n314,n315,n173);
nand (n315,n316,n393,n396);
nand (n316,n317,n319);
xor (n317,n318,n207);
xor (n318,n177,n196);
nand (n319,n320,n353,n392);
nand (n320,n321,n351);
nand (n321,n322,n328,n350);
nand (n322,n323,n23);
xor (n323,n324,n23);
or (n324,n325,n326);
and (n325,n191,n188);
and (n326,n327,n192);
nand (n328,n329,n23);
nand (n329,n330,n338,n349);
nand (n330,n331,n334);
xor (n331,n332,n121);
or (n332,n217,n333);
and (n333,n41,n222);
xor (n334,n335,n44);
or (n335,n336,n337);
and (n336,n46,n119);
and (n337,n54,n123);
nand (n338,n339,n334);
not (n339,n340);
xor (n340,n341,n220);
or (n341,n342,n346);
and (n342,n145,n343);
xor (n343,n344,n345);
and (n346,n145,n347);
nor (n347,n343,n348);
xnor (n348,n220,n344);
nand (n349,n331,n339);
nand (n350,n323,n329);
xor (n351,n352,n23);
xor (n352,n179,n184);
nand (n353,n354,n351);
nand (n354,n355,n374,n391);
nand (n355,n356,n372);
nand (n356,n357,n366,n371);
nand (n357,n358,n362);
xor (n358,n359,n49);
or (n359,n360,n361);
and (n360,n58,n42);
and (n361,n29,n47);
xor (n362,n363,n32);
or (n363,n364,n365);
and (n364,n34,n55);
and (n365,n70,n59);
nand (n366,n367,n362);
xor (n367,n368,n37);
or (n368,n369,n370);
and (n369,n79,n30);
and (n370,n83,n35);
nand (n371,n358,n367);
xor (n372,n373,n264);
xor (n373,n215,n259);
nand (n374,n375,n372);
nand (n375,n376,n385,n390);
nand (n376,n377,n381);
xor (n377,n378,n17);
or (n378,n379,n380);
and (n379,n133,n97);
and (n380,n105,n100);
xor (n381,n382,n121);
or (n382,n383,n384);
and (n383,n41,n218);
and (n384,n46,n222);
nand (n385,n386,n381);
xor (n386,n387,n86);
or (n387,n388,n389);
and (n388,n14,n80);
and (n389,n19,n84);
nand (n390,n377,n386);
nand (n391,n356,n375);
nand (n392,n321,n354);
nand (n393,n394,n319);
xor (n394,n395,n311);
xor (n395,n255,n275);
nand (n396,n317,n394);
nand (n397,n7,n315);
xor (n398,n399,n474);
xor (n399,n400,n404);
nand (n400,n401,n402,n403);
nand (n401,n9,n62);
nand (n402,n137,n62);
nand (n403,n9,n137);
xor (n404,n405,n444);
xor (n405,n406,n410);
nand (n406,n407,n408,n409);
nand (n407,n235,n239);
nand (n408,n249,n239);
nand (n409,n235,n249);
xor (n410,n411,n430);
xor (n411,n412,n416);
nand (n412,n413,n414,n415);
nand (n413,n241,n245);
nand (n414,n142,n245);
nand (n415,n241,n142);
xor (n416,n417,n426);
xor (n417,n418,n422);
xor (n418,n419,n22);
or (n419,n420,n421);
and (n420,n83,n15);
and (n421,n14,n20);
xor (n422,n423,n112);
or (n423,n424,n425);
and (n424,n19,n106);
and (n425,n133,n110);
nand (n426,n427,n428,n429);
nand (n427,n141,n147);
nand (n428,n151,n147);
nand (n429,n141,n151);
xor (n430,n431,n440);
xor (n431,n432,n436);
xor (n432,n433,n17);
or (n433,n434,n435);
and (n434,n70,n97);
and (n435,n79,n100);
xor (n436,n437,n23);
or (n437,n438,n439);
and (n438,n105,n188);
and (n439,n109,n192);
not (n440,n441);
xor (n441,n442,n49);
or (n442,n149,n443);
and (n443,n145,n47);
xor (n444,n445,n470);
xor (n445,n446,n450);
nand (n446,n447,n448,n449);
nand (n447,n11,n23);
nand (n448,n24,n23);
nand (n449,n11,n24);
xor (n450,n451,n466);
xor (n451,n23,n452);
xor (n452,n453,n462);
xor (n453,n454,n458);
xor (n454,n455,n32);
or (n455,n456,n457);
and (n456,n41,n55);
and (n457,n46,n59);
xor (n458,n459,n37);
or (n459,n460,n461);
and (n460,n54,n30);
and (n461,n58,n35);
xor (n462,n463,n86);
or (n463,n464,n465);
and (n464,n29,n80);
and (n465,n34,n84);
nand (n466,n467,n468,n469);
nand (n467,n157,n161);
nand (n468,n165,n161);
nand (n469,n157,n165);
nand (n470,n471,n472,n473);
nand (n471,n139,n155);
nand (n472,n169,n155);
nand (n473,n139,n169);
nand (n474,n475,n476,n477);
nand (n475,n175,n233);
nand (n476,n253,n233);
nand (n477,n175,n253);
nor (n478,n479,n483);
nand (n479,n480,n481,n482);
nand (n480,n400,n404);
nand (n481,n474,n404);
nand (n482,n400,n474);
xor (n483,n484,n551);
xor (n484,n485,n511);
xor (n485,n486,n495);
xor (n486,n487,n491);
nand (n487,n488,n489,n490);
nand (n488,n418,n422);
nand (n489,n426,n422);
nand (n490,n418,n426);
nand (n491,n492,n493,n494);
nand (n492,n23,n452);
nand (n493,n466,n452);
nand (n494,n23,n466);
xor (n495,n496,n507);
xor (n496,n23,n497);
xor (n497,n498,n503);
xor (n498,n440,n499);
xor (n499,n500,n32);
or (n500,n501,n502);
and (n501,n145,n55);
and (n502,n41,n59);
xor (n503,n504,n37);
or (n504,n505,n506);
and (n505,n46,n30);
and (n506,n54,n35);
nand (n507,n508,n509,n510);
nand (n508,n454,n458);
nand (n509,n462,n458);
nand (n510,n454,n462);
xor (n511,n512,n547);
xor (n512,n513,n543);
xor (n513,n514,n533);
xor (n514,n515,n519);
nand (n515,n516,n517,n518);
nand (n516,n432,n436);
nand (n517,n440,n436);
nand (n518,n432,n440);
xor (n519,n520,n529);
xor (n520,n521,n525);
xor (n521,n522,n86);
or (n522,n523,n524);
and (n523,n58,n80);
and (n524,n29,n84);
xor (n525,n526,n17);
or (n526,n527,n528);
and (n527,n34,n97);
and (n528,n70,n100);
xor (n529,n530,n23);
or (n530,n531,n532);
and (n531,n133,n188);
and (n532,n105,n192);
xor (n533,n534,n539);
xor (n534,n441,n535);
xor (n535,n536,n22);
or (n536,n537,n538);
and (n537,n79,n15);
and (n538,n83,n20);
xor (n539,n540,n112);
or (n540,n541,n542);
and (n541,n14,n106);
and (n542,n19,n110);
nand (n543,n544,n545,n546);
nand (n544,n412,n416);
nand (n545,n430,n416);
nand (n546,n412,n430);
nand (n547,n548,n549,n550);
nand (n548,n446,n450);
nand (n549,n470,n450);
nand (n550,n446,n470);
nand (n551,n552,n553,n554);
nand (n552,n406,n410);
nand (n553,n444,n410);
nand (n554,n406,n444);
not (n555,n556);
nand (n556,n479,n483);
nand (n557,n558,n560);
nor (n558,n559,n478);
nor (n559,n5,n398);
nand (n560,n561,n2091);
nor (n561,n562,n2059);
nor (n562,n563,n1532);
nor (n563,n564,n1517);
nor (n564,n565,n1238);
nand (n565,n566,n1021);
nor (n566,n567,n920);
nor (n567,n568,n830);
nand (n568,n569,n745,n829);
nand (n569,n570,n647);
xor (n570,n571,n623);
xor (n571,n572,n597);
xor (n572,n573,n585);
xor (n573,n574,n579);
xor (n574,n575,n86);
or (n575,n576,n577);
and (n576,n327,n80);
and (n577,n578,n84);
xor (n579,n580,n17);
or (n580,n581,n583);
and (n581,n582,n97);
and (n583,n584,n100);
xor (n585,n586,n590);
xor (n586,n587,n220);
or (n587,n588,n589);
and (n588,n34,n343);
and (n589,n70,n347);
xnor (n590,n591,n345);
nor (n591,n592,n596);
and (n592,n29,n593);
and (n593,n594,n345);
not (n594,n595);
and (n596,n58,n595);
nand (n597,n598,n608,n622);
nand (n598,n599,n603);
xor (n599,n600,n86);
or (n600,n601,n602);
and (n601,n578,n80);
and (n602,n582,n84);
xor (n603,n604,n17);
or (n604,n605,n606);
and (n605,n584,n97);
and (n606,n607,n100);
nand (n608,n609,n603);
xor (n609,n610,n619);
xor (n610,n611,n615);
xor (n611,n612,n220);
or (n612,n613,n614);
and (n613,n70,n343);
and (n614,n79,n347);
xor (n615,n616,n44);
or (n616,n617,n618);
and (n617,n19,n119);
and (n618,n133,n123);
xnor (n619,n620,n22);
nand (n620,n621,n15);
nand (n622,n599,n609);
xor (n623,n624,n633);
xor (n624,n625,n629);
xor (n625,n626,n22);
or (n626,n627,n628);
and (n627,n607,n15);
and (n628,n621,n20);
nand (n629,n630,n631,n632);
nand (n630,n611,n615);
nand (n631,n619,n615);
nand (n632,n611,n619);
xor (n633,n634,n643);
xor (n634,n635,n639);
xor (n635,n636,n44);
or (n636,n637,n638);
and (n637,n14,n119);
and (n638,n19,n123);
xor (n639,n640,n121);
or (n640,n641,n642);
and (n641,n79,n218);
and (n642,n83,n222);
xor (n643,n644,n49);
or (n644,n645,n646);
and (n645,n133,n42);
and (n646,n105,n47);
nand (n647,n648,n702,n744);
nand (n648,n649,n651);
xor (n649,n650,n609);
xor (n650,n599,n603);
xor (n651,n652,n691);
xor (n652,n653,n669);
nand (n653,n654,n663,n668);
nand (n654,n655,n659);
xor (n655,n656,n44);
or (n656,n657,n658);
and (n657,n133,n119);
and (n658,n105,n123);
xor (n659,n660,n121);
or (n660,n661,n662);
and (n661,n14,n218);
and (n662,n19,n222);
nand (n663,n664,n659);
xor (n664,n665,n49);
or (n665,n666,n667);
and (n666,n109,n42);
and (n667,n183,n47);
nand (n668,n655,n664);
nand (n669,n670,n685,n690);
nand (n670,n671,n680);
xor (n671,n672,n676);
xnor (n672,n673,n345);
nor (n673,n674,n675);
and (n674,n70,n593);
and (n675,n34,n595);
xor (n676,n677,n220);
or (n677,n678,n679);
and (n678,n79,n343);
and (n679,n83,n347);
and (n680,n681,n17);
xnor (n681,n682,n345);
nor (n682,n683,n684);
and (n683,n79,n593);
and (n684,n70,n595);
nand (n685,n686,n680);
xor (n686,n687,n32);
or (n687,n688,n689);
and (n688,n187,n55);
and (n689,n191,n59);
nand (n690,n671,n686);
xor (n691,n692,n698);
xor (n692,n693,n697);
xor (n693,n694,n32);
or (n694,n695,n696);
and (n695,n183,n55);
and (n696,n187,n59);
and (n697,n672,n676);
xor (n698,n699,n37);
or (n699,n700,n701);
and (n700,n191,n30);
and (n701,n327,n35);
nand (n702,n703,n651);
nand (n703,n704,n728,n743);
nand (n704,n705,n726);
nand (n705,n706,n720,n725);
nand (n706,n707,n716);
and (n707,n708,n712);
xnor (n708,n709,n345);
nor (n709,n710,n711);
and (n710,n83,n593);
and (n711,n79,n595);
xor (n712,n713,n220);
or (n713,n714,n715);
and (n714,n14,n343);
and (n715,n19,n347);
xor (n716,n717,n32);
or (n717,n718,n719);
and (n718,n191,n55);
and (n719,n327,n59);
nand (n720,n721,n716);
xor (n721,n722,n37);
or (n722,n723,n724);
and (n723,n578,n30);
and (n724,n582,n35);
nand (n725,n707,n721);
xor (n726,n727,n686);
xor (n727,n671,n680);
nand (n728,n729,n726);
xor (n729,n730,n739);
xor (n730,n731,n735);
xor (n731,n732,n37);
or (n732,n733,n734);
and (n733,n327,n30);
and (n734,n578,n35);
xor (n735,n736,n86);
or (n736,n737,n738);
and (n737,n582,n80);
and (n738,n584,n84);
xor (n739,n740,n17);
or (n740,n741,n742);
and (n741,n607,n97);
and (n742,n621,n100);
nand (n743,n705,n729);
nand (n744,n649,n703);
nand (n745,n746,n647);
xor (n746,n747,n786);
xor (n747,n748,n752);
nand (n748,n749,n750,n751);
nand (n749,n653,n669);
nand (n750,n691,n669);
nand (n751,n653,n691);
xor (n752,n753,n775);
xor (n753,n754,n771);
nand (n754,n755,n765,n770);
nand (n755,n756,n760);
xor (n756,n757,n121);
or (n757,n758,n759);
and (n758,n83,n218);
and (n759,n14,n222);
xor (n760,n761,n22);
xnor (n761,n762,n345);
nor (n762,n763,n764);
and (n763,n34,n593);
and (n764,n29,n595);
nand (n765,n766,n760);
xor (n766,n767,n49);
or (n767,n768,n769);
and (n768,n105,n42);
and (n769,n109,n47);
nand (n770,n756,n766);
nand (n771,n772,n773,n774);
nand (n772,n693,n697);
nand (n773,n698,n697);
nand (n774,n693,n698);
xor (n775,n776,n782);
xor (n776,n777,n778);
and (n777,n761,n22);
xor (n778,n779,n32);
or (n779,n780,n781);
and (n780,n109,n55);
and (n781,n183,n59);
xor (n782,n783,n37);
or (n783,n784,n785);
and (n784,n187,n30);
and (n785,n191,n35);
nand (n786,n787,n794,n828);
nand (n787,n788,n792);
nand (n788,n789,n790,n791);
nand (n789,n731,n735);
nand (n790,n739,n735);
nand (n791,n731,n739);
xor (n792,n793,n766);
xor (n793,n756,n760);
nand (n794,n795,n792);
nand (n795,n796,n813,n827);
nand (n796,n797,n811);
nand (n797,n798,n807,n810);
nand (n798,n799,n803);
xor (n799,n800,n220);
or (n800,n801,n802);
and (n801,n83,n343);
and (n802,n14,n347);
xor (n803,n804,n44);
or (n804,n805,n806);
and (n805,n105,n119);
and (n806,n109,n123);
nand (n807,n808,n803);
xnor (n808,n809,n17);
nand (n809,n621,n97);
nand (n810,n799,n808);
xor (n811,n812,n664);
xor (n812,n655,n659);
nand (n813,n814,n811);
nand (n814,n815,n821,n826);
nand (n815,n816,n820);
xor (n816,n817,n121);
or (n817,n818,n819);
and (n818,n19,n218);
and (n819,n133,n222);
xor (n820,n681,n17);
nand (n821,n822,n820);
xor (n822,n823,n49);
or (n823,n824,n825);
and (n824,n183,n42);
and (n825,n187,n47);
nand (n826,n816,n822);
nand (n827,n797,n814);
nand (n828,n788,n795);
nand (n829,n570,n746);
xor (n830,n831,n916);
xor (n831,n832,n853);
xor (n832,n833,n849);
xor (n833,n834,n845);
xor (n834,n835,n841);
xor (n835,n836,n840);
xor (n836,n837,n17);
or (n837,n838,n839);
and (n838,n578,n97);
and (n839,n582,n100);
and (n840,n586,n590);
xor (n841,n842,n22);
or (n842,n843,n844);
and (n843,n584,n15);
and (n844,n607,n20);
nand (n845,n846,n847,n848);
nand (n846,n625,n629);
nand (n847,n633,n629);
nand (n848,n625,n633);
nand (n849,n850,n851,n852);
nand (n850,n754,n771);
nand (n851,n775,n771);
nand (n852,n754,n775);
xor (n853,n854,n912);
xor (n854,n855,n879);
xor (n855,n856,n875);
xor (n856,n857,n861);
nand (n857,n858,n859,n860);
nand (n858,n777,n778);
nand (n859,n782,n778);
nand (n860,n777,n782);
xor (n861,n862,n871);
xor (n862,n863,n867);
xnor (n863,n864,n345);
nor (n864,n865,n866);
and (n865,n58,n593);
and (n866,n54,n595);
xor (n867,n868,n44);
or (n868,n869,n870);
and (n869,n83,n119);
and (n870,n14,n123);
xor (n871,n872,n121);
or (n872,n873,n874);
and (n873,n70,n218);
and (n874,n79,n222);
nand (n875,n876,n877,n878);
nand (n876,n635,n639);
nand (n877,n643,n639);
nand (n878,n635,n643);
xor (n879,n880,n898);
xor (n880,n881,n885);
nand (n881,n882,n883,n884);
nand (n882,n574,n579);
nand (n883,n585,n579);
nand (n884,n574,n585);
xor (n885,n886,n896);
xor (n886,n887,n891);
xor (n887,n888,n49);
or (n888,n889,n890);
and (n889,n19,n42);
and (n890,n133,n47);
xor (n891,n112,n892);
xor (n892,n893,n220);
or (n893,n894,n895);
and (n894,n29,n343);
and (n895,n34,n347);
xnor (n896,n897,n112);
nand (n897,n621,n106);
xor (n898,n899,n908);
xor (n899,n900,n904);
xor (n900,n901,n32);
or (n901,n902,n903);
and (n902,n105,n55);
and (n903,n109,n59);
xor (n904,n905,n37);
or (n905,n906,n907);
and (n906,n183,n30);
and (n907,n187,n35);
xor (n908,n909,n86);
or (n909,n910,n911);
and (n910,n191,n80);
and (n911,n327,n84);
nand (n912,n913,n914,n915);
nand (n913,n572,n597);
nand (n914,n623,n597);
nand (n915,n572,n623);
nand (n916,n917,n918,n919);
nand (n917,n748,n752);
nand (n918,n786,n752);
nand (n919,n748,n786);
nor (n920,n921,n925);
nand (n921,n922,n923,n924);
nand (n922,n832,n853);
nand (n923,n916,n853);
nand (n924,n832,n916);
xor (n925,n926,n935);
xor (n926,n927,n931);
nand (n927,n928,n929,n930);
nand (n928,n834,n845);
nand (n929,n849,n845);
nand (n930,n834,n849);
nand (n931,n932,n933,n934);
nand (n932,n855,n879);
nand (n933,n912,n879);
nand (n934,n855,n912);
xor (n935,n936,n997);
xor (n936,n937,n968);
xor (n937,n938,n957);
xor (n938,n939,n953);
xor (n939,n940,n949);
xor (n940,n941,n945);
xor (n941,n942,n44);
or (n942,n943,n944);
and (n943,n79,n119);
and (n944,n83,n123);
xor (n945,n946,n121);
or (n946,n947,n948);
and (n947,n34,n218);
and (n948,n70,n222);
xor (n949,n950,n49);
or (n950,n951,n952);
and (n951,n14,n42);
and (n952,n19,n47);
nand (n953,n954,n955,n956);
nand (n954,n887,n891);
nand (n955,n896,n891);
nand (n956,n887,n896);
xor (n957,n958,n964);
xor (n958,n959,n963);
xor (n959,n960,n32);
or (n960,n961,n962);
and (n961,n133,n55);
and (n962,n105,n59);
and (n963,n112,n892);
xor (n964,n965,n37);
or (n965,n966,n967);
and (n966,n109,n30);
and (n967,n183,n35);
xor (n968,n969,n993);
xor (n969,n970,n974);
nand (n970,n971,n972,n973);
nand (n971,n900,n904);
nand (n972,n908,n904);
nand (n973,n900,n908);
xor (n974,n975,n984);
xor (n975,n976,n980);
xor (n976,n977,n86);
or (n977,n978,n979);
and (n978,n187,n80);
and (n979,n191,n84);
xor (n980,n981,n17);
or (n981,n982,n983);
and (n982,n327,n97);
and (n983,n578,n100);
xor (n984,n985,n989);
xnor (n985,n986,n345);
nor (n986,n987,n988);
and (n987,n54,n593);
and (n988,n46,n595);
xor (n989,n990,n220);
or (n990,n991,n992);
and (n991,n58,n343);
and (n992,n29,n347);
nand (n993,n994,n995,n996);
nand (n994,n836,n840);
nand (n995,n841,n840);
nand (n996,n836,n841);
xor (n997,n998,n1017);
xor (n998,n999,n1013);
xor (n999,n1000,n1009);
xor (n1000,n1001,n1005);
xor (n1001,n1002,n22);
or (n1002,n1003,n1004);
and (n1003,n582,n15);
and (n1004,n584,n20);
xor (n1005,n1006,n112);
or (n1006,n1007,n1008);
and (n1007,n607,n106);
and (n1008,n621,n110);
nand (n1009,n1010,n1011,n1012);
nand (n1010,n863,n867);
nand (n1011,n871,n867);
nand (n1012,n863,n871);
nand (n1013,n1014,n1015,n1016);
nand (n1014,n857,n861);
nand (n1015,n875,n861);
nand (n1016,n857,n875);
nand (n1017,n1018,n1019,n1020);
nand (n1018,n881,n885);
nand (n1019,n898,n885);
nand (n1020,n881,n898);
nor (n1021,n1022,n1127);
nor (n1022,n1023,n1027);
nand (n1023,n1024,n1025,n1026);
nand (n1024,n927,n931);
nand (n1025,n935,n931);
nand (n1026,n927,n935);
xor (n1027,n1028,n1123);
xor (n1028,n1029,n1063);
xor (n1029,n1030,n1059);
xor (n1030,n1031,n1035);
nand (n1031,n1032,n1033,n1034);
nand (n1032,n939,n953);
nand (n1033,n957,n953);
nand (n1034,n939,n957);
xor (n1035,n1036,n1045);
xor (n1036,n1037,n1041);
xor (n1037,n1038,n112);
or (n1038,n1039,n1040);
and (n1039,n584,n106);
and (n1040,n607,n110);
nand (n1041,n1042,n1043,n1044);
nand (n1042,n959,n963);
nand (n1043,n964,n963);
nand (n1044,n959,n964);
xor (n1045,n1046,n1055);
xor (n1046,n1047,n1051);
xor (n1047,n1048,n44);
or (n1048,n1049,n1050);
and (n1049,n70,n119);
and (n1050,n79,n123);
xnor (n1051,n1052,n345);
nor (n1052,n1053,n1054);
and (n1053,n46,n593);
and (n1054,n41,n595);
xor (n1055,n1056,n121);
or (n1056,n1057,n1058);
and (n1057,n29,n218);
and (n1058,n34,n222);
nand (n1059,n1060,n1061,n1062);
nand (n1060,n970,n974);
nand (n1061,n993,n974);
nand (n1062,n970,n993);
xor (n1063,n1064,n1119);
xor (n1064,n1065,n1087);
xor (n1065,n1066,n1075);
xor (n1066,n1067,n1071);
nand (n1067,n1068,n1069,n1070);
nand (n1068,n941,n945);
nand (n1069,n949,n945);
nand (n1070,n941,n949);
nand (n1071,n1072,n1073,n1074);
nand (n1072,n976,n980);
nand (n1073,n984,n980);
nand (n1074,n976,n984);
xor (n1075,n1076,n1083);
xor (n1076,n1077,n1081);
xor (n1077,n1078,n49);
or (n1078,n1079,n1080);
and (n1079,n83,n42);
and (n1080,n14,n47);
xnor (n1081,n1082,n23);
nand (n1082,n621,n188);
xor (n1083,n1084,n32);
or (n1084,n1085,n1086);
and (n1085,n19,n55);
and (n1086,n133,n59);
xor (n1087,n1088,n1107);
xor (n1088,n1089,n1093);
nand (n1089,n1090,n1091,n1092);
nand (n1090,n1001,n1005);
nand (n1091,n1009,n1005);
nand (n1092,n1001,n1009);
xor (n1093,n1094,n1103);
xor (n1094,n1095,n1099);
xor (n1095,n1096,n37);
or (n1096,n1097,n1098);
and (n1097,n105,n30);
and (n1098,n109,n35);
xor (n1099,n1100,n86);
or (n1100,n1101,n1102);
and (n1101,n183,n80);
and (n1102,n187,n84);
xor (n1103,n1104,n17);
or (n1104,n1105,n1106);
and (n1105,n191,n97);
and (n1106,n327,n100);
xor (n1107,n1108,n1115);
xor (n1108,n1109,n1114);
xor (n1109,n23,n1110);
xor (n1110,n1111,n220);
or (n1111,n1112,n1113);
and (n1112,n54,n343);
and (n1113,n58,n347);
and (n1114,n985,n989);
xor (n1115,n1116,n22);
or (n1116,n1117,n1118);
and (n1117,n578,n15);
and (n1118,n582,n20);
nand (n1119,n1120,n1121,n1122);
nand (n1120,n999,n1013);
nand (n1121,n1017,n1013);
nand (n1122,n999,n1017);
nand (n1123,n1124,n1125,n1126);
nand (n1124,n937,n968);
nand (n1125,n997,n968);
nand (n1126,n937,n997);
nor (n1127,n1128,n1132);
nand (n1128,n1129,n1130,n1131);
nand (n1129,n1029,n1063);
nand (n1130,n1123,n1063);
nand (n1131,n1029,n1123);
xor (n1132,n1133,n1142);
xor (n1133,n1134,n1138);
nand (n1134,n1135,n1136,n1137);
nand (n1135,n1031,n1035);
nand (n1136,n1059,n1035);
nand (n1137,n1031,n1059);
nand (n1138,n1139,n1140,n1141);
nand (n1139,n1065,n1087);
nand (n1140,n1119,n1087);
nand (n1141,n1065,n1119);
xor (n1142,n1143,n1204);
xor (n1143,n1144,n1168);
xor (n1144,n1145,n1164);
xor (n1145,n1146,n1150);
nand (n1146,n1147,n1148,n1149);
nand (n1147,n1095,n1099);
nand (n1148,n1103,n1099);
nand (n1149,n1095,n1103);
xor (n1150,n1151,n1160);
xor (n1151,n1152,n1156);
xor (n1152,n1153,n32);
or (n1153,n1154,n1155);
and (n1154,n14,n55);
and (n1155,n19,n59);
xor (n1156,n1157,n37);
or (n1157,n1158,n1159);
and (n1158,n133,n30);
and (n1159,n105,n35);
xor (n1160,n1161,n86);
or (n1161,n1162,n1163);
and (n1162,n109,n80);
and (n1163,n183,n84);
nand (n1164,n1165,n1166,n1167);
nand (n1165,n1109,n1114);
nand (n1166,n1115,n1114);
nand (n1167,n1109,n1115);
xor (n1168,n1169,n1190);
xor (n1169,n1170,n1186);
xor (n1170,n1171,n1185);
xor (n1171,n1172,n1176);
xor (n1172,n1173,n17);
or (n1173,n1174,n1175);
and (n1174,n187,n97);
and (n1175,n191,n100);
xor (n1176,n1177,n1181);
xnor (n1177,n1178,n345);
nor (n1178,n1179,n1180);
and (n1179,n41,n593);
and (n1180,n145,n595);
xor (n1181,n1182,n220);
or (n1182,n1183,n1184);
and (n1183,n46,n343);
and (n1184,n54,n347);
and (n1185,n23,n1110);
nand (n1186,n1187,n1188,n1189);
nand (n1187,n1037,n1041);
nand (n1188,n1045,n1041);
nand (n1189,n1037,n1045);
xor (n1190,n1191,n1200);
xor (n1191,n1192,n1196);
xor (n1192,n1193,n22);
or (n1193,n1194,n1195);
and (n1194,n327,n15);
and (n1195,n578,n20);
xor (n1196,n1197,n23);
or (n1197,n1198,n1199);
and (n1198,n607,n188);
and (n1199,n621,n192);
xor (n1200,n1201,n112);
or (n1201,n1202,n1203);
and (n1202,n582,n106);
and (n1203,n584,n110);
xor (n1204,n1205,n1234);
xor (n1205,n1206,n1230);
xor (n1206,n1207,n1226);
xor (n1207,n1208,n1212);
nand (n1208,n1209,n1210,n1211);
nand (n1209,n1047,n1051);
nand (n1210,n1055,n1051);
nand (n1211,n1047,n1055);
xor (n1212,n1213,n1222);
xor (n1213,n1214,n1218);
xor (n1214,n1215,n44);
or (n1215,n1216,n1217);
and (n1216,n34,n119);
and (n1217,n70,n123);
xor (n1218,n1219,n121);
or (n1219,n1220,n1221);
and (n1220,n58,n218);
and (n1221,n29,n222);
xor (n1222,n1223,n49);
or (n1223,n1224,n1225);
and (n1224,n79,n42);
and (n1225,n83,n47);
nand (n1226,n1227,n1228,n1229);
nand (n1227,n1077,n1081);
nand (n1228,n1083,n1081);
nand (n1229,n1077,n1083);
nand (n1230,n1231,n1232,n1233);
nand (n1231,n1067,n1071);
nand (n1232,n1075,n1071);
nand (n1233,n1067,n1075);
nand (n1234,n1235,n1236,n1237);
nand (n1235,n1089,n1093);
nand (n1236,n1107,n1093);
nand (n1237,n1089,n1107);
nor (n1238,n1239,n1511);
nor (n1239,n1240,n1487);
nor (n1240,n1241,n1485);
nor (n1241,n1242,n1460);
nand (n1242,n1243,n1422);
nand (n1243,n1244,n1369,n1421);
nand (n1244,n1245,n1296);
xor (n1245,n1246,n1283);
xor (n1246,n1247,n1268);
nand (n1247,n1248,n1262,n1267);
nand (n1248,n1249,n1258);
and (n1249,n1250,n1254);
xnor (n1250,n1251,n345);
nor (n1251,n1252,n1253);
and (n1252,n19,n593);
and (n1253,n14,n595);
xor (n1254,n1255,n220);
or (n1255,n1256,n1257);
and (n1256,n133,n343);
and (n1257,n105,n347);
xor (n1258,n1259,n32);
or (n1259,n1260,n1261);
and (n1260,n578,n55);
and (n1261,n582,n59);
nand (n1262,n1263,n1258);
xor (n1263,n1264,n37);
or (n1264,n1265,n1266);
and (n1265,n584,n30);
and (n1266,n607,n35);
nand (n1267,n1249,n1263);
xor (n1268,n1269,n1278);
xor (n1269,n1270,n1274);
xor (n1270,n1271,n44);
or (n1271,n1272,n1273);
and (n1272,n109,n119);
and (n1273,n183,n123);
xor (n1274,n1275,n121);
or (n1275,n1276,n1277);
and (n1276,n133,n218);
and (n1277,n105,n222);
and (n1278,n1279,n86);
xnor (n1279,n1280,n345);
nor (n1280,n1281,n1282);
and (n1281,n14,n593);
and (n1282,n83,n595);
nand (n1283,n1284,n1290,n1295);
nand (n1284,n1285,n1289);
xor (n1285,n1286,n121);
or (n1286,n1287,n1288);
and (n1287,n105,n218);
and (n1288,n109,n222);
xor (n1289,n1279,n86);
nand (n1290,n1291,n1289);
xor (n1291,n1292,n49);
or (n1292,n1293,n1294);
and (n1293,n191,n42);
and (n1294,n327,n47);
nand (n1295,n1285,n1291);
xor (n1296,n1297,n1333);
xor (n1297,n1298,n1309);
xor (n1298,n1299,n1305);
xor (n1299,n1300,n1304);
xor (n1300,n1301,n49);
or (n1301,n1302,n1303);
and (n1302,n187,n42);
and (n1303,n191,n47);
xor (n1304,n708,n712);
xor (n1305,n1306,n32);
or (n1306,n1307,n1308);
and (n1307,n327,n55);
and (n1308,n578,n59);
xor (n1309,n1310,n1319);
xor (n1310,n1311,n1315);
xor (n1311,n1312,n37);
or (n1312,n1313,n1314);
and (n1313,n582,n30);
and (n1314,n584,n35);
xor (n1315,n1316,n86);
or (n1316,n1317,n1318);
and (n1317,n607,n80);
and (n1318,n621,n84);
nand (n1319,n1320,n1327,n1332);
nand (n1320,n1321,n1325);
xor (n1321,n1322,n220);
or (n1322,n1323,n1324);
and (n1323,n19,n343);
and (n1324,n133,n347);
xnor (n1325,n1326,n86);
nand (n1326,n621,n80);
nand (n1327,n1328,n1325);
xor (n1328,n1329,n44);
or (n1329,n1330,n1331);
and (n1330,n183,n119);
and (n1331,n187,n123);
nand (n1332,n1321,n1328);
nand (n1333,n1334,n1354,n1368);
nand (n1334,n1335,n1337);
xor (n1335,n1336,n1328);
xor (n1336,n1321,n1325);
nand (n1337,n1338,n1347,n1353);
nand (n1338,n1339,n1343);
xor (n1339,n1340,n44);
or (n1340,n1341,n1342);
and (n1341,n187,n119);
and (n1342,n191,n123);
xor (n1343,n1344,n121);
or (n1344,n1345,n1346);
and (n1345,n109,n218);
and (n1346,n183,n222);
nand (n1347,n1348,n1343);
and (n1348,n1349,n37);
xnor (n1349,n1350,n345);
nor (n1350,n1351,n1352);
and (n1351,n133,n593);
and (n1352,n19,n595);
nand (n1353,n1339,n1348);
nand (n1354,n1355,n1337);
nand (n1355,n1356,n1362,n1367);
nand (n1356,n1357,n1361);
xor (n1357,n1358,n49);
or (n1358,n1359,n1360);
and (n1359,n327,n42);
and (n1360,n578,n47);
xor (n1361,n1250,n1254);
nand (n1362,n1363,n1361);
xor (n1363,n1364,n32);
or (n1364,n1365,n1366);
and (n1365,n582,n55);
and (n1366,n584,n59);
nand (n1367,n1357,n1363);
nand (n1368,n1335,n1355);
nand (n1369,n1370,n1296);
nand (n1370,n1371,n1376,n1420);
nand (n1371,n1372,n1374);
xor (n1372,n1373,n1263);
xor (n1373,n1249,n1258);
xor (n1374,n1375,n1291);
xor (n1375,n1285,n1289);
nand (n1376,n1377,n1374);
nand (n1377,n1378,n1397,n1419);
nand (n1378,n1379,n1383);
xor (n1379,n1380,n37);
or (n1380,n1381,n1382);
and (n1381,n607,n30);
and (n1382,n621,n35);
nand (n1383,n1384,n1391,n1396);
nand (n1384,n1385,n1389);
xor (n1385,n1386,n220);
or (n1386,n1387,n1388);
and (n1387,n105,n343);
and (n1388,n109,n347);
xnor (n1389,n1390,n37);
nand (n1390,n621,n30);
nand (n1391,n1392,n1389);
xor (n1392,n1393,n44);
or (n1393,n1394,n1395);
and (n1394,n191,n119);
and (n1395,n327,n123);
nand (n1396,n1385,n1392);
nand (n1397,n1398,n1383);
nand (n1398,n1399,n1413,n1418);
nand (n1399,n1400,n1404);
xor (n1400,n1401,n121);
or (n1401,n1402,n1403);
and (n1402,n183,n218);
and (n1403,n187,n222);
and (n1404,n1405,n1409);
xnor (n1405,n1406,n345);
nor (n1406,n1407,n1408);
and (n1407,n105,n593);
and (n1408,n133,n595);
xor (n1409,n1410,n220);
or (n1410,n1411,n1412);
and (n1411,n109,n343);
and (n1412,n183,n347);
nand (n1413,n1414,n1404);
xor (n1414,n1415,n49);
or (n1415,n1416,n1417);
and (n1416,n578,n42);
and (n1417,n582,n47);
nand (n1418,n1400,n1414);
nand (n1419,n1379,n1398);
nand (n1420,n1372,n1377);
nand (n1421,n1245,n1370);
xor (n1422,n1423,n1438);
xor (n1423,n1424,n1434);
xor (n1424,n1425,n1432);
xor (n1425,n1426,n1430);
nand (n1426,n1427,n1428,n1429);
nand (n1427,n1270,n1274);
nand (n1428,n1278,n1274);
nand (n1429,n1270,n1278);
xor (n1430,n1431,n721);
xor (n1431,n707,n716);
xor (n1432,n1433,n822);
xor (n1433,n816,n820);
nand (n1434,n1435,n1436,n1437);
nand (n1435,n1298,n1309);
nand (n1436,n1333,n1309);
nand (n1437,n1298,n1333);
xor (n1438,n1439,n1448);
xor (n1439,n1440,n1444);
nand (n1440,n1441,n1442,n1443);
nand (n1441,n1311,n1315);
nand (n1442,n1319,n1315);
nand (n1443,n1311,n1319);
nand (n1444,n1445,n1446,n1447);
nand (n1445,n1247,n1268);
nand (n1446,n1283,n1268);
nand (n1447,n1247,n1283);
xor (n1448,n1449,n1458);
xor (n1449,n1450,n1454);
xor (n1450,n1451,n86);
or (n1451,n1452,n1453);
and (n1452,n584,n80);
and (n1453,n607,n84);
nand (n1454,n1455,n1456,n1457);
nand (n1455,n1300,n1304);
nand (n1456,n1305,n1304);
nand (n1457,n1300,n1305);
xor (n1458,n1459,n808);
xor (n1459,n799,n803);
nor (n1460,n1461,n1465);
nand (n1461,n1462,n1463,n1464);
nand (n1462,n1424,n1434);
nand (n1463,n1438,n1434);
nand (n1464,n1424,n1438);
xor (n1465,n1466,n1473);
xor (n1466,n1467,n1469);
xor (n1467,n1468,n729);
xor (n1468,n705,n726);
nand (n1469,n1470,n1471,n1472);
nand (n1470,n1440,n1444);
nand (n1471,n1448,n1444);
nand (n1472,n1440,n1448);
xor (n1473,n1474,n1483);
xor (n1474,n1475,n1479);
nand (n1475,n1476,n1477,n1478);
nand (n1476,n1450,n1454);
nand (n1477,n1458,n1454);
nand (n1478,n1450,n1458);
nand (n1479,n1480,n1481,n1482);
nand (n1480,n1426,n1430);
nand (n1481,n1432,n1430);
nand (n1482,n1426,n1432);
xor (n1483,n1484,n814);
xor (n1484,n797,n811);
not (n1485,n1486);
nand (n1486,n1461,n1465);
not (n1487,n1488);
nor (n1488,n1489,n1504);
nor (n1489,n1490,n1494);
nand (n1490,n1491,n1492,n1493);
nand (n1491,n1467,n1469);
nand (n1492,n1473,n1469);
nand (n1493,n1467,n1473);
xor (n1494,n1495,n1502);
xor (n1495,n1496,n1498);
xor (n1496,n1497,n795);
xor (n1497,n788,n792);
nand (n1498,n1499,n1500,n1501);
nand (n1499,n1475,n1479);
nand (n1500,n1483,n1479);
nand (n1501,n1475,n1483);
xor (n1502,n1503,n703);
xor (n1503,n649,n651);
nor (n1504,n1505,n1509);
nand (n1505,n1506,n1507,n1508);
nand (n1506,n1496,n1498);
nand (n1507,n1502,n1498);
nand (n1508,n1496,n1502);
xor (n1509,n1510,n746);
xor (n1510,n570,n647);
not (n1511,n1512);
nor (n1512,n1513,n1515);
nor (n1513,n1514,n1504);
nand (n1514,n1490,n1494);
not (n1515,n1516);
nand (n1516,n1505,n1509);
not (n1517,n1518);
nor (n1518,n1519,n1526);
nor (n1519,n1520,n1525);
nor (n1520,n1521,n1523);
nor (n1521,n1522,n920);
nand (n1522,n568,n830);
not (n1523,n1524);
nand (n1524,n921,n925);
not (n1525,n1021);
not (n1526,n1527);
nor (n1527,n1528,n1530);
nor (n1528,n1529,n1127);
nand (n1529,n1023,n1027);
not (n1530,n1531);
nand (n1531,n1128,n1132);
not (n1532,n1533);
nor (n1533,n1534,n1949);
nand (n1534,n1535,n1762);
nor (n1535,n1536,n1648);
nor (n1536,n1537,n1541);
nand (n1537,n1538,n1539,n1540);
nand (n1538,n1134,n1138);
nand (n1539,n1142,n1138);
nand (n1540,n1134,n1142);
xor (n1541,n1542,n1644);
xor (n1542,n1543,n1576);
xor (n1543,n1544,n1572);
xor (n1544,n1545,n1568);
xor (n1545,n1546,n1564);
xor (n1546,n1547,n1560);
xor (n1547,n1548,n1557);
xor (n1548,n1549,n1553);
xor (n1549,n1550,n220);
or (n1550,n1551,n1552);
and (n1551,n41,n343);
and (n1552,n46,n347);
xor (n1553,n1554,n121);
or (n1554,n1555,n1556);
and (n1555,n54,n218);
and (n1556,n58,n222);
xnor (n1557,n1558,n345);
nor (n1558,n1559,n1180);
and (n1559,n145,n593);
nand (n1560,n1561,n1562,n1563);
nand (n1561,n1152,n1156);
nand (n1562,n1160,n1156);
nand (n1563,n1152,n1160);
nand (n1564,n1565,n1566,n1567);
nand (n1565,n1172,n1176);
nand (n1566,n1185,n1176);
nand (n1567,n1172,n1185);
nand (n1568,n1569,n1570,n1571);
nand (n1569,n1146,n1150);
nand (n1570,n1164,n1150);
nand (n1571,n1146,n1164);
nand (n1572,n1573,n1574,n1575);
nand (n1573,n1170,n1186);
nand (n1574,n1190,n1186);
nand (n1575,n1170,n1190);
xor (n1576,n1577,n1640);
xor (n1577,n1578,n1616);
xor (n1578,n1579,n1601);
xor (n1579,n1580,n1594);
xor (n1580,n1581,n1590);
xor (n1581,n1582,n1586);
xor (n1582,n1583,n49);
or (n1583,n1584,n1585);
and (n1584,n70,n42);
and (n1585,n79,n47);
xor (n1586,n1587,n32);
or (n1587,n1588,n1589);
and (n1588,n83,n55);
and (n1589,n14,n59);
xor (n1590,n1591,n37);
or (n1591,n1592,n1593);
and (n1592,n19,n30);
and (n1593,n133,n35);
xor (n1594,n1595,n1597);
xor (n1595,n23,n1596);
and (n1596,n1177,n1181);
xor (n1597,n1598,n22);
or (n1598,n1599,n1600);
and (n1599,n191,n15);
and (n1600,n327,n20);
xor (n1601,n1602,n1611);
xor (n1602,n1603,n1607);
xor (n1603,n1604,n86);
or (n1604,n1605,n1606);
and (n1605,n105,n80);
and (n1606,n109,n84);
xor (n1607,n1608,n17);
or (n1608,n1609,n1610);
and (n1609,n183,n97);
and (n1610,n187,n100);
xor (n1611,n23,n1612);
xor (n1612,n1613,n44);
or (n1613,n1614,n1615);
and (n1614,n29,n119);
and (n1615,n34,n123);
xor (n1616,n1617,n1626);
xor (n1617,n1618,n1622);
nand (n1618,n1619,n1620,n1621);
nand (n1619,n1192,n1196);
nand (n1620,n1200,n1196);
nand (n1621,n1192,n1200);
nand (n1622,n1623,n1624,n1625);
nand (n1623,n1208,n1212);
nand (n1624,n1226,n1212);
nand (n1625,n1208,n1226);
xor (n1626,n1627,n1636);
xor (n1627,n1628,n1632);
xor (n1628,n1629,n112);
or (n1629,n1630,n1631);
and (n1630,n578,n106);
and (n1631,n582,n110);
xor (n1632,n1633,n23);
or (n1633,n1634,n1635);
and (n1634,n584,n188);
and (n1635,n607,n192);
nand (n1636,n1637,n1638,n1639);
nand (n1637,n1214,n1218);
nand (n1638,n1222,n1218);
nand (n1639,n1214,n1222);
nand (n1640,n1641,n1642,n1643);
nand (n1641,n1206,n1230);
nand (n1642,n1234,n1230);
nand (n1643,n1206,n1234);
nand (n1644,n1645,n1646,n1647);
nand (n1645,n1144,n1168);
nand (n1646,n1204,n1168);
nand (n1647,n1144,n1204);
nor (n1648,n1649,n1653);
nand (n1649,n1650,n1651,n1652);
nand (n1650,n1543,n1576);
nand (n1651,n1644,n1576);
nand (n1652,n1543,n1644);
xor (n1653,n1654,n1663);
xor (n1654,n1655,n1659);
nand (n1655,n1656,n1657,n1658);
nand (n1656,n1545,n1568);
nand (n1657,n1572,n1568);
nand (n1658,n1545,n1572);
nand (n1659,n1660,n1661,n1662);
nand (n1660,n1578,n1616);
nand (n1661,n1640,n1616);
nand (n1662,n1578,n1640);
xor (n1663,n1664,n1721);
xor (n1664,n1665,n1696);
xor (n1665,n1666,n1682);
xor (n1666,n1667,n1671);
nand (n1667,n1668,n1669,n1670);
nand (n1668,n23,n1596);
nand (n1669,n1597,n1596);
nand (n1670,n23,n1597);
xor (n1671,n1672,n1678);
xor (n1672,n1673,n1677);
xor (n1673,n1674,n17);
or (n1674,n1675,n1676);
and (n1675,n109,n97);
and (n1676,n183,n100);
and (n1677,n23,n1612);
xor (n1678,n1679,n22);
or (n1679,n1680,n1681);
and (n1680,n187,n15);
and (n1681,n191,n20);
xor (n1682,n1683,n1692);
xor (n1683,n1684,n1688);
xor (n1684,n1685,n112);
or (n1685,n1686,n1687);
and (n1686,n327,n106);
and (n1687,n578,n110);
xor (n1688,n1689,n23);
or (n1689,n1690,n1691);
and (n1690,n582,n188);
and (n1691,n584,n192);
nand (n1692,n1693,n1694,n1695);
nand (n1693,n1549,n1553);
nand (n1694,n1557,n1553);
nand (n1695,n1549,n1557);
xor (n1696,n1697,n1706);
xor (n1697,n1698,n1702);
nand (n1698,n1699,n1700,n1701);
nand (n1699,n1628,n1632);
nand (n1700,n1636,n1632);
nand (n1701,n1628,n1636);
nand (n1702,n1703,n1704,n1705);
nand (n1703,n1547,n1560);
nand (n1704,n1564,n1560);
nand (n1705,n1547,n1564);
xor (n1706,n1707,n23);
xor (n1707,n1708,n1712);
nand (n1708,n1709,n1710,n1711);
nand (n1709,n1582,n1586);
nand (n1710,n1590,n1586);
nand (n1711,n1582,n1590);
xor (n1712,n1713,n1718);
not (n1713,n1714);
xor (n1714,n1715,n44);
or (n1715,n1716,n1717);
and (n1716,n58,n119);
and (n1717,n29,n123);
xor (n1718,n1719,n220);
or (n1719,n342,n1720);
and (n1720,n41,n347);
xor (n1721,n1722,n1758);
xor (n1722,n1723,n1727);
nand (n1723,n1724,n1725,n1726);
nand (n1724,n1580,n1594);
nand (n1725,n1601,n1594);
nand (n1726,n1580,n1601);
xor (n1727,n1728,n1747);
xor (n1728,n1729,n1733);
nand (n1729,n1730,n1731,n1732);
nand (n1730,n1603,n1607);
nand (n1731,n1611,n1607);
nand (n1732,n1603,n1611);
xor (n1733,n1734,n1743);
xor (n1734,n1735,n1739);
xor (n1735,n1736,n32);
or (n1736,n1737,n1738);
and (n1737,n79,n55);
and (n1738,n83,n59);
xor (n1739,n1740,n37);
or (n1740,n1741,n1742);
and (n1741,n14,n30);
and (n1742,n19,n35);
xor (n1743,n1744,n86);
or (n1744,n1745,n1746);
and (n1745,n133,n80);
and (n1746,n105,n84);
xor (n1747,n1748,n1754);
xor (n1748,n1749,n1753);
xor (n1749,n1750,n121);
or (n1750,n1751,n1752);
and (n1751,n46,n218);
and (n1752,n54,n222);
not (n1753,n1557);
xor (n1754,n1755,n49);
or (n1755,n1756,n1757);
and (n1756,n34,n42);
and (n1757,n70,n47);
nand (n1758,n1759,n1760,n1761);
nand (n1759,n1618,n1622);
nand (n1760,n1626,n1622);
nand (n1761,n1618,n1626);
nor (n1762,n1763,n1870);
nor (n1763,n1764,n1768);
nand (n1764,n1765,n1766,n1767);
nand (n1765,n1655,n1659);
nand (n1766,n1663,n1659);
nand (n1767,n1655,n1663);
xor (n1768,n1769,n1866);
xor (n1769,n1770,n1810);
xor (n1770,n1771,n1806);
xor (n1771,n1772,n1802);
xor (n1772,n1773,n1798);
xor (n1773,n1774,n1788);
xor (n1774,n1775,n1784);
xor (n1775,n1776,n1780);
xor (n1776,n1777,n32);
or (n1777,n1778,n1779);
and (n1778,n70,n55);
and (n1779,n79,n59);
xor (n1780,n1781,n37);
or (n1781,n1782,n1783);
and (n1782,n83,n30);
and (n1783,n14,n35);
xor (n1784,n1785,n17);
or (n1785,n1786,n1787);
and (n1786,n105,n97);
and (n1787,n109,n100);
xor (n1788,n1789,n1794);
xor (n1789,n1790,n340);
xor (n1790,n1791,n44);
or (n1791,n1792,n1793);
and (n1792,n54,n119);
and (n1793,n58,n123);
xor (n1794,n1795,n49);
or (n1795,n1796,n1797);
and (n1796,n29,n42);
and (n1797,n34,n47);
nand (n1798,n1799,n1800,n1801);
nand (n1799,n1673,n1677);
nand (n1800,n1678,n1677);
nand (n1801,n1673,n1678);
nand (n1802,n1803,n1804,n1805);
nand (n1803,n1667,n1671);
nand (n1804,n1682,n1671);
nand (n1805,n1667,n1682);
nand (n1806,n1807,n1808,n1809);
nand (n1807,n1698,n1702);
nand (n1808,n1706,n1702);
nand (n1809,n1698,n1706);
xor (n1810,n1811,n1862);
xor (n1811,n1812,n1833);
xor (n1812,n1813,n1829);
xor (n1813,n1814,n1825);
xor (n1814,n1815,n1821);
xor (n1815,n1816,n1817);
not (n1816,n381);
xor (n1817,n1818,n86);
or (n1818,n1819,n1820);
and (n1819,n19,n80);
and (n1820,n133,n84);
xor (n1821,n1822,n22);
or (n1822,n1823,n1824);
and (n1823,n183,n15);
and (n1824,n187,n20);
nand (n1825,n1826,n1827,n1828);
nand (n1826,n1684,n1688);
nand (n1827,n1692,n1688);
nand (n1828,n1684,n1692);
nand (n1829,n1830,n1831,n1832);
nand (n1830,n1708,n1712);
nand (n1831,n23,n1712);
nand (n1832,n1708,n23);
xor (n1833,n1834,n1858);
xor (n1834,n1835,n1848);
xor (n1835,n1836,n1845);
xor (n1836,n1837,n1841);
xor (n1837,n1838,n112);
or (n1838,n1839,n1840);
and (n1839,n191,n106);
and (n1840,n327,n110);
xor (n1841,n1842,n23);
or (n1842,n1843,n1844);
and (n1843,n578,n188);
and (n1844,n582,n192);
nand (n1845,n1713,n1846,n1847);
nand (n1846,n1718,n1714);
not (n1847,n1718);
xor (n1848,n1849,n1854);
xor (n1849,n23,n1850);
nand (n1850,n1851,n1852,n1853);
nand (n1851,n1749,n1753);
nand (n1852,n1754,n1753);
nand (n1853,n1749,n1754);
nand (n1854,n1855,n1856,n1857);
nand (n1855,n1735,n1739);
nand (n1856,n1743,n1739);
nand (n1857,n1735,n1743);
nand (n1858,n1859,n1860,n1861);
nand (n1859,n1729,n1733);
nand (n1860,n1747,n1733);
nand (n1861,n1729,n1747);
nand (n1862,n1863,n1864,n1865);
nand (n1863,n1723,n1727);
nand (n1864,n1758,n1727);
nand (n1865,n1723,n1758);
nand (n1866,n1867,n1868,n1869);
nand (n1867,n1665,n1696);
nand (n1868,n1721,n1696);
nand (n1869,n1665,n1721);
nor (n1870,n1871,n1875);
nand (n1871,n1872,n1873,n1874);
nand (n1872,n1770,n1810);
nand (n1873,n1866,n1810);
nand (n1874,n1770,n1866);
xor (n1875,n1876,n1885);
xor (n1876,n1877,n1881);
nand (n1877,n1878,n1879,n1880);
nand (n1878,n1772,n1802);
nand (n1879,n1806,n1802);
nand (n1880,n1772,n1806);
nand (n1881,n1882,n1883,n1884);
nand (n1882,n1812,n1833);
nand (n1883,n1862,n1833);
nand (n1884,n1812,n1862);
xor (n1885,n1886,n1917);
xor (n1886,n1887,n1891);
nand (n1887,n1888,n1889,n1890);
nand (n1888,n1835,n1848);
nand (n1889,n1858,n1848);
nand (n1890,n1835,n1858);
xor (n1891,n1892,n1905);
xor (n1892,n1893,n1897);
nand (n1893,n1894,n1895,n1896);
nand (n1894,n23,n1850);
nand (n1895,n1854,n1850);
nand (n1896,n23,n1854);
xor (n1897,n1898,n1901);
xor (n1898,n1899,n23);
xor (n1899,n1900,n339);
xor (n1900,n331,n334);
nand (n1901,n1902,n1903,n1904);
nand (n1902,n1790,n340);
nand (n1903,n1794,n340);
nand (n1904,n1790,n1794);
xor (n1905,n1906,n1913);
xor (n1906,n1907,n1909);
xor (n1907,n1908,n367);
xor (n1908,n358,n362);
nand (n1909,n1910,n1911,n1912);
nand (n1910,n1776,n1780);
nand (n1911,n1784,n1780);
nand (n1912,n1776,n1784);
nand (n1913,n1914,n1915,n1916);
nand (n1914,n1837,n1841);
nand (n1915,n1845,n1841);
nand (n1916,n1837,n1845);
xor (n1917,n1918,n1927);
xor (n1918,n1919,n1923);
nand (n1919,n1920,n1921,n1922);
nand (n1920,n1774,n1788);
nand (n1921,n1798,n1788);
nand (n1922,n1774,n1798);
nand (n1923,n1924,n1925,n1926);
nand (n1924,n1814,n1825);
nand (n1925,n1829,n1825);
nand (n1926,n1814,n1829);
xor (n1927,n1928,n1935);
xor (n1928,n1929,n1933);
nand (n1929,n1930,n1931,n1932);
nand (n1930,n1816,n1817);
nand (n1931,n1821,n1817);
nand (n1932,n1816,n1821);
xor (n1933,n1934,n386);
xor (n1934,n377,n381);
xor (n1935,n1936,n1945);
xor (n1936,n1937,n1941);
xor (n1937,n1938,n22);
or (n1938,n1939,n1940);
and (n1939,n109,n15);
and (n1940,n183,n20);
xor (n1941,n1942,n112);
or (n1942,n1943,n1944);
and (n1943,n187,n106);
and (n1944,n191,n110);
xor (n1945,n1946,n23);
or (n1946,n1947,n1948);
and (n1947,n327,n188);
and (n1948,n578,n192);
nand (n1949,n1950,n2034);
nor (n1950,n1951,n2001);
nor (n1951,n1952,n1956);
nand (n1952,n1953,n1954,n1955);
nand (n1953,n1877,n1881);
nand (n1954,n1885,n1881);
nand (n1955,n1877,n1885);
xor (n1956,n1957,n1997);
xor (n1957,n1958,n1978);
xor (n1958,n1959,n1966);
xor (n1959,n1960,n1962);
xor (n1960,n1961,n375);
xor (n1961,n356,n372);
nand (n1962,n1963,n1964,n1965);
nand (n1963,n1929,n1933);
nand (n1964,n1935,n1933);
nand (n1965,n1929,n1935);
xor (n1966,n1967,n1974);
xor (n1967,n1968,n1972);
nand (n1968,n1969,n1970,n1971);
nand (n1969,n1937,n1941);
nand (n1970,n1945,n1941);
nand (n1971,n1937,n1945);
xor (n1972,n1973,n285);
xor (n1973,n279,n283);
nand (n1974,n1975,n1976,n1977);
nand (n1975,n1899,n23);
nand (n1976,n1901,n23);
nand (n1977,n1899,n1901);
xor (n1978,n1979,n1993);
xor (n1979,n1980,n1984);
nand (n1980,n1981,n1982,n1983);
nand (n1981,n1893,n1897);
nand (n1982,n1905,n1897);
nand (n1983,n1893,n1905);
xor (n1984,n1985,n1989);
xor (n1985,n1986,n1988);
xor (n1986,n1987,n301);
xor (n1987,n292,n296);
xor (n1988,n324,n329);
nand (n1989,n1990,n1991,n1992);
nand (n1990,n1907,n1909);
nand (n1991,n1913,n1909);
nand (n1992,n1907,n1913);
nand (n1993,n1994,n1995,n1996);
nand (n1994,n1919,n1923);
nand (n1995,n1927,n1923);
nand (n1996,n1919,n1927);
nand (n1997,n1998,n1999,n2000);
nand (n1998,n1887,n1891);
nand (n1999,n1917,n1891);
nand (n2000,n1887,n1917);
nor (n2001,n2002,n2006);
nand (n2002,n2003,n2004,n2005);
nand (n2003,n1958,n1978);
nand (n2004,n1997,n1978);
nand (n2005,n1958,n1997);
xor (n2006,n2007,n2030);
xor (n2007,n2008,n2018);
xor (n2008,n2009,n2016);
xor (n2009,n2010,n2012);
xor (n2010,n2011,n272);
xor (n2011,n257,n269);
nand (n2012,n2013,n2014,n2015);
nand (n2013,n1968,n1972);
nand (n2014,n1974,n1972);
nand (n2015,n1968,n1974);
xor (n2016,n2017,n307);
xor (n2017,n277,n290);
xor (n2018,n2019,n2026);
xor (n2019,n2020,n2022);
xor (n2020,n2021,n354);
xor (n2021,n321,n351);
nand (n2022,n2023,n2024,n2025);
nand (n2023,n1986,n1988);
nand (n2024,n1989,n1988);
nand (n2025,n1986,n1989);
nand (n2026,n2027,n2028,n2029);
nand (n2027,n1960,n1962);
nand (n2028,n1966,n1962);
nand (n2029,n1960,n1966);
nand (n2030,n2031,n2032,n2033);
nand (n2031,n1980,n1984);
nand (n2032,n1993,n1984);
nand (n2033,n1980,n1993);
nor (n2034,n2035,n2052);
nor (n2035,n2036,n2040);
nand (n2036,n2037,n2038,n2039);
nand (n2037,n2008,n2018);
nand (n2038,n2030,n2018);
nand (n2039,n2008,n2030);
xor (n2040,n2041,n2048);
xor (n2041,n2042,n2046);
nand (n2042,n2043,n2044,n2045);
nand (n2043,n2010,n2012);
nand (n2044,n2016,n2012);
nand (n2045,n2010,n2016);
xor (n2046,n2047,n394);
xor (n2047,n317,n319);
nand (n2048,n2049,n2050,n2051);
nand (n2049,n2020,n2022);
nand (n2050,n2026,n2022);
nand (n2051,n2020,n2026);
nor (n2052,n2053,n2057);
nand (n2053,n2054,n2055,n2056);
nand (n2054,n2042,n2046);
nand (n2055,n2048,n2046);
nand (n2056,n2042,n2048);
xor (n2057,n2058,n315);
xor (n2058,n7,n173);
not (n2059,n2060);
nor (n2060,n2061,n2076);
nor (n2061,n1949,n2062);
nor (n2062,n2063,n2070);
nor (n2063,n2064,n2069);
nor (n2064,n2065,n2067);
nor (n2065,n2066,n1648);
nand (n2066,n1537,n1541);
not (n2067,n2068);
nand (n2068,n1649,n1653);
not (n2069,n1762);
not (n2070,n2071);
nor (n2071,n2072,n2074);
nor (n2072,n2073,n1870);
nand (n2073,n1764,n1768);
not (n2074,n2075);
nand (n2075,n1871,n1875);
not (n2076,n2077);
nor (n2077,n2078,n2085);
nor (n2078,n2079,n2084);
nor (n2079,n2080,n2082);
nor (n2080,n2081,n2001);
nand (n2081,n1952,n1956);
not (n2082,n2083);
nand (n2083,n2002,n2006);
not (n2084,n2034);
not (n2085,n2086);
nor (n2086,n2087,n2089);
nor (n2087,n2088,n2052);
nand (n2088,n2036,n2040);
not (n2089,n2090);
nand (n2090,n2053,n2057);
nand (n2091,n2092,n2511);
nand (n2092,n2093,n2404);
nor (n2093,n2094,n2389);
nor (n2094,n2095,n2260);
nand (n2095,n2096,n2237);
nor (n2096,n2097,n2214);
nor (n2097,n2098,n2187);
nand (n2098,n2099,n2144,n2186);
nand (n2099,n2100,n2112);
xor (n2100,n2101,n2107);
xor (n2101,n2102,n2103);
xor (n2102,n1405,n1409);
xor (n2103,n2104,n32);
or (n2104,n2105,n2106);
and (n2105,n607,n55);
and (n2106,n621,n59);
and (n2107,n32,n2108);
xor (n2108,n2109,n220);
or (n2109,n2110,n2111);
and (n2110,n183,n343);
and (n2111,n187,n347);
nand (n2112,n2113,n2130,n2143);
nand (n2113,n2114,n2115);
xor (n2114,n32,n2108);
nand (n2115,n2116,n2125,n2129);
nand (n2116,n2117,n2121);
xor (n2117,n2118,n44);
or (n2118,n2119,n2120);
and (n2119,n582,n119);
and (n2120,n584,n123);
xor (n2121,n2122,n121);
or (n2122,n2123,n2124);
and (n2123,n327,n218);
and (n2124,n578,n222);
nand (n2125,n2126,n2121);
and (n2126,n49,n2127);
xnor (n2127,n2128,n49);
nand (n2128,n621,n42);
nand (n2129,n2117,n2126);
nand (n2130,n2131,n2115);
xor (n2131,n2132,n2139);
xor (n2132,n2133,n2137);
xnor (n2133,n2134,n345);
nor (n2134,n2135,n2136);
and (n2135,n109,n593);
and (n2136,n105,n595);
xnor (n2137,n2138,n32);
nand (n2138,n621,n55);
xor (n2139,n2140,n44);
or (n2140,n2141,n2142);
and (n2141,n578,n119);
and (n2142,n582,n123);
nand (n2143,n2114,n2131);
nand (n2144,n2145,n2112);
xor (n2145,n2146,n2165);
xor (n2146,n2147,n2151);
nand (n2147,n2148,n2149,n2150);
nand (n2148,n2133,n2137);
nand (n2149,n2139,n2137);
nand (n2150,n2133,n2139);
xor (n2151,n2152,n2161);
xor (n2152,n2153,n2157);
xor (n2153,n2154,n44);
or (n2154,n2155,n2156);
and (n2155,n327,n119);
and (n2156,n578,n123);
xor (n2157,n2158,n121);
or (n2158,n2159,n2160);
and (n2159,n187,n218);
and (n2160,n191,n222);
xor (n2161,n2162,n49);
or (n2162,n2163,n2164);
and (n2163,n582,n42);
and (n2164,n584,n47);
nand (n2165,n2166,n2180,n2185);
nand (n2166,n2167,n2171);
xor (n2167,n2168,n121);
or (n2168,n2169,n2170);
and (n2169,n191,n218);
and (n2170,n327,n222);
and (n2171,n2172,n2176);
xnor (n2172,n2173,n345);
nor (n2173,n2174,n2175);
and (n2174,n183,n593);
and (n2175,n109,n595);
xor (n2176,n2177,n220);
or (n2177,n2178,n2179);
and (n2178,n187,n343);
and (n2179,n191,n347);
nand (n2180,n2181,n2171);
xor (n2181,n2182,n49);
or (n2182,n2183,n2184);
and (n2183,n584,n42);
and (n2184,n607,n47);
nand (n2185,n2167,n2181);
nand (n2186,n2100,n2145);
xor (n2187,n2188,n2202);
xor (n2188,n2189,n2198);
xor (n2189,n2190,n2196);
xor (n2190,n2191,n2195);
xor (n2191,n2192,n32);
or (n2192,n2193,n2194);
and (n2193,n584,n55);
and (n2194,n607,n59);
xor (n2195,n1349,n37);
xor (n2196,n2197,n1392);
xor (n2197,n1385,n1389);
nand (n2198,n2199,n2200,n2201);
nand (n2199,n2147,n2151);
nand (n2200,n2165,n2151);
nand (n2201,n2147,n2165);
xor (n2202,n2203,n2212);
xor (n2203,n2204,n2208);
nand (n2204,n2205,n2206,n2207);
nand (n2205,n2102,n2103);
nand (n2206,n2107,n2103);
nand (n2207,n2102,n2107);
nand (n2208,n2209,n2210,n2211);
nand (n2209,n2153,n2157);
nand (n2210,n2161,n2157);
nand (n2211,n2153,n2161);
xor (n2212,n2213,n1414);
xor (n2213,n1400,n1404);
nor (n2214,n2215,n2219);
nand (n2215,n2216,n2217,n2218);
nand (n2216,n2189,n2198);
nand (n2217,n2202,n2198);
nand (n2218,n2189,n2202);
xor (n2219,n2220,n2227);
xor (n2220,n2221,n2223);
xor (n2221,n2222,n1398);
xor (n2222,n1379,n1383);
nand (n2223,n2224,n2225,n2226);
nand (n2224,n2204,n2208);
nand (n2225,n2212,n2208);
nand (n2226,n2204,n2212);
xor (n2227,n2228,n2233);
xor (n2228,n2229,n2231);
xor (n2229,n2230,n1348);
xor (n2230,n1339,n1343);
xor (n2231,n2232,n1363);
xor (n2232,n1357,n1361);
nand (n2233,n2234,n2235,n2236);
nand (n2234,n2191,n2195);
nand (n2235,n2196,n2195);
nand (n2236,n2191,n2196);
nor (n2237,n2238,n2253);
nor (n2238,n2239,n2243);
nand (n2239,n2240,n2241,n2242);
nand (n2240,n2221,n2223);
nand (n2241,n2227,n2223);
nand (n2242,n2221,n2227);
xor (n2243,n2244,n2251);
xor (n2244,n2245,n2247);
xor (n2245,n2246,n1355);
xor (n2246,n1335,n1337);
nand (n2247,n2248,n2249,n2250);
nand (n2248,n2229,n2231);
nand (n2249,n2233,n2231);
nand (n2250,n2229,n2233);
xor (n2251,n2252,n1377);
xor (n2252,n1372,n1374);
nor (n2253,n2254,n2258);
nand (n2254,n2255,n2256,n2257);
nand (n2255,n2245,n2247);
nand (n2256,n2251,n2247);
nand (n2257,n2245,n2251);
xor (n2258,n2259,n1370);
xor (n2259,n1245,n1296);
nor (n2260,n2261,n2383);
nor (n2261,n2262,n2359);
nor (n2262,n2263,n2356);
nor (n2263,n2264,n2332);
nand (n2264,n2265,n2304);
or (n2265,n2266,n2290,n2303);
and (n2266,n2267,n2276);
xor (n2267,n2268,n2272);
xnor (n2268,n2269,n345);
nor (n2269,n2270,n2271);
and (n2270,n191,n593);
and (n2271,n187,n595);
xnor (n2272,n2273,n220);
nor (n2273,n2274,n2275);
and (n2274,n578,n347);
and (n2275,n327,n343);
or (n2276,n2277,n2284,n2289);
and (n2277,n2278,n2280);
not (n2278,n2279);
nand (n2279,n621,n119);
xnor (n2280,n2281,n345);
nor (n2281,n2282,n2283);
and (n2282,n327,n593);
and (n2283,n191,n595);
and (n2284,n2280,n2285);
xnor (n2285,n2286,n220);
nor (n2286,n2287,n2288);
and (n2287,n582,n347);
and (n2288,n578,n343);
and (n2289,n2278,n2285);
and (n2290,n2276,n2291);
xor (n2291,n2292,n2299);
xor (n2292,n2293,n2295);
and (n2293,n44,n2294);
xnor (n2294,n2279,n44);
xnor (n2295,n2296,n121);
nor (n2296,n2297,n2298);
and (n2297,n584,n222);
and (n2298,n582,n218);
xnor (n2299,n2300,n44);
nor (n2300,n2301,n2302);
and (n2301,n621,n123);
and (n2302,n607,n119);
and (n2303,n2267,n2291);
xor (n2304,n2305,n2321);
xor (n2305,n2306,n2310);
or (n2306,n2307,n2308,n2309);
and (n2307,n2293,n2295);
and (n2308,n2295,n2299);
and (n2309,n2293,n2299);
xor (n2310,n2311,n2317);
xor (n2311,n2312,n2313);
and (n2312,n2268,n2272);
xnor (n2313,n2314,n121);
nor (n2314,n2315,n2316);
and (n2315,n582,n222);
and (n2316,n578,n218);
xnor (n2317,n2318,n44);
nor (n2318,n2319,n2320);
and (n2319,n607,n123);
and (n2320,n584,n119);
xor (n2321,n2322,n2328);
xor (n2322,n2323,n2324);
not (n2323,n2128);
xnor (n2324,n2325,n345);
nor (n2325,n2326,n2327);
and (n2326,n187,n593);
and (n2327,n183,n595);
xnor (n2328,n2329,n220);
nor (n2329,n2330,n2331);
and (n2330,n327,n347);
and (n2331,n191,n343);
nor (n2332,n2333,n2337);
or (n2333,n2334,n2335,n2336);
and (n2334,n2306,n2310);
and (n2335,n2310,n2321);
and (n2336,n2306,n2321);
xor (n2337,n2338,n2345);
xor (n2338,n2339,n2343);
or (n2339,n2340,n2341,n2342);
and (n2340,n2312,n2313);
and (n2341,n2313,n2317);
and (n2342,n2312,n2317);
xor (n2343,n2344,n2126);
xor (n2344,n2117,n2121);
xor (n2345,n2346,n2352);
xor (n2346,n2347,n2351);
xor (n2347,n2348,n49);
or (n2348,n2349,n2350);
and (n2349,n607,n42);
and (n2350,n621,n47);
xor (n2351,n2172,n2176);
or (n2352,n2353,n2354,n2355);
and (n2353,n2323,n2324);
and (n2354,n2324,n2328);
and (n2355,n2323,n2328);
not (n2356,n2357);
not (n2357,n2358);
and (n2358,n2333,n2337);
not (n2359,n2360);
nor (n2360,n2361,n2376);
nor (n2361,n2362,n2366);
nand (n2362,n2363,n2364,n2365);
nand (n2363,n2339,n2343);
nand (n2364,n2345,n2343);
nand (n2365,n2339,n2345);
xor (n2366,n2367,n2374);
xor (n2367,n2368,n2370);
xor (n2368,n2369,n2181);
xor (n2369,n2167,n2171);
nand (n2370,n2371,n2372,n2373);
nand (n2371,n2347,n2351);
nand (n2372,n2352,n2351);
nand (n2373,n2347,n2352);
xor (n2374,n2375,n2131);
xor (n2375,n2114,n2115);
nor (n2376,n2377,n2381);
nand (n2377,n2378,n2379,n2380);
nand (n2378,n2368,n2370);
nand (n2379,n2374,n2370);
nand (n2380,n2368,n2374);
xor (n2381,n2382,n2145);
xor (n2382,n2100,n2112);
not (n2383,n2384);
nor (n2384,n2385,n2387);
nor (n2385,n2386,n2376);
nand (n2386,n2362,n2366);
not (n2387,n2388);
nand (n2388,n2377,n2381);
not (n2389,n2390);
nor (n2390,n2391,n2398);
nor (n2391,n2392,n2397);
nor (n2392,n2393,n2395);
nor (n2393,n2394,n2214);
nand (n2394,n2098,n2187);
not (n2395,n2396);
nand (n2396,n2215,n2219);
not (n2397,n2237);
not (n2398,n2399);
nor (n2399,n2400,n2402);
nor (n2400,n2401,n2253);
nand (n2401,n2239,n2243);
not (n2402,n2403);
nand (n2403,n2254,n2258);
nand (n2404,n2405,n2409);
nor (n2405,n2406,n2095);
nand (n2406,n2407,n2360);
nor (n2407,n2408,n2332);
nor (n2408,n2265,n2304);
or (n2409,n2410,n2432);
and (n2410,n2411,n2413);
xor (n2411,n2412,n2291);
xor (n2412,n2267,n2276);
or (n2413,n2414,n2428,n2431);
and (n2414,n2415,n2424);
and (n2415,n2416,n2420);
xnor (n2416,n2417,n345);
nor (n2417,n2418,n2419);
and (n2418,n578,n593);
and (n2419,n327,n595);
xnor (n2420,n2421,n220);
nor (n2421,n2422,n2423);
and (n2422,n584,n347);
and (n2423,n582,n343);
xnor (n2424,n2425,n121);
nor (n2425,n2426,n2427);
and (n2426,n607,n222);
and (n2427,n584,n218);
and (n2428,n2424,n2429);
xor (n2429,n2430,n2285);
xor (n2430,n2278,n2280);
and (n2431,n2415,n2429);
and (n2432,n2433,n2434);
xor (n2433,n2411,n2413);
or (n2434,n2435,n2450);
and (n2435,n2436,n2448);
or (n2436,n2437,n2442,n2447);
and (n2437,n2438,n2439);
xor (n2438,n2416,n2420);
and (n2439,n121,n2440);
xnor (n2440,n2441,n121);
nand (n2441,n621,n218);
and (n2442,n2439,n2443);
xnor (n2443,n2444,n121);
nor (n2444,n2445,n2446);
and (n2445,n621,n222);
and (n2446,n607,n218);
and (n2447,n2438,n2443);
xor (n2448,n2449,n2429);
xor (n2449,n2415,n2424);
and (n2450,n2451,n2452);
xor (n2451,n2436,n2448);
or (n2452,n2453,n2469);
and (n2453,n2454,n2456);
xor (n2454,n2455,n2443);
xor (n2455,n2438,n2439);
or (n2456,n2457,n2463,n2468);
and (n2457,n2458,n2459);
not (n2458,n2441);
xnor (n2459,n2460,n345);
nor (n2460,n2461,n2462);
and (n2461,n582,n593);
and (n2462,n578,n595);
and (n2463,n2459,n2464);
xnor (n2464,n2465,n220);
nor (n2465,n2466,n2467);
and (n2466,n607,n347);
and (n2467,n584,n343);
and (n2468,n2458,n2464);
and (n2469,n2470,n2471);
xor (n2470,n2454,n2456);
or (n2471,n2472,n2483);
and (n2472,n2473,n2475);
xor (n2473,n2474,n2464);
xor (n2474,n2458,n2459);
and (n2475,n2476,n2479);
and (n2476,n220,n2477);
xnor (n2477,n2478,n220);
nand (n2478,n621,n343);
xnor (n2479,n2480,n345);
nor (n2480,n2481,n2482);
and (n2481,n584,n593);
and (n2482,n582,n595);
and (n2483,n2484,n2485);
xor (n2484,n2473,n2475);
or (n2485,n2486,n2492);
and (n2486,n2487,n2491);
xnor (n2487,n2488,n220);
nor (n2488,n2489,n2490);
and (n2489,n621,n347);
and (n2490,n607,n343);
xor (n2491,n2476,n2479);
and (n2492,n2493,n2494);
xor (n2493,n2487,n2491);
or (n2494,n2495,n2501);
and (n2495,n2496,n2500);
xnor (n2496,n2497,n345);
nor (n2497,n2498,n2499);
and (n2498,n607,n593);
and (n2499,n584,n595);
not (n2500,n2478);
and (n2501,n2502,n2503);
xor (n2502,n2496,n2500);
and (n2503,n2504,n2508);
xnor (n2504,n2505,n345);
nor (n2505,n2506,n2507);
and (n2506,n621,n593);
and (n2507,n607,n595);
and (n2508,n2509,n345);
xnor (n2509,n2510,n345);
nand (n2510,n621,n595);
not (n2511,n2512);
nand (n2512,n2513,n1533);
nor (n2513,n2514,n565);
nand (n2514,n2515,n1488);
nor (n2515,n2516,n1460);
nor (n2516,n1243,n1422);
nand (n2517,n2518,n2592);
not (n2518,n2519);
nor (n2519,n2520,n2524);
nand (n2520,n2521,n2522,n2523);
nand (n2521,n485,n511);
nand (n2522,n551,n511);
nand (n2523,n485,n551);
xor (n2524,n2525,n2588);
xor (n2525,n2526,n2554);
xor (n2526,n2527,n2550);
xor (n2527,n2528,n2542);
xor (n2528,n2529,n2538);
xor (n2529,n2530,n2534);
not (n2530,n2531);
xor (n2531,n2532,n32);
or (n2532,n501,n2533);
and (n2533,n145,n59);
xor (n2534,n2535,n22);
or (n2535,n2536,n2537);
and (n2536,n70,n15);
and (n2537,n79,n20);
xor (n2538,n2539,n112);
or (n2539,n2540,n2541);
and (n2540,n83,n106);
and (n2541,n14,n110);
xor (n2542,n2543,n2546);
or (n2543,n2544,n2545);
and (n2544,n19,n188);
and (n2545,n133,n192);
nand (n2546,n2547,n2548,n2549);
nand (n2547,n440,n499);
nand (n2548,n503,n499);
nand (n2549,n440,n503);
nand (n2550,n2551,n2552,n2553);
nand (n2551,n23,n497);
nand (n2552,n507,n497);
nand (n2553,n23,n507);
xor (n2554,n2555,n2584);
xor (n2555,n2556,n2580);
xor (n2556,n2557,n2576);
xor (n2557,n2558,n2572);
xor (n2558,n2559,n2568);
xor (n2559,n2560,n2564);
xor (n2560,n2561,n37);
or (n2561,n2562,n2563);
and (n2562,n41,n30);
and (n2563,n46,n35);
xor (n2564,n2565,n17);
or (n2565,n2566,n2567);
and (n2566,n29,n97);
and (n2567,n34,n100);
xor (n2568,n2569,n86);
or (n2569,n2570,n2571);
and (n2570,n54,n80);
and (n2571,n58,n84);
nand (n2572,n2573,n2574,n2575);
nand (n2573,n521,n525);
nand (n2574,n529,n525);
nand (n2575,n521,n529);
nand (n2576,n2577,n2578,n2579);
nand (n2577,n441,n535);
nand (n2578,n539,n535);
nand (n2579,n441,n539);
nand (n2580,n2581,n2582,n2583);
nand (n2581,n515,n519);
nand (n2582,n533,n519);
nand (n2583,n515,n533);
nand (n2584,n2585,n2586,n2587);
nand (n2585,n487,n491);
nand (n2586,n495,n491);
nand (n2587,n487,n495);
nand (n2588,n2589,n2590,n2591);
nand (n2589,n513,n543);
nand (n2590,n547,n543);
nand (n2591,n513,n547);
nand (n2592,n2520,n2524);
xor (n2593,n2594,n2736);
xnor (n2594,n2595,n2662);
xor (n2595,n2596,n2648);
xor (n2596,n2597,n2608);
xor (n2597,n2598,n2604);
xor (n2598,n2557,n2599);
and (n2599,n2600,n519);
or (n2600,n2601,n2602,n2603);
and (n2601,n441,n432);
not (n2602,n516);
and (n2603,n441,n436);
or (n2604,n2605,n2606,n2607);
not (n2605,n2578);
and (n2606,n539,n507);
and (n2607,n535,n507);
or (n2608,n2609,n2633,n2647);
and (n2609,n2610,n2629);
or (n2610,n2611,n2624,n2628);
and (n2611,n2612,n2616);
or (n2612,n2613,n2614,n2615);
and (n2613,n11,n155);
and (n2614,n155,n240);
and (n2615,n11,n240);
or (n2616,n2617,n2618,n2623);
and (n2617,n24,n169);
and (n2618,n169,n2619);
or (n2619,n2620,n2621,n2622);
and (n2620,n142,n202);
not (n2621,n238);
and (n2622,n142,n198);
and (n2623,n24,n2619);
and (n2624,n2616,n2625);
xor (n2625,n2626,n417);
xor (n2626,n452,n2627);
not (n2627,n430);
and (n2628,n2612,n2625);
xor (n2629,n2630,n2632);
xor (n2630,n2631,n497);
not (n2631,n488);
xor (n2632,n2600,n519);
and (n2633,n2629,n2634);
xor (n2634,n2635,n2645);
xor (n2635,n2636,n2640);
or (n2636,n2637,n2638,n2639);
and (n2637,n452,n2627);
and (n2638,n2627,n417);
and (n2639,n452,n417);
or (n2640,n2641,n2643,n2644);
and (n2641,n466,n2642);
not (n2642,n413);
and (n2643,n2642,n426);
and (n2644,n466,n426);
xor (n2645,n2646,n507);
xor (n2646,n535,n539);
and (n2647,n2610,n2634);
xor (n2648,n2649,n2658);
xor (n2649,n2650,n2654);
xor (n2650,n2651,n2546);
xor (n2651,n2652,n2653);
xor (n2652,n2543,n23);
not (n2653,n2528);
or (n2654,n2655,n2656,n2657);
and (n2655,n2631,n497);
and (n2656,n497,n2632);
and (n2657,n2631,n2632);
or (n2658,n2659,n2660,n2661);
and (n2659,n2636,n2640);
and (n2660,n2640,n2645);
and (n2661,n2636,n2645);
or (n2662,n2663,n2686,n2735);
and (n2663,n2664,n2684);
or (n2664,n2665,n2680,n2683);
and (n2665,n2666,n2668);
xor (n2666,n2667,n426);
xor (n2667,n466,n2642);
or (n2668,n2669,n2676,n2679);
and (n2669,n139,n2670);
or (n2670,n2671,n2673,n2675);
and (n2671,n230,n2672);
not (n2672,n196);
and (n2673,n2672,n2674);
not (n2674,n178);
and (n2675,n230,n2674);
and (n2676,n2670,n2677);
xor (n2677,n2678,n240);
xor (n2678,n11,n155);
and (n2679,n139,n2677);
and (n2680,n2668,n2681);
xor (n2681,n2682,n2625);
xor (n2682,n2612,n2616);
and (n2683,n2666,n2681);
xor (n2684,n2685,n2634);
xor (n2685,n2610,n2629);
and (n2686,n2684,n2687);
or (n2687,n2688,n2699,n2734);
and (n2688,n2689,n2697);
or (n2689,n2690,n2693,n2696);
and (n2690,n2691,n62);
xor (n2691,n2692,n2619);
xor (n2692,n24,n169);
and (n2693,n62,n2694);
xor (n2694,n2695,n2677);
xor (n2695,n139,n2670);
and (n2696,n2691,n2694);
xor (n2697,n2698,n2681);
xor (n2698,n2666,n2668);
and (n2699,n2697,n2700);
or (n2700,n2701,n2730,n2733);
and (n2701,n2702,n2715);
or (n2702,n2703,n2713,n2714);
and (n2703,n2704,n275);
or (n2704,n2705,n2710,n2712);
and (n2705,n2706,n269);
or (n2706,n2707,n2708,n2709);
and (n2707,n214,n259);
not (n2708,n263);
and (n2709,n214,n264);
and (n2710,n269,n2711);
not (n2711,n272);
and (n2712,n2706,n2711);
not (n2713,n310);
and (n2714,n2704,n311);
or (n2715,n2716,n2723,n2729);
and (n2716,n2717,n2721);
or (n2717,n2718,n2719,n2720);
and (n2718,n215,n211);
not (n2719,n229);
and (n2720,n215,n225);
xor (n2721,n2722,n2674);
xor (n2722,n230,n2672);
and (n2723,n2721,n2724);
or (n2724,n2725,n2726,n2728);
and (n2725,n214,n352);
and (n2726,n352,n2727);
not (n2727,n2013);
and (n2728,n214,n2727);
and (n2729,n2717,n2724);
and (n2730,n2715,n2731);
xor (n2731,n2732,n2694);
xor (n2732,n2691,n62);
and (n2733,n2702,n2731);
and (n2734,n2689,n2700);
and (n2735,n2664,n2687);
or (n2736,n2737,n2822);
and (n2737,n2738,n2740);
xor (n2738,n2739,n2687);
xor (n2739,n2664,n2684);
or (n2740,n2741,n2743);
xor (n2741,n2742,n2700);
xor (n2742,n2689,n2697);
or (n2743,n2744,n2766,n2821);
and (n2744,n2745,n2764);
or (n2745,n2746,n2760,n2763);
and (n2746,n2747,n2749);
xor (n2747,n2748,n311);
xor (n2748,n2704,n275);
or (n2749,n2750,n2753,n2759);
and (n2750,n2751,n2016);
xor (n2751,n2752,n2711);
xor (n2752,n2706,n269);
and (n2753,n2016,n2754);
or (n2754,n2755,n2756,n2758);
not (n2755,n391);
and (n2756,n375,n2757);
not (n2757,n372);
and (n2758,n356,n2757);
and (n2759,n2751,n2754);
and (n2760,n2749,n2761);
xor (n2761,n2762,n2724);
xor (n2762,n2717,n2721);
and (n2763,n2747,n2761);
xor (n2764,n2765,n2731);
xor (n2765,n2702,n2715);
and (n2766,n2764,n2767);
or (n2767,n2768,n2783,n2820);
and (n2768,n2769,n2781);
or (n2769,n2770,n2777,n2780);
and (n2770,n2771,n2775);
or (n2771,n2772,n2773,n2774);
and (n2772,n323,n1986);
and (n2773,n1986,n1967);
and (n2774,n323,n1967);
xor (n2775,n2776,n2727);
xor (n2776,n214,n352);
and (n2777,n2775,n2778);
and (n2778,n1962,n2779);
not (n2779,n1960);
and (n2780,n2771,n2778);
xor (n2781,n2782,n2761);
xor (n2782,n2747,n2749);
and (n2783,n2781,n2784);
or (n2784,n2785,n2805,n2819);
and (n2785,n2786,n2803);
or (n2786,n2787,n2792,n2802);
and (n2787,n2788,n1989);
or (n2788,n2789,n2790,n2791);
and (n2789,n340,n331);
not (n2790,n330);
and (n2791,n340,n334);
and (n2792,n1989,n2793);
or (n2793,n2794,n2799,n2801);
and (n2794,n339,n2795);
or (n2795,n2796,n2797,n2798);
and (n2796,n339,n1790);
not (n2797,n1904);
and (n2798,n339,n1794);
and (n2799,n2795,n2800);
not (n2800,n1899);
and (n2801,n339,n2800);
and (n2802,n2788,n2793);
xor (n2803,n2804,n2754);
xor (n2804,n2751,n2016);
and (n2805,n2803,n2806);
or (n2806,n2807,n2811,n2818);
and (n2807,n2808,n2810);
xor (n2808,n2809,n1967);
xor (n2809,n323,n1986);
not (n2810,n1959);
and (n2811,n2810,n2812);
or (n2812,n2813,n2816,n2817);
and (n2813,n2814,n1905);
and (n2814,n1774,n2815);
not (n2815,n1788);
and (n2816,n1905,n1927);
and (n2817,n2814,n1927);
and (n2818,n2808,n2812);
and (n2819,n2786,n2806);
and (n2820,n2769,n2784);
and (n2821,n2745,n2767);
and (n2822,n2823,n2824);
xor (n2823,n2738,n2740);
and (n2824,n2825,n2826);
xnor (n2825,n2741,n2743);
or (n2826,n2827,n3031);
and (n2827,n2828,n2830);
xor (n2828,n2829,n2767);
xor (n2829,n2745,n2764);
or (n2830,n2831,n2906,n3030);
and (n2831,n2832,n2904);
or (n2832,n2833,n2900,n2903);
and (n2833,n2834,n2836);
xor (n2834,n2835,n2778);
xor (n2835,n2771,n2775);
or (n2836,n2837,n2871,n2899);
and (n2837,n2838,n2869);
or (n2838,n2839,n2857,n2868);
and (n2839,n2840,n2849);
and (n2840,n2841,n1814);
or (n2841,n2842,n2847,n2848);
and (n2842,n2843,n1684);
or (n2843,n2844,n2845,n2846);
and (n2844,n1753,n1549);
not (n2845,n1693);
and (n2846,n1753,n1553);
not (n2847,n1826);
and (n2848,n2843,n1688);
or (n2849,n2850,n2855,n2856);
and (n2850,n1854,n2851);
or (n2851,n2852,n2853,n2854);
and (n2852,n1753,n1673);
not (n2853,n1801);
and (n2854,n1753,n1678);
and (n2855,n2851,n1835);
and (n2856,n1854,n1835);
and (n2857,n2849,n2858);
or (n2858,n2859,n2865,n2867);
and (n2859,n2860,n2861);
not (n2860,n1773);
or (n2861,n2862,n2863,n2864);
and (n2862,n1557,n1749);
not (n2863,n1853);
and (n2864,n1557,n1754);
and (n2865,n2861,n2866);
not (n2866,n1830);
and (n2867,n2860,n2866);
and (n2868,n2840,n2858);
xor (n2869,n2870,n2793);
xor (n2870,n2788,n1989);
and (n2871,n2869,n2872);
or (n2872,n2873,n2895,n2898);
and (n2873,n2874,n2876);
xor (n2874,n2875,n2800);
xor (n2875,n339,n2795);
or (n2876,n2877,n2886,n2894);
and (n2877,n2878,n2885);
or (n2878,n2879,n2881,n2884);
and (n2879,n1733,n2880);
not (n2880,n1730);
and (n2881,n2880,n2882);
xor (n2882,n2883,n1678);
xor (n2883,n1753,n1673);
and (n2884,n1733,n2882);
xor (n2885,n2841,n1814);
and (n2886,n2885,n2887);
or (n2887,n2888,n2892,n2893);
and (n2888,n2889,n2890);
not (n2889,n1747);
xor (n2890,n2891,n1688);
xor (n2891,n2843,n1684);
and (n2892,n2890,n1707);
and (n2893,n2889,n1707);
and (n2894,n2878,n2887);
and (n2895,n2876,n2896);
xor (n2896,n2897,n1927);
xor (n2897,n2814,n1905);
and (n2898,n2874,n2896);
and (n2899,n2838,n2872);
and (n2900,n2836,n2901);
xor (n2901,n2902,n2806);
xor (n2902,n2786,n2803);
and (n2903,n2834,n2901);
xor (n2904,n2905,n2784);
xor (n2905,n2769,n2781);
and (n2906,n2904,n2907);
or (n2907,n2908,n2941,n3029);
and (n2908,n2909,n2939);
or (n2909,n2910,n2935,n2938);
and (n2910,n2911,n2913);
xor (n2911,n2912,n2812);
xor (n2912,n2808,n2810);
or (n2913,n2914,n2931,n2934);
and (n2914,n2915,n2917);
xor (n2915,n2916,n2858);
xor (n2916,n2840,n2849);
or (n2917,n2918,n2923,n2930);
and (n2918,n2919,n2921);
xor (n2919,n2920,n1835);
xor (n2920,n1854,n2851);
xor (n2921,n2922,n2866);
xor (n2922,n2860,n2861);
and (n2923,n2921,n2924);
and (n2924,n1698,n2925);
or (n2925,n2926,n2927,n2929);
not (n2926,n1704);
and (n2927,n1564,n2928);
not (n2928,n1547);
and (n2929,n1560,n2928);
and (n2930,n2919,n2924);
and (n2931,n2917,n2932);
xor (n2932,n2933,n2896);
xor (n2933,n2874,n2876);
and (n2934,n2915,n2932);
and (n2935,n2913,n2936);
xor (n2936,n2937,n2872);
xor (n2937,n2838,n2869);
and (n2938,n2911,n2936);
xor (n2939,n2940,n2901);
xor (n2940,n2834,n2836);
and (n2941,n2939,n2942);
or (n2942,n2943,n3000,n3028);
and (n2943,n2944,n2946);
xor (n2944,n2945,n2936);
xor (n2945,n2911,n2913);
or (n2946,n2947,n2979,n2999);
and (n2947,n2948,n2977);
or (n2948,n2949,n2962,n2976);
and (n2949,n2950,n2960);
or (n2950,n2951,n2958,n2959);
and (n2951,n2952,n2956);
or (n2952,n2953,n2954,n2955);
and (n2953,n1612,n1597);
and (n2954,n1597,n1580);
and (n2955,n1612,n1580);
xor (n2956,n2957,n2882);
xor (n2957,n1733,n2880);
and (n2958,n2956,n1758);
and (n2959,n2952,n1758);
xor (n2960,n2961,n2887);
xor (n2961,n2878,n2885);
and (n2962,n2960,n2963);
or (n2963,n2964,n2973,n2975);
and (n2964,n2965,n2971);
or (n2965,n2966,n2967,n2970);
and (n2966,n1602,n1596);
and (n2967,n1596,n2968);
xor (n2968,n2969,n1580);
xor (n2969,n1612,n1597);
and (n2970,n1602,n2968);
xor (n2971,n2972,n1707);
xor (n2972,n2889,n2890);
and (n2973,n2971,n2974);
xor (n2974,n1698,n2925);
and (n2975,n2965,n2974);
and (n2976,n2950,n2963);
xor (n2977,n2978,n2932);
xor (n2978,n2915,n2917);
and (n2979,n2977,n2980);
or (n2980,n2981,n2995,n2998);
and (n2981,n2982,n2984);
xor (n2982,n2983,n2924);
xor (n2983,n2919,n2921);
or (n2984,n2985,n2993,n2994);
and (n2985,n2986,n2988);
xor (n2986,n2987,n1758);
xor (n2987,n2952,n2956);
or (n2988,n2989,n2990,n2992);
not (n2989,n1657);
and (n2990,n1572,n2991);
not (n2991,n1545);
and (n2992,n1568,n2991);
and (n2993,n2988,n1659);
and (n2994,n2986,n1659);
and (n2995,n2984,n2996);
xor (n2996,n2997,n2963);
xor (n2997,n2950,n2960);
and (n2998,n2982,n2996);
and (n2999,n2948,n2980);
and (n3000,n2946,n3001);
or (n3001,n3002,n3004);
xor (n3002,n3003,n2980);
xor (n3003,n2948,n2977);
or (n3004,n3005,n3021,n3027);
and (n3005,n3006,n3019);
or (n3006,n3007,n3015,n3018);
and (n3007,n3008,n3010);
xor (n3008,n3009,n2974);
xor (n3009,n2965,n2971);
or (n3010,n3011,n3013,n3014);
and (n3011,n3012,n1644);
not (n3012,n1543);
not (n3013,n1651);
and (n3014,n3012,n1576);
and (n3015,n3010,n3016);
xor (n3016,n3017,n1659);
xor (n3017,n2986,n2988);
and (n3018,n3008,n3016);
xor (n3019,n3020,n2996);
xor (n3020,n2982,n2984);
and (n3021,n3019,n3022);
or (n3022,n3023,n3025);
or (n3023,n1537,n3024);
not (n3024,n1541);
xor (n3025,n3026,n3016);
xor (n3026,n3008,n3010);
and (n3027,n3006,n3022);
and (n3028,n2944,n3001);
and (n3029,n2909,n2942);
and (n3030,n2832,n2907);
and (n3031,n3032,n3033);
xor (n3032,n2828,n2830);
and (n3033,n3034,n3036);
xor (n3034,n3035,n2907);
xor (n3035,n2832,n2904);
or (n3036,n3037,n3039);
xor (n3037,n3038,n2942);
xor (n3038,n2909,n2939);
and (n3039,n3040,n3041);
not (n3040,n3037);
and (n3041,n3042,n3044);
xor (n3042,n3043,n3001);
xor (n3043,n2944,n2946);
and (n3044,n3045,n3046);
xnor (n3045,n3002,n3004);
and (n3046,n3047,n3049);
xor (n3047,n3048,n3022);
xor (n3048,n3006,n3019);
and (n3049,n3050,n3051);
xnor (n3050,n3023,n3025);
and (n3051,n3052,n3055);
not (n3052,n3053);
nand (n3053,n3054,n2066);
not (n3054,n1536);
nand (n3055,n563,n3056);
nand (n3056,n2513,n2092);
endmodule
