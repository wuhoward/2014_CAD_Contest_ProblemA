module top (out,n12,n15,n17,n18,n23,n24,n32,n34,n35
        ,n38,n78,n82,n128,n158,n211,n320,n323,n328,n336
        ,n339,n381,n454,n506);
output out;
input n12;
input n15;
input n17;
input n18;
input n23;
input n24;
input n32;
input n34;
input n35;
input n38;
input n78;
input n82;
input n128;
input n158;
input n211;
input n320;
input n323;
input n328;
input n336;
input n339;
input n381;
input n454;
input n506;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n13;
wire n14;
wire n16;
wire n19;
wire n20;
wire n21;
wire n22;
wire n25;
wire n26;
wire n27;
wire n28;
wire n29;
wire n30;
wire n31;
wire n33;
wire n36;
wire n37;
wire n39;
wire n40;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n79;
wire n80;
wire n81;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n321;
wire n322;
wire n324;
wire n325;
wire n326;
wire n327;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n337;
wire n338;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
xor (out,n0,n672);
xor (n0,n1,n605);
xor (n1,n2,n310);
xor (n2,n3,n101);
xor (n3,n4,n66);
xor (n4,n5,n56);
xor (n5,n6,n53);
or (n6,n7,n44,n52);
and (n7,n8,n27);
or (n8,n9,n19,n26);
and (n9,n10,n16);
nor (n10,n11,n13);
not (n11,n12);
and (n13,n14,n12);
not (n14,n15);
and (n16,n17,n18);
and (n19,n16,n20);
nor (n20,n21,n25);
and (n21,n22,n24);
not (n22,n23);
not (n25,n24);
and (n26,n10,n20);
or (n27,n28,n41,n43);
and (n28,n29,n40);
or (n29,n30,n36,n39);
and (n30,n31,n33);
and (n31,n17,n32);
and (n33,n34,n35);
and (n36,n33,n37);
and (n37,n38,n24);
and (n39,n31,n37);
and (n40,n34,n32);
and (n41,n40,n42);
and (n42,n38,n35);
and (n43,n29,n42);
and (n44,n27,n45);
xor (n45,n46,n51);
xor (n46,n47,n50);
nor (n47,n48,n49);
not (n48,n17);
and (n49,n14,n17);
and (n50,n34,n18);
and (n51,n38,n32);
and (n52,n8,n45);
nor (n53,n54,n55);
and (n54,n22,n32);
not (n55,n32);
xor (n56,n57,n65);
xor (n57,n58,n62);
or (n58,n59,n60,n61);
and (n59,n47,n50);
and (n60,n50,n51);
and (n61,n47,n51);
nor (n62,n63,n64);
not (n63,n34);
and (n64,n14,n34);
and (n65,n38,n18);
or (n66,n67,n97,n100);
and (n67,n68,n94);
or (n68,n69,n90,n93);
and (n69,n70,n88);
or (n70,n71,n84,n87);
and (n71,n72,n80);
or (n72,n73,n76,n79);
and (n73,n74,n75);
and (n74,n17,n35);
and (n75,n34,n24);
and (n76,n75,n77);
and (n77,n38,n78);
and (n79,n74,n77);
and (n80,n81,n83);
and (n81,n82,n18);
and (n83,n12,n32);
and (n84,n80,n85);
xor (n85,n86,n37);
xor (n86,n31,n33);
and (n87,n72,n85);
xor (n88,n89,n20);
xor (n89,n10,n16);
and (n90,n88,n91);
xor (n91,n92,n42);
xor (n92,n29,n40);
and (n93,n70,n91);
nor (n94,n95,n96);
and (n95,n22,n35);
not (n96,n35);
and (n97,n94,n98);
xor (n98,n99,n45);
xor (n99,n8,n27);
and (n100,n68,n98);
or (n101,n102,n145);
and (n102,n103,n105);
xor (n103,n104,n98);
xor (n104,n68,n94);
or (n105,n106,n141,n144);
and (n106,n107,n118);
or (n107,n108,n113,n117);
and (n108,n109,n112);
nor (n109,n110,n111);
not (n110,n82);
and (n111,n14,n82);
and (n112,n12,n18);
and (n113,n112,n114);
nor (n114,n115,n116);
and (n115,n22,n78);
not (n116,n78);
and (n117,n109,n114);
or (n118,n119,n137,n140);
and (n119,n120,n135);
or (n120,n121,n132,n134);
and (n121,n122,n130);
or (n122,n123,n126,n129);
and (n123,n124,n125);
and (n124,n17,n24);
and (n125,n34,n78);
and (n126,n125,n127);
and (n127,n38,n128);
and (n129,n124,n127);
xor (n130,n131,n77);
xor (n131,n74,n75);
and (n132,n130,n133);
xor (n133,n81,n83);
and (n134,n122,n133);
xor (n135,n136,n114);
xor (n136,n109,n112);
and (n137,n135,n138);
xor (n138,n139,n85);
xor (n139,n72,n80);
and (n140,n120,n138);
and (n141,n118,n142);
xor (n142,n143,n91);
xor (n143,n70,n88);
and (n144,n107,n142);
and (n145,n146,n147);
xor (n146,n103,n105);
or (n147,n148,n194);
and (n148,n149,n151);
xor (n149,n150,n142);
xor (n150,n107,n118);
or (n151,n152,n190,n193);
and (n152,n153,n171);
or (n153,n154,n166,n170);
and (n154,n155,n163);
or (n155,n156,n160,n162);
and (n156,n157,n159);
and (n157,n158,n18);
and (n159,n82,n32);
and (n160,n159,n161);
and (n161,n12,n35);
and (n162,n157,n161);
nor (n163,n164,n165);
not (n164,n158);
and (n165,n14,n158);
and (n166,n163,n167);
nor (n167,n168,n169);
and (n168,n22,n128);
not (n169,n128);
and (n170,n155,n167);
or (n171,n172,n186,n189);
and (n172,n173,n184);
or (n173,n174,n180,n183);
and (n174,n175,n178);
and (n175,n176,n177);
and (n176,n17,n78);
and (n177,n34,n128);
xor (n178,n179,n161);
xor (n179,n157,n159);
and (n180,n178,n181);
xor (n181,n182,n127);
xor (n182,n124,n125);
and (n183,n175,n181);
xor (n184,n185,n167);
xor (n185,n155,n163);
and (n186,n184,n187);
xor (n187,n188,n133);
xor (n188,n122,n130);
and (n189,n173,n187);
and (n190,n171,n191);
xor (n191,n192,n138);
xor (n192,n120,n135);
and (n193,n153,n191);
and (n194,n195,n196);
xor (n195,n149,n151);
or (n196,n197,n216);
and (n197,n198,n200);
xor (n198,n199,n191);
xor (n199,n153,n171);
and (n200,n201,n214);
or (n201,n202,n208,n213);
and (n202,n203,n206);
and (n203,n204,n205);
and (n204,n12,n24);
xor (n205,n176,n177);
xor (n206,n207,n181);
xor (n207,n175,n178);
and (n208,n206,n209);
nor (n209,n210,n212);
not (n210,n211);
and (n212,n14,n211);
and (n213,n203,n209);
xor (n214,n215,n187);
xor (n215,n173,n184);
and (n216,n217,n218);
xor (n217,n198,n200);
or (n218,n219,n249);
and (n219,n220,n221);
xor (n220,n201,n214);
or (n221,n222,n245,n248);
and (n222,n223,n230);
or (n223,n224,n227,n229);
and (n224,n225,n226);
and (n225,n211,n18);
and (n226,n158,n32);
and (n227,n226,n228);
and (n228,n82,n35);
and (n229,n225,n228);
or (n230,n231,n242,n244);
and (n231,n232,n240);
or (n232,n233,n236,n239);
and (n233,n234,n235);
and (n234,n82,n78);
and (n235,n12,n128);
and (n236,n237,n238);
and (n237,n12,n78);
and (n238,n17,n128);
and (n239,n233,n238);
xor (n240,n241,n228);
xor (n241,n225,n226);
and (n242,n240,n243);
xor (n243,n204,n205);
and (n244,n232,n243);
and (n245,n230,n246);
xor (n246,n247,n209);
xor (n247,n203,n206);
and (n248,n223,n246);
and (n249,n250,n251);
xor (n250,n220,n221);
or (n251,n252,n280);
and (n252,n253,n255);
xor (n253,n254,n246);
xor (n254,n223,n230);
or (n255,n256,n276,n279);
and (n256,n257,n260);
and (n257,n258,n259);
and (n258,n158,n35);
and (n259,n82,n24);
or (n260,n261,n272,n275);
and (n261,n262,n271);
or (n262,n263,n268,n270);
and (n263,n264,n267);
and (n264,n265,n266);
and (n265,n158,n78);
and (n266,n82,n128);
and (n267,n158,n24);
and (n268,n267,n269);
xor (n269,n234,n235);
and (n270,n264,n269);
xor (n271,n258,n259);
and (n272,n271,n273);
xor (n273,n274,n238);
xor (n274,n233,n237);
and (n275,n262,n273);
and (n276,n260,n277);
xor (n277,n278,n243);
xor (n278,n232,n240);
and (n279,n257,n277);
and (n280,n281,n282);
xor (n281,n253,n255);
or (n282,n283,n305);
and (n283,n284,n286);
xor (n284,n285,n277);
xor (n285,n257,n260);
and (n286,n287,n303);
or (n287,n288,n299,n302);
and (n288,n289,n298);
or (n289,n290,n295,n297);
and (n290,n291,n294);
and (n291,n292,n293);
and (n292,n211,n78);
and (n293,n158,n128);
and (n294,n211,n24);
and (n295,n294,n296);
xor (n296,n265,n266);
and (n297,n291,n296);
and (n298,n211,n35);
and (n299,n298,n300);
xor (n300,n301,n269);
xor (n301,n264,n267);
and (n302,n289,n300);
xor (n303,n304,n273);
xor (n304,n262,n271);
and (n305,n306,n307);
xor (n306,n284,n286);
and (n307,n308,n309);
and (n308,n211,n32);
xor (n309,n287,n303);
xor (n310,n311,n399);
xor (n311,n312,n366);
xor (n312,n313,n356);
xor (n313,n314,n354);
or (n314,n315,n345,n353);
and (n315,n316,n330);
or (n316,n317,n324,n329);
and (n317,n318,n322);
nor (n318,n319,n321);
not (n319,n320);
and (n321,n14,n320);
and (n322,n323,n18);
and (n324,n322,n325);
nor (n325,n326,n25);
and (n326,n327,n24);
not (n327,n328);
and (n329,n318,n325);
or (n330,n331,n342,n344);
and (n331,n332,n341);
or (n332,n333,n337,n340);
and (n333,n334,n335);
and (n334,n323,n32);
and (n335,n336,n35);
and (n337,n335,n338);
and (n338,n339,n24);
and (n340,n334,n338);
and (n341,n336,n32);
and (n342,n341,n343);
and (n343,n339,n35);
and (n344,n332,n343);
and (n345,n330,n346);
xor (n346,n347,n352);
xor (n347,n348,n351);
nor (n348,n349,n350);
not (n349,n323);
and (n350,n14,n323);
and (n351,n336,n18);
and (n352,n339,n32);
and (n353,n316,n346);
nor (n354,n355,n55);
and (n355,n327,n32);
xor (n356,n357,n365);
xor (n357,n358,n362);
or (n358,n359,n360,n361);
and (n359,n348,n351);
and (n360,n351,n352);
and (n361,n348,n352);
nor (n362,n363,n364);
not (n363,n336);
and (n364,n14,n336);
and (n365,n339,n18);
or (n366,n367,n395,n398);
and (n367,n368,n393);
or (n368,n369,n389,n392);
and (n369,n370,n387);
or (n370,n371,n383,n386);
and (n371,n372,n379);
or (n372,n373,n376,n378);
and (n373,n374,n375);
and (n374,n323,n35);
and (n375,n336,n24);
and (n376,n375,n377);
and (n377,n339,n78);
and (n378,n374,n377);
and (n379,n380,n382);
and (n380,n381,n18);
and (n382,n320,n32);
and (n383,n379,n384);
xor (n384,n385,n338);
xor (n385,n334,n335);
and (n386,n372,n384);
xor (n387,n388,n325);
xor (n388,n318,n322);
and (n389,n387,n390);
xor (n390,n391,n343);
xor (n391,n332,n341);
and (n392,n370,n390);
nor (n393,n394,n96);
and (n394,n327,n35);
and (n395,n393,n396);
xor (n396,n397,n346);
xor (n397,n316,n330);
and (n398,n368,n396);
or (n399,n400,n441);
and (n400,n401,n403);
xor (n401,n402,n396);
xor (n402,n368,n393);
or (n403,n404,n437,n440);
and (n404,n405,n415);
or (n405,n406,n411,n414);
and (n406,n407,n410);
nor (n407,n408,n409);
not (n408,n381);
and (n409,n14,n381);
and (n410,n320,n18);
and (n411,n410,n412);
nor (n412,n413,n116);
and (n413,n327,n78);
and (n414,n407,n412);
or (n415,n416,n433,n436);
and (n416,n417,n431);
or (n417,n418,n428,n430);
and (n418,n419,n426);
or (n419,n420,n423,n425);
and (n420,n421,n422);
and (n421,n323,n24);
and (n422,n336,n78);
and (n423,n422,n424);
and (n424,n339,n128);
and (n425,n421,n424);
xor (n426,n427,n377);
xor (n427,n374,n375);
and (n428,n426,n429);
xor (n429,n380,n382);
and (n430,n419,n429);
xor (n431,n432,n412);
xor (n432,n407,n410);
and (n433,n431,n434);
xor (n434,n435,n384);
xor (n435,n372,n379);
and (n436,n417,n434);
and (n437,n415,n438);
xor (n438,n439,n390);
xor (n439,n370,n387);
and (n440,n405,n438);
and (n441,n442,n443);
xor (n442,n401,n403);
or (n443,n444,n489);
and (n444,n445,n447);
xor (n445,n446,n438);
xor (n446,n405,n415);
or (n447,n448,n485,n488);
and (n448,n449,n466);
or (n449,n450,n462,n465);
and (n450,n451,n459);
or (n451,n452,n456,n458);
and (n452,n453,n455);
and (n453,n454,n18);
and (n455,n381,n32);
and (n456,n455,n457);
and (n457,n320,n35);
and (n458,n453,n457);
nor (n459,n460,n461);
not (n460,n454);
and (n461,n14,n454);
and (n462,n459,n463);
nor (n463,n464,n169);
and (n464,n327,n128);
and (n465,n451,n463);
or (n466,n467,n481,n484);
and (n467,n468,n479);
or (n468,n469,n475,n478);
and (n469,n470,n473);
and (n470,n471,n472);
and (n471,n323,n78);
and (n472,n336,n128);
xor (n473,n474,n457);
xor (n474,n453,n455);
and (n475,n473,n476);
xor (n476,n477,n424);
xor (n477,n421,n422);
and (n478,n470,n476);
xor (n479,n480,n463);
xor (n480,n451,n459);
and (n481,n479,n482);
xor (n482,n483,n429);
xor (n483,n419,n426);
and (n484,n468,n482);
and (n485,n466,n486);
xor (n486,n487,n434);
xor (n487,n417,n431);
and (n488,n449,n486);
and (n489,n490,n491);
xor (n490,n445,n447);
or (n491,n492,n511);
and (n492,n493,n495);
xor (n493,n494,n486);
xor (n494,n449,n466);
and (n495,n496,n509);
or (n496,n497,n503,n508);
and (n497,n498,n501);
and (n498,n499,n500);
and (n499,n320,n24);
xor (n500,n471,n472);
xor (n501,n502,n476);
xor (n502,n470,n473);
and (n503,n501,n504);
nor (n504,n505,n507);
not (n505,n506);
and (n507,n14,n506);
and (n508,n498,n504);
xor (n509,n510,n482);
xor (n510,n468,n479);
and (n511,n512,n513);
xor (n512,n493,n495);
or (n513,n514,n544);
and (n514,n515,n516);
xor (n515,n496,n509);
or (n516,n517,n540,n543);
and (n517,n518,n525);
or (n518,n519,n522,n524);
and (n519,n520,n521);
and (n520,n506,n18);
and (n521,n454,n32);
and (n522,n521,n523);
and (n523,n381,n35);
and (n524,n520,n523);
or (n525,n526,n537,n539);
and (n526,n527,n535);
or (n527,n528,n531,n534);
and (n528,n529,n530);
and (n529,n381,n78);
and (n530,n320,n128);
and (n531,n532,n533);
and (n532,n320,n78);
and (n533,n323,n128);
and (n534,n528,n533);
xor (n535,n536,n523);
xor (n536,n520,n521);
and (n537,n535,n538);
xor (n538,n499,n500);
and (n539,n527,n538);
and (n540,n525,n541);
xor (n541,n542,n504);
xor (n542,n498,n501);
and (n543,n518,n541);
and (n544,n545,n546);
xor (n545,n515,n516);
or (n546,n547,n575);
and (n547,n548,n550);
xor (n548,n549,n541);
xor (n549,n518,n525);
or (n550,n551,n571,n574);
and (n551,n552,n555);
and (n552,n553,n554);
and (n553,n454,n35);
and (n554,n381,n24);
or (n555,n556,n567,n570);
and (n556,n557,n566);
or (n557,n558,n563,n565);
and (n558,n559,n562);
and (n559,n560,n561);
and (n560,n454,n78);
and (n561,n381,n128);
and (n562,n454,n24);
and (n563,n562,n564);
xor (n564,n529,n530);
and (n565,n559,n564);
xor (n566,n553,n554);
and (n567,n566,n568);
xor (n568,n569,n533);
xor (n569,n528,n532);
and (n570,n557,n568);
and (n571,n555,n572);
xor (n572,n573,n538);
xor (n573,n527,n535);
and (n574,n552,n572);
and (n575,n576,n577);
xor (n576,n548,n550);
or (n577,n578,n600);
and (n578,n579,n581);
xor (n579,n580,n572);
xor (n580,n552,n555);
and (n581,n582,n598);
or (n582,n583,n594,n597);
and (n583,n584,n593);
or (n584,n585,n590,n592);
and (n585,n586,n589);
and (n586,n587,n588);
and (n587,n506,n78);
and (n588,n454,n128);
and (n589,n506,n24);
and (n590,n589,n591);
xor (n591,n560,n561);
and (n592,n586,n591);
and (n593,n506,n35);
and (n594,n593,n595);
xor (n595,n596,n564);
xor (n596,n559,n562);
and (n597,n584,n595);
xor (n598,n599,n568);
xor (n599,n557,n566);
and (n600,n601,n602);
xor (n601,n579,n581);
and (n602,n603,n604);
and (n603,n506,n32);
xor (n604,n582,n598);
or (n605,n606,n609,n671);
and (n606,n607,n608);
xor (n607,n146,n147);
xor (n608,n442,n443);
and (n609,n608,n610);
or (n610,n611,n614,n670);
and (n611,n612,n613);
xor (n612,n195,n196);
xor (n613,n490,n491);
and (n614,n613,n615);
or (n615,n616,n619,n669);
and (n616,n617,n618);
xor (n617,n217,n218);
xor (n618,n512,n513);
and (n619,n618,n620);
or (n620,n621,n624,n668);
and (n621,n622,n623);
xor (n622,n250,n251);
xor (n623,n545,n546);
and (n624,n623,n625);
or (n625,n626,n629,n667);
and (n626,n627,n628);
xor (n627,n281,n282);
xor (n628,n576,n577);
and (n629,n628,n630);
or (n630,n631,n634,n666);
and (n631,n632,n633);
xor (n632,n306,n307);
xor (n633,n601,n602);
and (n634,n633,n635);
or (n635,n636,n639,n665);
and (n636,n637,n638);
xor (n637,n308,n309);
xor (n638,n603,n604);
and (n639,n638,n640);
or (n640,n641,n646,n664);
and (n641,n642,n644);
xor (n642,n643,n300);
xor (n643,n289,n298);
xor (n644,n645,n595);
xor (n645,n584,n593);
and (n646,n644,n647);
or (n647,n648,n653,n663);
and (n648,n649,n651);
xor (n649,n650,n296);
xor (n650,n291,n294);
xor (n651,n652,n591);
xor (n652,n586,n589);
and (n653,n651,n654);
or (n654,n655,n658,n662);
and (n655,n656,n657);
xor (n656,n292,n293);
xor (n657,n587,n588);
and (n658,n657,n659);
and (n659,n660,n661);
and (n660,n211,n128);
and (n661,n506,n128);
and (n662,n656,n659);
and (n663,n649,n654);
and (n664,n642,n647);
and (n665,n637,n640);
and (n666,n632,n635);
and (n667,n627,n630);
and (n668,n622,n625);
and (n669,n617,n620);
and (n670,n612,n615);
and (n671,n607,n610);
xor (n672,n673,n821);
xor (n673,n674,n782);
xor (n674,n675,n765);
xor (n675,n676,n763);
or (n676,n677,n753,n762);
and (n677,n678,n740);
or (n678,n679,n733,n739);
and (n679,n680,n718);
or (n680,n681,n709,n717);
and (n681,n682,n702);
and (n682,n683,n35);
xor (n683,n684,n685);
xor (n684,n34,n336);
or (n685,n686,n687,n701);
and (n686,n17,n323);
and (n687,n323,n688);
or (n688,n689,n690,n700);
and (n689,n12,n320);
and (n690,n320,n691);
or (n691,n692,n693,n699);
and (n692,n82,n381);
and (n693,n381,n694);
or (n694,n695,n696,n698);
and (n695,n158,n454);
and (n696,n454,n697);
and (n697,n211,n506);
and (n698,n158,n697);
and (n699,n82,n694);
and (n700,n12,n691);
and (n701,n17,n688);
and (n702,n703,n24);
xor (n703,n704,n705);
xor (n704,n38,n339);
or (n705,n706,n707,n708);
and (n706,n34,n336);
and (n707,n336,n685);
and (n708,n34,n685);
and (n709,n702,n710);
and (n710,n711,n78);
xor (n711,n712,n713);
xor (n712,n23,n328);
or (n713,n714,n715,n716);
and (n714,n38,n339);
and (n715,n339,n705);
and (n716,n38,n705);
and (n717,n682,n710);
or (n718,n719,n728,n732);
and (n719,n720,n725);
nor (n720,n721,n724);
not (n721,n722);
xor (n722,n723,n694);
xor (n723,n82,n381);
and (n724,n14,n722);
and (n725,n726,n18);
xor (n726,n727,n691);
xor (n727,n12,n320);
and (n728,n725,n729);
and (n729,n730,n32);
xor (n730,n731,n688);
xor (n731,n17,n323);
and (n732,n720,n729);
and (n733,n718,n734);
xor (n734,n735,n738);
xor (n735,n736,n737);
and (n736,n683,n32);
and (n737,n703,n35);
and (n738,n711,n24);
and (n739,n680,n734);
xor (n740,n741,n746);
xor (n741,n742,n745);
nor (n742,n743,n744);
not (n743,n730);
and (n744,n14,n730);
and (n745,n683,n18);
nor (n746,n747,n25);
and (n747,n748,n24);
not (n748,n749);
or (n749,n750,n751,n752);
and (n750,n23,n328);
and (n751,n328,n713);
and (n752,n23,n713);
and (n753,n740,n754);
xor (n754,n755,n761);
xor (n755,n756,n760);
or (n756,n757,n758,n759);
and (n757,n736,n737);
and (n758,n737,n738);
and (n759,n736,n738);
and (n760,n703,n32);
and (n761,n711,n35);
and (n762,n678,n754);
nor (n763,n764,n96);
and (n764,n748,n35);
xor (n765,n766,n775);
xor (n766,n767,n771);
or (n767,n768,n769,n770);
and (n768,n742,n745);
and (n769,n745,n746);
and (n770,n742,n746);
or (n771,n772,n773,n774);
and (n772,n756,n760);
and (n773,n760,n761);
and (n774,n756,n761);
xor (n775,n776,n781);
xor (n776,n777,n780);
nor (n777,n778,n779);
not (n778,n683);
and (n779,n14,n683);
and (n780,n703,n18);
and (n781,n711,n32);
or (n782,n783,n817,n820);
and (n783,n784,n794);
or (n784,n785,n790,n793);
and (n785,n786,n789);
nor (n786,n787,n788);
not (n787,n726);
and (n788,n14,n726);
and (n789,n730,n18);
and (n790,n789,n791);
nor (n791,n792,n116);
and (n792,n748,n78);
and (n793,n786,n791);
or (n794,n795,n813,n816);
and (n795,n796,n811);
or (n796,n797,n807,n810);
and (n797,n798,n805);
or (n798,n799,n802,n804);
and (n799,n800,n801);
and (n800,n683,n24);
and (n801,n703,n78);
and (n802,n801,n803);
and (n803,n711,n128);
and (n804,n800,n803);
xor (n805,n806,n710);
xor (n806,n682,n702);
and (n807,n805,n808);
xor (n808,n809,n729);
xor (n809,n720,n725);
and (n810,n798,n808);
xor (n811,n812,n791);
xor (n812,n786,n789);
and (n813,n811,n814);
xor (n814,n815,n734);
xor (n815,n680,n718);
and (n816,n796,n814);
and (n817,n794,n818);
xor (n818,n819,n754);
xor (n819,n678,n740);
and (n820,n784,n818);
or (n821,n822,n861);
and (n822,n823,n825);
xor (n823,n824,n818);
xor (n824,n784,n794);
or (n825,n826,n857,n860);
and (n826,n827,n837);
and (n827,n828,n835);
or (n828,n829,n832,n834);
and (n829,n830,n831);
and (n830,n722,n18);
and (n831,n726,n32);
and (n832,n831,n833);
and (n833,n730,n35);
and (n834,n830,n833);
nor (n835,n836,n169);
and (n836,n748,n128);
or (n837,n838,n854,n856);
and (n838,n839,n852);
or (n839,n840,n848,n851);
and (n840,n841,n846);
nor (n841,n842,n845);
not (n842,n843);
xor (n843,n844,n697);
xor (n844,n158,n454);
and (n845,n14,n843);
xor (n846,n847,n803);
xor (n847,n800,n801);
and (n848,n846,n849);
xor (n849,n850,n833);
xor (n850,n830,n831);
and (n851,n841,n849);
xor (n852,n853,n808);
xor (n853,n798,n805);
and (n854,n852,n855);
xor (n855,n828,n835);
and (n856,n839,n855);
and (n857,n837,n858);
xor (n858,n859,n814);
xor (n859,n796,n811);
and (n860,n827,n858);
and (n861,n862,n863);
xor (n862,n823,n825);
or (n863,n864,n901);
and (n864,n865,n867);
xor (n865,n866,n858);
xor (n866,n827,n837);
or (n867,n868,n897,n900);
and (n868,n869,n880);
and (n869,n870,n877);
or (n870,n871,n874,n876);
and (n871,n872,n873);
and (n872,n722,n32);
and (n873,n726,n35);
and (n874,n873,n875);
and (n875,n730,n24);
and (n876,n872,n875);
and (n877,n878,n879);
and (n878,n683,n78);
and (n879,n703,n128);
or (n880,n881,n893,n896);
and (n881,n882,n892);
or (n882,n883,n889,n891);
and (n883,n884,n887);
and (n884,n885,n886);
and (n885,n730,n78);
and (n886,n683,n128);
xor (n887,n888,n875);
xor (n888,n872,n873);
and (n889,n887,n890);
xor (n890,n878,n879);
and (n891,n884,n890);
xor (n892,n870,n877);
and (n893,n892,n894);
xor (n894,n895,n849);
xor (n895,n841,n846);
and (n896,n882,n894);
and (n897,n880,n898);
xor (n898,n899,n855);
xor (n899,n839,n852);
and (n900,n869,n898);
and (n901,n902,n903);
xor (n902,n865,n867);
or (n903,n904,n929);
and (n904,n905,n907);
xor (n905,n906,n898);
xor (n906,n869,n880);
or (n907,n908,n925,n928);
and (n908,n909,n915);
and (n909,n910,n914);
nor (n910,n911,n913);
not (n911,n912);
xor (n912,n211,n506);
and (n913,n14,n912);
and (n914,n843,n18);
or (n915,n916,n922,n924);
and (n916,n917,n920);
and (n917,n918,n919);
and (n918,n726,n24);
xor (n919,n885,n886);
xor (n920,n921,n890);
xor (n921,n884,n887);
and (n922,n920,n923);
xor (n923,n910,n914);
and (n924,n917,n923);
and (n925,n915,n926);
xor (n926,n927,n894);
xor (n927,n882,n892);
and (n928,n909,n926);
and (n929,n930,n931);
xor (n930,n905,n907);
or (n931,n932,n963);
and (n932,n933,n935);
xor (n933,n934,n926);
xor (n934,n909,n915);
or (n935,n936,n959,n962);
and (n936,n937,n944);
or (n937,n938,n941,n943);
and (n938,n939,n940);
and (n939,n912,n18);
and (n940,n843,n32);
and (n941,n940,n942);
and (n942,n722,n35);
and (n943,n939,n942);
or (n944,n945,n956,n958);
and (n945,n946,n954);
or (n946,n947,n950,n953);
and (n947,n948,n949);
and (n948,n722,n78);
and (n949,n726,n128);
and (n950,n951,n952);
and (n951,n726,n78);
and (n952,n730,n128);
and (n953,n947,n952);
xor (n954,n955,n942);
xor (n955,n939,n940);
and (n956,n954,n957);
xor (n957,n918,n919);
and (n958,n946,n957);
and (n959,n944,n960);
xor (n960,n961,n923);
xor (n961,n917,n920);
and (n962,n937,n960);
and (n963,n964,n965);
xor (n964,n933,n935);
or (n965,n966,n994);
and (n966,n967,n969);
xor (n967,n968,n960);
xor (n968,n937,n944);
or (n969,n970,n990,n993);
and (n970,n971,n974);
and (n971,n972,n973);
and (n972,n843,n35);
and (n973,n722,n24);
or (n974,n975,n986,n989);
and (n975,n976,n985);
or (n976,n977,n982,n984);
and (n977,n978,n981);
and (n978,n979,n980);
and (n979,n843,n78);
and (n980,n722,n128);
and (n981,n843,n24);
and (n982,n981,n983);
xor (n983,n948,n949);
and (n984,n978,n983);
xor (n985,n972,n973);
and (n986,n985,n987);
xor (n987,n988,n952);
xor (n988,n947,n951);
and (n989,n976,n987);
and (n990,n974,n991);
xor (n991,n992,n957);
xor (n992,n946,n954);
and (n993,n971,n991);
and (n994,n995,n996);
xor (n995,n967,n969);
or (n996,n997,n1019);
and (n997,n998,n1000);
xor (n998,n999,n991);
xor (n999,n971,n974);
and (n1000,n1001,n1017);
or (n1001,n1002,n1013,n1016);
and (n1002,n1003,n1012);
or (n1003,n1004,n1009,n1011);
and (n1004,n1005,n1008);
and (n1005,n1006,n1007);
and (n1006,n912,n78);
and (n1007,n843,n128);
and (n1008,n912,n24);
and (n1009,n1008,n1010);
xor (n1010,n979,n980);
and (n1011,n1005,n1010);
and (n1012,n912,n35);
and (n1013,n1012,n1014);
xor (n1014,n1015,n983);
xor (n1015,n978,n981);
and (n1016,n1003,n1014);
xor (n1017,n1018,n987);
xor (n1018,n976,n985);
and (n1019,n1020,n1021);
xor (n1020,n998,n1000);
and (n1021,n1022,n1023);
and (n1022,n912,n32);
xor (n1023,n1001,n1017);
endmodule
