module top (out,n3,n4,n5,n23,n24,n29,n34,n43,n56
        ,n57,n68,n75,n76,n77,n79,n89,n91,n99,n106
        ,n115,n122,n131,n138,n142,n147,n186,n204,n227,n252);
output out;
input n3;
input n4;
input n5;
input n23;
input n24;
input n29;
input n34;
input n43;
input n56;
input n57;
input n68;
input n75;
input n76;
input n77;
input n79;
input n89;
input n91;
input n99;
input n106;
input n115;
input n122;
input n131;
input n138;
input n142;
input n147;
input n186;
input n204;
input n227;
input n252;
wire n0;
wire n1;
wire n2;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n25;
wire n26;
wire n27;
wire n28;
wire n30;
wire n31;
wire n32;
wire n33;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n78;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n90;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n139;
wire n140;
wire n141;
wire n143;
wire n144;
wire n145;
wire n146;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
xnor (out,n0,n627);
nor (n0,n1,n6);
and (n1,n2,n5);
nor (n2,n3,n4);
and (n6,n7,n624);
nand (n7,n8,n623);
or (n8,n9,n334);
not (n9,n10);
nand (n10,n11,n333);
or (n11,n12,n284);
xor (n12,n13,n210);
xor (n13,n14,n151);
xor (n14,n15,n80);
xor (n15,n16,n45);
nand (n16,n17,n37);
or (n17,n18,n31);
not (n18,n19);
nor (n19,n20,n26);
nor (n20,n21,n25);
and (n21,n22,n24);
not (n22,n23);
nor (n25,n24,n22);
nand (n26,n27,n30);
or (n27,n28,n23);
not (n28,n29);
nand (n30,n28,n23);
nor (n31,n32,n35);
and (n32,n33,n34);
not (n33,n24);
and (n35,n24,n36);
not (n36,n34);
or (n37,n38,n39);
not (n38,n26);
not (n39,n40);
nor (n40,n41,n44);
and (n41,n42,n33);
not (n42,n43);
and (n44,n24,n43);
and (n45,n46,n70);
nand (n46,n47,n63);
or (n47,n48,n52);
not (n48,n49);
nor (n49,n50,n51);
and (n50,n42,n28);
and (n51,n29,n43);
nand (n52,n53,n60);
nor (n53,n54,n58);
and (n54,n55,n57);
not (n55,n56);
and (n58,n56,n59);
not (n59,n57);
nand (n60,n61,n62);
or (n61,n59,n29);
nand (n62,n29,n59);
nand (n63,n64,n65);
not (n64,n53);
nor (n65,n66,n69);
and (n66,n67,n28);
not (n67,n68);
and (n69,n29,n68);
not (n70,n71);
nand (n71,n72,n79);
nand (n72,n73,n78);
or (n73,n74,n77);
and (n74,n75,n76);
or (n78,n75,n76);
or (n80,n81,n150);
and (n81,n82,n133);
xor (n82,n83,n109);
nand (n83,n84,n102);
or (n84,n85,n97);
not (n85,n86);
nor (n86,n87,n94);
nor (n87,n88,n92);
and (n88,n89,n90);
not (n90,n91);
and (n92,n91,n93);
not (n93,n89);
nand (n94,n95,n96);
or (n95,n33,n89);
nand (n96,n33,n89);
nor (n97,n98,n100);
and (n98,n90,n99);
and (n100,n91,n101);
not (n101,n99);
or (n102,n103,n104);
not (n103,n94);
nor (n104,n105,n107);
and (n105,n90,n106);
and (n107,n91,n108);
not (n108,n106);
nand (n109,n110,n127);
or (n110,n111,n118);
not (n111,n112);
nor (n112,n113,n117);
and (n113,n114,n116);
not (n114,n115);
not (n116,n75);
and (n117,n75,n115);
nand (n118,n119,n124);
not (n119,n120);
nand (n120,n121,n123);
or (n121,n90,n122);
nand (n123,n122,n90);
nand (n124,n125,n126);
or (n125,n122,n116);
nand (n126,n116,n122);
nand (n127,n120,n128);
nor (n128,n129,n132);
and (n129,n130,n116);
not (n130,n131);
and (n132,n75,n131);
nand (n133,n134,n143);
or (n134,n135,n140);
nor (n135,n136,n139);
and (n136,n137,n56);
not (n137,n138);
and (n139,n138,n55);
nand (n140,n56,n141);
not (n141,n142);
or (n143,n144,n141);
not (n144,n145);
nor (n145,n146,n148);
and (n146,n56,n147);
and (n148,n149,n55);
not (n149,n147);
and (n150,n83,n109);
or (n151,n152,n209);
and (n152,n153,n208);
xor (n153,n154,n178);
or (n154,n155,n177);
and (n155,n156,n169);
xor (n156,n157,n162);
and (n157,n158,n77);
nand (n158,n159,n161);
or (n159,n160,n75);
not (n160,n76);
or (n161,n116,n76);
nand (n162,n163,n168);
or (n163,n164,n52);
not (n164,n165);
nor (n165,n166,n167);
and (n166,n36,n28);
and (n167,n29,n34);
nand (n168,n64,n49);
nand (n169,n170,n175);
or (n170,n171,n85);
not (n171,n172);
nor (n172,n173,n174);
and (n173,n91,n131);
and (n174,n130,n90);
nand (n175,n176,n94);
not (n176,n97);
and (n177,n157,n162);
or (n178,n179,n207);
and (n179,n180,n196);
xor (n180,n181,n190);
nand (n181,n182,n189);
or (n182,n183,n118);
not (n183,n184);
nor (n184,n185,n187);
and (n185,n75,n186);
and (n187,n188,n116);
not (n188,n186);
nand (n189,n120,n112);
nand (n190,n191,n195);
or (n191,n192,n140);
nor (n192,n193,n194);
and (n193,n55,n68);
and (n194,n56,n67);
or (n195,n135,n141);
nand (n196,n197,n201);
or (n197,n198,n18);
nor (n198,n199,n200);
and (n199,n33,n106);
and (n200,n24,n108);
or (n201,n202,n38);
nor (n202,n203,n205);
and (n203,n33,n204);
and (n205,n24,n206);
not (n206,n204);
and (n207,n181,n190);
xor (n208,n82,n133);
and (n209,n154,n178);
xor (n210,n211,n268);
xor (n211,n212,n247);
xor (n212,n213,n231);
xor (n213,n214,n221);
nand (n214,n215,n217);
or (n215,n216,n118);
not (n216,n128);
nand (n217,n120,n218);
nor (n218,n219,n220);
and (n219,n101,n116);
and (n220,n75,n99);
nand (n221,n222,n229);
or (n222,n141,n223);
not (n223,n224);
nor (n224,n225,n228);
and (n225,n226,n55);
not (n226,n227);
and (n228,n56,n227);
nand (n229,n145,n230);
not (n230,n140);
nand (n231,n232,n243);
or (n232,n233,n238);
not (n233,n234);
nor (n234,n235,n237);
and (n235,n188,n236);
not (n236,n79);
and (n237,n79,n186);
not (n238,n239);
nor (n239,n158,n240);
nor (n240,n241,n242);
and (n241,n236,n76);
and (n242,n79,n160);
nand (n243,n158,n244);
nor (n244,n245,n246);
and (n245,n114,n236);
and (n246,n79,n115);
xor (n247,n248,n261);
xor (n248,n249,n254);
and (n249,n250,n77);
nand (n250,n251,n253);
or (n251,n236,n252);
nand (n253,n236,n252);
nand (n254,n255,n257);
or (n255,n256,n52);
not (n256,n65);
nand (n257,n64,n258);
nand (n258,n259,n260);
or (n259,n137,n29);
nand (n260,n29,n137);
nand (n261,n262,n267);
or (n262,n263,n103);
not (n263,n264);
nand (n264,n265,n266);
or (n265,n206,n91);
or (n266,n90,n204);
or (n267,n85,n104);
or (n268,n269,n283);
and (n269,n270,n282);
xor (n270,n271,n279);
nand (n271,n272,n277);
or (n272,n238,n273);
nor (n273,n274,n275);
and (n274,n77,n236);
and (n275,n276,n79);
not (n276,n77);
or (n277,n278,n233);
not (n278,n158);
nand (n279,n280,n281);
or (n280,n18,n202);
or (n281,n38,n31);
xnor (n282,n71,n46);
and (n283,n271,n279);
or (n284,n285,n332);
and (n285,n286,n289);
xor (n286,n287,n288);
xor (n287,n270,n282);
xor (n288,n153,n208);
or (n289,n290,n331);
and (n290,n291,n330);
xor (n291,n292,n306);
and (n292,n293,n299);
and (n293,n294,n75);
nand (n294,n295,n296);
or (n295,n91,n122);
nand (n296,n297,n276);
or (n297,n298,n90);
not (n298,n122);
nand (n299,n300,n305);
or (n300,n301,n52);
not (n301,n302);
nand (n302,n303,n304);
or (n303,n29,n206);
or (n304,n28,n204);
nand (n305,n64,n165);
or (n306,n307,n329);
and (n307,n308,n323);
xor (n308,n309,n316);
nand (n309,n310,n315);
or (n310,n311,n85);
not (n311,n312);
nor (n312,n313,n314);
and (n313,n114,n90);
and (n314,n91,n115);
nand (n315,n94,n172);
nand (n316,n317,n322);
or (n317,n318,n118);
not (n318,n319);
nand (n319,n320,n321);
or (n320,n75,n276);
or (n321,n116,n77);
nand (n322,n120,n184);
nand (n323,n324,n328);
or (n324,n140,n325);
nor (n325,n326,n327);
and (n326,n55,n43);
and (n327,n56,n42);
or (n328,n192,n141);
and (n329,n309,n316);
xor (n330,n156,n169);
and (n331,n292,n306);
and (n332,n287,n288);
nand (n333,n12,n284);
not (n334,n335);
nand (n335,n336,n481,n622);
nand (n336,n337,n474);
nand (n337,n338,n473);
or (n338,n339,n460);
not (n339,n340);
nand (n340,n341,n459);
or (n341,n342,n433);
nor (n342,n343,n403);
xor (n343,n344,n383);
xor (n344,n345,n346);
xor (n345,n308,n323);
or (n346,n347,n382);
and (n347,n348,n365);
xor (n348,n349,n356);
nand (n349,n350,n355);
or (n350,n351,n52);
not (n351,n352);
nand (n352,n353,n354);
or (n353,n29,n108);
or (n354,n28,n106);
nand (n355,n64,n302);
nand (n356,n357,n361);
or (n357,n18,n358);
nor (n358,n359,n360);
and (n359,n33,n131);
and (n360,n24,n130);
or (n361,n362,n38);
nor (n362,n363,n364);
and (n363,n33,n99);
and (n364,n24,n101);
and (n365,n366,n371);
nor (n366,n367,n90);
nor (n367,n368,n370);
and (n368,n369,n276);
nand (n369,n24,n89);
and (n370,n33,n93);
nand (n371,n372,n377);
or (n372,n140,n373);
not (n373,n374);
nor (n374,n375,n376);
and (n375,n206,n55);
and (n376,n56,n204);
or (n377,n378,n141);
not (n378,n379);
nor (n379,n380,n381);
and (n380,n36,n55);
and (n381,n56,n34);
and (n382,n349,n356);
xor (n383,n384,n389);
xor (n384,n385,n388);
nand (n385,n386,n387);
or (n386,n18,n362);
or (n387,n38,n198);
xor (n388,n293,n299);
or (n389,n390,n402);
and (n390,n391,n396);
xor (n391,n392,n393);
and (n392,n120,n77);
nand (n393,n394,n395);
or (n394,n140,n378);
or (n395,n325,n141);
nand (n396,n397,n398);
or (n397,n311,n103);
or (n398,n85,n399);
nor (n399,n400,n401);
and (n400,n186,n90);
and (n401,n188,n91);
and (n402,n392,n393);
or (n403,n404,n432);
and (n404,n405,n431);
xor (n405,n406,n430);
or (n406,n407,n429);
and (n407,n408,n423);
xor (n408,n409,n417);
nand (n409,n410,n415);
or (n410,n411,n85);
not (n411,n412);
nand (n412,n413,n414);
or (n413,n91,n276);
or (n414,n90,n77);
nand (n415,n416,n94);
not (n416,n399);
nand (n417,n418,n422);
or (n418,n419,n52);
nor (n419,n420,n421);
and (n420,n101,n29);
and (n421,n99,n28);
nand (n422,n64,n352);
nand (n423,n424,n428);
or (n424,n18,n425);
nor (n425,n426,n427);
and (n426,n33,n115);
and (n427,n24,n114);
or (n428,n358,n38);
and (n429,n409,n417);
xor (n430,n391,n396);
xor (n431,n348,n365);
and (n432,n406,n430);
nand (n433,n434,n435);
xor (n434,n405,n431);
or (n435,n436,n458);
and (n436,n437,n457);
xor (n437,n438,n439);
xor (n438,n366,n371);
or (n439,n440,n456);
and (n440,n441,n450);
xor (n441,n442,n443);
and (n442,n94,n77);
nand (n443,n444,n445);
or (n444,n141,n373);
or (n445,n446,n140);
not (n446,n447);
nand (n447,n448,n449);
or (n448,n108,n56);
nand (n449,n56,n108);
nand (n450,n451,n455);
or (n451,n52,n452);
nor (n452,n453,n454);
and (n453,n28,n131);
and (n454,n29,n130);
or (n455,n53,n419);
and (n456,n442,n443);
xor (n457,n408,n423);
and (n458,n438,n439);
nand (n459,n343,n403);
not (n460,n461);
not (n461,n462);
nor (n462,n463,n470);
xor (n463,n464,n469);
xor (n464,n465,n466);
xor (n465,n180,n196);
or (n466,n467,n468);
and (n467,n384,n389);
and (n468,n385,n388);
xor (n469,n291,n330);
or (n470,n471,n472);
and (n471,n344,n383);
and (n472,n345,n346);
nand (n473,n463,n470);
nand (n474,n475,n477);
not (n475,n476);
xor (n476,n286,n289);
not (n477,n478);
or (n478,n479,n480);
and (n479,n464,n469);
and (n480,n465,n466);
nand (n481,n474,n482,n486);
nor (n482,n462,n483);
nand (n483,n484,n485);
not (n484,n342);
or (n485,n434,n435);
or (n486,n487,n621);
and (n487,n488,n514);
xor (n488,n489,n513);
or (n489,n490,n512);
and (n490,n491,n511);
xor (n491,n492,n498);
nand (n492,n493,n497);
or (n493,n18,n494);
nor (n494,n495,n496);
and (n495,n33,n186);
and (n496,n24,n188);
or (n497,n425,n38);
and (n498,n499,n504);
and (n499,n500,n24);
nand (n500,n501,n502);
or (n501,n29,n23);
nand (n502,n503,n276);
or (n503,n22,n28);
nand (n504,n505,n510);
or (n505,n140,n506);
not (n506,n507);
nor (n507,n508,n509);
and (n508,n101,n55);
and (n509,n56,n99);
nand (n510,n447,n142);
xor (n511,n441,n450);
and (n512,n492,n498);
xor (n513,n437,n457);
or (n514,n515,n620);
and (n515,n516,n539);
xor (n516,n517,n538);
or (n517,n518,n537);
and (n518,n519,n536);
xor (n519,n520,n528);
nand (n520,n521,n526);
or (n521,n522,n52);
not (n522,n523);
nor (n523,n524,n525);
and (n524,n114,n28);
and (n525,n29,n115);
nand (n526,n527,n64);
not (n527,n452);
nand (n528,n529,n534);
or (n529,n530,n18);
not (n530,n531);
nand (n531,n532,n533);
or (n532,n24,n276);
or (n533,n33,n77);
nand (n534,n535,n26);
not (n535,n494);
xor (n536,n499,n504);
and (n537,n520,n528);
xor (n538,n491,n511);
nand (n539,n540,n619);
or (n540,n541,n614);
nor (n541,n542,n613);
and (n542,n543,n575);
nand (n543,n544,n562);
not (n544,n545);
xor (n545,n546,n555);
xor (n546,n547,n548);
and (n547,n26,n77);
nand (n548,n549,n554);
or (n549,n550,n52);
not (n550,n551);
nor (n551,n552,n553);
and (n552,n29,n186);
and (n553,n188,n28);
nand (n554,n64,n523);
nand (n555,n556,n557);
or (n556,n141,n506);
or (n557,n140,n558);
not (n558,n559);
nor (n559,n560,n561);
and (n560,n130,n55);
and (n561,n56,n131);
nand (n562,n563,n569);
nand (n563,n564,n565);
or (n564,n141,n558);
nand (n565,n566,n230);
nand (n566,n567,n568);
or (n567,n115,n55);
nand (n568,n55,n115);
not (n569,n570);
nand (n570,n571,n29);
nand (n571,n572,n574);
or (n572,n573,n77);
nor (n573,n55,n59);
or (n574,n56,n57);
or (n575,n576,n612);
and (n576,n577,n589);
xor (n577,n578,n585);
nand (n578,n579,n584);
or (n579,n580,n52);
not (n580,n581);
nand (n581,n582,n583);
or (n582,n29,n276);
or (n583,n28,n77);
nand (n584,n64,n551);
nand (n585,n586,n588);
or (n586,n569,n587);
not (n587,n563);
nand (n588,n587,n569);
or (n589,n590,n611);
and (n590,n591,n601);
xor (n591,n592,n593);
nor (n592,n53,n276);
nand (n593,n594,n599);
or (n594,n140,n595);
not (n595,n596);
nand (n596,n597,n598);
or (n597,n186,n55);
nand (n598,n55,n186);
or (n599,n600,n141);
not (n600,n566);
nor (n601,n602,n609);
nor (n602,n603,n608);
and (n603,n604,n230);
not (n604,n605);
nor (n605,n606,n607);
and (n606,n55,n77);
and (n607,n56,n276);
and (n608,n596,n142);
or (n609,n610,n55);
nor (n610,n276,n141);
and (n611,n592,n593);
and (n612,n578,n585);
nor (n613,n544,n562);
nor (n614,n615,n616);
xor (n615,n519,n536);
or (n616,n617,n618);
and (n617,n546,n555);
and (n618,n547,n548);
nand (n619,n615,n616);
and (n620,n517,n538);
and (n621,n489,n513);
nand (n622,n476,n478);
or (n623,n335,n10);
not (n624,n625);
nand (n625,n626,n3);
not (n626,n4);
wire s0n627,s1n627,notn627;
or (n627,s0n627,s1n627);
not(notn627,n4);
and (s0n627,notn627,n628);
and (s1n627,n4,1'b0);
wire s0n628,s1n628,notn628;
or (n628,s0n628,s1n628);
not(notn628,n3);
and (s0n628,notn628,n5);
and (s1n628,n3,n629);
xor (n629,n630,n1011);
xor (n630,n631,n1008);
xor (n631,n632,n146);
xor (n632,n633,n999);
xor (n633,n634,n998);
xor (n634,n635,n983);
xor (n635,n636,n69);
xor (n636,n637,n963);
xor (n637,n638,n962);
xor (n638,n639,n937);
xor (n639,n640,n936);
xor (n640,n641,n904);
xor (n641,n642,n903);
xor (n642,n643,n864);
xor (n643,n644,n863);
xor (n644,n645,n819);
xor (n645,n646,n818);
xor (n646,n647,n769);
xor (n647,n648,n132);
xor (n648,n649,n715);
xor (n649,n650,n714);
xor (n650,n651,n653);
xor (n651,n652,n237);
and (n652,n252,n77);
or (n653,n654,n657);
and (n654,n655,n656);
and (n655,n79,n77);
and (n656,n76,n186);
and (n657,n658,n659);
xor (n658,n655,n656);
or (n659,n660,n662);
and (n660,n661,n185);
and (n661,n76,n77);
and (n662,n663,n664);
xor (n663,n661,n185);
or (n664,n665,n668);
and (n665,n666,n667);
and (n666,n75,n77);
and (n667,n122,n186);
and (n668,n669,n670);
xor (n669,n666,n667);
or (n670,n671,n674);
and (n671,n672,n673);
and (n672,n122,n77);
and (n673,n91,n186);
and (n674,n675,n676);
xor (n675,n672,n673);
or (n676,n677,n680);
and (n677,n678,n679);
and (n678,n91,n77);
and (n679,n89,n186);
and (n680,n681,n682);
xor (n681,n678,n679);
or (n682,n683,n686);
and (n683,n684,n685);
and (n684,n89,n77);
and (n685,n24,n186);
and (n686,n687,n688);
xor (n687,n684,n685);
or (n688,n689,n692);
and (n689,n690,n691);
and (n690,n24,n77);
and (n691,n23,n186);
and (n692,n693,n694);
xor (n693,n690,n691);
or (n694,n695,n697);
and (n695,n696,n552);
and (n696,n23,n77);
and (n697,n698,n699);
xor (n698,n696,n552);
or (n699,n700,n703);
and (n700,n701,n702);
and (n701,n29,n77);
and (n702,n57,n186);
and (n703,n704,n705);
xor (n704,n701,n702);
or (n705,n706,n709);
and (n706,n707,n708);
and (n707,n57,n77);
and (n708,n56,n186);
and (n709,n710,n711);
xor (n710,n707,n708);
and (n711,n712,n713);
and (n712,n56,n77);
and (n713,n142,n186);
and (n714,n76,n115);
or (n715,n716,n718);
and (n716,n717,n117);
xor (n717,n658,n659);
and (n718,n719,n720);
xor (n719,n717,n117);
or (n720,n721,n724);
and (n721,n722,n723);
xor (n722,n663,n664);
and (n723,n122,n115);
and (n724,n725,n726);
xor (n725,n722,n723);
or (n726,n727,n729);
and (n727,n728,n314);
xor (n728,n669,n670);
and (n729,n730,n731);
xor (n730,n728,n314);
or (n731,n732,n735);
and (n732,n733,n734);
xor (n733,n675,n676);
and (n734,n89,n115);
and (n735,n736,n737);
xor (n736,n733,n734);
or (n737,n738,n741);
and (n738,n739,n740);
xor (n739,n681,n682);
and (n740,n24,n115);
and (n741,n742,n743);
xor (n742,n739,n740);
or (n743,n744,n747);
and (n744,n745,n746);
xor (n745,n687,n688);
and (n746,n23,n115);
and (n747,n748,n749);
xor (n748,n745,n746);
or (n749,n750,n752);
and (n750,n751,n525);
xor (n751,n693,n694);
and (n752,n753,n754);
xor (n753,n751,n525);
or (n754,n755,n758);
and (n755,n756,n757);
xor (n756,n698,n699);
and (n757,n57,n115);
and (n758,n759,n760);
xor (n759,n756,n757);
or (n760,n761,n764);
and (n761,n762,n763);
xor (n762,n704,n705);
and (n763,n56,n115);
and (n764,n765,n766);
xor (n765,n762,n763);
and (n766,n767,n768);
xor (n767,n710,n711);
and (n768,n142,n115);
or (n769,n770,n773);
and (n770,n771,n772);
xor (n771,n719,n720);
and (n772,n122,n131);
and (n773,n774,n775);
xor (n774,n771,n772);
or (n775,n776,n778);
and (n776,n777,n173);
xor (n777,n725,n726);
and (n778,n779,n780);
xor (n779,n777,n173);
or (n780,n781,n784);
and (n781,n782,n783);
xor (n782,n730,n731);
and (n783,n89,n131);
and (n784,n785,n786);
xor (n785,n782,n783);
or (n786,n787,n790);
and (n787,n788,n789);
xor (n788,n736,n737);
and (n789,n24,n131);
and (n790,n791,n792);
xor (n791,n788,n789);
or (n792,n793,n796);
and (n793,n794,n795);
xor (n794,n742,n743);
and (n795,n23,n131);
and (n796,n797,n798);
xor (n797,n794,n795);
or (n798,n799,n802);
and (n799,n800,n801);
xor (n800,n748,n749);
and (n801,n29,n131);
and (n802,n803,n804);
xor (n803,n800,n801);
or (n804,n805,n808);
and (n805,n806,n807);
xor (n806,n753,n754);
and (n807,n57,n131);
and (n808,n809,n810);
xor (n809,n806,n807);
or (n810,n811,n813);
and (n811,n812,n561);
xor (n812,n759,n760);
and (n813,n814,n815);
xor (n814,n812,n561);
and (n815,n816,n817);
xor (n816,n765,n766);
and (n817,n142,n131);
and (n818,n122,n99);
or (n819,n820,n823);
and (n820,n821,n822);
xor (n821,n774,n775);
and (n822,n91,n99);
and (n823,n824,n825);
xor (n824,n821,n822);
or (n825,n826,n829);
and (n826,n827,n828);
xor (n827,n779,n780);
and (n828,n89,n99);
and (n829,n830,n831);
xor (n830,n827,n828);
or (n831,n832,n835);
and (n832,n833,n834);
xor (n833,n785,n786);
and (n834,n24,n99);
and (n835,n836,n837);
xor (n836,n833,n834);
or (n837,n838,n841);
and (n838,n839,n840);
xor (n839,n791,n792);
and (n840,n23,n99);
and (n841,n842,n843);
xor (n842,n839,n840);
or (n843,n844,n847);
and (n844,n845,n846);
xor (n845,n797,n798);
and (n846,n29,n99);
and (n847,n848,n849);
xor (n848,n845,n846);
or (n849,n850,n853);
and (n850,n851,n852);
xor (n851,n803,n804);
and (n852,n57,n99);
and (n853,n854,n855);
xor (n854,n851,n852);
or (n855,n856,n858);
and (n856,n857,n509);
xor (n857,n809,n810);
and (n858,n859,n860);
xor (n859,n857,n509);
and (n860,n861,n862);
xor (n861,n814,n815);
and (n862,n142,n99);
and (n863,n91,n106);
or (n864,n865,n868);
and (n865,n866,n867);
xor (n866,n824,n825);
and (n867,n89,n106);
and (n868,n869,n870);
xor (n869,n866,n867);
or (n870,n871,n874);
and (n871,n872,n873);
xor (n872,n830,n831);
and (n873,n24,n106);
and (n874,n875,n876);
xor (n875,n872,n873);
or (n876,n877,n880);
and (n877,n878,n879);
xor (n878,n836,n837);
and (n879,n23,n106);
and (n880,n881,n882);
xor (n881,n878,n879);
or (n882,n883,n886);
and (n883,n884,n885);
xor (n884,n842,n843);
and (n885,n29,n106);
and (n886,n887,n888);
xor (n887,n884,n885);
or (n888,n889,n892);
and (n889,n890,n891);
xor (n890,n848,n849);
and (n891,n57,n106);
and (n892,n893,n894);
xor (n893,n890,n891);
or (n894,n895,n898);
and (n895,n896,n897);
xor (n896,n854,n855);
and (n897,n56,n106);
and (n898,n899,n900);
xor (n899,n896,n897);
and (n900,n901,n902);
xor (n901,n859,n860);
and (n902,n142,n106);
and (n903,n89,n204);
or (n904,n905,n908);
and (n905,n906,n907);
xor (n906,n869,n870);
and (n907,n24,n204);
and (n908,n909,n910);
xor (n909,n906,n907);
or (n910,n911,n914);
and (n911,n912,n913);
xor (n912,n875,n876);
and (n913,n23,n204);
and (n914,n915,n916);
xor (n915,n912,n913);
or (n916,n917,n920);
and (n917,n918,n919);
xor (n918,n881,n882);
and (n919,n29,n204);
and (n920,n921,n922);
xor (n921,n918,n919);
or (n922,n923,n926);
and (n923,n924,n925);
xor (n924,n887,n888);
and (n925,n57,n204);
and (n926,n927,n928);
xor (n927,n924,n925);
or (n928,n929,n931);
and (n929,n930,n376);
xor (n930,n893,n894);
and (n931,n932,n933);
xor (n932,n930,n376);
and (n933,n934,n935);
xor (n934,n899,n900);
and (n935,n142,n204);
and (n936,n24,n34);
or (n937,n938,n941);
and (n938,n939,n940);
xor (n939,n909,n910);
and (n940,n23,n34);
and (n941,n942,n943);
xor (n942,n939,n940);
or (n943,n944,n946);
and (n944,n945,n167);
xor (n945,n915,n916);
and (n946,n947,n948);
xor (n947,n945,n167);
or (n948,n949,n952);
and (n949,n950,n951);
xor (n950,n921,n922);
and (n951,n57,n34);
and (n952,n953,n954);
xor (n953,n950,n951);
or (n954,n955,n957);
and (n955,n956,n381);
xor (n956,n927,n928);
and (n957,n958,n959);
xor (n958,n956,n381);
and (n959,n960,n961);
xor (n960,n932,n933);
and (n961,n142,n34);
and (n962,n23,n43);
or (n963,n964,n966);
and (n964,n965,n51);
xor (n965,n942,n943);
and (n966,n967,n968);
xor (n967,n965,n51);
or (n968,n969,n972);
and (n969,n970,n971);
xor (n970,n947,n948);
and (n971,n57,n43);
and (n972,n973,n974);
xor (n973,n970,n971);
or (n974,n975,n978);
and (n975,n976,n977);
xor (n976,n953,n954);
and (n977,n56,n43);
and (n978,n979,n980);
xor (n979,n976,n977);
and (n980,n981,n982);
xor (n981,n958,n959);
and (n982,n142,n43);
or (n983,n984,n987);
and (n984,n985,n986);
xor (n985,n967,n968);
and (n986,n57,n68);
and (n987,n988,n989);
xor (n988,n985,n986);
or (n989,n990,n993);
and (n990,n991,n992);
xor (n991,n973,n974);
and (n992,n56,n68);
and (n993,n994,n995);
xor (n994,n991,n992);
and (n995,n996,n997);
xor (n996,n979,n980);
and (n997,n142,n68);
and (n998,n57,n138);
or (n999,n1000,n1003);
and (n1000,n1001,n1002);
xor (n1001,n988,n989);
and (n1002,n56,n138);
and (n1003,n1004,n1005);
xor (n1004,n1001,n1002);
and (n1005,n1006,n1007);
xor (n1006,n994,n995);
and (n1007,n142,n138);
and (n1008,n1009,n1010);
xor (n1009,n1004,n1005);
and (n1010,n142,n147);
and (n1011,n142,n227);
endmodule
