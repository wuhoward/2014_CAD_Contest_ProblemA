module top (out,n17,n18,n24,n30,n36,n43,n45,n53,n54
        ,n63,n68,n72,n77,n86,n88,n95,n96,n105,n112
        ,n114,n121,n131,n139,n149,n155,n166,n168,n175,n184
        ,n193,n199,n205,n212,n217);
output out;
input n17;
input n18;
input n24;
input n30;
input n36;
input n43;
input n45;
input n53;
input n54;
input n63;
input n68;
input n72;
input n77;
input n86;
input n88;
input n95;
input n96;
input n105;
input n112;
input n114;
input n121;
input n131;
input n139;
input n149;
input n155;
input n166;
input n168;
input n175;
input n184;
input n193;
input n199;
input n205;
input n212;
input n217;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n25;
wire n26;
wire n27;
wire n28;
wire n29;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n37;
wire n38;
wire n39;
wire n40;
wire n41;
wire n42;
wire n44;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n64;
wire n65;
wire n66;
wire n67;
wire n69;
wire n70;
wire n71;
wire n73;
wire n74;
wire n75;
wire n76;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n87;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n113;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n167;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n213;
wire n214;
wire n215;
wire n216;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
xor (out,n0,n1104);
nand (n0,n1,n1103);
or (n1,n2,n521);
not (n2,n3);
nor (n3,n4,n520);
not (n4,n5);
nand (n5,n6,n428);
xor (n6,n7,n374);
xor (n7,n8,n221);
xor (n8,n9,n158);
xor (n9,n10,n78);
xor (n10,n11,n65);
xor (n11,n12,n38);
nand (n12,n13,n32);
or (n13,n14,n21);
nor (n14,n15,n19);
and (n15,n16,n18);
not (n16,n17);
and (n19,n17,n20);
not (n20,n18);
nand (n21,n22,n26);
nand (n22,n23,n25);
or (n23,n24,n20);
nand (n25,n20,n24);
not (n26,n27);
nand (n27,n28,n31);
or (n28,n29,n24);
not (n29,n30);
nand (n31,n24,n29);
nand (n32,n33,n27);
nor (n33,n34,n37);
and (n34,n35,n20);
not (n35,n36);
and (n37,n36,n18);
nand (n38,n39,n59);
or (n39,n40,n48);
not (n40,n41);
nand (n41,n42,n46);
or (n42,n43,n44);
not (n44,n45);
or (n46,n47,n45);
not (n47,n43);
nand (n48,n49,n56);
not (n49,n50);
nand (n50,n51,n55);
or (n51,n52,n54);
not (n52,n53);
nand (n55,n52,n54);
nand (n56,n57,n58);
or (n57,n54,n47);
nand (n58,n47,n54);
nand (n59,n50,n60);
nor (n60,n61,n64);
and (n61,n62,n47);
not (n62,n63);
and (n64,n63,n43);
nand (n65,n66,n76);
or (n66,n67,n69);
not (n67,n68);
not (n69,n70);
nor (n70,n71,n73);
not (n71,n72);
nand (n73,n74,n75);
or (n74,n47,n72);
nand (n75,n72,n47);
nand (n76,n73,n77);
xor (n78,n79,n133);
xor (n79,n80,n107);
nand (n80,n81,n101);
or (n81,n82,n90);
not (n82,n83);
nor (n83,n84,n89);
and (n84,n85,n87);
not (n85,n86);
not (n87,n88);
and (n89,n86,n88);
nand (n90,n91,n98);
not (n91,n92);
nand (n92,n93,n97);
or (n93,n94,n96);
not (n94,n95);
nand (n97,n94,n96);
nand (n98,n99,n100);
or (n99,n88,n94);
nand (n100,n94,n88);
nand (n101,n92,n102);
or (n102,n103,n106);
and (n103,n104,n88);
not (n104,n105);
and (n106,n105,n87);
nand (n107,n108,n127);
or (n108,n109,n117);
not (n109,n110);
nand (n110,n111,n115);
or (n111,n112,n113);
not (n113,n114);
or (n115,n116,n114);
not (n116,n112);
not (n117,n118);
nor (n118,n119,n124);
nor (n119,n120,n122);
and (n120,n121,n116);
and (n122,n112,n123);
not (n123,n121);
nand (n124,n125,n126);
or (n125,n20,n121);
nand (n126,n121,n20);
nand (n127,n124,n128);
nor (n128,n129,n132);
and (n129,n130,n116);
not (n130,n131);
and (n132,n131,n112);
nand (n133,n134,n151);
or (n134,n135,n145);
not (n135,n136);
nor (n136,n137,n141);
nand (n137,n138,n140);
or (n138,n87,n139);
nand (n140,n139,n87);
nor (n141,n142,n144);
and (n142,n143,n30);
not (n143,n139);
and (n144,n139,n29);
not (n145,n146);
nor (n146,n147,n150);
and (n147,n29,n148);
not (n148,n149);
and (n150,n149,n30);
or (n151,n152,n157);
nor (n152,n153,n156);
and (n153,n154,n30);
not (n154,n155);
and (n156,n155,n29);
not (n157,n137);
xor (n158,n159,n208);
xor (n159,n160,n187);
nand (n160,n161,n180);
or (n161,n162,n170);
not (n162,n163);
nor (n163,n164,n169);
and (n164,n165,n167);
not (n165,n166);
not (n167,n168);
and (n169,n166,n168);
nand (n170,n171,n177);
not (n171,n172);
nand (n172,n173,n176);
or (n173,n174,n112);
not (n174,n175);
nand (n176,n112,n174);
nand (n177,n178,n179);
nand (n178,n174,n168);
nand (n179,n175,n167);
nand (n180,n181,n172);
not (n181,n182);
nor (n182,n183,n185);
and (n183,n167,n184);
and (n185,n168,n186);
not (n186,n184);
nand (n187,n188,n202);
or (n188,n189,n195);
not (n189,n190);
nand (n190,n191,n194);
or (n191,n53,n192);
not (n192,n193);
or (n194,n52,n193);
nand (n195,n196,n201);
nor (n196,n197,n200);
and (n197,n198,n168);
not (n198,n199);
and (n200,n199,n167);
xor (n201,n198,n52);
or (n202,n196,n203);
nor (n203,n204,n206);
and (n204,n52,n205);
and (n206,n53,n207);
not (n207,n205);
nand (n208,n209,n220);
or (n209,n210,n213);
nand (n210,n211,n96);
not (n211,n212);
not (n213,n214);
nor (n214,n215,n219);
and (n215,n216,n218);
not (n216,n217);
not (n218,n96);
and (n219,n217,n96);
or (n220,n218,n211);
or (n221,n222,n373);
and (n222,n223,n344);
xor (n223,n224,n277);
or (n224,n225,n276);
and (n225,n226,n252);
xor (n226,n227,n236);
nand (n227,n228,n232);
or (n228,n195,n229);
nor (n229,n230,n231);
and (n230,n52,n45);
and (n231,n53,n44);
or (n232,n196,n233);
nor (n233,n234,n235);
and (n234,n63,n52);
and (n235,n53,n62);
xor (n236,n237,n243);
nor (n237,n238,n47);
nor (n238,n239,n241);
and (n239,n240,n52);
nand (n240,n68,n54);
and (n241,n67,n242);
not (n242,n54);
nand (n243,n244,n248);
or (n244,n245,n210);
nor (n245,n246,n247);
and (n246,n85,n96);
and (n247,n86,n218);
or (n248,n249,n211);
nor (n249,n250,n251);
and (n250,n218,n105);
and (n251,n96,n104);
or (n252,n253,n275);
and (n253,n254,n264);
xor (n254,n255,n256);
nor (n255,n49,n67);
nand (n256,n257,n262);
or (n257,n210,n258);
not (n258,n259);
nor (n259,n260,n261);
and (n260,n154,n218);
and (n261,n155,n96);
nand (n262,n263,n212);
not (n263,n245);
nand (n264,n265,n270);
or (n265,n90,n266);
not (n266,n267);
nand (n267,n268,n269);
or (n268,n88,n35);
or (n269,n87,n36);
or (n270,n91,n271);
not (n271,n272);
nand (n272,n273,n274);
or (n273,n88,n148);
or (n274,n87,n149);
and (n275,n255,n256);
and (n276,n227,n236);
xor (n277,n278,n311);
xor (n278,n279,n280);
and (n279,n237,n243);
or (n280,n281,n310);
and (n281,n282,n300);
xor (n282,n283,n289);
nand (n283,n284,n285);
or (n284,n271,n90);
nand (n285,n92,n286);
nor (n286,n287,n288);
and (n287,n154,n87);
and (n288,n155,n88);
nand (n289,n290,n295);
or (n290,n291,n48);
not (n291,n292);
nand (n292,n293,n294);
or (n293,n47,n68);
or (n294,n43,n67);
nand (n295,n296,n50);
nand (n296,n297,n299);
or (n297,n43,n298);
not (n298,n77);
or (n299,n47,n77);
nand (n300,n301,n306);
or (n301,n21,n302);
not (n302,n303);
nor (n303,n304,n305);
and (n304,n113,n20);
and (n305,n114,n18);
or (n306,n26,n307);
nor (n307,n308,n309);
and (n308,n130,n18);
and (n309,n131,n20);
and (n310,n283,n289);
or (n311,n312,n343);
and (n312,n313,n334);
xor (n313,n314,n325);
nand (n314,n315,n320);
or (n315,n316,n117);
not (n316,n317);
nor (n317,n318,n319);
and (n318,n165,n116);
and (n319,n166,n112);
or (n320,n321,n324);
nor (n321,n322,n323);
and (n322,n186,n112);
and (n323,n184,n116);
not (n324,n124);
nand (n325,n326,n330);
or (n326,n327,n135);
nor (n327,n328,n329);
and (n328,n29,n17);
and (n329,n30,n16);
nand (n330,n137,n331);
nand (n331,n332,n333);
or (n332,n30,n35);
or (n333,n29,n36);
nand (n334,n335,n339);
or (n335,n170,n336);
nor (n336,n337,n338);
and (n337,n167,n193);
and (n338,n168,n192);
or (n339,n171,n340);
nor (n340,n341,n342);
and (n341,n207,n168);
and (n342,n205,n167);
and (n343,n314,n325);
or (n344,n345,n372);
and (n345,n346,n371);
xor (n346,n347,n370);
or (n347,n348,n369);
and (n348,n349,n363);
xor (n349,n350,n357);
nand (n350,n351,n356);
or (n351,n352,n21);
not (n352,n353);
nand (n353,n354,n355);
or (n354,n18,n186);
or (n355,n20,n184);
nand (n356,n27,n303);
nand (n357,n358,n362);
or (n358,n117,n359);
nor (n359,n360,n361);
and (n360,n116,n205);
and (n361,n112,n207);
nand (n362,n124,n317);
nand (n363,n364,n368);
or (n364,n135,n365);
nor (n365,n366,n367);
and (n366,n29,n131);
and (n367,n30,n130);
or (n368,n327,n157);
and (n369,n350,n357);
xor (n370,n313,n334);
xor (n371,n282,n300);
and (n372,n347,n370);
and (n373,n224,n277);
xor (n374,n375,n421);
xor (n375,n376,n379);
or (n376,n377,n378);
and (n377,n278,n311);
and (n378,n279,n280);
xor (n379,n380,n407);
xor (n380,n381,n393);
or (n381,n382,n392);
and (n382,n383,n388);
xor (n383,n384,n385);
and (n384,n73,n68);
nand (n385,n386,n387);
or (n386,n211,n213);
or (n387,n249,n210);
nand (n388,n389,n391);
or (n389,n90,n390);
not (n390,n286);
nand (n391,n92,n83);
and (n392,n384,n385);
or (n393,n394,n406);
and (n394,n395,n403);
xor (n395,n396,n400);
nand (n396,n397,n399);
or (n397,n398,n135);
not (n398,n331);
nand (n399,n146,n137);
nand (n400,n401,n402);
or (n401,n340,n170);
nand (n402,n163,n172);
nand (n403,n404,n405);
or (n404,n189,n196);
or (n405,n195,n233);
and (n406,n396,n400);
or (n407,n408,n420);
and (n408,n409,n417);
xor (n409,n410,n414);
nand (n410,n411,n413);
or (n411,n412,n48);
not (n412,n296);
nand (n413,n41,n50);
nand (n414,n415,n416);
or (n415,n21,n307);
or (n416,n26,n14);
nand (n417,n418,n419);
or (n418,n117,n321);
or (n419,n324,n109);
and (n420,n410,n414);
or (n421,n422,n427);
and (n422,n423,n426);
xor (n423,n424,n425);
xor (n424,n395,n403);
xor (n425,n383,n388);
xor (n426,n409,n417);
and (n427,n424,n425);
or (n428,n429,n519);
and (n429,n430,n518);
xor (n430,n431,n432);
xor (n431,n423,n426);
or (n432,n433,n517);
and (n433,n434,n465);
xor (n434,n435,n464);
or (n435,n436,n463);
and (n436,n437,n451);
xor (n437,n438,n445);
nand (n438,n439,n443);
or (n439,n440,n170);
nor (n440,n441,n442);
and (n441,n62,n168);
and (n442,n63,n167);
nand (n443,n444,n172);
not (n444,n336);
nand (n445,n446,n450);
or (n446,n447,n195);
nor (n447,n448,n449);
and (n448,n52,n77);
and (n449,n53,n298);
or (n450,n196,n229);
and (n451,n452,n457);
nor (n452,n453,n52);
nor (n453,n454,n456);
and (n454,n455,n167);
nand (n455,n68,n199);
and (n456,n67,n198);
nand (n457,n458,n459);
or (n458,n211,n258);
or (n459,n460,n210);
nor (n460,n461,n462);
and (n461,n148,n96);
and (n462,n149,n218);
and (n463,n438,n445);
xor (n464,n226,n252);
or (n465,n466,n516);
and (n466,n467,n515);
xor (n467,n468,n493);
or (n468,n469,n492);
and (n469,n470,n485);
xor (n470,n471,n478);
nand (n471,n472,n477);
or (n472,n473,n90);
not (n473,n474);
nor (n474,n475,n476);
and (n475,n16,n87);
and (n476,n17,n88);
nand (n477,n267,n92);
nand (n478,n479,n484);
or (n479,n480,n21);
not (n480,n481);
nand (n481,n482,n483);
or (n482,n18,n165);
or (n483,n20,n166);
nand (n484,n27,n353);
nand (n485,n486,n491);
or (n486,n117,n487);
not (n487,n488);
nand (n488,n489,n490);
or (n489,n112,n192);
or (n490,n116,n193);
or (n491,n324,n359);
and (n492,n471,n478);
or (n493,n494,n514);
and (n494,n495,n508);
xor (n495,n496,n502);
nand (n496,n497,n501);
or (n497,n135,n498);
nor (n498,n499,n500);
and (n499,n29,n114);
and (n500,n30,n113);
or (n501,n365,n157);
nand (n502,n503,n507);
or (n503,n170,n504);
nor (n504,n505,n506);
and (n505,n167,n45);
and (n506,n168,n44);
or (n507,n440,n171);
nand (n508,n509,n513);
or (n509,n195,n510);
nor (n510,n511,n512);
and (n511,n67,n53);
and (n512,n68,n52);
or (n513,n447,n196);
and (n514,n496,n502);
xor (n515,n254,n264);
and (n516,n468,n493);
and (n517,n435,n464);
xor (n518,n223,n344);
and (n519,n431,n432);
nor (n520,n6,n428);
not (n521,n522);
nor (n522,n523,n1101);
and (n523,n524,n1095);
nand (n524,n525,n1082);
or (n525,n526,n978);
not (n526,n527);
nand (n527,n528,n967,n977);
nand (n528,n529,n722,n826);
nand (n529,n530,n686);
not (n530,n531);
xor (n531,n532,n645);
xor (n532,n533,n574);
xor (n533,n534,n553);
xor (n534,n535,n544);
nand (n535,n536,n540);
or (n536,n170,n537);
nor (n537,n538,n539);
and (n538,n67,n168);
and (n539,n167,n68);
or (n540,n171,n541);
nor (n541,n542,n543);
and (n542,n167,n77);
and (n543,n168,n298);
nand (n544,n545,n549);
or (n545,n135,n546);
nor (n546,n547,n548);
and (n547,n29,n166);
and (n548,n30,n165);
or (n549,n550,n157);
nor (n550,n551,n552);
and (n551,n29,n184);
and (n552,n30,n186);
nand (n553,n554,n573);
or (n554,n555,n562);
not (n555,n556);
nand (n556,n557,n168);
nand (n557,n558,n559);
or (n558,n68,n175);
nand (n559,n560,n116);
not (n560,n561);
and (n561,n68,n175);
not (n562,n563);
nand (n563,n564,n569);
or (n564,n565,n90);
not (n565,n566);
nand (n566,n567,n568);
or (n567,n88,n113);
or (n568,n87,n114);
nand (n569,n92,n570);
nand (n570,n571,n572);
or (n571,n88,n130);
or (n572,n87,n131);
or (n573,n563,n556);
xor (n574,n575,n625);
xor (n575,n576,n597);
or (n576,n577,n596);
and (n577,n578,n586);
xor (n578,n579,n580);
and (n579,n172,n68);
nand (n580,n581,n585);
or (n581,n582,n90);
nor (n582,n583,n584);
and (n583,n186,n88);
and (n584,n184,n87);
nand (n585,n92,n566);
nand (n586,n587,n592);
or (n587,n21,n588);
not (n588,n589);
nor (n589,n590,n591);
and (n590,n62,n20);
and (n591,n63,n18);
or (n592,n26,n593);
nor (n593,n594,n595);
and (n594,n193,n20);
and (n595,n192,n18);
and (n596,n579,n580);
or (n597,n598,n624);
and (n598,n599,n618);
xor (n599,n600,n609);
nand (n600,n601,n605);
or (n601,n117,n602);
nor (n602,n603,n604);
and (n603,n298,n112);
and (n604,n77,n116);
or (n605,n324,n606);
nor (n606,n607,n608);
and (n607,n45,n116);
and (n608,n44,n112);
nand (n609,n610,n614);
or (n610,n611,n210);
nor (n611,n612,n613);
and (n612,n218,n131);
and (n613,n96,n130);
or (n614,n615,n211);
nor (n615,n616,n617);
and (n616,n218,n17);
and (n617,n96,n16);
nand (n618,n619,n623);
or (n619,n135,n620);
nor (n620,n621,n622);
and (n621,n29,n205);
and (n622,n30,n207);
or (n623,n546,n157);
and (n624,n600,n609);
xor (n625,n626,n639);
xor (n626,n627,n633);
nand (n627,n628,n629);
or (n628,n21,n593);
or (n629,n630,n26);
nor (n630,n631,n632);
and (n631,n207,n18);
and (n632,n205,n20);
nand (n633,n634,n635);
or (n634,n117,n606);
or (n635,n324,n636);
nor (n636,n637,n638);
and (n637,n62,n112);
and (n638,n63,n116);
nand (n639,n640,n641);
or (n640,n615,n210);
or (n641,n642,n211);
nor (n642,n643,n644);
and (n643,n218,n36);
and (n644,n96,n35);
or (n645,n646,n685);
and (n646,n647,n684);
xor (n647,n648,n661);
and (n648,n649,n655);
and (n649,n650,n112);
nand (n650,n651,n652);
or (n651,n68,n121);
nand (n652,n653,n20);
not (n653,n654);
and (n654,n68,n121);
nand (n655,n656,n660);
or (n656,n90,n657);
nor (n657,n658,n659);
and (n658,n87,n166);
and (n659,n88,n165);
or (n660,n91,n582);
or (n661,n662,n683);
and (n662,n663,n677);
xor (n663,n664,n671);
nand (n664,n665,n670);
or (n665,n666,n21);
not (n666,n667);
nor (n667,n668,n669);
and (n668,n45,n18);
and (n669,n44,n20);
nand (n670,n27,n589);
nand (n671,n672,n676);
or (n672,n117,n673);
nor (n673,n674,n675);
and (n674,n112,n67);
and (n675,n116,n68);
or (n676,n324,n602);
nand (n677,n678,n682);
or (n678,n210,n679);
nor (n679,n680,n681);
and (n680,n218,n114);
and (n681,n96,n113);
or (n682,n611,n211);
and (n683,n664,n671);
xor (n684,n578,n586);
and (n685,n648,n661);
not (n686,n687);
or (n687,n688,n721);
and (n688,n689,n720);
xor (n689,n690,n691);
xor (n690,n599,n618);
or (n691,n692,n719);
and (n692,n693,n701);
xor (n693,n694,n700);
nand (n694,n695,n699);
or (n695,n135,n696);
nor (n696,n697,n698);
and (n697,n29,n193);
and (n698,n30,n192);
or (n699,n620,n157);
xor (n700,n649,n655);
or (n701,n702,n718);
and (n702,n703,n711);
xor (n703,n704,n705);
and (n704,n124,n68);
nand (n705,n706,n710);
or (n706,n707,n210);
nor (n707,n708,n709);
and (n708,n218,n184);
and (n709,n96,n186);
or (n710,n679,n211);
nand (n711,n712,n717);
or (n712,n21,n713);
not (n713,n714);
nand (n714,n715,n716);
or (n715,n18,n298);
or (n716,n20,n77);
or (n717,n26,n666);
and (n718,n704,n705);
and (n719,n694,n700);
xor (n720,n647,n684);
and (n721,n690,n691);
nor (n722,n723,n763);
not (n723,n724);
or (n724,n725,n726);
xor (n725,n689,n720);
or (n726,n727,n762);
and (n727,n728,n761);
xor (n728,n729,n730);
xor (n729,n663,n677);
or (n730,n731,n760);
and (n731,n732,n745);
xor (n732,n733,n739);
nand (n733,n734,n738);
or (n734,n90,n735);
nor (n735,n736,n737);
and (n736,n87,n205);
and (n737,n88,n207);
or (n738,n91,n657);
nand (n739,n740,n744);
or (n740,n135,n741);
nor (n741,n742,n743);
and (n742,n29,n63);
and (n743,n30,n62);
or (n744,n696,n157);
and (n745,n746,n753);
nor (n746,n747,n20);
nor (n747,n748,n751);
and (n748,n749,n29);
not (n749,n750);
and (n750,n68,n24);
and (n751,n67,n752);
not (n752,n24);
nand (n753,n754,n759);
or (n754,n210,n755);
not (n755,n756);
nor (n756,n757,n758);
and (n757,n166,n96);
and (n758,n165,n218);
or (n759,n707,n211);
and (n760,n733,n739);
xor (n761,n693,n701);
and (n762,n729,n730);
nand (n763,n764,n820);
not (n764,n765);
nor (n765,n766,n795);
xor (n766,n767,n794);
xor (n767,n768,n793);
or (n768,n769,n792);
and (n769,n770,n786);
xor (n770,n771,n778);
nand (n771,n772,n777);
or (n772,n773,n21);
not (n773,n774);
nand (n774,n775,n776);
or (n775,n20,n68);
or (n776,n18,n67);
nand (n777,n27,n714);
nand (n778,n779,n784);
or (n779,n780,n90);
not (n780,n781);
nand (n781,n782,n783);
or (n782,n88,n192);
or (n783,n87,n193);
nand (n784,n785,n92);
not (n785,n735);
nand (n786,n787,n791);
or (n787,n135,n788);
nor (n788,n789,n790);
and (n789,n29,n45);
and (n790,n30,n44);
or (n791,n741,n157);
and (n792,n771,n778);
xor (n793,n703,n711);
xor (n794,n732,n745);
or (n795,n796,n819);
and (n796,n797,n818);
xor (n797,n798,n799);
xor (n798,n746,n753);
or (n799,n800,n817);
and (n800,n801,n810);
xor (n801,n802,n803);
and (n802,n27,n68);
nand (n803,n804,n805);
or (n804,n211,n755);
or (n805,n806,n210);
not (n806,n807);
nand (n807,n808,n809);
or (n808,n205,n218);
nand (n809,n218,n205);
nand (n810,n811,n816);
or (n811,n812,n90);
not (n812,n813);
nand (n813,n814,n815);
or (n814,n88,n62);
or (n815,n87,n63);
nand (n816,n92,n781);
and (n817,n802,n803);
xor (n818,n770,n786);
and (n819,n798,n799);
not (n820,n821);
nor (n821,n822,n823);
xor (n822,n728,n761);
or (n823,n824,n825);
and (n824,n767,n794);
and (n825,n768,n793);
or (n826,n827,n966);
and (n827,n828,n855);
xor (n828,n829,n854);
or (n829,n830,n853);
and (n830,n831,n852);
xor (n831,n832,n838);
nand (n832,n833,n837);
or (n833,n135,n834);
nor (n834,n835,n836);
and (n835,n29,n77);
and (n836,n30,n298);
or (n837,n788,n157);
nor (n838,n839,n847);
not (n839,n840);
nand (n840,n841,n846);
or (n841,n210,n842);
not (n842,n843);
nor (n843,n844,n845);
and (n844,n193,n96);
and (n845,n192,n218);
nand (n846,n807,n212);
nand (n847,n848,n30);
nand (n848,n849,n851);
or (n849,n850,n88);
and (n850,n68,n139);
or (n851,n68,n139);
xor (n852,n801,n810);
and (n853,n832,n838);
xor (n854,n797,n818);
or (n855,n856,n965);
and (n856,n857,n881);
xor (n857,n858,n880);
or (n858,n859,n879);
and (n859,n860,n875);
xor (n860,n861,n868);
nand (n861,n862,n867);
or (n862,n863,n90);
not (n863,n864);
nor (n864,n865,n866);
and (n865,n44,n87);
and (n866,n45,n88);
nand (n867,n92,n813);
nand (n868,n869,n874);
or (n869,n870,n135);
not (n870,n871);
nand (n871,n872,n873);
or (n872,n29,n68);
or (n873,n67,n30);
or (n874,n834,n157);
nand (n875,n876,n878);
or (n876,n877,n839);
not (n877,n847);
or (n878,n840,n847);
and (n879,n861,n868);
xor (n880,n831,n852);
or (n881,n882,n964);
and (n882,n883,n904);
xor (n883,n884,n903);
or (n884,n885,n902);
and (n885,n886,n895);
xor (n886,n887,n888);
and (n887,n137,n68);
nand (n888,n889,n894);
or (n889,n890,n90);
not (n890,n891);
nor (n891,n892,n893);
and (n892,n298,n87);
and (n893,n77,n88);
nand (n894,n92,n864);
nand (n895,n896,n897);
or (n896,n211,n842);
or (n897,n210,n898);
not (n898,n899);
nor (n899,n900,n901);
and (n900,n62,n218);
and (n901,n63,n96);
and (n902,n887,n888);
xor (n903,n860,n875);
nand (n904,n905,n963);
or (n905,n906,n922);
nor (n906,n907,n908);
xor (n907,n886,n895);
and (n908,n909,n916);
nand (n909,n910,n911);
nand (n910,n899,n212);
nand (n911,n912,n915);
nor (n912,n913,n914);
and (n913,n44,n218);
and (n914,n45,n96);
not (n915,n210);
not (n916,n917);
nand (n917,n918,n88);
nand (n918,n919,n921);
or (n919,n920,n96);
and (n920,n68,n95);
or (n921,n68,n95);
nor (n922,n923,n962);
and (n923,n924,n936);
nand (n924,n925,n929);
nor (n925,n926,n928);
and (n926,n927,n916);
not (n927,n909);
and (n928,n909,n917);
nor (n929,n930,n931);
and (n930,n92,n891);
and (n931,n932,n933);
not (n932,n90);
nand (n933,n934,n935);
or (n934,n87,n68);
or (n935,n67,n88);
nand (n936,n937,n960);
or (n937,n938,n952);
not (n938,n939);
and (n939,n940,n950);
nand (n940,n941,n946);
or (n941,n211,n942);
not (n942,n943);
nor (n943,n944,n945);
and (n944,n298,n218);
and (n945,n77,n96);
nand (n946,n947,n915);
nand (n947,n948,n949);
or (n948,n218,n68);
or (n949,n96,n67);
nor (n950,n951,n218);
and (n951,n68,n212);
not (n952,n953);
nand (n953,n954,n959);
not (n954,n955);
nand (n955,n956,n958);
or (n956,n211,n957);
not (n957,n912);
nand (n958,n943,n915);
nand (n959,n92,n68);
nand (n960,n961,n955);
not (n961,n959);
nor (n962,n925,n929);
nand (n963,n907,n908);
and (n964,n884,n903);
and (n965,n858,n880);
and (n966,n829,n854);
nand (n967,n968,n529);
or (n968,n969,n971);
not (n969,n970);
nand (n970,n725,n726);
not (n971,n972);
nand (n972,n724,n973);
nand (n973,n974,n976);
or (n974,n821,n975);
nand (n975,n766,n795);
nand (n976,n822,n823);
nand (n977,n531,n687);
not (n978,n979);
nor (n979,n980,n1045);
nor (n980,n981,n1022);
xor (n981,n982,n1021);
xor (n982,n983,n984);
xor (n983,n346,n371);
or (n984,n985,n1020);
and (n985,n986,n989);
xor (n986,n987,n988);
xor (n987,n349,n363);
xor (n988,n437,n451);
or (n989,n990,n1019);
and (n990,n991,n1006);
xor (n991,n992,n993);
xor (n992,n452,n457);
or (n993,n994,n1005);
and (n994,n995,n1002);
xor (n995,n996,n998);
and (n996,n997,n68);
not (n997,n196);
nand (n998,n999,n1001);
or (n999,n1000,n90);
not (n1000,n570);
nand (n1001,n92,n474);
nand (n1002,n1003,n1004);
or (n1003,n480,n26);
or (n1004,n21,n630);
and (n1005,n996,n998);
or (n1006,n1007,n1018);
and (n1007,n1008,n1015);
xor (n1008,n1009,n1012);
nand (n1009,n1010,n1011);
or (n1010,n636,n117);
nand (n1011,n488,n124);
nand (n1012,n1013,n1014);
or (n1013,n642,n210);
or (n1014,n460,n211);
nand (n1015,n1016,n1017);
or (n1016,n541,n170);
or (n1017,n504,n171);
and (n1018,n1009,n1012);
and (n1019,n992,n993);
and (n1020,n987,n988);
xor (n1021,n434,n465);
or (n1022,n1023,n1044);
and (n1023,n1024,n1027);
xor (n1024,n1025,n1026);
xor (n1025,n467,n515);
xor (n1026,n986,n989);
or (n1027,n1028,n1043);
and (n1028,n1029,n1032);
xor (n1029,n1030,n1031);
xor (n1030,n495,n508);
xor (n1031,n470,n485);
or (n1032,n1033,n1042);
and (n1033,n1034,n1039);
xor (n1034,n1035,n1038);
nand (n1035,n1036,n1037);
or (n1036,n135,n550);
or (n1037,n498,n157);
and (n1038,n563,n555);
or (n1039,n1040,n1041);
and (n1040,n626,n639);
and (n1041,n627,n633);
and (n1042,n1035,n1038);
and (n1043,n1030,n1031);
and (n1044,n1025,n1026);
nand (n1045,n1046,n1075);
nor (n1046,n1047,n1070);
nor (n1047,n1048,n1061);
xor (n1048,n1049,n1060);
xor (n1049,n1050,n1051);
xor (n1050,n991,n1006);
or (n1051,n1052,n1059);
and (n1052,n1053,n1056);
xor (n1053,n1054,n1055);
xor (n1054,n1008,n1015);
xor (n1055,n995,n1002);
or (n1056,n1057,n1058);
and (n1057,n534,n553);
and (n1058,n535,n544);
and (n1059,n1054,n1055);
xor (n1060,n1029,n1032);
or (n1061,n1062,n1069);
and (n1062,n1063,n1068);
xor (n1063,n1064,n1065);
xor (n1064,n1034,n1039);
or (n1065,n1066,n1067);
and (n1066,n575,n625);
and (n1067,n576,n597);
xor (n1068,n1053,n1056);
and (n1069,n1064,n1065);
nor (n1070,n1071,n1074);
or (n1071,n1072,n1073);
and (n1072,n532,n645);
and (n1073,n533,n574);
xor (n1074,n1063,n1068);
nand (n1075,n1076,n1078);
not (n1076,n1077);
xor (n1077,n1024,n1027);
not (n1078,n1079);
or (n1079,n1080,n1081);
and (n1080,n1049,n1060);
and (n1081,n1050,n1051);
nor (n1082,n1083,n1094);
and (n1083,n1084,n1085);
not (n1084,n980);
nand (n1085,n1086,n1093);
or (n1086,n1087,n1088);
not (n1087,n1075);
not (n1088,n1089);
nand (n1089,n1090,n1092);
or (n1090,n1047,n1091);
nand (n1091,n1071,n1074);
nand (n1092,n1048,n1061);
nand (n1093,n1077,n1079);
and (n1094,n981,n1022);
not (n1095,n1096);
nor (n1096,n1097,n1098);
xor (n1097,n430,n518);
or (n1098,n1099,n1100);
and (n1099,n982,n1021);
and (n1100,n983,n984);
not (n1101,n1102);
nand (n1102,n1097,n1098);
or (n1103,n522,n3);
xor (n1104,n1105,n1893);
xor (n1105,n1106,n1892);
xor (n1106,n1107,n1883);
xor (n1107,n1108,n1882);
xor (n1108,n1109,n1867);
xor (n1109,n1110,n1866);
xor (n1110,n1111,n1845);
xor (n1111,n1112,n1844);
xor (n1112,n1113,n1817);
xor (n1113,n1114,n1816);
xor (n1114,n1115,n1783);
xor (n1115,n1116,n169);
xor (n1116,n1117,n1745);
xor (n1117,n1118,n1744);
xor (n1118,n1119,n1700);
xor (n1119,n1120,n1699);
xor (n1120,n1121,n1649);
xor (n1121,n1122,n1648);
xor (n1122,n1123,n1594);
xor (n1123,n1124,n1593);
xor (n1124,n1125,n1531);
xor (n1125,n1126,n1530);
xor (n1126,n1127,n1461);
xor (n1127,n1128,n150);
xor (n1128,n1129,n1387);
xor (n1129,n1130,n1386);
xor (n1130,n1131,n1309);
xor (n1131,n1132,n89);
xor (n1132,n1133,n1223);
xor (n1133,n1134,n1222);
xor (n1134,n219,n1135);
or (n1135,n1136,n1139);
and (n1136,n1137,n1138);
and (n1137,n217,n212);
and (n1138,n105,n96);
and (n1139,n1140,n1141);
xor (n1140,n1137,n1138);
or (n1141,n1142,n1145);
and (n1142,n1143,n1144);
and (n1143,n105,n212);
and (n1144,n86,n96);
and (n1145,n1146,n1147);
xor (n1146,n1143,n1144);
or (n1147,n1148,n1150);
and (n1148,n1149,n261);
and (n1149,n86,n212);
and (n1150,n1151,n1152);
xor (n1151,n1149,n261);
or (n1152,n1153,n1156);
and (n1153,n1154,n1155);
and (n1154,n155,n212);
and (n1155,n149,n96);
and (n1156,n1157,n1158);
xor (n1157,n1154,n1155);
or (n1158,n1159,n1162);
and (n1159,n1160,n1161);
and (n1160,n149,n212);
and (n1161,n36,n96);
and (n1162,n1163,n1164);
xor (n1163,n1160,n1161);
or (n1164,n1165,n1168);
and (n1165,n1166,n1167);
and (n1166,n36,n212);
and (n1167,n17,n96);
and (n1168,n1169,n1170);
xor (n1169,n1166,n1167);
or (n1170,n1171,n1174);
and (n1171,n1172,n1173);
and (n1172,n17,n212);
and (n1173,n131,n96);
and (n1174,n1175,n1176);
xor (n1175,n1172,n1173);
or (n1176,n1177,n1180);
and (n1177,n1178,n1179);
and (n1178,n131,n212);
and (n1179,n114,n96);
and (n1180,n1181,n1182);
xor (n1181,n1178,n1179);
or (n1182,n1183,n1186);
and (n1183,n1184,n1185);
and (n1184,n114,n212);
and (n1185,n184,n96);
and (n1186,n1187,n1188);
xor (n1187,n1184,n1185);
or (n1188,n1189,n1191);
and (n1189,n1190,n757);
and (n1190,n184,n212);
and (n1191,n1192,n1193);
xor (n1192,n1190,n757);
or (n1193,n1194,n1197);
and (n1194,n1195,n1196);
and (n1195,n166,n212);
and (n1196,n205,n96);
and (n1197,n1198,n1199);
xor (n1198,n1195,n1196);
or (n1199,n1200,n1202);
and (n1200,n1201,n844);
and (n1201,n205,n212);
and (n1202,n1203,n1204);
xor (n1203,n1201,n844);
or (n1204,n1205,n1207);
and (n1205,n1206,n901);
and (n1206,n193,n212);
and (n1207,n1208,n1209);
xor (n1208,n1206,n901);
or (n1209,n1210,n1212);
and (n1210,n1211,n914);
and (n1211,n63,n212);
and (n1212,n1213,n1214);
xor (n1213,n1211,n914);
or (n1214,n1215,n1217);
and (n1215,n1216,n945);
and (n1216,n45,n212);
and (n1217,n1218,n1219);
xor (n1218,n1216,n945);
and (n1219,n1220,n1221);
and (n1220,n77,n212);
and (n1221,n68,n96);
and (n1222,n105,n95);
or (n1223,n1224,n1227);
and (n1224,n1225,n1226);
xor (n1225,n1140,n1141);
and (n1226,n86,n95);
and (n1227,n1228,n1229);
xor (n1228,n1225,n1226);
or (n1229,n1230,n1233);
and (n1230,n1231,n1232);
xor (n1231,n1146,n1147);
and (n1232,n155,n95);
and (n1233,n1234,n1235);
xor (n1234,n1231,n1232);
or (n1235,n1236,n1239);
and (n1236,n1237,n1238);
xor (n1237,n1151,n1152);
and (n1238,n149,n95);
and (n1239,n1240,n1241);
xor (n1240,n1237,n1238);
or (n1241,n1242,n1245);
and (n1242,n1243,n1244);
xor (n1243,n1157,n1158);
and (n1244,n36,n95);
and (n1245,n1246,n1247);
xor (n1246,n1243,n1244);
or (n1247,n1248,n1251);
and (n1248,n1249,n1250);
xor (n1249,n1163,n1164);
and (n1250,n17,n95);
and (n1251,n1252,n1253);
xor (n1252,n1249,n1250);
or (n1253,n1254,n1257);
and (n1254,n1255,n1256);
xor (n1255,n1169,n1170);
and (n1256,n131,n95);
and (n1257,n1258,n1259);
xor (n1258,n1255,n1256);
or (n1259,n1260,n1263);
and (n1260,n1261,n1262);
xor (n1261,n1175,n1176);
and (n1262,n114,n95);
and (n1263,n1264,n1265);
xor (n1264,n1261,n1262);
or (n1265,n1266,n1269);
and (n1266,n1267,n1268);
xor (n1267,n1181,n1182);
and (n1268,n184,n95);
and (n1269,n1270,n1271);
xor (n1270,n1267,n1268);
or (n1271,n1272,n1275);
and (n1272,n1273,n1274);
xor (n1273,n1187,n1188);
and (n1274,n166,n95);
and (n1275,n1276,n1277);
xor (n1276,n1273,n1274);
or (n1277,n1278,n1281);
and (n1278,n1279,n1280);
xor (n1279,n1192,n1193);
and (n1280,n205,n95);
and (n1281,n1282,n1283);
xor (n1282,n1279,n1280);
or (n1283,n1284,n1287);
and (n1284,n1285,n1286);
xor (n1285,n1198,n1199);
and (n1286,n193,n95);
and (n1287,n1288,n1289);
xor (n1288,n1285,n1286);
or (n1289,n1290,n1293);
and (n1290,n1291,n1292);
xor (n1291,n1203,n1204);
and (n1292,n63,n95);
and (n1293,n1294,n1295);
xor (n1294,n1291,n1292);
or (n1295,n1296,n1299);
and (n1296,n1297,n1298);
xor (n1297,n1208,n1209);
and (n1298,n45,n95);
and (n1299,n1300,n1301);
xor (n1300,n1297,n1298);
or (n1301,n1302,n1305);
and (n1302,n1303,n1304);
xor (n1303,n1213,n1214);
and (n1304,n77,n95);
and (n1305,n1306,n1307);
xor (n1306,n1303,n1304);
and (n1307,n1308,n920);
xor (n1308,n1218,n1219);
or (n1309,n1310,n1312);
and (n1310,n1311,n288);
xor (n1311,n1228,n1229);
and (n1312,n1313,n1314);
xor (n1313,n1311,n288);
or (n1314,n1315,n1318);
and (n1315,n1316,n1317);
xor (n1316,n1234,n1235);
and (n1317,n149,n88);
and (n1318,n1319,n1320);
xor (n1319,n1316,n1317);
or (n1320,n1321,n1324);
and (n1321,n1322,n1323);
xor (n1322,n1240,n1241);
and (n1323,n36,n88);
and (n1324,n1325,n1326);
xor (n1325,n1322,n1323);
or (n1326,n1327,n1329);
and (n1327,n1328,n476);
xor (n1328,n1246,n1247);
and (n1329,n1330,n1331);
xor (n1330,n1328,n476);
or (n1331,n1332,n1335);
and (n1332,n1333,n1334);
xor (n1333,n1252,n1253);
and (n1334,n131,n88);
and (n1335,n1336,n1337);
xor (n1336,n1333,n1334);
or (n1337,n1338,n1341);
and (n1338,n1339,n1340);
xor (n1339,n1258,n1259);
and (n1340,n114,n88);
and (n1341,n1342,n1343);
xor (n1342,n1339,n1340);
or (n1343,n1344,n1347);
and (n1344,n1345,n1346);
xor (n1345,n1264,n1265);
and (n1346,n184,n88);
and (n1347,n1348,n1349);
xor (n1348,n1345,n1346);
or (n1349,n1350,n1353);
and (n1350,n1351,n1352);
xor (n1351,n1270,n1271);
and (n1352,n166,n88);
and (n1353,n1354,n1355);
xor (n1354,n1351,n1352);
or (n1355,n1356,n1359);
and (n1356,n1357,n1358);
xor (n1357,n1276,n1277);
and (n1358,n205,n88);
and (n1359,n1360,n1361);
xor (n1360,n1357,n1358);
or (n1361,n1362,n1365);
and (n1362,n1363,n1364);
xor (n1363,n1282,n1283);
and (n1364,n193,n88);
and (n1365,n1366,n1367);
xor (n1366,n1363,n1364);
or (n1367,n1368,n1371);
and (n1368,n1369,n1370);
xor (n1369,n1288,n1289);
and (n1370,n63,n88);
and (n1371,n1372,n1373);
xor (n1372,n1369,n1370);
or (n1373,n1374,n1376);
and (n1374,n1375,n866);
xor (n1375,n1294,n1295);
and (n1376,n1377,n1378);
xor (n1377,n1375,n866);
or (n1378,n1379,n1381);
and (n1379,n1380,n893);
xor (n1380,n1300,n1301);
and (n1381,n1382,n1383);
xor (n1382,n1380,n893);
and (n1383,n1384,n1385);
xor (n1384,n1306,n1307);
and (n1385,n68,n88);
and (n1386,n155,n139);
or (n1387,n1388,n1391);
and (n1388,n1389,n1390);
xor (n1389,n1313,n1314);
and (n1390,n149,n139);
and (n1391,n1392,n1393);
xor (n1392,n1389,n1390);
or (n1393,n1394,n1397);
and (n1394,n1395,n1396);
xor (n1395,n1319,n1320);
and (n1396,n36,n139);
and (n1397,n1398,n1399);
xor (n1398,n1395,n1396);
or (n1399,n1400,n1403);
and (n1400,n1401,n1402);
xor (n1401,n1325,n1326);
and (n1402,n17,n139);
and (n1403,n1404,n1405);
xor (n1404,n1401,n1402);
or (n1405,n1406,n1409);
and (n1406,n1407,n1408);
xor (n1407,n1330,n1331);
and (n1408,n131,n139);
and (n1409,n1410,n1411);
xor (n1410,n1407,n1408);
or (n1411,n1412,n1415);
and (n1412,n1413,n1414);
xor (n1413,n1336,n1337);
and (n1414,n114,n139);
and (n1415,n1416,n1417);
xor (n1416,n1413,n1414);
or (n1417,n1418,n1421);
and (n1418,n1419,n1420);
xor (n1419,n1342,n1343);
and (n1420,n184,n139);
and (n1421,n1422,n1423);
xor (n1422,n1419,n1420);
or (n1423,n1424,n1427);
and (n1424,n1425,n1426);
xor (n1425,n1348,n1349);
and (n1426,n166,n139);
and (n1427,n1428,n1429);
xor (n1428,n1425,n1426);
or (n1429,n1430,n1433);
and (n1430,n1431,n1432);
xor (n1431,n1354,n1355);
and (n1432,n205,n139);
and (n1433,n1434,n1435);
xor (n1434,n1431,n1432);
or (n1435,n1436,n1439);
and (n1436,n1437,n1438);
xor (n1437,n1360,n1361);
and (n1438,n193,n139);
and (n1439,n1440,n1441);
xor (n1440,n1437,n1438);
or (n1441,n1442,n1445);
and (n1442,n1443,n1444);
xor (n1443,n1366,n1367);
and (n1444,n63,n139);
and (n1445,n1446,n1447);
xor (n1446,n1443,n1444);
or (n1447,n1448,n1451);
and (n1448,n1449,n1450);
xor (n1449,n1372,n1373);
and (n1450,n45,n139);
and (n1451,n1452,n1453);
xor (n1452,n1449,n1450);
or (n1453,n1454,n1457);
and (n1454,n1455,n1456);
xor (n1455,n1377,n1378);
and (n1456,n77,n139);
and (n1457,n1458,n1459);
xor (n1458,n1455,n1456);
and (n1459,n1460,n850);
xor (n1460,n1382,n1383);
or (n1461,n1462,n1465);
and (n1462,n1463,n1464);
xor (n1463,n1392,n1393);
and (n1464,n36,n30);
and (n1465,n1466,n1467);
xor (n1466,n1463,n1464);
or (n1467,n1468,n1471);
and (n1468,n1469,n1470);
xor (n1469,n1398,n1399);
and (n1470,n17,n30);
and (n1471,n1472,n1473);
xor (n1472,n1469,n1470);
or (n1473,n1474,n1477);
and (n1474,n1475,n1476);
xor (n1475,n1404,n1405);
and (n1476,n131,n30);
and (n1477,n1478,n1479);
xor (n1478,n1475,n1476);
or (n1479,n1480,n1483);
and (n1480,n1481,n1482);
xor (n1481,n1410,n1411);
and (n1482,n114,n30);
and (n1483,n1484,n1485);
xor (n1484,n1481,n1482);
or (n1485,n1486,n1489);
and (n1486,n1487,n1488);
xor (n1487,n1416,n1417);
and (n1488,n184,n30);
and (n1489,n1490,n1491);
xor (n1490,n1487,n1488);
or (n1491,n1492,n1495);
and (n1492,n1493,n1494);
xor (n1493,n1422,n1423);
and (n1494,n166,n30);
and (n1495,n1496,n1497);
xor (n1496,n1493,n1494);
or (n1497,n1498,n1501);
and (n1498,n1499,n1500);
xor (n1499,n1428,n1429);
and (n1500,n205,n30);
and (n1501,n1502,n1503);
xor (n1502,n1499,n1500);
or (n1503,n1504,n1507);
and (n1504,n1505,n1506);
xor (n1505,n1434,n1435);
and (n1506,n193,n30);
and (n1507,n1508,n1509);
xor (n1508,n1505,n1506);
or (n1509,n1510,n1513);
and (n1510,n1511,n1512);
xor (n1511,n1440,n1441);
and (n1512,n63,n30);
and (n1513,n1514,n1515);
xor (n1514,n1511,n1512);
or (n1515,n1516,n1519);
and (n1516,n1517,n1518);
xor (n1517,n1446,n1447);
and (n1518,n45,n30);
and (n1519,n1520,n1521);
xor (n1520,n1517,n1518);
or (n1521,n1522,n1525);
and (n1522,n1523,n1524);
xor (n1523,n1452,n1453);
and (n1524,n77,n30);
and (n1525,n1526,n1527);
xor (n1526,n1523,n1524);
and (n1527,n1528,n1529);
xor (n1528,n1458,n1459);
and (n1529,n68,n30);
and (n1530,n36,n24);
or (n1531,n1532,n1535);
and (n1532,n1533,n1534);
xor (n1533,n1466,n1467);
and (n1534,n17,n24);
and (n1535,n1536,n1537);
xor (n1536,n1533,n1534);
or (n1537,n1538,n1541);
and (n1538,n1539,n1540);
xor (n1539,n1472,n1473);
and (n1540,n131,n24);
and (n1541,n1542,n1543);
xor (n1542,n1539,n1540);
or (n1543,n1544,n1547);
and (n1544,n1545,n1546);
xor (n1545,n1478,n1479);
and (n1546,n114,n24);
and (n1547,n1548,n1549);
xor (n1548,n1545,n1546);
or (n1549,n1550,n1553);
and (n1550,n1551,n1552);
xor (n1551,n1484,n1485);
and (n1552,n184,n24);
and (n1553,n1554,n1555);
xor (n1554,n1551,n1552);
or (n1555,n1556,n1559);
and (n1556,n1557,n1558);
xor (n1557,n1490,n1491);
and (n1558,n166,n24);
and (n1559,n1560,n1561);
xor (n1560,n1557,n1558);
or (n1561,n1562,n1565);
and (n1562,n1563,n1564);
xor (n1563,n1496,n1497);
and (n1564,n205,n24);
and (n1565,n1566,n1567);
xor (n1566,n1563,n1564);
or (n1567,n1568,n1571);
and (n1568,n1569,n1570);
xor (n1569,n1502,n1503);
and (n1570,n193,n24);
and (n1571,n1572,n1573);
xor (n1572,n1569,n1570);
or (n1573,n1574,n1577);
and (n1574,n1575,n1576);
xor (n1575,n1508,n1509);
and (n1576,n63,n24);
and (n1577,n1578,n1579);
xor (n1578,n1575,n1576);
or (n1579,n1580,n1583);
and (n1580,n1581,n1582);
xor (n1581,n1514,n1515);
and (n1582,n45,n24);
and (n1583,n1584,n1585);
xor (n1584,n1581,n1582);
or (n1585,n1586,n1589);
and (n1586,n1587,n1588);
xor (n1587,n1520,n1521);
and (n1588,n77,n24);
and (n1589,n1590,n1591);
xor (n1590,n1587,n1588);
and (n1591,n1592,n750);
xor (n1592,n1526,n1527);
and (n1593,n17,n18);
or (n1594,n1595,n1598);
and (n1595,n1596,n1597);
xor (n1596,n1536,n1537);
and (n1597,n131,n18);
and (n1598,n1599,n1600);
xor (n1599,n1596,n1597);
or (n1600,n1601,n1603);
and (n1601,n1602,n305);
xor (n1602,n1542,n1543);
and (n1603,n1604,n1605);
xor (n1604,n1602,n305);
or (n1605,n1606,n1609);
and (n1606,n1607,n1608);
xor (n1607,n1548,n1549);
and (n1608,n184,n18);
and (n1609,n1610,n1611);
xor (n1610,n1607,n1608);
or (n1611,n1612,n1615);
and (n1612,n1613,n1614);
xor (n1613,n1554,n1555);
and (n1614,n166,n18);
and (n1615,n1616,n1617);
xor (n1616,n1613,n1614);
or (n1617,n1618,n1621);
and (n1618,n1619,n1620);
xor (n1619,n1560,n1561);
and (n1620,n205,n18);
and (n1621,n1622,n1623);
xor (n1622,n1619,n1620);
or (n1623,n1624,n1627);
and (n1624,n1625,n1626);
xor (n1625,n1566,n1567);
and (n1626,n193,n18);
and (n1627,n1628,n1629);
xor (n1628,n1625,n1626);
or (n1629,n1630,n1632);
and (n1630,n1631,n591);
xor (n1631,n1572,n1573);
and (n1632,n1633,n1634);
xor (n1633,n1631,n591);
or (n1634,n1635,n1637);
and (n1635,n1636,n668);
xor (n1636,n1578,n1579);
and (n1637,n1638,n1639);
xor (n1638,n1636,n668);
or (n1639,n1640,n1643);
and (n1640,n1641,n1642);
xor (n1641,n1584,n1585);
and (n1642,n77,n18);
and (n1643,n1644,n1645);
xor (n1644,n1641,n1642);
and (n1645,n1646,n1647);
xor (n1646,n1590,n1591);
and (n1647,n68,n18);
and (n1648,n131,n121);
or (n1649,n1650,n1653);
and (n1650,n1651,n1652);
xor (n1651,n1599,n1600);
and (n1652,n114,n121);
and (n1653,n1654,n1655);
xor (n1654,n1651,n1652);
or (n1655,n1656,n1659);
and (n1656,n1657,n1658);
xor (n1657,n1604,n1605);
and (n1658,n184,n121);
and (n1659,n1660,n1661);
xor (n1660,n1657,n1658);
or (n1661,n1662,n1665);
and (n1662,n1663,n1664);
xor (n1663,n1610,n1611);
and (n1664,n166,n121);
and (n1665,n1666,n1667);
xor (n1666,n1663,n1664);
or (n1667,n1668,n1671);
and (n1668,n1669,n1670);
xor (n1669,n1616,n1617);
and (n1670,n205,n121);
and (n1671,n1672,n1673);
xor (n1672,n1669,n1670);
or (n1673,n1674,n1677);
and (n1674,n1675,n1676);
xor (n1675,n1622,n1623);
and (n1676,n193,n121);
and (n1677,n1678,n1679);
xor (n1678,n1675,n1676);
or (n1679,n1680,n1683);
and (n1680,n1681,n1682);
xor (n1681,n1628,n1629);
and (n1682,n63,n121);
and (n1683,n1684,n1685);
xor (n1684,n1681,n1682);
or (n1685,n1686,n1689);
and (n1686,n1687,n1688);
xor (n1687,n1633,n1634);
and (n1688,n45,n121);
and (n1689,n1690,n1691);
xor (n1690,n1687,n1688);
or (n1691,n1692,n1695);
and (n1692,n1693,n1694);
xor (n1693,n1638,n1639);
and (n1694,n77,n121);
and (n1695,n1696,n1697);
xor (n1696,n1693,n1694);
and (n1697,n1698,n654);
xor (n1698,n1644,n1645);
and (n1699,n114,n112);
or (n1700,n1701,n1704);
and (n1701,n1702,n1703);
xor (n1702,n1654,n1655);
and (n1703,n184,n112);
and (n1704,n1705,n1706);
xor (n1705,n1702,n1703);
or (n1706,n1707,n1709);
and (n1707,n1708,n319);
xor (n1708,n1660,n1661);
and (n1709,n1710,n1711);
xor (n1710,n1708,n319);
or (n1711,n1712,n1715);
and (n1712,n1713,n1714);
xor (n1713,n1666,n1667);
and (n1714,n205,n112);
and (n1715,n1716,n1717);
xor (n1716,n1713,n1714);
or (n1717,n1718,n1721);
and (n1718,n1719,n1720);
xor (n1719,n1672,n1673);
and (n1720,n193,n112);
and (n1721,n1722,n1723);
xor (n1722,n1719,n1720);
or (n1723,n1724,n1727);
and (n1724,n1725,n1726);
xor (n1725,n1678,n1679);
and (n1726,n63,n112);
and (n1727,n1728,n1729);
xor (n1728,n1725,n1726);
or (n1729,n1730,n1733);
and (n1730,n1731,n1732);
xor (n1731,n1684,n1685);
and (n1732,n45,n112);
and (n1733,n1734,n1735);
xor (n1734,n1731,n1732);
or (n1735,n1736,n1739);
and (n1736,n1737,n1738);
xor (n1737,n1690,n1691);
and (n1738,n77,n112);
and (n1739,n1740,n1741);
xor (n1740,n1737,n1738);
and (n1741,n1742,n1743);
xor (n1742,n1696,n1697);
and (n1743,n68,n112);
and (n1744,n184,n175);
or (n1745,n1746,n1749);
and (n1746,n1747,n1748);
xor (n1747,n1705,n1706);
and (n1748,n166,n175);
and (n1749,n1750,n1751);
xor (n1750,n1747,n1748);
or (n1751,n1752,n1755);
and (n1752,n1753,n1754);
xor (n1753,n1710,n1711);
and (n1754,n205,n175);
and (n1755,n1756,n1757);
xor (n1756,n1753,n1754);
or (n1757,n1758,n1761);
and (n1758,n1759,n1760);
xor (n1759,n1716,n1717);
and (n1760,n193,n175);
and (n1761,n1762,n1763);
xor (n1762,n1759,n1760);
or (n1763,n1764,n1767);
and (n1764,n1765,n1766);
xor (n1765,n1722,n1723);
and (n1766,n63,n175);
and (n1767,n1768,n1769);
xor (n1768,n1765,n1766);
or (n1769,n1770,n1773);
and (n1770,n1771,n1772);
xor (n1771,n1728,n1729);
and (n1772,n45,n175);
and (n1773,n1774,n1775);
xor (n1774,n1771,n1772);
or (n1775,n1776,n1779);
and (n1776,n1777,n1778);
xor (n1777,n1734,n1735);
and (n1778,n77,n175);
and (n1779,n1780,n1781);
xor (n1780,n1777,n1778);
and (n1781,n1782,n561);
xor (n1782,n1740,n1741);
or (n1783,n1784,n1787);
and (n1784,n1785,n1786);
xor (n1785,n1750,n1751);
and (n1786,n205,n168);
and (n1787,n1788,n1789);
xor (n1788,n1785,n1786);
or (n1789,n1790,n1793);
and (n1790,n1791,n1792);
xor (n1791,n1756,n1757);
and (n1792,n193,n168);
and (n1793,n1794,n1795);
xor (n1794,n1791,n1792);
or (n1795,n1796,n1799);
and (n1796,n1797,n1798);
xor (n1797,n1762,n1763);
and (n1798,n63,n168);
and (n1799,n1800,n1801);
xor (n1800,n1797,n1798);
or (n1801,n1802,n1805);
and (n1802,n1803,n1804);
xor (n1803,n1768,n1769);
and (n1804,n45,n168);
and (n1805,n1806,n1807);
xor (n1806,n1803,n1804);
or (n1807,n1808,n1811);
and (n1808,n1809,n1810);
xor (n1809,n1774,n1775);
and (n1810,n77,n168);
and (n1811,n1812,n1813);
xor (n1812,n1809,n1810);
and (n1813,n1814,n1815);
xor (n1814,n1780,n1781);
and (n1815,n68,n168);
and (n1816,n205,n199);
or (n1817,n1818,n1821);
and (n1818,n1819,n1820);
xor (n1819,n1788,n1789);
and (n1820,n193,n199);
and (n1821,n1822,n1823);
xor (n1822,n1819,n1820);
or (n1823,n1824,n1827);
and (n1824,n1825,n1826);
xor (n1825,n1794,n1795);
and (n1826,n63,n199);
and (n1827,n1828,n1829);
xor (n1828,n1825,n1826);
or (n1829,n1830,n1833);
and (n1830,n1831,n1832);
xor (n1831,n1800,n1801);
and (n1832,n45,n199);
and (n1833,n1834,n1835);
xor (n1834,n1831,n1832);
or (n1835,n1836,n1839);
and (n1836,n1837,n1838);
xor (n1837,n1806,n1807);
and (n1838,n77,n199);
and (n1839,n1840,n1841);
xor (n1840,n1837,n1838);
and (n1841,n1842,n1843);
xor (n1842,n1812,n1813);
not (n1843,n455);
and (n1844,n193,n53);
or (n1845,n1846,n1849);
and (n1846,n1847,n1848);
xor (n1847,n1822,n1823);
and (n1848,n63,n53);
and (n1849,n1850,n1851);
xor (n1850,n1847,n1848);
or (n1851,n1852,n1855);
and (n1852,n1853,n1854);
xor (n1853,n1828,n1829);
and (n1854,n45,n53);
and (n1855,n1856,n1857);
xor (n1856,n1853,n1854);
or (n1857,n1858,n1861);
and (n1858,n1859,n1860);
xor (n1859,n1834,n1835);
and (n1860,n77,n53);
and (n1861,n1862,n1863);
xor (n1862,n1859,n1860);
and (n1863,n1864,n1865);
xor (n1864,n1840,n1841);
and (n1865,n68,n53);
and (n1866,n63,n54);
or (n1867,n1868,n1871);
and (n1868,n1869,n1870);
xor (n1869,n1850,n1851);
and (n1870,n45,n54);
and (n1871,n1872,n1873);
xor (n1872,n1869,n1870);
or (n1873,n1874,n1877);
and (n1874,n1875,n1876);
xor (n1875,n1856,n1857);
and (n1876,n77,n54);
and (n1877,n1878,n1879);
xor (n1878,n1875,n1876);
and (n1879,n1880,n1881);
xor (n1880,n1862,n1863);
not (n1881,n240);
and (n1882,n45,n43);
or (n1883,n1884,n1887);
and (n1884,n1885,n1886);
xor (n1885,n1872,n1873);
and (n1886,n77,n43);
and (n1887,n1888,n1889);
xor (n1888,n1885,n1886);
and (n1889,n1890,n1891);
xor (n1890,n1878,n1879);
and (n1891,n68,n43);
and (n1892,n77,n72);
and (n1893,n1894,n1895);
xor (n1894,n1888,n1889);
and (n1895,n68,n72);
endmodule
