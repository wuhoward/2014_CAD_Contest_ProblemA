module top (out,n16,n18,n19,n21,n24,n28,n30,n32,n35
        ,n39,n41,n42,n44,n47,n53,n55,n56,n58,n61
        ,n65,n67,n68,n72,n76,n78,n80,n89,n91,n100
        ,n102,n104,n107,n117,n120,n125,n132,n143,n145,n148
        ,n152,n154,n156,n169,n192,n221,n225,n232,n405);
output out;
input n16;
input n18;
input n19;
input n21;
input n24;
input n28;
input n30;
input n32;
input n35;
input n39;
input n41;
input n42;
input n44;
input n47;
input n53;
input n55;
input n56;
input n58;
input n61;
input n65;
input n67;
input n68;
input n72;
input n76;
input n78;
input n80;
input n89;
input n91;
input n100;
input n102;
input n104;
input n107;
input n117;
input n120;
input n125;
input n132;
input n143;
input n145;
input n148;
input n152;
input n154;
input n156;
input n169;
input n192;
input n221;
input n225;
input n232;
input n405;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n17;
wire n20;
wire n22;
wire n23;
wire n25;
wire n26;
wire n27;
wire n29;
wire n31;
wire n33;
wire n34;
wire n36;
wire n37;
wire n38;
wire n40;
wire n43;
wire n45;
wire n46;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n54;
wire n57;
wire n59;
wire n60;
wire n62;
wire n63;
wire n64;
wire n66;
wire n69;
wire n70;
wire n71;
wire n73;
wire n74;
wire n75;
wire n77;
wire n79;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n90;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n101;
wire n103;
wire n105;
wire n106;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n118;
wire n119;
wire n121;
wire n122;
wire n123;
wire n124;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n144;
wire n146;
wire n147;
wire n149;
wire n150;
wire n151;
wire n153;
wire n155;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n193;
wire n194;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n222;
wire n223;
wire n224;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
xor (out,n0,n2247);
xnor (n0,n1,n2149);
nand (n1,n2,n748);
nor (n2,n3,n746);
nor (n3,n4,n647);
nand (n4,n5,n549);
nand (n5,n6,n454,n548);
nand (n6,n7,n283);
nand (n7,n8,n179,n282);
nand (n8,n9,n109);
xor (n9,n10,n83);
xor (n10,n11,n48);
xor (n11,n12,n36);
xor (n12,n13,n25);
xor (n13,n14,n24);
or (n14,n15,n20);
and (n15,n16,n17);
xor (n17,n18,n19);
and (n20,n21,n22);
nor (n22,n17,n23);
xnor (n23,n24,n18);
xor (n25,n26,n35);
or (n26,n27,n31);
and (n27,n28,n29);
xor (n29,n30,n24);
and (n31,n32,n33);
nor (n33,n29,n34);
xnor (n34,n35,n30);
xor (n36,n37,n47);
or (n37,n38,n43);
and (n38,n39,n40);
xor (n40,n41,n42);
and (n43,n44,n45);
nor (n45,n40,n46);
xnor (n46,n47,n41);
xor (n48,n49,n73);
xor (n49,n50,n62);
xor (n50,n51,n61);
or (n51,n52,n57);
and (n52,n53,n54);
xor (n54,n55,n56);
and (n57,n58,n59);
nor (n59,n54,n60);
xnor (n60,n61,n55);
xor (n62,n63,n72);
or (n63,n64,n69);
and (n64,n65,n66);
xor (n66,n67,n68);
and (n69,n65,n70);
nor (n70,n66,n71);
xnor (n71,n72,n67);
xor (n73,n74,n19);
or (n74,n75,n79);
and (n75,n76,n77);
xor (n77,n78,n61);
and (n79,n80,n81);
nor (n81,n77,n82);
xnor (n82,n19,n78);
nand (n83,n84,n96,n108);
nand (n84,n85,n90);
xor (n85,n86,n47);
or (n86,n87,n88);
and (n87,n44,n40);
and (n88,n89,n45);
and (n90,n91,n92);
xor (n92,n93,n61);
or (n93,n94,n95);
and (n94,n76,n54);
and (n95,n80,n59);
nand (n96,n97,n90);
xor (n97,n98,n107);
or (n98,n99,n103);
and (n99,n100,n101);
xor (n101,n102,n47);
and (n103,n104,n105);
nor (n105,n101,n106);
xnor (n106,n107,n102);
nand (n108,n85,n97);
nand (n109,n110,n136,n178);
nand (n110,n111,n134);
nand (n111,n112,n127,n133);
nand (n112,n91,n113);
and (n113,n114,n122);
xnor (n114,n115,n68);
nor (n115,n116,n121);
and (n116,n117,n118);
and (n118,n119,n68);
not (n119,n120);
and (n121,n65,n120);
xor (n122,n123,n72);
or (n123,n124,n126);
and (n124,n125,n66);
and (n126,n53,n70);
nand (n127,n128,n113);
xor (n128,n129,n107);
or (n129,n130,n131);
and (n130,n104,n101);
and (n131,n132,n105);
nand (n133,n91,n128);
xor (n134,n135,n97);
xor (n135,n85,n90);
nand (n136,n137,n134);
xor (n137,n138,n159);
xor (n138,n139,n149);
xor (n139,n140,n148);
or (n140,n141,n144);
and (n141,n132,n142);
xor (n142,n143,n107);
and (n144,n145,n146);
nor (n146,n142,n147);
xnor (n147,n148,n143);
xor (n149,n150,n91);
or (n150,n151,n155);
and (n151,n152,n153);
xor (n153,n154,n148);
and (n155,n156,n157);
nor (n157,n153,n158);
xnor (n158,n91,n154);
nand (n159,n160,n173,n177);
nand (n160,n161,n165);
xor (n161,n162,n72);
or (n162,n163,n164);
and (n163,n117,n66);
and (n164,n125,n70);
xor (n165,n166,n56);
or (n166,n167,n170);
and (n167,n53,n168);
xor (n168,n169,n72);
and (n170,n58,n171);
nor (n171,n168,n172);
xnor (n172,n56,n169);
nand (n173,n174,n165);
xnor (n174,n175,n68);
nor (n175,n176,n121);
and (n176,n65,n118);
nand (n177,n161,n174);
nand (n178,n111,n137);
nand (n179,n180,n109);
nand (n180,n181,n253,n281);
nand (n181,n182,n211);
nand (n182,n183,n193,n210);
nand (n183,n184,n188);
xor (n184,n185,n148);
or (n185,n186,n187);
and (n186,n145,n142);
and (n187,n152,n146);
xor (n188,n189,n91);
or (n189,n190,n191);
and (n190,n156,n153);
and (n191,n192,n157);
nand (n193,n194,n188);
nand (n194,n195,n204,n209);
nand (n195,n196,n200);
xor (n196,n197,n61);
or (n197,n198,n199);
and (n198,n80,n54);
and (n199,n16,n59);
xor (n200,n201,n56);
or (n201,n202,n203);
and (n202,n58,n168);
and (n203,n76,n171);
nand (n204,n205,n200);
xor (n205,n206,n19);
or (n206,n207,n208);
and (n207,n21,n77);
and (n208,n28,n81);
nand (n209,n196,n205);
nand (n210,n184,n194);
nand (n211,n212,n237,n252);
nand (n212,n213,n215);
xor (n213,n214,n174);
xor (n214,n161,n165);
nand (n215,n216,n227,n236);
nand (n216,n217,n222);
xor (n217,n218,n24);
or (n218,n219,n220);
and (n219,n32,n17);
and (n220,n221,n22);
xor (n222,n223,n35);
or (n223,n224,n226);
and (n224,n225,n29);
and (n226,n39,n33);
nand (n227,n228,n222);
xor (n228,n229,n42);
or (n229,n230,n233);
and (n230,n44,n231);
xor (n231,n232,n35);
and (n233,n89,n234);
nor (n234,n231,n235);
xnor (n235,n42,n232);
nand (n236,n217,n228);
nand (n237,n238,n215);
nand (n238,n239,n245,n251);
nand (n239,n240,n244);
xor (n240,n241,n47);
or (n241,n242,n243);
and (n242,n100,n40);
and (n243,n104,n45);
xor (n244,n114,n122);
nand (n245,n246,n244);
and (n246,n91,n247);
xor (n247,n248,n72);
or (n248,n249,n250);
and (n249,n53,n66);
and (n250,n58,n70);
nand (n251,n240,n246);
nand (n252,n213,n238);
nand (n253,n254,n211);
xor (n254,n255,n91);
xor (n255,n256,n272);
nand (n256,n257,n266,n271);
nand (n257,n258,n262);
xor (n258,n259,n19);
or (n259,n260,n261);
and (n260,n16,n77);
and (n261,n21,n81);
xor (n262,n263,n24);
or (n263,n264,n265);
and (n264,n28,n17);
and (n265,n32,n22);
nand (n266,n267,n262);
xor (n267,n268,n35);
or (n268,n269,n270);
and (n269,n221,n29);
and (n270,n225,n33);
nand (n271,n258,n267);
xor (n272,n273,n278);
not (n273,n274);
xor (n274,n275,n61);
or (n275,n276,n277);
and (n276,n58,n54);
and (n277,n76,n59);
xor (n278,n279,n72);
or (n279,n64,n280);
and (n280,n117,n70);
nand (n281,n182,n254);
nand (n282,n9,n180);
nand (n283,n284,n377,n453);
nand (n284,n285,n310);
xor (n285,n286,n306);
xor (n286,n287,n302);
xor (n287,n288,n298);
xor (n288,n289,n294);
not (n289,n290);
xor (n290,n291,n56);
or (n291,n292,n293);
and (n292,n117,n168);
and (n293,n125,n171);
xor (n294,n295,n42);
or (n295,n296,n297);
and (n296,n221,n231);
and (n297,n225,n234);
xor (n298,n299,n107);
or (n299,n300,n301);
and (n300,n89,n101);
and (n301,n100,n105);
nand (n302,n303,n304,n305);
nand (n303,n139,n149);
nand (n304,n159,n149);
nand (n305,n139,n159);
nand (n306,n307,n308,n309);
nand (n307,n256,n272);
nand (n308,n91,n272);
nand (n309,n256,n91);
xor (n310,n311,n356);
xor (n311,n312,n325);
xor (n312,n313,n322);
xor (n313,n314,n318);
xor (n314,n315,n148);
or (n315,n316,n317);
and (n316,n104,n142);
and (n317,n132,n146);
xor (n318,n319,n91);
or (n319,n320,n321);
and (n320,n145,n153);
and (n321,n152,n157);
nand (n322,n273,n323,n324);
nand (n323,n278,n274);
not (n324,n278);
xor (n325,n326,n340);
xor (n326,n91,n327);
nand (n327,n328,n334,n339);
nand (n328,n329,n333);
xor (n329,n330,n56);
or (n330,n331,n332);
and (n331,n125,n168);
and (n332,n53,n171);
not (n333,n174);
nand (n334,n335,n333);
xor (n335,n336,n19);
or (n336,n337,n338);
and (n337,n80,n77);
and (n338,n16,n81);
nand (n339,n329,n335);
nand (n340,n341,n350,n355);
nand (n341,n342,n346);
xor (n342,n343,n24);
or (n343,n344,n345);
and (n344,n21,n17);
and (n345,n28,n22);
xor (n346,n347,n35);
or (n347,n348,n349);
and (n348,n32,n29);
and (n349,n221,n33);
nand (n350,n351,n346);
xor (n351,n352,n42);
or (n352,n353,n354);
and (n353,n225,n231);
and (n354,n39,n234);
nand (n355,n342,n351);
nand (n356,n357,n373,n376);
nand (n357,n358,n371);
nand (n358,n359,n368,n370);
nand (n359,n360,n364);
xor (n360,n361,n42);
or (n361,n362,n363);
and (n362,n39,n231);
and (n363,n44,n234);
xor (n364,n365,n47);
or (n365,n366,n367);
and (n366,n89,n40);
and (n367,n100,n45);
nand (n368,n369,n364);
xor (n369,n91,n92);
nand (n370,n360,n369);
xor (n371,n372,n351);
xor (n372,n342,n346);
nand (n373,n374,n371);
xor (n374,n375,n335);
xor (n375,n329,n333);
nand (n376,n358,n374);
nand (n377,n378,n310);
nand (n378,n379,n392,n452);
nand (n379,n380,n390);
nand (n380,n381,n386,n389);
nand (n381,n382,n384);
xor (n382,n383,n267);
xor (n383,n258,n262);
xor (n384,n385,n128);
xor (n385,n91,n113);
nand (n386,n387,n384);
xor (n387,n388,n369);
xor (n388,n360,n364);
nand (n389,n382,n387);
xor (n390,n391,n374);
xor (n391,n358,n371);
nand (n392,n393,n390);
nand (n393,n394,n448,n451);
nand (n394,n395,n412);
nand (n395,n396,n406,n411);
nand (n396,n397,n401);
xor (n397,n398,n107);
or (n398,n399,n400);
and (n399,n132,n101);
and (n400,n145,n105);
xor (n401,n402,n91);
or (n402,n403,n404);
and (n403,n192,n153);
and (n404,n405,n157);
nand (n406,n407,n401);
xor (n407,n408,n148);
or (n408,n409,n410);
and (n409,n152,n142);
and (n410,n156,n146);
nand (n411,n397,n407);
nand (n412,n413,n432,n447);
nand (n413,n414,n430);
nand (n414,n415,n424,n429);
nand (n415,n416,n420);
xor (n416,n417,n61);
or (n417,n418,n419);
and (n418,n16,n54);
and (n419,n21,n59);
xnor (n420,n421,n68);
nor (n421,n422,n423);
and (n422,n125,n118);
and (n423,n117,n120);
nand (n424,n425,n420);
xor (n425,n426,n56);
or (n426,n427,n428);
and (n427,n76,n168);
and (n428,n80,n171);
nand (n429,n416,n425);
xor (n430,n431,n205);
xor (n431,n196,n200);
nand (n432,n433,n430);
nand (n433,n434,n441,n446);
nand (n434,n435,n439);
xor (n435,n436,n19);
or (n436,n437,n438);
and (n437,n28,n77);
and (n438,n32,n81);
xnor (n439,n440,n91);
nand (n440,n405,n153);
nand (n441,n442,n439);
xor (n442,n443,n24);
or (n443,n444,n445);
and (n444,n221,n17);
and (n445,n225,n22);
nand (n446,n435,n442);
nand (n447,n414,n433);
nand (n448,n449,n412);
xor (n449,n450,n194);
xor (n450,n184,n188);
nand (n451,n395,n449);
nand (n452,n380,n393);
nand (n453,n285,n378);
nand (n454,n455,n283);
xor (n455,n456,n508);
xor (n456,n457,n461);
nand (n457,n458,n459,n460);
nand (n458,n312,n325);
nand (n459,n356,n325);
nand (n460,n312,n356);
xor (n461,n462,n484);
xor (n462,n463,n467);
nand (n463,n464,n465,n466);
nand (n464,n91,n327);
nand (n465,n340,n327);
nand (n466,n91,n340);
xor (n467,n468,n480);
xor (n468,n469,n91);
xor (n469,n470,n479);
xor (n470,n471,n475);
xor (n471,n472,n56);
or (n472,n473,n474);
and (n473,n65,n168);
and (n474,n117,n171);
xor (n475,n476,n61);
or (n476,n477,n478);
and (n477,n125,n54);
and (n478,n53,n59);
not (n479,n62);
nand (n480,n481,n482,n483);
nand (n481,n50,n62);
nand (n482,n73,n62);
nand (n483,n50,n73);
xor (n484,n485,n504);
xor (n485,n486,n500);
xor (n486,n487,n496);
xor (n487,n488,n492);
xor (n488,n489,n19);
or (n489,n490,n491);
and (n490,n58,n77);
and (n491,n76,n81);
xor (n492,n493,n24);
or (n493,n494,n495);
and (n494,n80,n17);
and (n495,n16,n22);
xor (n496,n497,n35);
or (n497,n498,n499);
and (n498,n21,n29);
and (n499,n28,n33);
nand (n500,n501,n502,n503);
nand (n501,n13,n25);
nand (n502,n36,n25);
nand (n503,n13,n36);
nand (n504,n505,n506,n507);
nand (n505,n314,n318);
nand (n506,n322,n318);
nand (n507,n314,n322);
xor (n508,n509,n518);
xor (n509,n510,n514);
nand (n510,n511,n512,n513);
nand (n511,n11,n48);
nand (n512,n83,n48);
nand (n513,n11,n83);
nand (n514,n515,n516,n517);
nand (n515,n287,n302);
nand (n516,n306,n302);
nand (n517,n287,n306);
xor (n518,n519,n534);
xor (n519,n520,n524);
nand (n520,n521,n522,n523);
nand (n521,n289,n294);
nand (n522,n298,n294);
nand (n523,n289,n298);
xor (n524,n525,n530);
xor (n525,n526,n290);
xor (n526,n527,n47);
or (n527,n528,n529);
and (n528,n225,n40);
and (n529,n39,n45);
xor (n530,n531,n42);
or (n531,n532,n533);
and (n532,n32,n231);
and (n533,n221,n234);
xor (n534,n535,n544);
xor (n535,n536,n540);
xor (n536,n537,n107);
or (n537,n538,n539);
and (n538,n44,n101);
and (n539,n89,n105);
xor (n540,n541,n148);
or (n541,n542,n543);
and (n542,n100,n142);
and (n543,n104,n146);
xor (n544,n545,n91);
or (n545,n546,n547);
and (n546,n132,n153);
and (n547,n145,n157);
nand (n548,n7,n455);
xor (n549,n550,n643);
xor (n550,n551,n605);
xor (n551,n552,n580);
xor (n552,n553,n576);
xor (n553,n554,n572);
xor (n554,n555,n559);
nand (n555,n556,n557,n558);
nand (n556,n488,n492);
nand (n557,n496,n492);
nand (n558,n488,n496);
xor (n559,n560,n568);
xor (n560,n561,n564);
xor (n561,n562,n56);
or (n562,n473,n563);
and (n563,n65,n171);
xor (n564,n565,n24);
or (n565,n566,n567);
and (n566,n76,n17);
and (n567,n80,n22);
xor (n568,n569,n35);
or (n569,n570,n571);
and (n570,n16,n29);
and (n571,n21,n33);
nand (n572,n573,n574,n575);
nand (n573,n526,n290);
nand (n574,n530,n290);
nand (n575,n526,n530);
nand (n576,n577,n578,n579);
nand (n577,n520,n524);
nand (n578,n534,n524);
nand (n579,n520,n534);
xor (n580,n581,n601);
xor (n581,n582,n586);
nand (n582,n583,n584,n585);
nand (n583,n536,n540);
nand (n584,n544,n540);
nand (n585,n536,n544);
xor (n586,n587,n597);
xor (n587,n588,n592);
xor (n588,n589,n19);
or (n589,n590,n591);
and (n590,n53,n77);
and (n591,n58,n81);
not (n592,n593);
xor (n593,n594,n61);
or (n594,n595,n596);
and (n595,n117,n54);
and (n596,n125,n59);
xor (n597,n598,n42);
or (n598,n599,n600);
and (n599,n28,n231);
and (n600,n32,n234);
nand (n601,n602,n603,n604);
nand (n602,n469,n91);
nand (n603,n480,n91);
nand (n604,n469,n480);
xor (n605,n606,n639);
xor (n606,n607,n611);
nand (n607,n608,n609,n610);
nand (n608,n463,n467);
nand (n609,n484,n467);
nand (n610,n463,n484);
xor (n611,n612,n635);
xor (n612,n613,n627);
xor (n613,n614,n623);
xor (n614,n615,n619);
xor (n615,n616,n47);
or (n616,n617,n618);
and (n617,n221,n40);
and (n618,n225,n45);
xor (n619,n620,n107);
or (n620,n621,n622);
and (n621,n39,n101);
and (n622,n44,n105);
xor (n623,n624,n148);
or (n624,n625,n626);
and (n625,n89,n142);
and (n626,n100,n146);
xor (n627,n628,n631);
or (n628,n629,n630);
and (n629,n104,n153);
and (n630,n132,n157);
nand (n631,n632,n633,n634);
nand (n632,n471,n475);
nand (n633,n479,n475);
nand (n634,n471,n479);
nand (n635,n636,n637,n638);
nand (n636,n486,n500);
nand (n637,n504,n500);
nand (n638,n486,n504);
nand (n639,n640,n641,n642);
nand (n640,n510,n514);
nand (n641,n518,n514);
nand (n642,n510,n518);
nand (n643,n644,n645,n646);
nand (n644,n457,n461);
nand (n645,n508,n461);
nand (n646,n457,n508);
nor (n647,n648,n652);
nand (n648,n649,n650,n651);
nand (n649,n551,n605);
nand (n650,n643,n605);
nand (n651,n551,n643);
xor (n652,n653,n742);
xor (n653,n654,n711);
xor (n654,n655,n691);
xor (n655,n656,n687);
xor (n656,n657,n676);
xor (n657,n658,n662);
nand (n658,n659,n660,n661);
nand (n659,n561,n564);
nand (n660,n568,n564);
nand (n661,n561,n568);
xor (n662,n663,n672);
xor (n663,n664,n668);
xor (n664,n665,n35);
or (n665,n666,n667);
and (n666,n80,n29);
and (n667,n16,n33);
xor (n668,n669,n19);
or (n669,n670,n671);
and (n670,n125,n77);
and (n671,n53,n81);
xor (n672,n673,n42);
or (n673,n674,n675);
and (n674,n21,n231);
and (n675,n28,n234);
xor (n676,n677,n683);
xor (n677,n678,n682);
xor (n678,n679,n61);
or (n679,n680,n681);
and (n680,n65,n54);
and (n681,n117,n59);
not (n682,n561);
xor (n683,n684,n24);
or (n684,n685,n686);
and (n685,n58,n17);
and (n686,n76,n22);
nand (n687,n688,n689,n690);
nand (n688,n582,n586);
nand (n689,n601,n586);
nand (n690,n582,n601);
xor (n691,n692,n701);
xor (n692,n693,n697);
nand (n693,n694,n695,n696);
nand (n694,n588,n592);
nand (n695,n597,n592);
nand (n696,n588,n597);
nand (n697,n698,n699,n700);
nand (n698,n615,n619);
nand (n699,n623,n619);
nand (n700,n615,n623);
xor (n701,n702,n707);
xor (n702,n593,n703);
xor (n703,n704,n47);
or (n704,n705,n706);
and (n705,n32,n40);
and (n706,n221,n45);
xor (n707,n708,n107);
or (n708,n709,n710);
and (n709,n225,n101);
and (n710,n39,n105);
xor (n711,n712,n738);
xor (n712,n713,n734);
xor (n713,n714,n730);
xor (n714,n715,n720);
nand (n715,n716,n718,n719);
nand (n716,n717,n91);
xor (n717,n628,n91);
nand (n718,n631,n91);
nand (n719,n717,n631);
xor (n720,n721,n91);
xor (n721,n722,n726);
xor (n722,n723,n148);
or (n723,n724,n725);
and (n724,n44,n142);
and (n725,n89,n146);
xor (n726,n727,n91);
or (n727,n728,n729);
and (n728,n100,n153);
and (n729,n104,n157);
nand (n730,n731,n732,n733);
nand (n731,n555,n559);
nand (n732,n572,n559);
nand (n733,n555,n572);
nand (n734,n735,n736,n737);
nand (n735,n613,n627);
nand (n736,n635,n627);
nand (n737,n613,n635);
nand (n738,n739,n740,n741);
nand (n739,n553,n576);
nand (n740,n580,n576);
nand (n741,n553,n580);
nand (n742,n743,n744,n745);
nand (n743,n607,n611);
nand (n744,n639,n611);
nand (n745,n607,n639);
not (n746,n747);
nand (n747,n648,n652);
nand (n748,n749,n751);
nor (n749,n750,n647);
nor (n750,n5,n549);
nand (n751,n752,n1134);
nor (n752,n753,n1128);
nor (n753,n754,n1104);
nor (n754,n755,n1102);
nor (n755,n756,n1079);
nand (n756,n757,n1051);
nand (n757,n758,n1013,n1050);
nand (n758,n759,n879);
nand (n759,n760,n817,n878);
nand (n760,n761,n805);
nand (n761,n762,n792,n804);
nand (n762,n763,n777);
xor (n763,n764,n773);
xor (n764,n765,n769);
xor (n765,n766,n61);
or (n766,n767,n768);
and (n767,n21,n54);
and (n768,n28,n59);
xor (n769,n770,n56);
or (n770,n771,n772);
and (n771,n80,n168);
and (n772,n16,n171);
xor (n773,n774,n19);
or (n774,n775,n776);
and (n775,n32,n77);
and (n776,n221,n81);
nand (n777,n778,n788,n791);
nand (n778,n779,n783);
xor (n779,n780,n19);
or (n780,n781,n782);
and (n781,n221,n77);
and (n782,n225,n81);
xor (n783,n148,n784);
xor (n784,n785,n72);
or (n785,n786,n787);
and (n786,n76,n66);
and (n787,n80,n70);
nand (n788,n789,n783);
xnor (n789,n790,n148);
nand (n790,n405,n142);
nand (n791,n779,n789);
nand (n792,n793,n777);
xor (n793,n794,n800);
xor (n794,n795,n799);
xor (n795,n796,n24);
or (n796,n797,n798);
and (n797,n225,n17);
and (n798,n39,n22);
and (n799,n148,n784);
xor (n800,n801,n35);
or (n801,n802,n803);
and (n802,n44,n29);
and (n803,n89,n33);
nand (n804,n763,n793);
xor (n805,n806,n815);
xor (n806,n807,n811);
xor (n807,n808,n148);
or (n808,n809,n810);
and (n809,n156,n142);
and (n810,n192,n146);
nand (n811,n812,n813,n814);
nand (n812,n795,n799);
nand (n813,n800,n799);
nand (n814,n795,n800);
xor (n815,n816,n425);
xor (n816,n416,n420);
nand (n817,n818,n805);
nand (n818,n819,n855,n877);
nand (n819,n820,n836);
nand (n820,n821,n830,n835);
nand (n821,n822,n826);
xor (n822,n823,n24);
or (n823,n824,n825);
and (n824,n39,n17);
and (n825,n44,n22);
xor (n826,n827,n35);
or (n827,n828,n829);
and (n828,n89,n29);
and (n829,n100,n33);
nand (n830,n831,n826);
xor (n831,n832,n42);
or (n832,n833,n834);
and (n833,n104,n231);
and (n834,n132,n234);
nand (n835,n822,n831);
xor (n836,n837,n846);
xor (n837,n838,n842);
xor (n838,n839,n42);
or (n839,n840,n841);
and (n840,n100,n231);
and (n841,n104,n234);
xor (n842,n843,n47);
or (n843,n844,n845);
and (n844,n132,n40);
and (n845,n145,n45);
xor (n846,n847,n851);
xnor (n847,n848,n68);
nor (n848,n849,n850);
and (n849,n53,n118);
and (n850,n125,n120);
xor (n851,n852,n72);
or (n852,n853,n854);
and (n853,n58,n66);
and (n854,n76,n70);
nand (n855,n856,n836);
nand (n856,n857,n871,n876);
nand (n857,n858,n862);
xor (n858,n859,n47);
or (n859,n860,n861);
and (n860,n145,n40);
and (n861,n152,n45);
and (n862,n863,n867);
xor (n863,n864,n72);
or (n864,n865,n866);
and (n865,n80,n66);
and (n866,n16,n70);
xnor (n867,n868,n68);
nor (n868,n869,n870);
and (n869,n76,n118);
and (n870,n58,n120);
nand (n871,n872,n862);
xor (n872,n873,n107);
or (n873,n874,n875);
and (n874,n156,n101);
and (n875,n192,n105);
nand (n876,n858,n872);
nand (n877,n820,n856);
nand (n878,n761,n818);
nand (n879,n880,n945,n1012);
nand (n880,n881,n893);
xor (n881,n882,n891);
xor (n882,n883,n887);
nand (n883,n884,n885,n886);
nand (n884,n765,n769);
nand (n885,n773,n769);
nand (n886,n765,n773);
nand (n887,n888,n889,n890);
nand (n888,n838,n842);
nand (n889,n846,n842);
nand (n890,n838,n846);
xor (n891,n892,n442);
xor (n892,n435,n439);
xor (n893,n894,n937);
xor (n894,n895,n923);
nand (n895,n896,n905,n922);
nand (n896,n897,n901);
xor (n897,n898,n107);
or (n898,n899,n900);
and (n899,n152,n101);
and (n900,n156,n105);
xor (n901,n902,n148);
or (n902,n903,n904);
and (n903,n192,n142);
and (n904,n405,n146);
nand (n905,n906,n901);
nand (n906,n907,n916,n921);
nand (n907,n908,n912);
xnor (n908,n909,n68);
nor (n909,n910,n911);
and (n910,n58,n118);
and (n911,n53,n120);
xor (n912,n913,n61);
or (n913,n914,n915);
and (n914,n28,n54);
and (n915,n32,n59);
nand (n916,n917,n912);
xor (n917,n918,n56);
or (n918,n919,n920);
and (n919,n16,n168);
and (n920,n21,n171);
nand (n921,n908,n917);
nand (n922,n897,n906);
xor (n923,n924,n933);
xor (n924,n925,n929);
xor (n925,n926,n35);
or (n926,n927,n928);
and (n927,n39,n29);
and (n928,n44,n33);
xor (n929,n930,n42);
or (n930,n931,n932);
and (n931,n89,n231);
and (n932,n100,n234);
xor (n933,n934,n47);
or (n934,n935,n936);
and (n935,n104,n40);
and (n936,n132,n45);
xor (n937,n938,n941);
xor (n938,n939,n940);
xor (n939,n91,n247);
and (n940,n847,n851);
xor (n941,n942,n107);
or (n942,n943,n944);
and (n943,n145,n101);
and (n944,n152,n105);
nand (n945,n946,n893);
nand (n946,n947,n989,n1011);
nand (n947,n948,n950);
xor (n948,n949,n906);
xor (n949,n897,n901);
nand (n950,n951,n971,n988);
nand (n951,n952,n969);
nand (n952,n953,n963,n968);
nand (n953,n954,n959);
and (n954,n955,n107);
xnor (n955,n956,n68);
nor (n956,n957,n958);
and (n957,n80,n118);
and (n958,n76,n120);
xor (n959,n960,n24);
or (n960,n961,n962);
and (n961,n44,n17);
and (n962,n89,n22);
nand (n963,n964,n959);
xor (n964,n965,n35);
or (n965,n966,n967);
and (n966,n100,n29);
and (n967,n104,n33);
nand (n968,n954,n964);
xor (n969,n970,n917);
xor (n970,n908,n912);
nand (n971,n972,n969);
nand (n972,n973,n982,n987);
nand (n973,n974,n978);
xor (n974,n975,n61);
or (n975,n976,n977);
and (n976,n32,n54);
and (n977,n221,n59);
xor (n978,n979,n56);
or (n979,n980,n981);
and (n980,n21,n168);
and (n981,n28,n171);
nand (n982,n983,n978);
xor (n983,n984,n19);
or (n984,n985,n986);
and (n985,n225,n77);
and (n986,n39,n81);
nand (n987,n974,n983);
nand (n988,n952,n972);
nand (n989,n990,n950);
nand (n990,n991,n1007,n1010);
nand (n991,n992,n1005);
nand (n992,n993,n1002,n1004);
nand (n993,n994,n998);
xor (n994,n995,n42);
or (n995,n996,n997);
and (n996,n132,n231);
and (n997,n145,n234);
xor (n998,n999,n47);
or (n999,n1000,n1001);
and (n1000,n152,n40);
and (n1001,n156,n45);
nand (n1002,n1003,n998);
xor (n1003,n863,n867);
nand (n1004,n994,n1003);
xor (n1005,n1006,n789);
xor (n1006,n779,n783);
nand (n1007,n1008,n1005);
xor (n1008,n1009,n831);
xor (n1009,n822,n826);
nand (n1010,n992,n1008);
nand (n1011,n948,n990);
nand (n1012,n881,n946);
nand (n1013,n1014,n879);
xor (n1014,n1015,n1038);
xor (n1015,n1016,n1028);
xor (n1016,n1017,n1024);
xor (n1017,n1018,n1022);
nand (n1018,n1019,n1020,n1021);
nand (n1019,n925,n929);
nand (n1020,n933,n929);
nand (n1021,n925,n933);
xor (n1022,n1023,n228);
xor (n1023,n217,n222);
nand (n1024,n1025,n1026,n1027);
nand (n1025,n939,n940);
nand (n1026,n941,n940);
nand (n1027,n939,n941);
xor (n1028,n1029,n1036);
xor (n1029,n1030,n1032);
xor (n1030,n1031,n246);
xor (n1031,n240,n244);
nand (n1032,n1033,n1034,n1035);
nand (n1033,n807,n811);
nand (n1034,n815,n811);
nand (n1035,n807,n815);
xor (n1036,n1037,n407);
xor (n1037,n397,n401);
xor (n1038,n1039,n1046);
xor (n1039,n1040,n1042);
xor (n1040,n1041,n433);
xor (n1041,n414,n430);
nand (n1042,n1043,n1044,n1045);
nand (n1043,n883,n887);
nand (n1044,n891,n887);
nand (n1045,n883,n891);
nand (n1046,n1047,n1048,n1049);
nand (n1047,n895,n923);
nand (n1048,n937,n923);
nand (n1049,n895,n937);
nand (n1050,n759,n1014);
xor (n1051,n1052,n1075);
xor (n1052,n1053,n1065);
xor (n1053,n1054,n1061);
xor (n1054,n1055,n1057);
xor (n1055,n1056,n238);
xor (n1056,n213,n215);
nand (n1057,n1058,n1059,n1060);
nand (n1058,n1018,n1022);
nand (n1059,n1024,n1022);
nand (n1060,n1018,n1024);
nand (n1061,n1062,n1063,n1064);
nand (n1062,n1030,n1032);
nand (n1063,n1036,n1032);
nand (n1064,n1030,n1036);
xor (n1065,n1066,n1071);
xor (n1066,n1067,n1069);
xor (n1067,n1068,n387);
xor (n1068,n382,n384);
xor (n1069,n1070,n449);
xor (n1070,n395,n412);
nand (n1071,n1072,n1073,n1074);
nand (n1072,n1040,n1042);
nand (n1073,n1046,n1042);
nand (n1074,n1040,n1046);
nand (n1075,n1076,n1077,n1078);
nand (n1076,n1016,n1028);
nand (n1077,n1038,n1028);
nand (n1078,n1016,n1038);
nor (n1079,n1080,n1084);
nand (n1080,n1081,n1082,n1083);
nand (n1081,n1053,n1065);
nand (n1082,n1075,n1065);
nand (n1083,n1053,n1075);
xor (n1084,n1085,n1094);
xor (n1085,n1086,n1090);
nand (n1086,n1087,n1088,n1089);
nand (n1087,n1055,n1057);
nand (n1088,n1061,n1057);
nand (n1089,n1055,n1061);
nand (n1090,n1091,n1092,n1093);
nand (n1091,n1067,n1069);
nand (n1092,n1071,n1069);
nand (n1093,n1067,n1071);
xor (n1094,n1095,n1100);
xor (n1095,n1096,n1098);
xor (n1096,n1097,n137);
xor (n1097,n111,n134);
xor (n1098,n1099,n254);
xor (n1099,n182,n211);
xor (n1100,n1101,n393);
xor (n1101,n380,n390);
not (n1102,n1103);
nand (n1103,n1080,n1084);
not (n1104,n1105);
nor (n1105,n1106,n1121);
nor (n1106,n1107,n1111);
nand (n1107,n1108,n1109,n1110);
nand (n1108,n1086,n1090);
nand (n1109,n1094,n1090);
nand (n1110,n1086,n1094);
xor (n1111,n1112,n1117);
xor (n1112,n1113,n1115);
xor (n1113,n1114,n180);
xor (n1114,n9,n109);
xor (n1115,n1116,n378);
xor (n1116,n285,n310);
nand (n1117,n1118,n1119,n1120);
nand (n1118,n1096,n1098);
nand (n1119,n1100,n1098);
nand (n1120,n1096,n1100);
nor (n1121,n1122,n1126);
nand (n1122,n1123,n1124,n1125);
nand (n1123,n1113,n1115);
nand (n1124,n1117,n1115);
nand (n1125,n1113,n1117);
xor (n1126,n1127,n455);
xor (n1127,n7,n283);
not (n1128,n1129);
nor (n1129,n1130,n1132);
nor (n1130,n1131,n1121);
nand (n1131,n1107,n1111);
not (n1132,n1133);
nand (n1133,n1122,n1126);
nand (n1134,n1135,n2145);
nand (n1135,n1136,n1721);
nor (n1136,n1137,n1706);
nor (n1137,n1138,n1427);
nand (n1138,n1139,n1404);
nor (n1139,n1140,n1381);
nor (n1140,n1141,n1353);
nand (n1141,n1142,n1281,n1352);
nand (n1142,n1143,n1183);
xor (n1143,n1144,n1171);
xor (n1144,n1145,n1147);
xor (n1145,n1146,n1003);
xor (n1146,n994,n998);
nand (n1147,n1148,n1157,n1170);
nand (n1148,n1149,n1153);
xor (n1149,n1150,n42);
or (n1150,n1151,n1152);
and (n1151,n145,n231);
and (n1152,n152,n234);
xor (n1153,n1154,n47);
or (n1154,n1155,n1156);
and (n1155,n156,n40);
and (n1156,n192,n45);
nand (n1157,n1158,n1153);
xor (n1158,n1159,n1168);
xor (n1159,n1160,n1164);
xor (n1160,n1161,n72);
or (n1161,n1162,n1163);
and (n1162,n16,n66);
and (n1163,n21,n70);
xor (n1164,n1165,n61);
or (n1165,n1166,n1167);
and (n1166,n221,n54);
and (n1167,n225,n59);
xnor (n1168,n1169,n107);
nand (n1169,n405,n101);
nand (n1170,n1149,n1158);
xor (n1171,n1172,n1181);
xor (n1172,n1173,n1177);
xor (n1173,n1174,n107);
or (n1174,n1175,n1176);
and (n1175,n192,n101);
and (n1176,n405,n105);
nand (n1177,n1178,n1179,n1180);
nand (n1178,n1160,n1164);
nand (n1179,n1168,n1164);
nand (n1180,n1160,n1168);
xor (n1181,n1182,n983);
xor (n1182,n974,n978);
nand (n1183,n1184,n1238,n1280);
nand (n1184,n1185,n1187);
xor (n1185,n1186,n1158);
xor (n1186,n1149,n1153);
xor (n1187,n1188,n1227);
xor (n1188,n1189,n1205);
nand (n1189,n1190,n1199,n1204);
nand (n1190,n1191,n1195);
xor (n1191,n1192,n61);
or (n1192,n1193,n1194);
and (n1193,n225,n54);
and (n1194,n39,n59);
xor (n1195,n1196,n56);
or (n1196,n1197,n1198);
and (n1197,n32,n168);
and (n1198,n221,n171);
nand (n1199,n1200,n1195);
xor (n1200,n1201,n19);
or (n1201,n1202,n1203);
and (n1202,n44,n77);
and (n1203,n89,n81);
nand (n1204,n1191,n1200);
nand (n1205,n1206,n1221,n1226);
nand (n1206,n1207,n1216);
xor (n1207,n1208,n1212);
xnor (n1208,n1209,n68);
nor (n1209,n1210,n1211);
and (n1210,n16,n118);
and (n1211,n80,n120);
xor (n1212,n1213,n72);
or (n1213,n1214,n1215);
and (n1214,n21,n66);
and (n1215,n28,n70);
and (n1216,n1217,n47);
xnor (n1217,n1218,n68);
nor (n1218,n1219,n1220);
and (n1219,n21,n118);
and (n1220,n16,n120);
nand (n1221,n1222,n1216);
xor (n1222,n1223,n24);
or (n1223,n1224,n1225);
and (n1224,n100,n17);
and (n1225,n104,n22);
nand (n1226,n1207,n1222);
xor (n1227,n1228,n1234);
xor (n1228,n1229,n1233);
xor (n1229,n1230,n24);
or (n1230,n1231,n1232);
and (n1231,n89,n17);
and (n1232,n100,n22);
and (n1233,n1208,n1212);
xor (n1234,n1235,n35);
or (n1235,n1236,n1237);
and (n1236,n104,n29);
and (n1237,n132,n33);
nand (n1238,n1239,n1187);
nand (n1239,n1240,n1264,n1279);
nand (n1240,n1241,n1262);
nand (n1241,n1242,n1256,n1261);
nand (n1242,n1243,n1252);
and (n1243,n1244,n1248);
xnor (n1244,n1245,n68);
nor (n1245,n1246,n1247);
and (n1246,n28,n118);
and (n1247,n21,n120);
xor (n1248,n1249,n72);
or (n1249,n1250,n1251);
and (n1250,n32,n66);
and (n1251,n221,n70);
xor (n1252,n1253,n24);
or (n1253,n1254,n1255);
and (n1254,n104,n17);
and (n1255,n132,n22);
nand (n1256,n1257,n1252);
xor (n1257,n1258,n35);
or (n1258,n1259,n1260);
and (n1259,n145,n29);
and (n1260,n152,n33);
nand (n1261,n1243,n1257);
xor (n1262,n1263,n1222);
xor (n1263,n1207,n1216);
nand (n1264,n1265,n1262);
xor (n1265,n1266,n1275);
xor (n1266,n1267,n1271);
xor (n1267,n1268,n35);
or (n1268,n1269,n1270);
and (n1269,n132,n29);
and (n1270,n145,n33);
xor (n1271,n1272,n42);
or (n1272,n1273,n1274);
and (n1273,n152,n231);
and (n1274,n156,n234);
xor (n1275,n1276,n47);
or (n1276,n1277,n1278);
and (n1277,n192,n40);
and (n1278,n405,n45);
nand (n1279,n1241,n1265);
nand (n1280,n1185,n1239);
nand (n1281,n1282,n1183);
xor (n1282,n1283,n1309);
xor (n1283,n1284,n1288);
nand (n1284,n1285,n1286,n1287);
nand (n1285,n1189,n1205);
nand (n1286,n1227,n1205);
nand (n1287,n1189,n1227);
xor (n1288,n1289,n1307);
xor (n1289,n1290,n1303);
nand (n1290,n1291,n1297,n1302);
nand (n1291,n1292,n1296);
xor (n1292,n1293,n56);
or (n1293,n1294,n1295);
and (n1294,n28,n168);
and (n1295,n32,n171);
xor (n1296,n955,n107);
nand (n1297,n1298,n1296);
xor (n1298,n1299,n19);
or (n1299,n1300,n1301);
and (n1300,n39,n77);
and (n1301,n44,n81);
nand (n1302,n1292,n1298);
nand (n1303,n1304,n1305,n1306);
nand (n1304,n1229,n1233);
nand (n1305,n1234,n1233);
nand (n1306,n1229,n1234);
xor (n1307,n1308,n964);
xor (n1308,n954,n959);
nand (n1309,n1310,n1317,n1351);
nand (n1310,n1311,n1315);
nand (n1311,n1312,n1313,n1314);
nand (n1312,n1267,n1271);
nand (n1313,n1275,n1271);
nand (n1314,n1267,n1275);
xor (n1315,n1316,n1298);
xor (n1316,n1292,n1296);
nand (n1317,n1318,n1315);
nand (n1318,n1319,n1336,n1350);
nand (n1319,n1320,n1334);
nand (n1320,n1321,n1330,n1333);
nand (n1321,n1322,n1326);
xor (n1322,n1323,n72);
or (n1323,n1324,n1325);
and (n1324,n28,n66);
and (n1325,n32,n70);
xor (n1326,n1327,n61);
or (n1327,n1328,n1329);
and (n1328,n39,n54);
and (n1329,n44,n59);
nand (n1330,n1331,n1326);
xnor (n1331,n1332,n47);
nand (n1332,n405,n40);
nand (n1333,n1322,n1331);
xor (n1334,n1335,n1200);
xor (n1335,n1191,n1195);
nand (n1336,n1337,n1334);
nand (n1337,n1338,n1344,n1349);
nand (n1338,n1339,n1343);
xor (n1339,n1340,n56);
or (n1340,n1341,n1342);
and (n1341,n221,n168);
and (n1342,n225,n171);
xor (n1343,n1217,n47);
nand (n1344,n1345,n1343);
xor (n1345,n1346,n19);
or (n1346,n1347,n1348);
and (n1347,n89,n77);
and (n1348,n100,n81);
nand (n1349,n1339,n1345);
nand (n1350,n1320,n1337);
nand (n1351,n1311,n1318);
nand (n1352,n1143,n1282);
xor (n1353,n1354,n1377);
xor (n1354,n1355,n1367);
xor (n1355,n1356,n1363);
xor (n1356,n1357,n1359);
xor (n1357,n1358,n872);
xor (n1358,n858,n862);
nand (n1359,n1360,n1361,n1362);
nand (n1360,n1173,n1177);
nand (n1361,n1181,n1177);
nand (n1362,n1173,n1181);
nand (n1363,n1364,n1365,n1366);
nand (n1364,n1290,n1303);
nand (n1365,n1307,n1303);
nand (n1366,n1290,n1307);
xor (n1367,n1368,n1373);
xor (n1368,n1369,n1371);
xor (n1369,n1370,n972);
xor (n1370,n952,n969);
xor (n1371,n1372,n1008);
xor (n1372,n992,n1005);
nand (n1373,n1374,n1375,n1376);
nand (n1374,n1145,n1147);
nand (n1375,n1171,n1147);
nand (n1376,n1145,n1171);
nand (n1377,n1378,n1379,n1380);
nand (n1378,n1284,n1288);
nand (n1379,n1309,n1288);
nand (n1380,n1284,n1309);
nor (n1381,n1382,n1386);
nand (n1382,n1383,n1384,n1385);
nand (n1383,n1355,n1367);
nand (n1384,n1377,n1367);
nand (n1385,n1355,n1377);
xor (n1386,n1387,n1396);
xor (n1387,n1388,n1392);
nand (n1388,n1389,n1390,n1391);
nand (n1389,n1357,n1359);
nand (n1390,n1363,n1359);
nand (n1391,n1357,n1363);
nand (n1392,n1393,n1394,n1395);
nand (n1393,n1369,n1371);
nand (n1394,n1373,n1371);
nand (n1395,n1369,n1373);
xor (n1396,n1397,n1402);
xor (n1397,n1398,n1400);
xor (n1398,n1399,n793);
xor (n1399,n763,n777);
xor (n1400,n1401,n856);
xor (n1401,n820,n836);
xor (n1402,n1403,n990);
xor (n1403,n948,n950);
nor (n1404,n1405,n1420);
nor (n1405,n1406,n1410);
nand (n1406,n1407,n1408,n1409);
nand (n1407,n1388,n1392);
nand (n1408,n1396,n1392);
nand (n1409,n1388,n1396);
xor (n1410,n1411,n1416);
xor (n1411,n1412,n1414);
xor (n1412,n1413,n818);
xor (n1413,n761,n805);
xor (n1414,n1415,n946);
xor (n1415,n881,n893);
nand (n1416,n1417,n1418,n1419);
nand (n1417,n1398,n1400);
nand (n1418,n1402,n1400);
nand (n1419,n1398,n1402);
nor (n1420,n1421,n1425);
nand (n1421,n1422,n1423,n1424);
nand (n1422,n1412,n1414);
nand (n1423,n1416,n1414);
nand (n1424,n1412,n1416);
xor (n1425,n1426,n1014);
xor (n1426,n759,n879);
nor (n1427,n1428,n1700);
nor (n1428,n1429,n1676);
nor (n1429,n1430,n1674);
nor (n1430,n1431,n1649);
nand (n1431,n1432,n1611);
nand (n1432,n1433,n1558,n1610);
nand (n1433,n1434,n1485);
xor (n1434,n1435,n1472);
xor (n1435,n1436,n1457);
nand (n1436,n1437,n1451,n1456);
nand (n1437,n1438,n1447);
and (n1438,n1439,n1443);
xnor (n1439,n1440,n68);
nor (n1440,n1441,n1442);
and (n1441,n221,n118);
and (n1442,n32,n120);
xor (n1443,n1444,n72);
or (n1444,n1445,n1446);
and (n1445,n225,n66);
and (n1446,n39,n70);
xor (n1447,n1448,n24);
or (n1448,n1449,n1450);
and (n1449,n145,n17);
and (n1450,n152,n22);
nand (n1451,n1452,n1447);
xor (n1452,n1453,n35);
or (n1453,n1454,n1455);
and (n1454,n156,n29);
and (n1455,n192,n33);
nand (n1456,n1438,n1452);
xor (n1457,n1458,n1467);
xor (n1458,n1459,n1463);
xor (n1459,n1460,n61);
or (n1460,n1461,n1462);
and (n1461,n44,n54);
and (n1462,n89,n59);
xor (n1463,n1464,n56);
or (n1464,n1465,n1466);
and (n1465,n225,n168);
and (n1466,n39,n171);
and (n1467,n1468,n42);
xnor (n1468,n1469,n68);
nor (n1469,n1470,n1471);
and (n1470,n32,n118);
and (n1471,n28,n120);
nand (n1472,n1473,n1479,n1484);
nand (n1473,n1474,n1478);
xor (n1474,n1475,n56);
or (n1475,n1476,n1477);
and (n1476,n39,n168);
and (n1477,n44,n171);
xor (n1478,n1468,n42);
nand (n1479,n1480,n1478);
xor (n1480,n1481,n19);
or (n1481,n1482,n1483);
and (n1482,n104,n77);
and (n1483,n132,n81);
nand (n1484,n1474,n1480);
xor (n1485,n1486,n1522);
xor (n1486,n1487,n1498);
xor (n1487,n1488,n1494);
xor (n1488,n1489,n1493);
xor (n1489,n1490,n19);
or (n1490,n1491,n1492);
and (n1491,n100,n77);
and (n1492,n104,n81);
xor (n1493,n1244,n1248);
xor (n1494,n1495,n24);
or (n1495,n1496,n1497);
and (n1496,n132,n17);
and (n1497,n145,n22);
xor (n1498,n1499,n1508);
xor (n1499,n1500,n1504);
xor (n1500,n1501,n35);
or (n1501,n1502,n1503);
and (n1502,n152,n29);
and (n1503,n156,n33);
xor (n1504,n1505,n42);
or (n1505,n1506,n1507);
and (n1506,n192,n231);
and (n1507,n405,n234);
nand (n1508,n1509,n1516,n1521);
nand (n1509,n1510,n1514);
xor (n1510,n1511,n72);
or (n1511,n1512,n1513);
and (n1512,n221,n66);
and (n1513,n225,n70);
xnor (n1514,n1515,n42);
nand (n1515,n405,n231);
nand (n1516,n1517,n1514);
xor (n1517,n1518,n61);
or (n1518,n1519,n1520);
and (n1519,n89,n54);
and (n1520,n100,n59);
nand (n1521,n1510,n1517);
nand (n1522,n1523,n1543,n1557);
nand (n1523,n1524,n1526);
xor (n1524,n1525,n1517);
xor (n1525,n1510,n1514);
nand (n1526,n1527,n1536,n1542);
nand (n1527,n1528,n1532);
xor (n1528,n1529,n61);
or (n1529,n1530,n1531);
and (n1530,n100,n54);
and (n1531,n104,n59);
xor (n1532,n1533,n56);
or (n1533,n1534,n1535);
and (n1534,n44,n168);
and (n1535,n89,n171);
nand (n1536,n1537,n1532);
and (n1537,n1538,n35);
xnor (n1538,n1539,n68);
nor (n1539,n1540,n1541);
and (n1540,n225,n118);
and (n1541,n221,n120);
nand (n1542,n1528,n1537);
nand (n1543,n1544,n1526);
nand (n1544,n1545,n1551,n1556);
nand (n1545,n1546,n1550);
xor (n1546,n1547,n19);
or (n1547,n1548,n1549);
and (n1548,n132,n77);
and (n1549,n145,n81);
xor (n1550,n1439,n1443);
nand (n1551,n1552,n1550);
xor (n1552,n1553,n24);
or (n1553,n1554,n1555);
and (n1554,n152,n17);
and (n1555,n156,n22);
nand (n1556,n1546,n1552);
nand (n1557,n1524,n1544);
nand (n1558,n1559,n1485);
nand (n1559,n1560,n1565,n1609);
nand (n1560,n1561,n1563);
xor (n1561,n1562,n1452);
xor (n1562,n1438,n1447);
xor (n1563,n1564,n1480);
xor (n1564,n1474,n1478);
nand (n1565,n1566,n1563);
nand (n1566,n1567,n1586,n1608);
nand (n1567,n1568,n1572);
xor (n1568,n1569,n35);
or (n1569,n1570,n1571);
and (n1570,n192,n29);
and (n1571,n405,n33);
nand (n1572,n1573,n1580,n1585);
nand (n1573,n1574,n1578);
xor (n1574,n1575,n72);
or (n1575,n1576,n1577);
and (n1576,n39,n66);
and (n1577,n44,n70);
xnor (n1578,n1579,n35);
nand (n1579,n405,n29);
nand (n1580,n1581,n1578);
xor (n1581,n1582,n61);
or (n1582,n1583,n1584);
and (n1583,n104,n54);
and (n1584,n132,n59);
nand (n1585,n1574,n1581);
nand (n1586,n1587,n1572);
nand (n1587,n1588,n1602,n1607);
nand (n1588,n1589,n1593);
xor (n1589,n1590,n56);
or (n1590,n1591,n1592);
and (n1591,n89,n168);
and (n1592,n100,n171);
and (n1593,n1594,n1598);
xnor (n1594,n1595,n68);
nor (n1595,n1596,n1597);
and (n1596,n39,n118);
and (n1597,n225,n120);
xor (n1598,n1599,n72);
or (n1599,n1600,n1601);
and (n1600,n44,n66);
and (n1601,n89,n70);
nand (n1602,n1603,n1593);
xor (n1603,n1604,n19);
or (n1604,n1605,n1606);
and (n1605,n145,n77);
and (n1606,n152,n81);
nand (n1607,n1589,n1603);
nand (n1608,n1568,n1587);
nand (n1609,n1561,n1566);
nand (n1610,n1434,n1559);
xor (n1611,n1612,n1627);
xor (n1612,n1613,n1623);
xor (n1613,n1614,n1621);
xor (n1614,n1615,n1619);
nand (n1615,n1616,n1617,n1618);
nand (n1616,n1459,n1463);
nand (n1617,n1467,n1463);
nand (n1618,n1459,n1467);
xor (n1619,n1620,n1257);
xor (n1620,n1243,n1252);
xor (n1621,n1622,n1345);
xor (n1622,n1339,n1343);
nand (n1623,n1624,n1625,n1626);
nand (n1624,n1487,n1498);
nand (n1625,n1522,n1498);
nand (n1626,n1487,n1522);
xor (n1627,n1628,n1637);
xor (n1628,n1629,n1633);
nand (n1629,n1630,n1631,n1632);
nand (n1630,n1500,n1504);
nand (n1631,n1508,n1504);
nand (n1632,n1500,n1508);
nand (n1633,n1634,n1635,n1636);
nand (n1634,n1436,n1457);
nand (n1635,n1472,n1457);
nand (n1636,n1436,n1472);
xor (n1637,n1638,n1647);
xor (n1638,n1639,n1643);
xor (n1639,n1640,n42);
or (n1640,n1641,n1642);
and (n1641,n156,n231);
and (n1642,n192,n234);
nand (n1643,n1644,n1645,n1646);
nand (n1644,n1489,n1493);
nand (n1645,n1494,n1493);
nand (n1646,n1489,n1494);
xor (n1647,n1648,n1331);
xor (n1648,n1322,n1326);
nor (n1649,n1650,n1654);
nand (n1650,n1651,n1652,n1653);
nand (n1651,n1613,n1623);
nand (n1652,n1627,n1623);
nand (n1653,n1613,n1627);
xor (n1654,n1655,n1662);
xor (n1655,n1656,n1658);
xor (n1656,n1657,n1265);
xor (n1657,n1241,n1262);
nand (n1658,n1659,n1660,n1661);
nand (n1659,n1629,n1633);
nand (n1660,n1637,n1633);
nand (n1661,n1629,n1637);
xor (n1662,n1663,n1672);
xor (n1663,n1664,n1668);
nand (n1664,n1665,n1666,n1667);
nand (n1665,n1639,n1643);
nand (n1666,n1647,n1643);
nand (n1667,n1639,n1647);
nand (n1668,n1669,n1670,n1671);
nand (n1669,n1615,n1619);
nand (n1670,n1621,n1619);
nand (n1671,n1615,n1621);
xor (n1672,n1673,n1337);
xor (n1673,n1320,n1334);
not (n1674,n1675);
nand (n1675,n1650,n1654);
not (n1676,n1677);
nor (n1677,n1678,n1693);
nor (n1678,n1679,n1683);
nand (n1679,n1680,n1681,n1682);
nand (n1680,n1656,n1658);
nand (n1681,n1662,n1658);
nand (n1682,n1656,n1662);
xor (n1683,n1684,n1691);
xor (n1684,n1685,n1687);
xor (n1685,n1686,n1318);
xor (n1686,n1311,n1315);
nand (n1687,n1688,n1689,n1690);
nand (n1688,n1664,n1668);
nand (n1689,n1672,n1668);
nand (n1690,n1664,n1672);
xor (n1691,n1692,n1239);
xor (n1692,n1185,n1187);
nor (n1693,n1694,n1698);
nand (n1694,n1695,n1696,n1697);
nand (n1695,n1685,n1687);
nand (n1696,n1691,n1687);
nand (n1697,n1685,n1691);
xor (n1698,n1699,n1282);
xor (n1699,n1143,n1183);
not (n1700,n1701);
nor (n1701,n1702,n1704);
nor (n1702,n1703,n1693);
nand (n1703,n1679,n1683);
not (n1704,n1705);
nand (n1705,n1694,n1698);
not (n1706,n1707);
nor (n1707,n1708,n1715);
nor (n1708,n1709,n1714);
nor (n1709,n1710,n1712);
nor (n1710,n1711,n1381);
nand (n1711,n1141,n1353);
not (n1712,n1713);
nand (n1713,n1382,n1386);
not (n1714,n1404);
not (n1715,n1716);
nor (n1716,n1717,n1719);
nor (n1717,n1718,n1420);
nand (n1718,n1406,n1410);
not (n1719,n1720);
nand (n1720,n1421,n1425);
nand (n1721,n1722,n1726);
nor (n1722,n1723,n1138);
nand (n1723,n1724,n1677);
nor (n1724,n1725,n1649);
nor (n1725,n1432,n1611);
nand (n1726,n1727,n2038);
nor (n1727,n1728,n2023);
nor (n1728,n1729,n1894);
nand (n1729,n1730,n1871);
nor (n1730,n1731,n1848);
nor (n1731,n1732,n1821);
nand (n1732,n1733,n1778,n1820);
nand (n1733,n1734,n1746);
xor (n1734,n1735,n1741);
xor (n1735,n1736,n1737);
xor (n1736,n1594,n1598);
xor (n1737,n1738,n24);
or (n1738,n1739,n1740);
and (n1739,n192,n17);
and (n1740,n405,n22);
and (n1741,n24,n1742);
xor (n1742,n1743,n72);
or (n1743,n1744,n1745);
and (n1744,n89,n66);
and (n1745,n100,n70);
nand (n1746,n1747,n1764,n1777);
nand (n1747,n1748,n1749);
xor (n1748,n24,n1742);
nand (n1749,n1750,n1759,n1763);
nand (n1750,n1751,n1755);
xor (n1751,n1752,n61);
or (n1752,n1753,n1754);
and (n1753,n152,n54);
and (n1754,n156,n59);
xor (n1755,n1756,n56);
or (n1756,n1757,n1758);
and (n1757,n132,n168);
and (n1758,n145,n171);
nand (n1759,n1760,n1755);
and (n1760,n19,n1761);
xnor (n1761,n1762,n19);
nand (n1762,n405,n77);
nand (n1763,n1751,n1760);
nand (n1764,n1765,n1749);
xor (n1765,n1766,n1773);
xor (n1766,n1767,n1771);
xnor (n1767,n1768,n68);
nor (n1768,n1769,n1770);
and (n1769,n44,n118);
and (n1770,n39,n120);
xnor (n1771,n1772,n24);
nand (n1772,n405,n17);
xor (n1773,n1774,n61);
or (n1774,n1775,n1776);
and (n1775,n145,n54);
and (n1776,n152,n59);
nand (n1777,n1748,n1765);
nand (n1778,n1779,n1746);
xor (n1779,n1780,n1799);
xor (n1780,n1781,n1785);
nand (n1781,n1782,n1783,n1784);
nand (n1782,n1767,n1771);
nand (n1783,n1773,n1771);
nand (n1784,n1767,n1773);
xor (n1785,n1786,n1795);
xor (n1786,n1787,n1791);
xor (n1787,n1788,n61);
or (n1788,n1789,n1790);
and (n1789,n132,n54);
and (n1790,n145,n59);
xor (n1791,n1792,n56);
or (n1792,n1793,n1794);
and (n1793,n100,n168);
and (n1794,n104,n171);
xor (n1795,n1796,n19);
or (n1796,n1797,n1798);
and (n1797,n152,n77);
and (n1798,n156,n81);
nand (n1799,n1800,n1814,n1819);
nand (n1800,n1801,n1805);
xor (n1801,n1802,n56);
or (n1802,n1803,n1804);
and (n1803,n104,n168);
and (n1804,n132,n171);
and (n1805,n1806,n1810);
xnor (n1806,n1807,n68);
nor (n1807,n1808,n1809);
and (n1808,n89,n118);
and (n1809,n44,n120);
xor (n1810,n1811,n72);
or (n1811,n1812,n1813);
and (n1812,n100,n66);
and (n1813,n104,n70);
nand (n1814,n1815,n1805);
xor (n1815,n1816,n19);
or (n1816,n1817,n1818);
and (n1817,n156,n77);
and (n1818,n192,n81);
nand (n1819,n1801,n1815);
nand (n1820,n1734,n1779);
xor (n1821,n1822,n1836);
xor (n1822,n1823,n1832);
xor (n1823,n1824,n1830);
xor (n1824,n1825,n1829);
xor (n1825,n1826,n24);
or (n1826,n1827,n1828);
and (n1827,n156,n17);
and (n1828,n192,n22);
xor (n1829,n1538,n35);
xor (n1830,n1831,n1581);
xor (n1831,n1574,n1578);
nand (n1832,n1833,n1834,n1835);
nand (n1833,n1781,n1785);
nand (n1834,n1799,n1785);
nand (n1835,n1781,n1799);
xor (n1836,n1837,n1846);
xor (n1837,n1838,n1842);
nand (n1838,n1839,n1840,n1841);
nand (n1839,n1736,n1737);
nand (n1840,n1741,n1737);
nand (n1841,n1736,n1741);
nand (n1842,n1843,n1844,n1845);
nand (n1843,n1787,n1791);
nand (n1844,n1795,n1791);
nand (n1845,n1787,n1795);
xor (n1846,n1847,n1603);
xor (n1847,n1589,n1593);
nor (n1848,n1849,n1853);
nand (n1849,n1850,n1851,n1852);
nand (n1850,n1823,n1832);
nand (n1851,n1836,n1832);
nand (n1852,n1823,n1836);
xor (n1853,n1854,n1861);
xor (n1854,n1855,n1857);
xor (n1855,n1856,n1587);
xor (n1856,n1568,n1572);
nand (n1857,n1858,n1859,n1860);
nand (n1858,n1838,n1842);
nand (n1859,n1846,n1842);
nand (n1860,n1838,n1846);
xor (n1861,n1862,n1867);
xor (n1862,n1863,n1865);
xor (n1863,n1864,n1537);
xor (n1864,n1528,n1532);
xor (n1865,n1866,n1552);
xor (n1866,n1546,n1550);
nand (n1867,n1868,n1869,n1870);
nand (n1868,n1825,n1829);
nand (n1869,n1830,n1829);
nand (n1870,n1825,n1830);
nor (n1871,n1872,n1887);
nor (n1872,n1873,n1877);
nand (n1873,n1874,n1875,n1876);
nand (n1874,n1855,n1857);
nand (n1875,n1861,n1857);
nand (n1876,n1855,n1861);
xor (n1877,n1878,n1885);
xor (n1878,n1879,n1881);
xor (n1879,n1880,n1544);
xor (n1880,n1524,n1526);
nand (n1881,n1882,n1883,n1884);
nand (n1882,n1863,n1865);
nand (n1883,n1867,n1865);
nand (n1884,n1863,n1867);
xor (n1885,n1886,n1566);
xor (n1886,n1561,n1563);
nor (n1887,n1888,n1892);
nand (n1888,n1889,n1890,n1891);
nand (n1889,n1879,n1881);
nand (n1890,n1885,n1881);
nand (n1891,n1879,n1885);
xor (n1892,n1893,n1559);
xor (n1893,n1434,n1485);
nor (n1894,n1895,n2017);
nor (n1895,n1896,n1993);
nor (n1896,n1897,n1990);
nor (n1897,n1898,n1966);
nand (n1898,n1899,n1938);
or (n1899,n1900,n1924,n1937);
and (n1900,n1901,n1910);
xor (n1901,n1902,n1906);
xnor (n1902,n1903,n68);
nor (n1903,n1904,n1905);
and (n1904,n104,n118);
and (n1905,n100,n120);
xnor (n1906,n1907,n72);
nor (n1907,n1908,n1909);
and (n1908,n145,n70);
and (n1909,n132,n66);
or (n1910,n1911,n1918,n1923);
and (n1911,n1912,n1914);
not (n1912,n1913);
nand (n1913,n405,n54);
xnor (n1914,n1915,n68);
nor (n1915,n1916,n1917);
and (n1916,n132,n118);
and (n1917,n104,n120);
and (n1918,n1914,n1919);
xnor (n1919,n1920,n72);
nor (n1920,n1921,n1922);
and (n1921,n152,n70);
and (n1922,n145,n66);
and (n1923,n1912,n1919);
and (n1924,n1910,n1925);
xor (n1925,n1926,n1933);
xor (n1926,n1927,n1929);
and (n1927,n61,n1928);
xnor (n1928,n1913,n61);
xnor (n1929,n1930,n56);
nor (n1930,n1931,n1932);
and (n1931,n156,n171);
and (n1932,n152,n168);
xnor (n1933,n1934,n61);
nor (n1934,n1935,n1936);
and (n1935,n405,n59);
and (n1936,n192,n54);
and (n1937,n1901,n1925);
xor (n1938,n1939,n1955);
xor (n1939,n1940,n1944);
or (n1940,n1941,n1942,n1943);
and (n1941,n1927,n1929);
and (n1942,n1929,n1933);
and (n1943,n1927,n1933);
xor (n1944,n1945,n1951);
xor (n1945,n1946,n1947);
and (n1946,n1902,n1906);
xnor (n1947,n1948,n56);
nor (n1948,n1949,n1950);
and (n1949,n152,n171);
and (n1950,n145,n168);
xnor (n1951,n1952,n61);
nor (n1952,n1953,n1954);
and (n1953,n192,n59);
and (n1954,n156,n54);
xor (n1955,n1956,n1962);
xor (n1956,n1957,n1958);
not (n1957,n1762);
xnor (n1958,n1959,n68);
nor (n1959,n1960,n1961);
and (n1960,n100,n118);
and (n1961,n89,n120);
xnor (n1962,n1963,n72);
nor (n1963,n1964,n1965);
and (n1964,n132,n70);
and (n1965,n104,n66);
nor (n1966,n1967,n1971);
or (n1967,n1968,n1969,n1970);
and (n1968,n1940,n1944);
and (n1969,n1944,n1955);
and (n1970,n1940,n1955);
xor (n1971,n1972,n1979);
xor (n1972,n1973,n1977);
or (n1973,n1974,n1975,n1976);
and (n1974,n1946,n1947);
and (n1975,n1947,n1951);
and (n1976,n1946,n1951);
xor (n1977,n1978,n1760);
xor (n1978,n1751,n1755);
xor (n1979,n1980,n1986);
xor (n1980,n1981,n1985);
xor (n1981,n1982,n19);
or (n1982,n1983,n1984);
and (n1983,n192,n77);
and (n1984,n405,n81);
xor (n1985,n1806,n1810);
or (n1986,n1987,n1988,n1989);
and (n1987,n1957,n1958);
and (n1988,n1958,n1962);
and (n1989,n1957,n1962);
not (n1990,n1991);
not (n1991,n1992);
and (n1992,n1967,n1971);
not (n1993,n1994);
nor (n1994,n1995,n2010);
nor (n1995,n1996,n2000);
nand (n1996,n1997,n1998,n1999);
nand (n1997,n1973,n1977);
nand (n1998,n1979,n1977);
nand (n1999,n1973,n1979);
xor (n2000,n2001,n2008);
xor (n2001,n2002,n2004);
xor (n2002,n2003,n1815);
xor (n2003,n1801,n1805);
nand (n2004,n2005,n2006,n2007);
nand (n2005,n1981,n1985);
nand (n2006,n1986,n1985);
nand (n2007,n1981,n1986);
xor (n2008,n2009,n1765);
xor (n2009,n1748,n1749);
nor (n2010,n2011,n2015);
nand (n2011,n2012,n2013,n2014);
nand (n2012,n2002,n2004);
nand (n2013,n2008,n2004);
nand (n2014,n2002,n2008);
xor (n2015,n2016,n1779);
xor (n2016,n1734,n1746);
not (n2017,n2018);
nor (n2018,n2019,n2021);
nor (n2019,n2020,n2010);
nand (n2020,n1996,n2000);
not (n2021,n2022);
nand (n2022,n2011,n2015);
not (n2023,n2024);
nor (n2024,n2025,n2032);
nor (n2025,n2026,n2031);
nor (n2026,n2027,n2029);
nor (n2027,n2028,n1848);
nand (n2028,n1732,n1821);
not (n2029,n2030);
nand (n2030,n1849,n1853);
not (n2031,n1871);
not (n2032,n2033);
nor (n2033,n2034,n2036);
nor (n2034,n2035,n1887);
nand (n2035,n1873,n1877);
not (n2036,n2037);
nand (n2037,n1888,n1892);
nand (n2038,n2039,n2043);
nor (n2039,n2040,n1729);
nand (n2040,n2041,n1994);
nor (n2041,n2042,n1966);
nor (n2042,n1899,n1938);
or (n2043,n2044,n2066);
and (n2044,n2045,n2047);
xor (n2045,n2046,n1925);
xor (n2046,n1901,n1910);
or (n2047,n2048,n2062,n2065);
and (n2048,n2049,n2058);
and (n2049,n2050,n2054);
xnor (n2050,n2051,n68);
nor (n2051,n2052,n2053);
and (n2052,n145,n118);
and (n2053,n132,n120);
xnor (n2054,n2055,n72);
nor (n2055,n2056,n2057);
and (n2056,n156,n70);
and (n2057,n152,n66);
xnor (n2058,n2059,n56);
nor (n2059,n2060,n2061);
and (n2060,n192,n171);
and (n2061,n156,n168);
and (n2062,n2058,n2063);
xor (n2063,n2064,n1919);
xor (n2064,n1912,n1914);
and (n2065,n2049,n2063);
and (n2066,n2067,n2068);
xor (n2067,n2045,n2047);
or (n2068,n2069,n2084);
and (n2069,n2070,n2082);
or (n2070,n2071,n2076,n2081);
and (n2071,n2072,n2073);
xor (n2072,n2050,n2054);
and (n2073,n56,n2074);
xnor (n2074,n2075,n56);
nand (n2075,n405,n168);
and (n2076,n2073,n2077);
xnor (n2077,n2078,n56);
nor (n2078,n2079,n2080);
and (n2079,n405,n171);
and (n2080,n192,n168);
and (n2081,n2072,n2077);
xor (n2082,n2083,n2063);
xor (n2083,n2049,n2058);
and (n2084,n2085,n2086);
xor (n2085,n2070,n2082);
or (n2086,n2087,n2103);
and (n2087,n2088,n2090);
xor (n2088,n2089,n2077);
xor (n2089,n2072,n2073);
or (n2090,n2091,n2097,n2102);
and (n2091,n2092,n2093);
not (n2092,n2075);
xnor (n2093,n2094,n68);
nor (n2094,n2095,n2096);
and (n2095,n152,n118);
and (n2096,n145,n120);
and (n2097,n2093,n2098);
xnor (n2098,n2099,n72);
nor (n2099,n2100,n2101);
and (n2100,n192,n70);
and (n2101,n156,n66);
and (n2102,n2092,n2098);
and (n2103,n2104,n2105);
xor (n2104,n2088,n2090);
or (n2105,n2106,n2117);
and (n2106,n2107,n2109);
xor (n2107,n2108,n2098);
xor (n2108,n2092,n2093);
and (n2109,n2110,n2113);
and (n2110,n72,n2111);
xnor (n2111,n2112,n72);
nand (n2112,n405,n66);
xnor (n2113,n2114,n68);
nor (n2114,n2115,n2116);
and (n2115,n156,n118);
and (n2116,n152,n120);
and (n2117,n2118,n2119);
xor (n2118,n2107,n2109);
or (n2119,n2120,n2126);
and (n2120,n2121,n2125);
xnor (n2121,n2122,n72);
nor (n2122,n2123,n2124);
and (n2123,n405,n70);
and (n2124,n192,n66);
xor (n2125,n2110,n2113);
and (n2126,n2127,n2128);
xor (n2127,n2121,n2125);
or (n2128,n2129,n2135);
and (n2129,n2130,n2134);
xnor (n2130,n2131,n68);
nor (n2131,n2132,n2133);
and (n2132,n192,n118);
and (n2133,n156,n120);
not (n2134,n2112);
and (n2135,n2136,n2137);
xor (n2136,n2130,n2134);
and (n2137,n2138,n2142);
xnor (n2138,n2139,n68);
nor (n2139,n2140,n2141);
and (n2140,n405,n118);
and (n2141,n192,n120);
and (n2142,n2143,n68);
xnor (n2143,n2144,n68);
nand (n2144,n405,n120);
not (n2145,n2146);
nand (n2146,n2147,n1105);
nor (n2147,n2148,n1079);
nor (n2148,n757,n1051);
nand (n2149,n2150,n2246);
not (n2150,n2151);
nor (n2151,n2152,n2156);
nand (n2152,n2153,n2154,n2155);
nand (n2153,n654,n711);
nand (n2154,n742,n711);
nand (n2155,n654,n742);
xor (n2156,n2157,n2242);
xor (n2157,n2158,n2162);
nand (n2158,n2159,n2160,n2161);
nand (n2159,n656,n687);
nand (n2160,n691,n687);
nand (n2161,n656,n691);
xor (n2162,n2163,n2208);
xor (n2163,n2164,n2204);
xor (n2164,n2165,n2184);
xor (n2165,n2166,n2170);
nand (n2166,n2167,n2168,n2169);
nand (n2167,n722,n726);
nand (n2168,n91,n726);
nand (n2169,n722,n91);
xor (n2170,n2171,n2180);
xor (n2171,n2172,n2176);
xor (n2172,n2173,n91);
or (n2173,n2174,n2175);
and (n2174,n89,n153);
and (n2175,n100,n157);
not (n2176,n2177);
xor (n2177,n2178,n61);
or (n2178,n680,n2179);
and (n2179,n65,n59);
xor (n2180,n2181,n107);
or (n2181,n2182,n2183);
and (n2182,n221,n101);
and (n2183,n225,n105);
xor (n2184,n2185,n2190);
xor (n2185,n91,n2186);
nand (n2186,n2187,n2188,n2189);
nand (n2187,n678,n682);
nand (n2188,n683,n682);
nand (n2189,n678,n683);
xor (n2190,n2191,n2200);
xor (n2191,n2192,n2196);
xor (n2192,n2193,n35);
or (n2193,n2194,n2195);
and (n2194,n76,n29);
and (n2195,n80,n33);
xor (n2196,n2197,n19);
or (n2197,n2198,n2199);
and (n2198,n117,n77);
and (n2199,n125,n81);
xor (n2200,n2201,n24);
or (n2201,n2202,n2203);
and (n2202,n53,n17);
and (n2203,n58,n22);
nand (n2204,n2205,n2206,n2207);
nand (n2205,n715,n720);
nand (n2206,n730,n720);
nand (n2207,n715,n730);
xor (n2208,n2209,n2218);
xor (n2209,n2210,n2214);
nand (n2210,n2211,n2212,n2213);
nand (n2211,n658,n662);
nand (n2212,n676,n662);
nand (n2213,n658,n676);
nand (n2214,n2215,n2216,n2217);
nand (n2215,n693,n697);
nand (n2216,n701,n697);
nand (n2217,n693,n701);
xor (n2218,n2219,n2238);
xor (n2219,n2220,n2224);
nand (n2220,n2221,n2222,n2223);
nand (n2221,n664,n668);
nand (n2222,n672,n668);
nand (n2223,n664,n672);
xor (n2224,n2225,n2234);
xor (n2225,n2226,n2230);
xor (n2226,n2227,n42);
or (n2227,n2228,n2229);
and (n2228,n16,n231);
and (n2229,n21,n234);
xor (n2230,n2231,n47);
or (n2231,n2232,n2233);
and (n2232,n28,n40);
and (n2233,n32,n45);
xor (n2234,n2235,n148);
or (n2235,n2236,n2237);
and (n2236,n39,n142);
and (n2237,n44,n146);
nand (n2238,n2239,n2240,n2241);
nand (n2239,n593,n703);
nand (n2240,n707,n703);
nand (n2241,n593,n707);
nand (n2242,n2243,n2244,n2245);
nand (n2243,n713,n734);
nand (n2244,n738,n734);
nand (n2245,n713,n738);
nand (n2246,n2152,n2156);
xor (n2247,n2248,n2534);
xor (n2248,n2249,n2411);
xor (n2249,n2250,n2375);
or (n2250,n2251,n2342,n2374);
and (n2251,n2252,n2263);
xor (n2252,n2253,n2261);
xor (n2253,n2254,n2258);
or (n2254,n2255,n2256,n2257);
and (n2255,n717,n613);
and (n2256,n613,n581);
and (n2257,n717,n581);
xor (n2258,n2259,n2260);
xor (n2259,n682,n721);
not (n2260,n688);
and (n2261,n576,n2262);
not (n2262,n553);
or (n2263,n2264,n2311,n2341);
and (n2264,n2265,n2296);
or (n2265,n2266,n2284,n2295);
and (n2266,n2267,n2276);
and (n2267,n2268,n287);
or (n2268,n2269,n2274,n2275);
and (n2269,n2270,n139);
or (n2270,n2271,n2272,n2273);
and (n2271,n333,n161);
not (n2272,n160);
and (n2273,n333,n165);
not (n2274,n303);
and (n2275,n2270,n149);
or (n2276,n2277,n2282,n2283);
and (n2277,n340,n2278);
or (n2278,n2279,n2280,n2281);
and (n2279,n333,n85);
not (n2280,n108);
and (n2281,n333,n97);
and (n2282,n2278,n312);
and (n2283,n340,n312);
and (n2284,n2276,n2285);
or (n2285,n2286,n2292,n2294);
and (n2286,n2287,n2288);
not (n2287,n10);
or (n2288,n2289,n2290,n2291);
and (n2289,n174,n329);
not (n2290,n339);
and (n2291,n174,n335);
and (n2292,n2288,n2293);
not (n2293,n307);
and (n2294,n2287,n2293);
and (n2295,n2267,n2285);
xor (n2296,n2297,n2302);
xor (n2297,n2298,n635);
or (n2298,n2299,n2300,n2301);
and (n2299,n62,n471);
not (n2300,n632);
and (n2301,n62,n475);
or (n2302,n2303,n2308,n2310);
and (n2303,n479,n2304);
or (n2304,n2305,n2306,n2307);
and (n2305,n479,n50);
not (n2306,n483);
and (n2307,n479,n73);
and (n2308,n2304,n2309);
not (n2309,n469);
and (n2310,n479,n2309);
and (n2311,n2296,n2312);
or (n2312,n2313,n2335,n2340);
and (n2313,n2314,n2316);
xor (n2314,n2315,n2309);
xor (n2315,n479,n2304);
or (n2316,n2317,n2326,n2334);
and (n2317,n2318,n2325);
or (n2318,n2319,n2321,n2324);
and (n2319,n371,n2320);
not (n2320,n359);
and (n2321,n2320,n2322);
xor (n2322,n2323,n97);
xor (n2323,n333,n85);
and (n2324,n371,n2322);
xor (n2325,n2268,n287);
and (n2326,n2325,n2327);
or (n2327,n2328,n2332,n2333);
and (n2328,n2329,n2330);
not (n2329,n374);
xor (n2330,n2331,n149);
xor (n2331,n2270,n139);
and (n2332,n2330,n255);
and (n2333,n2329,n255);
and (n2334,n2318,n2327);
and (n2335,n2316,n2336);
xor (n2336,n2337,n518);
xor (n2337,n2338,n484);
and (n2338,n11,n2339);
not (n2339,n48);
and (n2340,n2314,n2336);
and (n2341,n2265,n2312);
and (n2342,n2263,n2343);
xor (n2343,n2344,n2363);
xor (n2344,n2345,n2349);
or (n2345,n2346,n2347,n2348);
and (n2346,n2298,n635);
and (n2347,n635,n2302);
and (n2348,n2298,n2302);
xor (n2349,n2350,n2358);
xor (n2350,n2351,n691);
xor (n2351,n2352,n2357);
xor (n2352,n2353,n662);
or (n2353,n2354,n2355,n2356);
and (n2354,n682,n564);
not (n2355,n660);
and (n2356,n682,n568);
not (n2357,n676);
or (n2358,n2359,n2360,n2362);
not (n2359,n733);
and (n2360,n572,n2361);
not (n2361,n559);
and (n2362,n555,n2361);
or (n2363,n2364,n2368,n2373);
and (n2364,n2365,n2367);
xor (n2365,n2366,n581);
xor (n2366,n717,n613);
not (n2367,n552);
and (n2368,n2367,n2369);
or (n2369,n2370,n2371,n2372);
and (n2370,n2338,n484);
and (n2371,n484,n518);
and (n2372,n2338,n518);
and (n2373,n2365,n2369);
and (n2374,n2252,n2343);
xor (n2375,n2376,n2407);
xor (n2376,n2377,n2381);
or (n2377,n2378,n2379,n2380);
and (n2378,n2254,n2258);
and (n2379,n2258,n2261);
and (n2380,n2254,n2261);
xor (n2381,n2382,n2393);
xor (n2382,n2383,n2389);
xor (n2383,n2384,n2218);
xor (n2384,n2385,n2214);
or (n2385,n2386,n2387,n2388);
and (n2386,n2353,n662);
and (n2387,n662,n2357);
and (n2388,n2353,n2357);
or (n2389,n2390,n2391,n2392);
and (n2390,n2351,n691);
and (n2391,n691,n2358);
and (n2392,n2351,n2358);
xor (n2393,n2394,n2403);
xor (n2394,n2395,n2399);
or (n2395,n2396,n2397,n2398);
and (n2396,n561,n678);
not (n2397,n2189);
and (n2398,n561,n683);
xor (n2399,n2400,n2402);
xor (n2400,n2190,n2401);
not (n2401,n2170);
not (n2402,n2167);
or (n2403,n2404,n2405,n2406);
and (n2404,n682,n721);
and (n2405,n721,n2260);
and (n2406,n682,n2260);
or (n2407,n2408,n2409,n2410);
and (n2408,n2345,n2349);
and (n2409,n2349,n2363);
and (n2410,n2345,n2363);
or (n2411,n2412,n2445,n2533);
and (n2412,n2413,n2443);
or (n2413,n2414,n2439,n2442);
and (n2414,n2415,n2417);
xor (n2415,n2416,n2369);
xor (n2416,n2365,n2367);
or (n2417,n2418,n2435,n2438);
and (n2418,n2419,n2421);
xor (n2419,n2420,n2285);
xor (n2420,n2267,n2276);
or (n2421,n2422,n2427,n2434);
and (n2422,n2423,n2425);
xor (n2423,n2424,n312);
xor (n2424,n340,n2278);
xor (n2425,n2426,n2293);
xor (n2426,n2287,n2288);
and (n2427,n2425,n2428);
and (n2428,n182,n2429);
or (n2429,n2430,n2431,n2433);
not (n2430,n237);
and (n2431,n238,n2432);
not (n2432,n213);
and (n2433,n215,n2432);
and (n2434,n2423,n2428);
and (n2435,n2421,n2436);
xor (n2436,n2437,n2336);
xor (n2437,n2314,n2316);
and (n2438,n2419,n2436);
and (n2439,n2417,n2440);
xor (n2440,n2441,n2312);
xor (n2441,n2265,n2296);
and (n2442,n2415,n2440);
xor (n2443,n2444,n2343);
xor (n2444,n2252,n2263);
and (n2445,n2443,n2446);
or (n2446,n2447,n2504,n2532);
and (n2447,n2448,n2450);
xor (n2448,n2449,n2440);
xor (n2449,n2415,n2417);
or (n2450,n2451,n2483,n2503);
and (n2451,n2452,n2481);
or (n2452,n2453,n2466,n2480);
and (n2453,n2454,n2464);
or (n2454,n2455,n2462,n2463);
and (n2455,n2456,n2460);
or (n2456,n2457,n2458,n2459);
and (n2457,n92,n128);
and (n2458,n128,n382);
and (n2459,n92,n382);
xor (n2460,n2461,n2322);
xor (n2461,n371,n2320);
and (n2462,n2460,n393);
and (n2463,n2456,n393);
xor (n2464,n2465,n2327);
xor (n2465,n2318,n2325);
and (n2466,n2464,n2467);
or (n2467,n2468,n2477,n2479);
and (n2468,n2469,n2475);
or (n2469,n2470,n2471,n2474);
and (n2470,n388,n113);
and (n2471,n113,n2472);
xor (n2472,n2473,n382);
xor (n2473,n92,n128);
and (n2474,n388,n2472);
xor (n2475,n2476,n255);
xor (n2476,n2329,n2330);
and (n2477,n2475,n2478);
xor (n2478,n182,n2429);
and (n2479,n2469,n2478);
and (n2480,n2454,n2467);
xor (n2481,n2482,n2436);
xor (n2482,n2419,n2421);
and (n2483,n2481,n2484);
or (n2484,n2485,n2499,n2502);
and (n2485,n2486,n2488);
xor (n2486,n2487,n2428);
xor (n2487,n2423,n2425);
or (n2488,n2489,n2497,n2498);
and (n2489,n2490,n2492);
xor (n2490,n2491,n393);
xor (n2491,n2456,n2460);
or (n2492,n2493,n2494,n2496);
not (n2493,n1088);
and (n2494,n1061,n2495);
not (n2495,n1055);
and (n2496,n1057,n2495);
and (n2497,n2492,n1090);
and (n2498,n2490,n1090);
and (n2499,n2488,n2500);
xor (n2500,n2501,n2467);
xor (n2501,n2454,n2464);
and (n2502,n2486,n2500);
and (n2503,n2452,n2484);
and (n2504,n2450,n2505);
or (n2505,n2506,n2508);
xor (n2506,n2507,n2484);
xor (n2507,n2452,n2481);
or (n2508,n2509,n2525,n2531);
and (n2509,n2510,n2523);
or (n2510,n2511,n2519,n2522);
and (n2511,n2512,n2514);
xor (n2512,n2513,n2478);
xor (n2513,n2469,n2475);
or (n2514,n2515,n2517,n2518);
and (n2515,n2516,n1075);
not (n2516,n1053);
not (n2517,n1082);
and (n2518,n2516,n1065);
and (n2519,n2514,n2520);
xor (n2520,n2521,n1090);
xor (n2521,n2490,n2492);
and (n2522,n2512,n2520);
xor (n2523,n2524,n2500);
xor (n2524,n2486,n2488);
and (n2525,n2523,n2526);
or (n2526,n2527,n2529);
or (n2527,n757,n2528);
not (n2528,n1051);
xor (n2529,n2530,n2520);
xor (n2530,n2512,n2514);
and (n2531,n2510,n2526);
and (n2532,n2448,n2505);
and (n2533,n2413,n2446);
or (n2534,n2535,n2537);
xor (n2535,n2536,n2446);
xor (n2536,n2413,n2443);
and (n2537,n2538,n2539);
not (n2538,n2535);
and (n2539,n2540,n2542);
xor (n2540,n2541,n2505);
xor (n2541,n2448,n2450);
and (n2542,n2543,n2544);
xnor (n2543,n2506,n2508);
and (n2544,n2545,n2547);
xor (n2545,n2546,n2526);
xor (n2546,n2510,n2523);
and (n2547,n2548,n2549);
xnor (n2548,n2527,n2529);
and (n2549,n2550,n1135);
not (n2550,n2551);
nand (n2551,n2552,n756);
not (n2552,n2148);
endmodule
