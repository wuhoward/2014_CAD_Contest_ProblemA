module top (out,n4,n19,n20,n25,n29,n39,n40,n42,n43
        ,n48,n49,n53,n60,n70,n71,n79,n85,n98,n106
        ,n107,n109,n110,n144,n149,n150,n194,n244,n296,n335
        ,n383,n389,n398,n408,n414,n1030);
output out;
input n4;
input n19;
input n20;
input n25;
input n29;
input n39;
input n40;
input n42;
input n43;
input n48;
input n49;
input n53;
input n60;
input n70;
input n71;
input n79;
input n85;
input n98;
input n106;
input n107;
input n109;
input n110;
input n144;
input n149;
input n150;
input n194;
input n244;
input n296;
input n335;
input n383;
input n389;
input n398;
input n408;
input n414;
input n1030;
wire n0;
wire n1;
wire n2;
wire n3;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n21;
wire n22;
wire n24;
wire n26;
wire n27;
wire n28;
wire n30;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n41;
wire n44;
wire n45;
wire n46;
wire n47;
wire n50;
wire n51;
wire n52;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n108;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n145;
wire n146;
wire n147;
wire n148;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n195;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
xnor (out,n0,n1031);
nand (n0,n1,n1030);
nand (n1,n2,n869);
or (n2,n3,n5);
not (n3,n4);
not (n5,n6);
nand (n6,n7,n868);
or (n7,n8,n257);
not (n8,n9);
nand (n9,n10,n256);
not (n10,n11);
nor (n11,n12,n208);
xor (n12,n13,n164);
xor (n13,n14,n88);
xor (n14,n15,n63);
xor (n15,n16,n31);
nor (n16,n17,n26);
nand (n17,n18,n21);
wire s0n18,s1n18,notn18;
or (n18,s0n18,s1n18);
not(notn18,n4);
and (s0n18,notn18,n19);
and (s1n18,n4,n20);
not (n21,n22);
wire s0n22,s1n22,notn22;
or (n22,s0n22,s1n22);
not(notn22,n4);
and (s0n22,notn22,1'b0);
and (s1n22,n4,n24);
and (n24,n25,n20);
nor (n26,n27,n30);
and (n27,n22,n28);
not (n28,n29);
and (n30,n21,n29);
nand (n31,n32,n57);
or (n32,n33,n51);
nand (n33,n34,n45);
not (n34,n35);
nand (n35,n36,n44);
or (n36,n37,n41);
not (n37,n38);
wire s0n38,s1n38,notn38;
or (n38,s0n38,s1n38);
not(notn38,n4);
and (s0n38,notn38,n39);
and (s1n38,n4,n40);
wire s0n41,s1n41,notn41;
or (n41,s0n41,s1n41);
not(notn41,n4);
and (s0n41,notn41,n42);
and (s1n41,n4,n43);
nand (n44,n41,n37);
nand (n45,n46,n50);
or (n46,n37,n47);
wire s0n47,s1n47,notn47;
or (n47,s0n47,s1n47);
not(notn47,n4);
and (s0n47,notn47,n48);
and (s1n47,n4,n49);
nand (n50,n47,n37);
nor (n51,n52,n55);
and (n52,n53,n54);
not (n54,n47);
and (n55,n56,n47);
not (n56,n53);
or (n57,n34,n58);
nor (n58,n59,n61);
and (n59,n54,n60);
and (n61,n47,n62);
not (n62,n60);
nand (n63,n64,n82);
or (n64,n65,n76);
nand (n65,n66,n73);
nor (n66,n67,n72);
and (n67,n68,n47);
not (n68,n69);
wire s0n69,s1n69,notn69;
or (n69,s0n69,s1n69);
not(notn69,n4);
and (s0n69,notn69,n70);
and (s1n69,n4,n71);
and (n72,n69,n54);
nand (n73,n74,n75);
or (n74,n68,n18);
nand (n75,n18,n68);
nor (n76,n77,n80);
and (n77,n78,n79);
not (n78,n18);
and (n80,n18,n81);
not (n81,n79);
or (n82,n66,n83);
nor (n83,n84,n86);
and (n84,n78,n85);
and (n86,n18,n87);
not (n87,n85);
xor (n88,n89,n137);
xor (n89,n90,n122);
not (n90,n91);
nand (n91,n92,n112);
or (n92,n93,n101);
not (n93,n94);
nand (n94,n95,n99);
or (n95,n41,n96);
not (n96,n97);
and (n97,n25,n98);
or (n99,n100,n97);
not (n100,n41);
not (n101,n102);
nand (n102,n103,n111);
or (n103,n104,n108);
not (n104,n105);
wire s0n105,s1n105,notn105;
or (n105,s0n105,s1n105);
not(notn105,n4);
and (s0n105,notn105,n106);
and (s1n105,n4,n107);
wire s0n108,s1n108,notn108;
or (n108,s0n108,s1n108);
not(notn108,n4);
and (s0n108,notn108,n109);
and (s1n108,n4,n110);
nand (n111,n108,n104);
nand (n112,n113,n118);
not (n113,n114);
nor (n114,n115,n116);
and (n115,n100,n98);
and (n116,n41,n117);
not (n117,n98);
and (n118,n119,n101);
nand (n119,n120,n121);
or (n120,n104,n41);
nand (n121,n41,n104);
or (n122,n123,n129);
nand (n123,n124,n128);
or (n124,n65,n125);
nor (n125,n126,n127);
and (n126,n78,n29);
and (n127,n18,n28);
or (n128,n66,n76);
nand (n129,n130,n136);
or (n130,n131,n132);
not (n131,n118);
not (n132,n133);
nand (n133,n134,n135);
or (n134,n41,n62);
or (n135,n100,n60);
or (n136,n101,n114);
or (n137,n138,n163);
and (n138,n139,n157);
xor (n139,n140,n146);
nor (n140,n17,n141);
nor (n141,n142,n145);
and (n142,n22,n143);
not (n143,n144);
and (n145,n21,n144);
nand (n146,n147,n153);
or (n147,n148,n151);
wire s0n148,s1n148,notn148;
or (n148,s0n148,s1n148);
not(notn148,n4);
and (s0n148,notn148,n149);
and (s1n148,n4,n150);
nor (n151,n152,n148);
not (n152,n108);
not (n153,n154);
nor (n154,n155,n156);
and (n155,n152,n97);
and (n156,n108,n96);
nand (n157,n158,n159);
or (n158,n51,n34);
or (n159,n33,n160);
nor (n160,n161,n162);
and (n161,n54,n85);
and (n162,n47,n87);
and (n163,n140,n146);
or (n164,n165,n207);
and (n165,n166,n203);
xor (n166,n167,n180);
and (n167,n168,n176);
nand (n168,n169,n174);
or (n169,n170,n171);
not (n170,n151);
nor (n171,n172,n173);
and (n172,n152,n98);
and (n173,n108,n117);
or (n174,n154,n175);
not (n175,n148);
nand (n176,n177,n179);
or (n177,n178,n131);
xor (n178,n53,n100);
nand (n179,n102,n133);
or (n180,n181,n202);
and (n181,n182,n196);
xor (n182,n183,n190);
nand (n183,n184,n189);
or (n184,n185,n65);
not (n185,n186);
nor (n186,n187,n188);
and (n187,n144,n18);
and (n188,n143,n78);
or (n189,n66,n125);
nor (n190,n17,n191);
nor (n191,n192,n195);
and (n192,n22,n193);
not (n193,n194);
and (n195,n21,n194);
nand (n196,n197,n201);
or (n197,n33,n198);
nor (n198,n199,n200);
and (n199,n54,n79);
and (n200,n47,n81);
or (n201,n34,n160);
and (n202,n183,n190);
nand (n203,n204,n122);
or (n204,n205,n206);
not (n205,n129);
not (n206,n123);
and (n207,n167,n180);
or (n208,n209,n255);
and (n209,n210,n254);
xor (n210,n211,n212);
xor (n211,n139,n157);
or (n212,n213,n253);
and (n213,n214,n229);
xor (n214,n215,n216);
xor (n215,n168,n176);
and (n216,n217,n223);
nand (n217,n218,n222);
or (n218,n170,n219);
nor (n219,n220,n221);
and (n220,n152,n60);
and (n221,n108,n62);
or (n222,n171,n175);
nand (n223,n224,n228);
or (n224,n131,n225);
nor (n225,n226,n227);
and (n226,n100,n85);
and (n227,n41,n87);
or (n228,n178,n101);
or (n229,n230,n252);
and (n230,n231,n246);
xor (n231,n232,n240);
nand (n232,n233,n238);
or (n233,n234,n65);
not (n234,n235);
nor (n235,n236,n237);
and (n236,n194,n18);
and (n237,n193,n78);
nand (n238,n239,n186);
not (n239,n66);
nor (n240,n17,n241);
nor (n241,n242,n245);
and (n242,n22,n243);
not (n243,n244);
and (n245,n21,n244);
nand (n246,n247,n251);
or (n247,n33,n248);
nor (n248,n249,n250);
and (n249,n54,n29);
and (n250,n47,n28);
or (n251,n34,n198);
and (n252,n232,n240);
and (n253,n215,n216);
xor (n254,n166,n203);
and (n255,n211,n212);
nand (n256,n12,n208);
not (n257,n258);
nand (n258,n259,n864);
or (n259,n260,n361);
not (n260,n261);
nor (n261,n262,n353);
nor (n262,n263,n346);
or (n263,n264,n345);
and (n264,n265,n305);
xor (n265,n266,n267);
xor (n266,n231,n246);
xor (n267,n268,n283);
xor (n268,n269,n270);
xor (n269,n217,n223);
and (n270,n271,n277);
nand (n271,n272,n276);
or (n272,n170,n273);
nor (n273,n274,n275);
and (n274,n152,n53);
and (n275,n108,n56);
or (n276,n219,n175);
nand (n277,n278,n282);
or (n278,n131,n279);
nor (n279,n280,n281);
and (n280,n100,n79);
and (n281,n41,n81);
or (n282,n101,n225);
or (n283,n284,n304);
and (n284,n285,n298);
xor (n285,n286,n292);
nand (n286,n287,n291);
or (n287,n288,n65);
nor (n288,n289,n290);
and (n289,n244,n78);
and (n290,n243,n18);
nand (n291,n239,n235);
nor (n292,n17,n293);
nor (n293,n294,n297);
and (n294,n22,n295);
not (n295,n296);
and (n297,n21,n296);
nand (n298,n299,n303);
or (n299,n33,n300);
nor (n300,n301,n302);
and (n301,n54,n144);
and (n302,n47,n143);
or (n303,n34,n248);
and (n304,n286,n292);
or (n305,n306,n344);
and (n306,n307,n322);
xor (n307,n308,n309);
xor (n308,n271,n277);
and (n309,n310,n316);
nand (n310,n311,n315);
or (n311,n170,n312);
nor (n312,n313,n314);
and (n313,n152,n85);
and (n314,n108,n87);
or (n315,n273,n175);
nand (n316,n317,n321);
or (n317,n131,n318);
nor (n318,n319,n320);
and (n319,n100,n29);
and (n320,n41,n28);
or (n321,n279,n101);
or (n322,n323,n343);
and (n323,n324,n337);
xor (n324,n325,n331);
nand (n325,n326,n330);
or (n326,n65,n327);
nor (n327,n328,n329);
and (n328,n78,n296);
and (n329,n18,n295);
or (n330,n66,n288);
nor (n331,n17,n332);
nor (n332,n333,n336);
and (n333,n22,n334);
not (n334,n335);
and (n336,n21,n335);
nand (n337,n338,n339);
or (n338,n300,n34);
or (n339,n33,n340);
nor (n340,n341,n342);
and (n341,n54,n194);
and (n342,n47,n193);
and (n343,n325,n331);
and (n344,n308,n309);
and (n345,n266,n267);
xor (n346,n347,n350);
xor (n347,n348,n349);
xor (n348,n182,n196);
xor (n349,n214,n229);
or (n350,n351,n352);
and (n351,n268,n283);
and (n352,n269,n270);
not (n353,n354);
nand (n354,n355,n357);
not (n355,n356);
xor (n356,n210,n254);
not (n357,n358);
or (n358,n359,n360);
and (n359,n347,n350);
and (n360,n348,n349);
not (n361,n362);
nand (n362,n363,n853,n863);
nand (n363,n364,n774);
nand (n364,n365,n629,n773);
nand (n365,n366,n582);
nand (n366,n367,n581);
or (n367,n368,n536);
nor (n368,n369,n535);
and (n369,n370,n507);
not (n370,n371);
nor (n371,n372,n467);
or (n372,n373,n466);
and (n373,n374,n437);
xor (n374,n375,n418);
or (n375,n376,n417);
and (n376,n377,n404);
xor (n377,n378,n392);
nand (n378,n379,n386);
or (n379,n380,n65);
not (n380,n381);
nand (n381,n382,n384);
or (n382,n78,n383);
or (n384,n18,n385);
not (n385,n383);
or (n386,n66,n387);
nor (n387,n388,n390);
and (n388,n389,n78);
and (n390,n391,n18);
not (n391,n389);
nand (n392,n393,n400);
or (n393,n394,n131);
not (n394,n395);
nand (n395,n396,n399);
or (n396,n41,n397);
not (n397,n398);
or (n399,n100,n398);
nand (n400,n102,n401);
nor (n401,n402,n403);
and (n402,n335,n41);
and (n403,n334,n100);
nand (n404,n405,n411);
or (n405,n33,n406);
nor (n406,n407,n409);
and (n407,n54,n408);
and (n409,n47,n410);
not (n410,n408);
or (n411,n34,n412);
nor (n412,n413,n415);
and (n413,n54,n414);
and (n415,n47,n416);
not (n416,n414);
and (n417,n378,n392);
xor (n418,n419,n431);
xor (n419,n420,n422);
and (n420,n421,n383);
not (n421,n17);
nand (n422,n423,n427);
or (n423,n170,n424);
nor (n424,n425,n426);
and (n425,n243,n108);
and (n426,n244,n152);
or (n427,n428,n175);
nor (n428,n429,n430);
and (n429,n152,n194);
and (n430,n108,n193);
nand (n431,n432,n433);
or (n432,n65,n387);
or (n433,n66,n434);
nor (n434,n435,n436);
and (n435,n408,n78);
and (n436,n410,n18);
xor (n437,n438,n452);
xor (n438,n439,n446);
nand (n439,n440,n442);
or (n440,n131,n441);
not (n441,n401);
or (n442,n101,n443);
nor (n443,n444,n445);
and (n444,n100,n296);
and (n445,n41,n295);
nand (n446,n447,n448);
or (n447,n33,n412);
or (n448,n34,n449);
nor (n449,n450,n451);
and (n450,n54,n398);
and (n451,n47,n397);
and (n452,n453,n458);
nor (n453,n454,n78);
nor (n454,n455,n457);
and (n455,n54,n456);
nand (n456,n69,n383);
and (n457,n68,n385);
nand (n458,n459,n464);
or (n459,n460,n170);
not (n460,n461);
nor (n461,n462,n463);
and (n462,n296,n108);
and (n463,n295,n152);
nand (n464,n465,n148);
not (n465,n424);
and (n466,n375,n418);
xor (n467,n468,n490);
xor (n468,n469,n487);
xor (n469,n470,n481);
xor (n470,n471,n477);
nand (n471,n472,n473);
or (n472,n434,n65);
nand (n473,n474,n239);
nor (n474,n475,n476);
and (n475,n414,n18);
and (n476,n416,n78);
nor (n477,n17,n478);
nor (n478,n479,n480);
and (n479,n22,n391);
and (n480,n21,n389);
nand (n481,n482,n483);
or (n482,n170,n428);
or (n483,n484,n175);
nor (n484,n485,n486);
and (n485,n152,n144);
and (n486,n108,n143);
or (n487,n488,n489);
and (n488,n438,n452);
and (n489,n439,n446);
xor (n490,n491,n504);
xor (n491,n492,n498);
nand (n492,n493,n494);
or (n493,n33,n449);
or (n494,n34,n495);
nor (n495,n496,n497);
and (n496,n54,n335);
and (n497,n47,n334);
nand (n498,n499,n500);
or (n499,n131,n443);
or (n500,n501,n101);
nor (n501,n502,n503);
and (n502,n100,n244);
and (n503,n41,n243);
or (n504,n505,n506);
and (n505,n419,n431);
and (n506,n420,n422);
not (n507,n508);
nand (n508,n509,n510);
xor (n509,n374,n437);
or (n510,n511,n534);
and (n511,n512,n533);
xor (n512,n513,n514);
xor (n513,n453,n458);
or (n514,n515,n532);
and (n515,n516,n525);
xor (n516,n517,n518);
and (n517,n239,n383);
nand (n518,n519,n520);
or (n519,n175,n460);
nand (n520,n521,n151);
not (n521,n522);
nor (n522,n523,n524);
and (n523,n335,n152);
and (n524,n334,n108);
nand (n525,n526,n531);
or (n526,n527,n131);
not (n527,n528);
nor (n528,n529,n530);
and (n529,n414,n41);
and (n530,n100,n416);
nand (n531,n102,n395);
and (n532,n517,n518);
xor (n533,n377,n404);
and (n534,n513,n514);
and (n535,n372,n467);
nor (n536,n537,n578);
xor (n537,n538,n575);
xor (n538,n539,n558);
xor (n539,n540,n552);
xor (n540,n541,n548);
nand (n541,n542,n544);
or (n542,n543,n65);
not (n543,n474);
nand (n544,n239,n545);
nor (n545,n546,n547);
and (n546,n398,n18);
and (n547,n397,n78);
nor (n548,n17,n549);
nor (n549,n550,n551);
and (n550,n22,n410);
and (n551,n21,n408);
nand (n552,n553,n554);
or (n553,n33,n495);
or (n554,n34,n555);
nor (n555,n556,n557);
and (n556,n54,n296);
and (n557,n47,n295);
xor (n558,n559,n572);
xor (n559,n560,n566);
nand (n560,n561,n562);
or (n561,n170,n484);
or (n562,n563,n175);
nor (n563,n564,n565);
and (n564,n152,n29);
and (n565,n108,n28);
nand (n566,n567,n568);
or (n567,n131,n501);
or (n568,n569,n101);
nor (n569,n570,n571);
and (n570,n100,n194);
and (n571,n41,n193);
or (n572,n573,n574);
and (n573,n470,n481);
and (n574,n471,n477);
or (n575,n576,n577);
and (n576,n491,n504);
and (n577,n492,n498);
or (n578,n579,n580);
and (n579,n468,n490);
and (n580,n469,n487);
nand (n581,n537,n578);
nand (n582,n583,n625);
not (n583,n584);
xor (n584,n585,n624);
xor (n585,n586,n605);
xor (n586,n587,n599);
xor (n587,n588,n595);
nand (n588,n589,n591);
or (n589,n590,n65);
not (n590,n545);
nand (n591,n239,n592);
nor (n592,n593,n594);
and (n593,n335,n18);
and (n594,n334,n78);
nor (n595,n17,n596);
nor (n596,n597,n598);
and (n597,n22,n416);
and (n598,n21,n414);
nand (n599,n600,n601);
or (n600,n33,n555);
or (n601,n34,n602);
nor (n602,n603,n604);
and (n603,n54,n244);
and (n604,n47,n243);
xor (n605,n606,n621);
xor (n606,n607,n620);
xor (n607,n608,n614);
nand (n608,n609,n610);
or (n609,n170,n563);
or (n610,n611,n175);
nor (n611,n612,n613);
and (n612,n152,n79);
and (n613,n108,n81);
nand (n614,n615,n616);
or (n615,n131,n569);
or (n616,n101,n617);
nor (n617,n618,n619);
and (n618,n100,n144);
and (n619,n41,n143);
and (n620,n560,n566);
or (n621,n622,n623);
and (n622,n540,n552);
and (n623,n541,n548);
and (n624,n559,n572);
not (n625,n626);
or (n626,n627,n628);
and (n627,n538,n575);
and (n628,n539,n558);
nand (n629,n582,n630,n772);
nor (n630,n631,n769);
nor (n631,n632,n767);
and (n632,n633,n762);
or (n633,n634,n761);
and (n634,n635,n677);
xor (n635,n636,n670);
or (n636,n637,n669);
and (n637,n638,n657);
xor (n638,n639,n646);
nand (n639,n640,n645);
or (n640,n641,n131);
not (n641,n642);
nor (n642,n643,n644);
and (n643,n410,n100);
and (n644,n408,n41);
nand (n645,n102,n528);
nand (n646,n647,n652);
or (n647,n648,n34);
not (n648,n649);
nor (n649,n650,n651);
and (n650,n389,n47);
and (n651,n391,n54);
nand (n652,n653,n654);
not (n653,n33);
nand (n654,n655,n656);
or (n655,n54,n383);
or (n656,n47,n385);
xor (n657,n658,n663);
and (n658,n659,n47);
nand (n659,n660,n662);
or (n660,n41,n661);
and (n661,n383,n38);
or (n662,n38,n383);
nand (n663,n664,n668);
or (n664,n170,n665);
nor (n665,n666,n667);
and (n666,n152,n398);
and (n667,n108,n397);
or (n668,n522,n175);
and (n669,n639,n646);
xor (n670,n671,n676);
xor (n671,n672,n675);
nand (n672,n673,n674);
or (n673,n648,n33);
or (n674,n34,n406);
and (n675,n658,n663);
xor (n676,n516,n525);
or (n677,n678,n760);
and (n678,n679,n700);
xor (n679,n680,n699);
or (n680,n681,n698);
and (n681,n682,n691);
xor (n682,n683,n684);
and (n683,n35,n383);
nand (n684,n685,n690);
or (n685,n686,n131);
not (n686,n687);
nor (n687,n688,n689);
and (n688,n389,n41);
and (n689,n391,n100);
nand (n690,n642,n102);
nand (n691,n692,n697);
or (n692,n170,n693);
not (n693,n694);
nor (n694,n695,n696);
and (n695,n416,n152);
and (n696,n414,n108);
or (n697,n665,n175);
and (n698,n683,n684);
xor (n699,n638,n657);
or (n700,n701,n759);
and (n701,n702,n758);
xor (n702,n703,n717);
nor (n703,n704,n712);
not (n704,n705);
nand (n705,n706,n711);
or (n706,n707,n170);
not (n707,n708);
nand (n708,n709,n710);
or (n709,n410,n108);
nand (n710,n108,n410);
nand (n711,n694,n148);
nand (n712,n713,n41);
nand (n713,n714,n716);
or (n714,n108,n715);
and (n715,n383,n105);
or (n716,n105,n383);
nand (n717,n718,n756);
or (n718,n719,n742);
not (n719,n720);
nand (n720,n721,n741);
or (n721,n722,n731);
nor (n722,n723,n730);
nand (n723,n724,n729);
or (n724,n725,n170);
not (n725,n726);
nand (n726,n727,n728);
or (n727,n391,n108);
nand (n728,n108,n391);
nand (n729,n708,n148);
nor (n730,n101,n385);
nand (n731,n732,n739);
nand (n732,n733,n738);
or (n733,n734,n170);
not (n734,n735);
nand (n735,n736,n737);
or (n736,n152,n383);
or (n737,n108,n385);
nand (n738,n726,n148);
nor (n739,n740,n152);
and (n740,n383,n148);
nand (n741,n723,n730);
not (n742,n743);
nand (n743,n744,n752);
not (n744,n745);
nand (n745,n746,n751);
or (n746,n747,n131);
not (n747,n748);
nand (n748,n749,n750);
or (n749,n100,n383);
or (n750,n41,n385);
nand (n751,n102,n687);
nor (n752,n753,n755);
and (n753,n704,n754);
not (n754,n712);
and (n755,n705,n712);
nand (n756,n757,n745);
not (n757,n752);
xor (n758,n682,n691);
and (n759,n703,n717);
and (n760,n680,n699);
and (n761,n636,n670);
or (n762,n763,n764);
xor (n763,n512,n533);
or (n764,n765,n766);
and (n765,n671,n676);
and (n766,n672,n675);
not (n767,n768);
nand (n768,n763,n764);
nand (n769,n770,n370);
not (n770,n771);
nor (n771,n509,n510);
not (n772,n536);
nand (n773,n584,n626);
nor (n774,n775,n832);
nand (n775,n776,n825);
not (n776,n777);
nor (n777,n778,n816);
xor (n778,n779,n807);
xor (n779,n780,n781);
xor (n780,n324,n337);
xor (n781,n782,n791);
xor (n782,n783,n784);
xor (n783,n310,n316);
and (n784,n785,n788);
nand (n785,n786,n787);
or (n786,n170,n611);
or (n787,n312,n175);
nand (n788,n789,n790);
or (n789,n131,n617);
or (n790,n318,n101);
or (n791,n792,n806);
and (n792,n793,n803);
xor (n793,n794,n799);
nand (n794,n795,n797);
or (n795,n796,n65);
not (n796,n592);
nand (n797,n798,n239);
not (n798,n327);
nor (n799,n17,n800);
nor (n800,n801,n802);
and (n801,n22,n397);
and (n802,n21,n398);
nand (n803,n804,n805);
or (n804,n33,n602);
or (n805,n34,n340);
and (n806,n794,n799);
or (n807,n808,n815);
and (n808,n809,n812);
xor (n809,n810,n811);
xor (n810,n785,n788);
and (n811,n608,n614);
or (n812,n813,n814);
and (n813,n587,n599);
and (n814,n588,n595);
and (n815,n810,n811);
or (n816,n817,n824);
and (n817,n818,n821);
xor (n818,n819,n820);
xor (n819,n793,n803);
xor (n820,n809,n812);
or (n821,n822,n823);
and (n822,n606,n621);
and (n823,n607,n620);
and (n824,n819,n820);
nand (n825,n826,n828);
not (n826,n827);
xor (n827,n818,n821);
not (n828,n829);
or (n829,n830,n831);
and (n830,n585,n624);
and (n831,n586,n605);
nand (n832,n833,n846);
nand (n833,n834,n842);
not (n834,n835);
xor (n835,n836,n839);
xor (n836,n837,n838);
xor (n837,n285,n298);
xor (n838,n307,n322);
or (n839,n840,n841);
and (n840,n782,n791);
and (n841,n783,n784);
not (n842,n843);
or (n843,n844,n845);
and (n844,n779,n807);
and (n845,n780,n781);
nand (n846,n847,n849);
not (n847,n848);
xor (n848,n265,n305);
not (n849,n850);
or (n850,n851,n852);
and (n851,n836,n839);
and (n852,n837,n838);
nand (n853,n854,n846);
nand (n854,n855,n862);
or (n855,n856,n857);
not (n856,n833);
not (n857,n858);
nand (n858,n859,n861);
or (n859,n777,n860);
nand (n860,n827,n829);
nand (n861,n778,n816);
nand (n862,n835,n843);
nand (n863,n850,n848);
nor (n864,n865,n867);
and (n865,n866,n354);
and (n866,n263,n346);
nor (n867,n355,n357);
or (n868,n258,n9);
not (n869,n870);
and (n870,n871,n3,n25);
nand (n871,n872,n1029);
or (n872,n873,n926);
not (n873,n874);
nor (n874,n875,n925);
and (n875,n876,n914);
not (n876,n877);
or (n877,n878,n913);
and (n878,n879,n894);
xor (n879,n880,n890);
nand (n880,n881,n886);
or (n881,n882,n66);
not (n882,n883);
nand (n883,n884,n885);
or (n884,n18,n96);
or (n885,n78,n97);
or (n886,n65,n887);
nor (n887,n888,n889);
and (n888,n78,n98);
and (n889,n18,n117);
nand (n890,n891,n892,n421);
or (n891,n22,n60);
not (n892,n893);
and (n893,n60,n22);
or (n894,n895,n912);
and (n895,n896,n908);
xor (n896,n897,n902);
nand (n897,n898,n899);
or (n898,n653,n35);
nand (n899,n900,n901);
or (n900,n47,n96);
or (n901,n54,n97);
nand (n902,n903,n907);
or (n903,n65,n904);
nor (n904,n905,n906);
and (n905,n78,n60);
and (n906,n18,n62);
or (n907,n66,n887);
nor (n908,n17,n909);
nor (n909,n910,n911);
and (n910,n22,n56);
and (n911,n21,n53);
and (n912,n897,n902);
and (n913,n880,n890);
not (n914,n915);
xor (n915,n916,n924);
xor (n916,n917,n920);
nand (n917,n918,n883);
or (n918,n919,n239);
not (n919,n65);
nor (n920,n17,n921);
nor (n921,n922,n923);
and (n922,n22,n117);
and (n923,n21,n98);
not (n924,n890);
and (n925,n877,n915);
nand (n926,n927,n1010,n1028);
nand (n927,n362,n928);
and (n928,n929,n966,n1005);
and (n929,n261,n930,n10);
nand (n930,n931,n962);
not (n931,n932);
xor (n932,n933,n959);
xor (n933,n934,n948);
xor (n934,n935,n944);
xor (n935,n936,n938);
nand (n936,n937,n94);
or (n937,n118,n102);
nand (n938,n939,n940);
or (n939,n33,n58);
or (n940,n34,n941);
nor (n941,n942,n943);
and (n942,n54,n98);
and (n943,n47,n117);
nor (n944,n17,n945);
nor (n945,n946,n947);
and (n946,n22,n81);
and (n947,n21,n79);
xor (n948,n949,n956);
xor (n949,n950,n91);
nand (n950,n951,n952);
or (n951,n65,n83);
or (n952,n66,n953);
nor (n953,n954,n955);
and (n954,n78,n53);
and (n955,n18,n56);
or (n956,n957,n958);
and (n957,n15,n63);
and (n958,n16,n31);
or (n959,n960,n961);
and (n960,n89,n137);
and (n961,n90,n122);
not (n962,n963);
or (n963,n964,n965);
and (n964,n13,n164);
and (n965,n14,n88);
nor (n966,n967,n992);
nor (n967,n968,n971);
or (n968,n969,n970);
and (n969,n933,n959);
and (n970,n934,n948);
xor (n971,n972,n989);
xor (n972,n973,n976);
or (n973,n974,n975);
and (n974,n935,n944);
and (n975,n936,n938);
xor (n976,n977,n985);
xor (n977,n978,n981);
nand (n978,n979,n980);
or (n979,n65,n953);
or (n980,n66,n904);
nor (n981,n17,n982);
nor (n982,n983,n984);
and (n983,n22,n87);
and (n984,n21,n85);
nor (n985,n986,n988);
and (n986,n653,n987);
not (n987,n941);
and (n988,n35,n899);
or (n989,n990,n991);
and (n990,n949,n956);
and (n991,n950,n91);
and (n992,n993,n997);
not (n993,n994);
or (n994,n995,n996);
and (n995,n972,n989);
and (n996,n973,n976);
not (n997,n998);
xor (n998,n999,n1002);
xor (n999,n1000,n1001);
not (n1000,n985);
xor (n1001,n896,n908);
or (n1002,n1003,n1004);
and (n1003,n977,n985);
and (n1004,n978,n981);
or (n1005,n1006,n1009);
or (n1006,n1007,n1008);
and (n1007,n999,n1002);
and (n1008,n1000,n1001);
xor (n1009,n879,n894);
nand (n1010,n1011,n1005);
nand (n1011,n1012,n1022);
or (n1012,n1013,n1014);
not (n1013,n966);
not (n1014,n1015);
nand (n1015,n1016,n1021);
or (n1016,n1017,n1018);
not (n1017,n930);
not (n1018,n1019);
nand (n1019,n1020,n256);
or (n1020,n864,n11);
or (n1021,n931,n962);
nor (n1022,n1023,n1027);
and (n1023,n1024,n1026);
not (n1024,n1025);
nand (n1025,n968,n971);
not (n1026,n992);
nor (n1027,n993,n997);
nand (n1028,n1006,n1009);
nand (n1029,n873,n926);
and (n1031,n1030,n1032);
wire s0n1032,s1n1032,notn1032;
or (n1032,s0n1032,s1n1032);
not(notn1032,n4);
and (s0n1032,notn1032,n1033);
and (s1n1032,n4,n2333);
and (n1033,n25,n1034);
xor (n1034,n1035,n1849);
xor (n1035,n1036,n2331);
xor (n1036,n1037,n1844);
xor (n1037,n1038,n2324);
xor (n1038,n1039,n1838);
xor (n1039,n1040,n2312);
xor (n1040,n1041,n1832);
xor (n1041,n1042,n2295);
xor (n1042,n1043,n1826);
xor (n1043,n1044,n2273);
xor (n1044,n1045,n1820);
xor (n1045,n1046,n2246);
xor (n1046,n1047,n1814);
xor (n1047,n1048,n2214);
xor (n1048,n1049,n1808);
xor (n1049,n1050,n2177);
xor (n1050,n1051,n1802);
xor (n1051,n1052,n2135);
xor (n1052,n1053,n1796);
xor (n1053,n1054,n2088);
xor (n1054,n1055,n1790);
xor (n1055,n1056,n2036);
xor (n1056,n1057,n1784);
xor (n1057,n1058,n1979);
xor (n1058,n1059,n1778);
xor (n1059,n1060,n1917);
xor (n1060,n1061,n1772);
xor (n1061,n1062,n1850);
xor (n1062,n1063,n893);
xor (n1063,n1064,n1764);
xor (n1064,n1065,n1763);
xor (n1065,n1066,n1675);
xor (n1066,n1067,n1674);
xor (n1067,n1068,n1576);
xor (n1068,n1069,n1575);
xor (n1069,n1070,n1473);
xor (n1070,n1071,n1472);
xor (n1071,n1072,n1365);
xor (n1072,n1073,n1364);
xor (n1073,n1074,n1085);
xor (n1074,n1075,n1084);
xor (n1075,n1076,n1083);
xor (n1076,n1077,n1082);
xor (n1077,n1078,n1081);
xor (n1078,n1079,n1080);
and (n1079,n97,n148);
and (n1080,n97,n108);
and (n1081,n1079,n1080);
and (n1082,n97,n105);
and (n1083,n1077,n1082);
and (n1084,n97,n41);
or (n1085,n1086,n1087);
and (n1086,n1075,n1084);
and (n1087,n1074,n1088);
or (n1088,n1086,n1089);
and (n1089,n1074,n1090);
or (n1090,n1086,n1091);
and (n1091,n1074,n1092);
or (n1092,n1086,n1093);
and (n1093,n1074,n1094);
or (n1094,n1095,n1279);
and (n1095,n1096,n1278);
xor (n1096,n1076,n1097);
or (n1097,n1098,n1190);
and (n1098,n1099,n1189);
xor (n1099,n1078,n1100);
or (n1100,n1081,n1101);
and (n1101,n1102,n1104);
xor (n1102,n1079,n1103);
and (n1103,n98,n108);
or (n1104,n1105,n1108);
and (n1105,n1106,n1107);
and (n1106,n98,n148);
and (n1107,n60,n108);
and (n1108,n1109,n1110);
xor (n1109,n1106,n1107);
or (n1110,n1111,n1114);
and (n1111,n1112,n1113);
and (n1112,n60,n148);
and (n1113,n53,n108);
and (n1114,n1115,n1116);
xor (n1115,n1112,n1113);
or (n1116,n1117,n1120);
and (n1117,n1118,n1119);
and (n1118,n53,n148);
and (n1119,n85,n108);
and (n1120,n1121,n1122);
xor (n1121,n1118,n1119);
or (n1122,n1123,n1126);
and (n1123,n1124,n1125);
and (n1124,n85,n148);
and (n1125,n79,n108);
and (n1126,n1127,n1128);
xor (n1127,n1124,n1125);
or (n1128,n1129,n1132);
and (n1129,n1130,n1131);
and (n1130,n79,n148);
and (n1131,n29,n108);
and (n1132,n1133,n1134);
xor (n1133,n1130,n1131);
or (n1134,n1135,n1138);
and (n1135,n1136,n1137);
and (n1136,n29,n148);
and (n1137,n144,n108);
and (n1138,n1139,n1140);
xor (n1139,n1136,n1137);
or (n1140,n1141,n1144);
and (n1141,n1142,n1143);
and (n1142,n144,n148);
and (n1143,n194,n108);
and (n1144,n1145,n1146);
xor (n1145,n1142,n1143);
or (n1146,n1147,n1150);
and (n1147,n1148,n1149);
and (n1148,n194,n148);
and (n1149,n244,n108);
and (n1150,n1151,n1152);
xor (n1151,n1148,n1149);
or (n1152,n1153,n1155);
and (n1153,n1154,n462);
and (n1154,n244,n148);
and (n1155,n1156,n1157);
xor (n1156,n1154,n462);
or (n1157,n1158,n1161);
and (n1158,n1159,n1160);
and (n1159,n296,n148);
and (n1160,n335,n108);
and (n1161,n1162,n1163);
xor (n1162,n1159,n1160);
or (n1163,n1164,n1167);
and (n1164,n1165,n1166);
and (n1165,n335,n148);
and (n1166,n398,n108);
and (n1167,n1168,n1169);
xor (n1168,n1165,n1166);
or (n1169,n1170,n1172);
and (n1170,n1171,n696);
and (n1171,n398,n148);
and (n1172,n1173,n1174);
xor (n1173,n1171,n696);
or (n1174,n1175,n1178);
and (n1175,n1176,n1177);
and (n1176,n414,n148);
and (n1177,n408,n108);
and (n1178,n1179,n1180);
xor (n1179,n1176,n1177);
or (n1180,n1181,n1184);
and (n1181,n1182,n1183);
and (n1182,n408,n148);
and (n1183,n389,n108);
and (n1184,n1185,n1186);
xor (n1185,n1182,n1183);
and (n1186,n1187,n1188);
and (n1187,n389,n148);
and (n1188,n383,n108);
and (n1189,n98,n105);
and (n1190,n1191,n1192);
xor (n1191,n1099,n1189);
or (n1192,n1193,n1196);
and (n1193,n1194,n1195);
xor (n1194,n1102,n1104);
and (n1195,n60,n105);
and (n1196,n1197,n1198);
xor (n1197,n1194,n1195);
or (n1198,n1199,n1202);
and (n1199,n1200,n1201);
xor (n1200,n1109,n1110);
and (n1201,n53,n105);
and (n1202,n1203,n1204);
xor (n1203,n1200,n1201);
or (n1204,n1205,n1208);
and (n1205,n1206,n1207);
xor (n1206,n1115,n1116);
and (n1207,n85,n105);
and (n1208,n1209,n1210);
xor (n1209,n1206,n1207);
or (n1210,n1211,n1214);
and (n1211,n1212,n1213);
xor (n1212,n1121,n1122);
and (n1213,n79,n105);
and (n1214,n1215,n1216);
xor (n1215,n1212,n1213);
or (n1216,n1217,n1220);
and (n1217,n1218,n1219);
xor (n1218,n1127,n1128);
and (n1219,n29,n105);
and (n1220,n1221,n1222);
xor (n1221,n1218,n1219);
or (n1222,n1223,n1226);
and (n1223,n1224,n1225);
xor (n1224,n1133,n1134);
and (n1225,n144,n105);
and (n1226,n1227,n1228);
xor (n1227,n1224,n1225);
or (n1228,n1229,n1232);
and (n1229,n1230,n1231);
xor (n1230,n1139,n1140);
and (n1231,n194,n105);
and (n1232,n1233,n1234);
xor (n1233,n1230,n1231);
or (n1234,n1235,n1238);
and (n1235,n1236,n1237);
xor (n1236,n1145,n1146);
and (n1237,n244,n105);
and (n1238,n1239,n1240);
xor (n1239,n1236,n1237);
or (n1240,n1241,n1244);
and (n1241,n1242,n1243);
xor (n1242,n1151,n1152);
and (n1243,n296,n105);
and (n1244,n1245,n1246);
xor (n1245,n1242,n1243);
or (n1246,n1247,n1250);
and (n1247,n1248,n1249);
xor (n1248,n1156,n1157);
and (n1249,n335,n105);
and (n1250,n1251,n1252);
xor (n1251,n1248,n1249);
or (n1252,n1253,n1256);
and (n1253,n1254,n1255);
xor (n1254,n1162,n1163);
and (n1255,n398,n105);
and (n1256,n1257,n1258);
xor (n1257,n1254,n1255);
or (n1258,n1259,n1262);
and (n1259,n1260,n1261);
xor (n1260,n1168,n1169);
and (n1261,n414,n105);
and (n1262,n1263,n1264);
xor (n1263,n1260,n1261);
or (n1264,n1265,n1268);
and (n1265,n1266,n1267);
xor (n1266,n1173,n1174);
and (n1267,n408,n105);
and (n1268,n1269,n1270);
xor (n1269,n1266,n1267);
or (n1270,n1271,n1274);
and (n1271,n1272,n1273);
xor (n1272,n1179,n1180);
and (n1273,n389,n105);
and (n1274,n1275,n1276);
xor (n1275,n1272,n1273);
and (n1276,n1277,n715);
xor (n1277,n1185,n1186);
and (n1278,n98,n41);
and (n1279,n1280,n1281);
xor (n1280,n1096,n1278);
or (n1281,n1282,n1285);
and (n1282,n1283,n1284);
xor (n1283,n1191,n1192);
and (n1284,n60,n41);
and (n1285,n1286,n1287);
xor (n1286,n1283,n1284);
or (n1287,n1288,n1291);
and (n1288,n1289,n1290);
xor (n1289,n1197,n1198);
and (n1290,n53,n41);
and (n1291,n1292,n1293);
xor (n1292,n1289,n1290);
or (n1293,n1294,n1297);
and (n1294,n1295,n1296);
xor (n1295,n1203,n1204);
and (n1296,n85,n41);
and (n1297,n1298,n1299);
xor (n1298,n1295,n1296);
or (n1299,n1300,n1303);
and (n1300,n1301,n1302);
xor (n1301,n1209,n1210);
and (n1302,n79,n41);
and (n1303,n1304,n1305);
xor (n1304,n1301,n1302);
or (n1305,n1306,n1309);
and (n1306,n1307,n1308);
xor (n1307,n1215,n1216);
and (n1308,n29,n41);
and (n1309,n1310,n1311);
xor (n1310,n1307,n1308);
or (n1311,n1312,n1315);
and (n1312,n1313,n1314);
xor (n1313,n1221,n1222);
and (n1314,n144,n41);
and (n1315,n1316,n1317);
xor (n1316,n1313,n1314);
or (n1317,n1318,n1321);
and (n1318,n1319,n1320);
xor (n1319,n1227,n1228);
and (n1320,n194,n41);
and (n1321,n1322,n1323);
xor (n1322,n1319,n1320);
or (n1323,n1324,n1327);
and (n1324,n1325,n1326);
xor (n1325,n1233,n1234);
and (n1326,n244,n41);
and (n1327,n1328,n1329);
xor (n1328,n1325,n1326);
or (n1329,n1330,n1333);
and (n1330,n1331,n1332);
xor (n1331,n1239,n1240);
and (n1332,n296,n41);
and (n1333,n1334,n1335);
xor (n1334,n1331,n1332);
or (n1335,n1336,n1338);
and (n1336,n1337,n402);
xor (n1337,n1245,n1246);
and (n1338,n1339,n1340);
xor (n1339,n1337,n402);
or (n1340,n1341,n1344);
and (n1341,n1342,n1343);
xor (n1342,n1251,n1252);
and (n1343,n398,n41);
and (n1344,n1345,n1346);
xor (n1345,n1342,n1343);
or (n1346,n1347,n1349);
and (n1347,n1348,n529);
xor (n1348,n1257,n1258);
and (n1349,n1350,n1351);
xor (n1350,n1348,n529);
or (n1351,n1352,n1354);
and (n1352,n1353,n644);
xor (n1353,n1263,n1264);
and (n1354,n1355,n1356);
xor (n1355,n1353,n644);
or (n1356,n1357,n1359);
and (n1357,n1358,n688);
xor (n1358,n1269,n1270);
and (n1359,n1360,n1361);
xor (n1360,n1358,n688);
and (n1361,n1362,n1363);
xor (n1362,n1275,n1276);
and (n1363,n383,n41);
and (n1364,n97,n38);
or (n1365,n1366,n1368);
and (n1366,n1367,n1364);
xor (n1367,n1074,n1088);
and (n1368,n1369,n1370);
xor (n1369,n1367,n1364);
or (n1370,n1371,n1373);
and (n1371,n1372,n1364);
xor (n1372,n1074,n1090);
and (n1373,n1374,n1375);
xor (n1374,n1372,n1364);
or (n1375,n1376,n1378);
and (n1376,n1377,n1364);
xor (n1377,n1074,n1092);
and (n1378,n1379,n1380);
xor (n1379,n1377,n1364);
or (n1380,n1381,n1384);
and (n1381,n1382,n1383);
xor (n1382,n1074,n1094);
and (n1383,n98,n38);
and (n1384,n1385,n1386);
xor (n1385,n1382,n1383);
or (n1386,n1387,n1390);
and (n1387,n1388,n1389);
xor (n1388,n1280,n1281);
and (n1389,n60,n38);
and (n1390,n1391,n1392);
xor (n1391,n1388,n1389);
or (n1392,n1393,n1396);
and (n1393,n1394,n1395);
xor (n1394,n1286,n1287);
and (n1395,n53,n38);
and (n1396,n1397,n1398);
xor (n1397,n1394,n1395);
or (n1398,n1399,n1402);
and (n1399,n1400,n1401);
xor (n1400,n1292,n1293);
and (n1401,n85,n38);
and (n1402,n1403,n1404);
xor (n1403,n1400,n1401);
or (n1404,n1405,n1408);
and (n1405,n1406,n1407);
xor (n1406,n1298,n1299);
and (n1407,n79,n38);
and (n1408,n1409,n1410);
xor (n1409,n1406,n1407);
or (n1410,n1411,n1414);
and (n1411,n1412,n1413);
xor (n1412,n1304,n1305);
and (n1413,n29,n38);
and (n1414,n1415,n1416);
xor (n1415,n1412,n1413);
or (n1416,n1417,n1420);
and (n1417,n1418,n1419);
xor (n1418,n1310,n1311);
and (n1419,n144,n38);
and (n1420,n1421,n1422);
xor (n1421,n1418,n1419);
or (n1422,n1423,n1426);
and (n1423,n1424,n1425);
xor (n1424,n1316,n1317);
and (n1425,n194,n38);
and (n1426,n1427,n1428);
xor (n1427,n1424,n1425);
or (n1428,n1429,n1432);
and (n1429,n1430,n1431);
xor (n1430,n1322,n1323);
and (n1431,n244,n38);
and (n1432,n1433,n1434);
xor (n1433,n1430,n1431);
or (n1434,n1435,n1438);
and (n1435,n1436,n1437);
xor (n1436,n1328,n1329);
and (n1437,n296,n38);
and (n1438,n1439,n1440);
xor (n1439,n1436,n1437);
or (n1440,n1441,n1444);
and (n1441,n1442,n1443);
xor (n1442,n1334,n1335);
and (n1443,n335,n38);
and (n1444,n1445,n1446);
xor (n1445,n1442,n1443);
or (n1446,n1447,n1450);
and (n1447,n1448,n1449);
xor (n1448,n1339,n1340);
and (n1449,n398,n38);
and (n1450,n1451,n1452);
xor (n1451,n1448,n1449);
or (n1452,n1453,n1456);
and (n1453,n1454,n1455);
xor (n1454,n1345,n1346);
and (n1455,n414,n38);
and (n1456,n1457,n1458);
xor (n1457,n1454,n1455);
or (n1458,n1459,n1462);
and (n1459,n1460,n1461);
xor (n1460,n1350,n1351);
and (n1461,n408,n38);
and (n1462,n1463,n1464);
xor (n1463,n1460,n1461);
or (n1464,n1465,n1468);
and (n1465,n1466,n1467);
xor (n1466,n1355,n1356);
and (n1467,n389,n38);
and (n1468,n1469,n1470);
xor (n1469,n1466,n1467);
and (n1470,n1471,n661);
xor (n1471,n1360,n1361);
and (n1472,n97,n47);
or (n1473,n1474,n1476);
and (n1474,n1475,n1472);
xor (n1475,n1369,n1370);
and (n1476,n1477,n1478);
xor (n1477,n1475,n1472);
or (n1478,n1479,n1481);
and (n1479,n1480,n1472);
xor (n1480,n1374,n1375);
and (n1481,n1482,n1483);
xor (n1482,n1480,n1472);
or (n1483,n1484,n1487);
and (n1484,n1485,n1486);
xor (n1485,n1379,n1380);
and (n1486,n98,n47);
and (n1487,n1488,n1489);
xor (n1488,n1485,n1486);
or (n1489,n1490,n1493);
and (n1490,n1491,n1492);
xor (n1491,n1385,n1386);
and (n1492,n60,n47);
and (n1493,n1494,n1495);
xor (n1494,n1491,n1492);
or (n1495,n1496,n1499);
and (n1496,n1497,n1498);
xor (n1497,n1391,n1392);
and (n1498,n53,n47);
and (n1499,n1500,n1501);
xor (n1500,n1497,n1498);
or (n1501,n1502,n1505);
and (n1502,n1503,n1504);
xor (n1503,n1397,n1398);
and (n1504,n85,n47);
and (n1505,n1506,n1507);
xor (n1506,n1503,n1504);
or (n1507,n1508,n1511);
and (n1508,n1509,n1510);
xor (n1509,n1403,n1404);
and (n1510,n79,n47);
and (n1511,n1512,n1513);
xor (n1512,n1509,n1510);
or (n1513,n1514,n1517);
and (n1514,n1515,n1516);
xor (n1515,n1409,n1410);
and (n1516,n29,n47);
and (n1517,n1518,n1519);
xor (n1518,n1515,n1516);
or (n1519,n1520,n1523);
and (n1520,n1521,n1522);
xor (n1521,n1415,n1416);
and (n1522,n144,n47);
and (n1523,n1524,n1525);
xor (n1524,n1521,n1522);
or (n1525,n1526,n1529);
and (n1526,n1527,n1528);
xor (n1527,n1421,n1422);
and (n1528,n194,n47);
and (n1529,n1530,n1531);
xor (n1530,n1527,n1528);
or (n1531,n1532,n1535);
and (n1532,n1533,n1534);
xor (n1533,n1427,n1428);
and (n1534,n244,n47);
and (n1535,n1536,n1537);
xor (n1536,n1533,n1534);
or (n1537,n1538,n1541);
and (n1538,n1539,n1540);
xor (n1539,n1433,n1434);
and (n1540,n296,n47);
and (n1541,n1542,n1543);
xor (n1542,n1539,n1540);
or (n1543,n1544,n1547);
and (n1544,n1545,n1546);
xor (n1545,n1439,n1440);
and (n1546,n335,n47);
and (n1547,n1548,n1549);
xor (n1548,n1545,n1546);
or (n1549,n1550,n1553);
and (n1550,n1551,n1552);
xor (n1551,n1445,n1446);
and (n1552,n398,n47);
and (n1553,n1554,n1555);
xor (n1554,n1551,n1552);
or (n1555,n1556,n1559);
and (n1556,n1557,n1558);
xor (n1557,n1451,n1452);
and (n1558,n414,n47);
and (n1559,n1560,n1561);
xor (n1560,n1557,n1558);
or (n1561,n1562,n1565);
and (n1562,n1563,n1564);
xor (n1563,n1457,n1458);
and (n1564,n408,n47);
and (n1565,n1566,n1567);
xor (n1566,n1563,n1564);
or (n1567,n1568,n1570);
and (n1568,n1569,n650);
xor (n1569,n1463,n1464);
and (n1570,n1571,n1572);
xor (n1571,n1569,n650);
and (n1572,n1573,n1574);
xor (n1573,n1469,n1470);
and (n1574,n383,n47);
and (n1575,n97,n69);
or (n1576,n1577,n1579);
and (n1577,n1578,n1575);
xor (n1578,n1477,n1478);
and (n1579,n1580,n1581);
xor (n1580,n1578,n1575);
or (n1581,n1582,n1585);
and (n1582,n1583,n1584);
xor (n1583,n1482,n1483);
and (n1584,n98,n69);
and (n1585,n1586,n1587);
xor (n1586,n1583,n1584);
or (n1587,n1588,n1591);
and (n1588,n1589,n1590);
xor (n1589,n1488,n1489);
and (n1590,n60,n69);
and (n1591,n1592,n1593);
xor (n1592,n1589,n1590);
or (n1593,n1594,n1597);
and (n1594,n1595,n1596);
xor (n1595,n1494,n1495);
and (n1596,n53,n69);
and (n1597,n1598,n1599);
xor (n1598,n1595,n1596);
or (n1599,n1600,n1603);
and (n1600,n1601,n1602);
xor (n1601,n1500,n1501);
and (n1602,n85,n69);
and (n1603,n1604,n1605);
xor (n1604,n1601,n1602);
or (n1605,n1606,n1609);
and (n1606,n1607,n1608);
xor (n1607,n1506,n1507);
and (n1608,n79,n69);
and (n1609,n1610,n1611);
xor (n1610,n1607,n1608);
or (n1611,n1612,n1615);
and (n1612,n1613,n1614);
xor (n1613,n1512,n1513);
and (n1614,n29,n69);
and (n1615,n1616,n1617);
xor (n1616,n1613,n1614);
or (n1617,n1618,n1621);
and (n1618,n1619,n1620);
xor (n1619,n1518,n1519);
and (n1620,n144,n69);
and (n1621,n1622,n1623);
xor (n1622,n1619,n1620);
or (n1623,n1624,n1627);
and (n1624,n1625,n1626);
xor (n1625,n1524,n1525);
and (n1626,n194,n69);
and (n1627,n1628,n1629);
xor (n1628,n1625,n1626);
or (n1629,n1630,n1633);
and (n1630,n1631,n1632);
xor (n1631,n1530,n1531);
and (n1632,n244,n69);
and (n1633,n1634,n1635);
xor (n1634,n1631,n1632);
or (n1635,n1636,n1639);
and (n1636,n1637,n1638);
xor (n1637,n1536,n1537);
and (n1638,n296,n69);
and (n1639,n1640,n1641);
xor (n1640,n1637,n1638);
or (n1641,n1642,n1645);
and (n1642,n1643,n1644);
xor (n1643,n1542,n1543);
and (n1644,n335,n69);
and (n1645,n1646,n1647);
xor (n1646,n1643,n1644);
or (n1647,n1648,n1651);
and (n1648,n1649,n1650);
xor (n1649,n1548,n1549);
and (n1650,n398,n69);
and (n1651,n1652,n1653);
xor (n1652,n1649,n1650);
or (n1653,n1654,n1657);
and (n1654,n1655,n1656);
xor (n1655,n1554,n1555);
and (n1656,n414,n69);
and (n1657,n1658,n1659);
xor (n1658,n1655,n1656);
or (n1659,n1660,n1663);
and (n1660,n1661,n1662);
xor (n1661,n1560,n1561);
and (n1662,n408,n69);
and (n1663,n1664,n1665);
xor (n1664,n1661,n1662);
or (n1665,n1666,n1669);
and (n1666,n1667,n1668);
xor (n1667,n1566,n1567);
and (n1668,n389,n69);
and (n1669,n1670,n1671);
xor (n1670,n1667,n1668);
and (n1671,n1672,n1673);
xor (n1672,n1571,n1572);
not (n1673,n456);
and (n1674,n97,n18);
or (n1675,n1676,n1679);
and (n1676,n1677,n1678);
xor (n1677,n1580,n1581);
and (n1678,n98,n18);
and (n1679,n1680,n1681);
xor (n1680,n1677,n1678);
or (n1681,n1682,n1685);
and (n1682,n1683,n1684);
xor (n1683,n1586,n1587);
and (n1684,n60,n18);
and (n1685,n1686,n1687);
xor (n1686,n1683,n1684);
or (n1687,n1688,n1691);
and (n1688,n1689,n1690);
xor (n1689,n1592,n1593);
and (n1690,n53,n18);
and (n1691,n1692,n1693);
xor (n1692,n1689,n1690);
or (n1693,n1694,n1697);
and (n1694,n1695,n1696);
xor (n1695,n1598,n1599);
and (n1696,n85,n18);
and (n1697,n1698,n1699);
xor (n1698,n1695,n1696);
or (n1699,n1700,n1703);
and (n1700,n1701,n1702);
xor (n1701,n1604,n1605);
and (n1702,n79,n18);
and (n1703,n1704,n1705);
xor (n1704,n1701,n1702);
or (n1705,n1706,n1709);
and (n1706,n1707,n1708);
xor (n1707,n1610,n1611);
and (n1708,n29,n18);
and (n1709,n1710,n1711);
xor (n1710,n1707,n1708);
or (n1711,n1712,n1714);
and (n1712,n1713,n187);
xor (n1713,n1616,n1617);
and (n1714,n1715,n1716);
xor (n1715,n1713,n187);
or (n1716,n1717,n1719);
and (n1717,n1718,n236);
xor (n1718,n1622,n1623);
and (n1719,n1720,n1721);
xor (n1720,n1718,n236);
or (n1721,n1722,n1725);
and (n1722,n1723,n1724);
xor (n1723,n1628,n1629);
and (n1724,n244,n18);
and (n1725,n1726,n1727);
xor (n1726,n1723,n1724);
or (n1727,n1728,n1731);
and (n1728,n1729,n1730);
xor (n1729,n1634,n1635);
and (n1730,n296,n18);
and (n1731,n1732,n1733);
xor (n1732,n1729,n1730);
or (n1733,n1734,n1736);
and (n1734,n1735,n593);
xor (n1735,n1640,n1641);
and (n1736,n1737,n1738);
xor (n1737,n1735,n593);
or (n1738,n1739,n1741);
and (n1739,n1740,n546);
xor (n1740,n1646,n1647);
and (n1741,n1742,n1743);
xor (n1742,n1740,n546);
or (n1743,n1744,n1746);
and (n1744,n1745,n475);
xor (n1745,n1652,n1653);
and (n1746,n1747,n1748);
xor (n1747,n1745,n475);
or (n1748,n1749,n1752);
and (n1749,n1750,n1751);
xor (n1750,n1658,n1659);
and (n1751,n408,n18);
and (n1752,n1753,n1754);
xor (n1753,n1750,n1751);
or (n1754,n1755,n1758);
and (n1755,n1756,n1757);
xor (n1756,n1664,n1665);
and (n1757,n389,n18);
and (n1758,n1759,n1760);
xor (n1759,n1756,n1757);
and (n1760,n1761,n1762);
xor (n1761,n1670,n1671);
and (n1762,n383,n18);
and (n1763,n98,n22);
or (n1764,n1765,n1767);
and (n1765,n1766,n893);
xor (n1766,n1680,n1681);
and (n1767,n1768,n1769);
xor (n1768,n1766,n893);
or (n1769,n1770,n1773);
and (n1770,n1771,n1772);
xor (n1771,n1686,n1687);
and (n1772,n53,n22);
and (n1773,n1774,n1775);
xor (n1774,n1771,n1772);
or (n1775,n1776,n1779);
and (n1776,n1777,n1778);
xor (n1777,n1692,n1693);
and (n1778,n85,n22);
and (n1779,n1780,n1781);
xor (n1780,n1777,n1778);
or (n1781,n1782,n1785);
and (n1782,n1783,n1784);
xor (n1783,n1698,n1699);
and (n1784,n79,n22);
and (n1785,n1786,n1787);
xor (n1786,n1783,n1784);
or (n1787,n1788,n1791);
and (n1788,n1789,n1790);
xor (n1789,n1704,n1705);
and (n1790,n29,n22);
and (n1791,n1792,n1793);
xor (n1792,n1789,n1790);
or (n1793,n1794,n1797);
and (n1794,n1795,n1796);
xor (n1795,n1710,n1711);
and (n1796,n144,n22);
and (n1797,n1798,n1799);
xor (n1798,n1795,n1796);
or (n1799,n1800,n1803);
and (n1800,n1801,n1802);
xor (n1801,n1715,n1716);
and (n1802,n194,n22);
and (n1803,n1804,n1805);
xor (n1804,n1801,n1802);
or (n1805,n1806,n1809);
and (n1806,n1807,n1808);
xor (n1807,n1720,n1721);
and (n1808,n244,n22);
and (n1809,n1810,n1811);
xor (n1810,n1807,n1808);
or (n1811,n1812,n1815);
and (n1812,n1813,n1814);
xor (n1813,n1726,n1727);
and (n1814,n296,n22);
and (n1815,n1816,n1817);
xor (n1816,n1813,n1814);
or (n1817,n1818,n1821);
and (n1818,n1819,n1820);
xor (n1819,n1732,n1733);
and (n1820,n335,n22);
and (n1821,n1822,n1823);
xor (n1822,n1819,n1820);
or (n1823,n1824,n1827);
and (n1824,n1825,n1826);
xor (n1825,n1737,n1738);
and (n1826,n398,n22);
and (n1827,n1828,n1829);
xor (n1828,n1825,n1826);
or (n1829,n1830,n1833);
and (n1830,n1831,n1832);
xor (n1831,n1742,n1743);
and (n1832,n414,n22);
and (n1833,n1834,n1835);
xor (n1834,n1831,n1832);
or (n1835,n1836,n1839);
and (n1836,n1837,n1838);
xor (n1837,n1747,n1748);
and (n1838,n408,n22);
and (n1839,n1840,n1841);
xor (n1840,n1837,n1838);
or (n1841,n1842,n1845);
and (n1842,n1843,n1844);
xor (n1843,n1753,n1754);
and (n1844,n389,n22);
and (n1845,n1846,n1847);
xor (n1846,n1843,n1844);
and (n1847,n1848,n1849);
xor (n1848,n1759,n1760);
and (n1849,n383,n22);
or (n1850,n1851,n1853);
and (n1851,n1852,n1772);
xor (n1852,n1768,n1769);
and (n1853,n1854,n1855);
xor (n1854,n1852,n1772);
or (n1855,n1856,n1858);
and (n1856,n1857,n1778);
xor (n1857,n1774,n1775);
and (n1858,n1859,n1860);
xor (n1859,n1857,n1778);
or (n1860,n1861,n1863);
and (n1861,n1862,n1784);
xor (n1862,n1780,n1781);
and (n1863,n1864,n1865);
xor (n1864,n1862,n1784);
or (n1865,n1866,n1868);
and (n1866,n1867,n1790);
xor (n1867,n1786,n1787);
and (n1868,n1869,n1870);
xor (n1869,n1867,n1790);
or (n1870,n1871,n1873);
and (n1871,n1872,n1796);
xor (n1872,n1792,n1793);
and (n1873,n1874,n1875);
xor (n1874,n1872,n1796);
or (n1875,n1876,n1878);
and (n1876,n1877,n1802);
xor (n1877,n1798,n1799);
and (n1878,n1879,n1880);
xor (n1879,n1877,n1802);
or (n1880,n1881,n1883);
and (n1881,n1882,n1808);
xor (n1882,n1804,n1805);
and (n1883,n1884,n1885);
xor (n1884,n1882,n1808);
or (n1885,n1886,n1888);
and (n1886,n1887,n1814);
xor (n1887,n1810,n1811);
and (n1888,n1889,n1890);
xor (n1889,n1887,n1814);
or (n1890,n1891,n1893);
and (n1891,n1892,n1820);
xor (n1892,n1816,n1817);
and (n1893,n1894,n1895);
xor (n1894,n1892,n1820);
or (n1895,n1896,n1898);
and (n1896,n1897,n1826);
xor (n1897,n1822,n1823);
and (n1898,n1899,n1900);
xor (n1899,n1897,n1826);
or (n1900,n1901,n1903);
and (n1901,n1902,n1832);
xor (n1902,n1828,n1829);
and (n1903,n1904,n1905);
xor (n1904,n1902,n1832);
or (n1905,n1906,n1908);
and (n1906,n1907,n1838);
xor (n1907,n1834,n1835);
and (n1908,n1909,n1910);
xor (n1909,n1907,n1838);
or (n1910,n1911,n1913);
and (n1911,n1912,n1844);
xor (n1912,n1840,n1841);
and (n1913,n1914,n1915);
xor (n1914,n1912,n1844);
and (n1915,n1916,n1849);
xor (n1916,n1846,n1847);
or (n1917,n1918,n1920);
and (n1918,n1919,n1778);
xor (n1919,n1854,n1855);
and (n1920,n1921,n1922);
xor (n1921,n1919,n1778);
or (n1922,n1923,n1925);
and (n1923,n1924,n1784);
xor (n1924,n1859,n1860);
and (n1925,n1926,n1927);
xor (n1926,n1924,n1784);
or (n1927,n1928,n1930);
and (n1928,n1929,n1790);
xor (n1929,n1864,n1865);
and (n1930,n1931,n1932);
xor (n1931,n1929,n1790);
or (n1932,n1933,n1935);
and (n1933,n1934,n1796);
xor (n1934,n1869,n1870);
and (n1935,n1936,n1937);
xor (n1936,n1934,n1796);
or (n1937,n1938,n1940);
and (n1938,n1939,n1802);
xor (n1939,n1874,n1875);
and (n1940,n1941,n1942);
xor (n1941,n1939,n1802);
or (n1942,n1943,n1945);
and (n1943,n1944,n1808);
xor (n1944,n1879,n1880);
and (n1945,n1946,n1947);
xor (n1946,n1944,n1808);
or (n1947,n1948,n1950);
and (n1948,n1949,n1814);
xor (n1949,n1884,n1885);
and (n1950,n1951,n1952);
xor (n1951,n1949,n1814);
or (n1952,n1953,n1955);
and (n1953,n1954,n1820);
xor (n1954,n1889,n1890);
and (n1955,n1956,n1957);
xor (n1956,n1954,n1820);
or (n1957,n1958,n1960);
and (n1958,n1959,n1826);
xor (n1959,n1894,n1895);
and (n1960,n1961,n1962);
xor (n1961,n1959,n1826);
or (n1962,n1963,n1965);
and (n1963,n1964,n1832);
xor (n1964,n1899,n1900);
and (n1965,n1966,n1967);
xor (n1966,n1964,n1832);
or (n1967,n1968,n1970);
and (n1968,n1969,n1838);
xor (n1969,n1904,n1905);
and (n1970,n1971,n1972);
xor (n1971,n1969,n1838);
or (n1972,n1973,n1975);
and (n1973,n1974,n1844);
xor (n1974,n1909,n1910);
and (n1975,n1976,n1977);
xor (n1976,n1974,n1844);
and (n1977,n1978,n1849);
xor (n1978,n1914,n1915);
or (n1979,n1980,n1982);
and (n1980,n1981,n1784);
xor (n1981,n1921,n1922);
and (n1982,n1983,n1984);
xor (n1983,n1981,n1784);
or (n1984,n1985,n1987);
and (n1985,n1986,n1790);
xor (n1986,n1926,n1927);
and (n1987,n1988,n1989);
xor (n1988,n1986,n1790);
or (n1989,n1990,n1992);
and (n1990,n1991,n1796);
xor (n1991,n1931,n1932);
and (n1992,n1993,n1994);
xor (n1993,n1991,n1796);
or (n1994,n1995,n1997);
and (n1995,n1996,n1802);
xor (n1996,n1936,n1937);
and (n1997,n1998,n1999);
xor (n1998,n1996,n1802);
or (n1999,n2000,n2002);
and (n2000,n2001,n1808);
xor (n2001,n1941,n1942);
and (n2002,n2003,n2004);
xor (n2003,n2001,n1808);
or (n2004,n2005,n2007);
and (n2005,n2006,n1814);
xor (n2006,n1946,n1947);
and (n2007,n2008,n2009);
xor (n2008,n2006,n1814);
or (n2009,n2010,n2012);
and (n2010,n2011,n1820);
xor (n2011,n1951,n1952);
and (n2012,n2013,n2014);
xor (n2013,n2011,n1820);
or (n2014,n2015,n2017);
and (n2015,n2016,n1826);
xor (n2016,n1956,n1957);
and (n2017,n2018,n2019);
xor (n2018,n2016,n1826);
or (n2019,n2020,n2022);
and (n2020,n2021,n1832);
xor (n2021,n1961,n1962);
and (n2022,n2023,n2024);
xor (n2023,n2021,n1832);
or (n2024,n2025,n2027);
and (n2025,n2026,n1838);
xor (n2026,n1966,n1967);
and (n2027,n2028,n2029);
xor (n2028,n2026,n1838);
or (n2029,n2030,n2032);
and (n2030,n2031,n1844);
xor (n2031,n1971,n1972);
and (n2032,n2033,n2034);
xor (n2033,n2031,n1844);
and (n2034,n2035,n1849);
xor (n2035,n1976,n1977);
or (n2036,n2037,n2039);
and (n2037,n2038,n1790);
xor (n2038,n1983,n1984);
and (n2039,n2040,n2041);
xor (n2040,n2038,n1790);
or (n2041,n2042,n2044);
and (n2042,n2043,n1796);
xor (n2043,n1988,n1989);
and (n2044,n2045,n2046);
xor (n2045,n2043,n1796);
or (n2046,n2047,n2049);
and (n2047,n2048,n1802);
xor (n2048,n1993,n1994);
and (n2049,n2050,n2051);
xor (n2050,n2048,n1802);
or (n2051,n2052,n2054);
and (n2052,n2053,n1808);
xor (n2053,n1998,n1999);
and (n2054,n2055,n2056);
xor (n2055,n2053,n1808);
or (n2056,n2057,n2059);
and (n2057,n2058,n1814);
xor (n2058,n2003,n2004);
and (n2059,n2060,n2061);
xor (n2060,n2058,n1814);
or (n2061,n2062,n2064);
and (n2062,n2063,n1820);
xor (n2063,n2008,n2009);
and (n2064,n2065,n2066);
xor (n2065,n2063,n1820);
or (n2066,n2067,n2069);
and (n2067,n2068,n1826);
xor (n2068,n2013,n2014);
and (n2069,n2070,n2071);
xor (n2070,n2068,n1826);
or (n2071,n2072,n2074);
and (n2072,n2073,n1832);
xor (n2073,n2018,n2019);
and (n2074,n2075,n2076);
xor (n2075,n2073,n1832);
or (n2076,n2077,n2079);
and (n2077,n2078,n1838);
xor (n2078,n2023,n2024);
and (n2079,n2080,n2081);
xor (n2080,n2078,n1838);
or (n2081,n2082,n2084);
and (n2082,n2083,n1844);
xor (n2083,n2028,n2029);
and (n2084,n2085,n2086);
xor (n2085,n2083,n1844);
and (n2086,n2087,n1849);
xor (n2087,n2033,n2034);
or (n2088,n2089,n2091);
and (n2089,n2090,n1796);
xor (n2090,n2040,n2041);
and (n2091,n2092,n2093);
xor (n2092,n2090,n1796);
or (n2093,n2094,n2096);
and (n2094,n2095,n1802);
xor (n2095,n2045,n2046);
and (n2096,n2097,n2098);
xor (n2097,n2095,n1802);
or (n2098,n2099,n2101);
and (n2099,n2100,n1808);
xor (n2100,n2050,n2051);
and (n2101,n2102,n2103);
xor (n2102,n2100,n1808);
or (n2103,n2104,n2106);
and (n2104,n2105,n1814);
xor (n2105,n2055,n2056);
and (n2106,n2107,n2108);
xor (n2107,n2105,n1814);
or (n2108,n2109,n2111);
and (n2109,n2110,n1820);
xor (n2110,n2060,n2061);
and (n2111,n2112,n2113);
xor (n2112,n2110,n1820);
or (n2113,n2114,n2116);
and (n2114,n2115,n1826);
xor (n2115,n2065,n2066);
and (n2116,n2117,n2118);
xor (n2117,n2115,n1826);
or (n2118,n2119,n2121);
and (n2119,n2120,n1832);
xor (n2120,n2070,n2071);
and (n2121,n2122,n2123);
xor (n2122,n2120,n1832);
or (n2123,n2124,n2126);
and (n2124,n2125,n1838);
xor (n2125,n2075,n2076);
and (n2126,n2127,n2128);
xor (n2127,n2125,n1838);
or (n2128,n2129,n2131);
and (n2129,n2130,n1844);
xor (n2130,n2080,n2081);
and (n2131,n2132,n2133);
xor (n2132,n2130,n1844);
and (n2133,n2134,n1849);
xor (n2134,n2085,n2086);
or (n2135,n2136,n2138);
and (n2136,n2137,n1802);
xor (n2137,n2092,n2093);
and (n2138,n2139,n2140);
xor (n2139,n2137,n1802);
or (n2140,n2141,n2143);
and (n2141,n2142,n1808);
xor (n2142,n2097,n2098);
and (n2143,n2144,n2145);
xor (n2144,n2142,n1808);
or (n2145,n2146,n2148);
and (n2146,n2147,n1814);
xor (n2147,n2102,n2103);
and (n2148,n2149,n2150);
xor (n2149,n2147,n1814);
or (n2150,n2151,n2153);
and (n2151,n2152,n1820);
xor (n2152,n2107,n2108);
and (n2153,n2154,n2155);
xor (n2154,n2152,n1820);
or (n2155,n2156,n2158);
and (n2156,n2157,n1826);
xor (n2157,n2112,n2113);
and (n2158,n2159,n2160);
xor (n2159,n2157,n1826);
or (n2160,n2161,n2163);
and (n2161,n2162,n1832);
xor (n2162,n2117,n2118);
and (n2163,n2164,n2165);
xor (n2164,n2162,n1832);
or (n2165,n2166,n2168);
and (n2166,n2167,n1838);
xor (n2167,n2122,n2123);
and (n2168,n2169,n2170);
xor (n2169,n2167,n1838);
or (n2170,n2171,n2173);
and (n2171,n2172,n1844);
xor (n2172,n2127,n2128);
and (n2173,n2174,n2175);
xor (n2174,n2172,n1844);
and (n2175,n2176,n1849);
xor (n2176,n2132,n2133);
or (n2177,n2178,n2180);
and (n2178,n2179,n1808);
xor (n2179,n2139,n2140);
and (n2180,n2181,n2182);
xor (n2181,n2179,n1808);
or (n2182,n2183,n2185);
and (n2183,n2184,n1814);
xor (n2184,n2144,n2145);
and (n2185,n2186,n2187);
xor (n2186,n2184,n1814);
or (n2187,n2188,n2190);
and (n2188,n2189,n1820);
xor (n2189,n2149,n2150);
and (n2190,n2191,n2192);
xor (n2191,n2189,n1820);
or (n2192,n2193,n2195);
and (n2193,n2194,n1826);
xor (n2194,n2154,n2155);
and (n2195,n2196,n2197);
xor (n2196,n2194,n1826);
or (n2197,n2198,n2200);
and (n2198,n2199,n1832);
xor (n2199,n2159,n2160);
and (n2200,n2201,n2202);
xor (n2201,n2199,n1832);
or (n2202,n2203,n2205);
and (n2203,n2204,n1838);
xor (n2204,n2164,n2165);
and (n2205,n2206,n2207);
xor (n2206,n2204,n1838);
or (n2207,n2208,n2210);
and (n2208,n2209,n1844);
xor (n2209,n2169,n2170);
and (n2210,n2211,n2212);
xor (n2211,n2209,n1844);
and (n2212,n2213,n1849);
xor (n2213,n2174,n2175);
or (n2214,n2215,n2217);
and (n2215,n2216,n1814);
xor (n2216,n2181,n2182);
and (n2217,n2218,n2219);
xor (n2218,n2216,n1814);
or (n2219,n2220,n2222);
and (n2220,n2221,n1820);
xor (n2221,n2186,n2187);
and (n2222,n2223,n2224);
xor (n2223,n2221,n1820);
or (n2224,n2225,n2227);
and (n2225,n2226,n1826);
xor (n2226,n2191,n2192);
and (n2227,n2228,n2229);
xor (n2228,n2226,n1826);
or (n2229,n2230,n2232);
and (n2230,n2231,n1832);
xor (n2231,n2196,n2197);
and (n2232,n2233,n2234);
xor (n2233,n2231,n1832);
or (n2234,n2235,n2237);
and (n2235,n2236,n1838);
xor (n2236,n2201,n2202);
and (n2237,n2238,n2239);
xor (n2238,n2236,n1838);
or (n2239,n2240,n2242);
and (n2240,n2241,n1844);
xor (n2241,n2206,n2207);
and (n2242,n2243,n2244);
xor (n2243,n2241,n1844);
and (n2244,n2245,n1849);
xor (n2245,n2211,n2212);
or (n2246,n2247,n2249);
and (n2247,n2248,n1820);
xor (n2248,n2218,n2219);
and (n2249,n2250,n2251);
xor (n2250,n2248,n1820);
or (n2251,n2252,n2254);
and (n2252,n2253,n1826);
xor (n2253,n2223,n2224);
and (n2254,n2255,n2256);
xor (n2255,n2253,n1826);
or (n2256,n2257,n2259);
and (n2257,n2258,n1832);
xor (n2258,n2228,n2229);
and (n2259,n2260,n2261);
xor (n2260,n2258,n1832);
or (n2261,n2262,n2264);
and (n2262,n2263,n1838);
xor (n2263,n2233,n2234);
and (n2264,n2265,n2266);
xor (n2265,n2263,n1838);
or (n2266,n2267,n2269);
and (n2267,n2268,n1844);
xor (n2268,n2238,n2239);
and (n2269,n2270,n2271);
xor (n2270,n2268,n1844);
and (n2271,n2272,n1849);
xor (n2272,n2243,n2244);
or (n2273,n2274,n2276);
and (n2274,n2275,n1826);
xor (n2275,n2250,n2251);
and (n2276,n2277,n2278);
xor (n2277,n2275,n1826);
or (n2278,n2279,n2281);
and (n2279,n2280,n1832);
xor (n2280,n2255,n2256);
and (n2281,n2282,n2283);
xor (n2282,n2280,n1832);
or (n2283,n2284,n2286);
and (n2284,n2285,n1838);
xor (n2285,n2260,n2261);
and (n2286,n2287,n2288);
xor (n2287,n2285,n1838);
or (n2288,n2289,n2291);
and (n2289,n2290,n1844);
xor (n2290,n2265,n2266);
and (n2291,n2292,n2293);
xor (n2292,n2290,n1844);
and (n2293,n2294,n1849);
xor (n2294,n2270,n2271);
or (n2295,n2296,n2298);
and (n2296,n2297,n1832);
xor (n2297,n2277,n2278);
and (n2298,n2299,n2300);
xor (n2299,n2297,n1832);
or (n2300,n2301,n2303);
and (n2301,n2302,n1838);
xor (n2302,n2282,n2283);
and (n2303,n2304,n2305);
xor (n2304,n2302,n1838);
or (n2305,n2306,n2308);
and (n2306,n2307,n1844);
xor (n2307,n2287,n2288);
and (n2308,n2309,n2310);
xor (n2309,n2307,n1844);
and (n2310,n2311,n1849);
xor (n2311,n2292,n2293);
or (n2312,n2313,n2315);
and (n2313,n2314,n1838);
xor (n2314,n2299,n2300);
and (n2315,n2316,n2317);
xor (n2316,n2314,n1838);
or (n2317,n2318,n2320);
and (n2318,n2319,n1844);
xor (n2319,n2304,n2305);
and (n2320,n2321,n2322);
xor (n2321,n2319,n1844);
and (n2322,n2323,n1849);
xor (n2323,n2309,n2310);
or (n2324,n2325,n2327);
and (n2325,n2326,n1844);
xor (n2326,n2316,n2317);
and (n2327,n2328,n2329);
xor (n2328,n2326,n1844);
and (n2329,n2330,n1849);
xor (n2330,n2321,n2322);
and (n2331,n2332,n1849);
xor (n2332,n2328,n2329);
xor (n2333,n2294,n1849);
endmodule
