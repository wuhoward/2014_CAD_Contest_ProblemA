module top (out,n15,n16,n21,n24,n30,n40,n46,n47,n57
        ,n68,n70,n76,n85,n96,n100,n107,n121,n133,n140
        ,n144,n189,n195,n262,n320,n321,n352,n412,n434,n435
        ,n464,n604,n637,n698,n777);
output out;
input n15;
input n16;
input n21;
input n24;
input n30;
input n40;
input n46;
input n47;
input n57;
input n68;
input n70;
input n76;
input n85;
input n96;
input n100;
input n107;
input n121;
input n133;
input n140;
input n144;
input n189;
input n195;
input n262;
input n320;
input n321;
input n352;
input n412;
input n434;
input n435;
input n464;
input n604;
input n637;
input n698;
input n777;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n17;
wire n18;
wire n19;
wire n20;
wire n22;
wire n23;
wire n25;
wire n26;
wire n27;
wire n28;
wire n29;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n36;
wire n37;
wire n38;
wire n39;
wire n41;
wire n42;
wire n43;
wire n44;
wire n45;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n65;
wire n66;
wire n67;
wire n69;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n97;
wire n98;
wire n99;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n141;
wire n142;
wire n143;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
wire n1181;
wire n1182;
wire n1183;
wire n1184;
wire n1185;
wire n1186;
wire n1187;
wire n1188;
wire n1189;
wire n1190;
wire n1191;
wire n1192;
wire n1193;
wire n1194;
wire n1195;
wire n1196;
wire n1197;
wire n1198;
wire n1199;
wire n1200;
wire n1201;
wire n1202;
wire n1203;
wire n1204;
wire n1205;
wire n1206;
wire n1207;
wire n1208;
wire n1209;
wire n1210;
wire n1211;
wire n1212;
wire n1213;
wire n1214;
wire n1215;
wire n1216;
wire n1217;
wire n1218;
wire n1219;
wire n1220;
wire n1221;
wire n1222;
wire n1223;
wire n1224;
wire n1225;
wire n1226;
wire n1227;
wire n1228;
wire n1229;
wire n1230;
wire n1231;
wire n1232;
wire n1233;
wire n1234;
wire n1235;
wire n1236;
wire n1237;
wire n1238;
wire n1239;
wire n1240;
wire n1241;
wire n1242;
wire n1243;
wire n1244;
wire n1245;
wire n1246;
wire n1247;
wire n1248;
wire n1249;
wire n1250;
wire n1251;
wire n1252;
wire n1253;
wire n1254;
wire n1255;
wire n1256;
wire n1257;
wire n1258;
wire n1259;
wire n1260;
wire n1261;
wire n1262;
wire n1263;
wire n1264;
wire n1265;
wire n1266;
wire n1267;
wire n1268;
wire n1269;
wire n1270;
wire n1271;
wire n1272;
wire n1273;
wire n1274;
wire n1275;
wire n1276;
wire n1277;
wire n1278;
wire n1279;
wire n1280;
wire n1281;
wire n1282;
wire n1283;
wire n1284;
wire n1285;
wire n1286;
wire n1287;
wire n1288;
wire n1289;
wire n1290;
wire n1291;
wire n1292;
wire n1293;
wire n1294;
wire n1295;
wire n1296;
wire n1297;
wire n1298;
wire n1299;
wire n1300;
wire n1301;
wire n1302;
wire n1303;
wire n1304;
wire n1305;
wire n1306;
wire n1307;
wire n1308;
wire n1309;
wire n1310;
wire n1311;
wire n1312;
wire n1313;
wire n1314;
wire n1315;
wire n1316;
wire n1317;
wire n1318;
wire n1319;
wire n1320;
wire n1321;
wire n1322;
wire n1323;
wire n1324;
wire n1325;
wire n1326;
wire n1327;
wire n1328;
wire n1329;
wire n1330;
wire n1331;
wire n1332;
wire n1333;
wire n1334;
wire n1335;
wire n1336;
wire n1337;
wire n1338;
wire n1339;
wire n1340;
wire n1341;
wire n1342;
wire n1343;
wire n1344;
wire n1345;
wire n1346;
wire n1347;
wire n1348;
wire n1349;
wire n1350;
wire n1351;
wire n1352;
wire n1353;
wire n1354;
wire n1355;
wire n1356;
wire n1357;
wire n1358;
wire n1359;
wire n1360;
wire n1361;
wire n1362;
wire n1363;
wire n1364;
wire n1365;
wire n1366;
wire n1367;
wire n1368;
wire n1369;
wire n1370;
wire n1371;
wire n1372;
wire n1373;
wire n1374;
wire n1375;
wire n1376;
wire n1377;
wire n1378;
wire n1379;
wire n1380;
wire n1381;
wire n1382;
wire n1383;
wire n1384;
wire n1385;
wire n1386;
wire n1387;
wire n1388;
wire n1389;
wire n1390;
wire n1391;
wire n1392;
wire n1393;
wire n1394;
wire n1395;
wire n1396;
wire n1397;
wire n1398;
wire n1399;
wire n1400;
wire n1401;
wire n1402;
wire n1403;
wire n1404;
wire n1405;
wire n1406;
wire n1407;
wire n1408;
wire n1409;
wire n1410;
wire n1411;
wire n1412;
wire n1413;
wire n1414;
wire n1415;
wire n1416;
wire n1417;
wire n1418;
wire n1419;
wire n1420;
wire n1421;
wire n1422;
wire n1423;
wire n1424;
wire n1425;
wire n1426;
wire n1427;
wire n1428;
wire n1429;
wire n1430;
wire n1431;
wire n1432;
wire n1433;
wire n1434;
wire n1435;
wire n1436;
wire n1437;
wire n1438;
wire n1439;
wire n1440;
wire n1441;
wire n1442;
wire n1443;
wire n1444;
wire n1445;
wire n1446;
wire n1447;
wire n1448;
wire n1449;
wire n1450;
wire n1451;
wire n1452;
wire n1453;
wire n1454;
wire n1455;
wire n1456;
wire n1457;
wire n1458;
wire n1459;
wire n1460;
wire n1461;
wire n1462;
wire n1463;
wire n1464;
wire n1465;
wire n1466;
wire n1467;
wire n1468;
wire n1469;
wire n1470;
wire n1471;
wire n1472;
wire n1473;
wire n1474;
wire n1475;
wire n1476;
wire n1477;
wire n1478;
wire n1479;
wire n1480;
wire n1481;
wire n1482;
wire n1483;
wire n1484;
wire n1485;
wire n1486;
wire n1487;
wire n1488;
wire n1489;
wire n1490;
wire n1491;
wire n1492;
wire n1493;
wire n1494;
wire n1495;
wire n1496;
wire n1497;
wire n1498;
wire n1499;
wire n1500;
wire n1501;
wire n1502;
wire n1503;
wire n1504;
wire n1505;
wire n1506;
wire n1507;
wire n1508;
wire n1509;
wire n1510;
wire n1511;
wire n1512;
wire n1513;
wire n1514;
wire n1515;
wire n1516;
wire n1517;
wire n1518;
wire n1519;
wire n1520;
wire n1521;
wire n1522;
wire n1523;
wire n1524;
wire n1525;
wire n1526;
wire n1527;
wire n1528;
wire n1529;
wire n1530;
wire n1531;
wire n1532;
wire n1533;
wire n1534;
wire n1535;
wire n1536;
wire n1537;
wire n1538;
wire n1539;
wire n1540;
wire n1541;
wire n1542;
wire n1543;
wire n1544;
wire n1545;
wire n1546;
wire n1547;
wire n1548;
wire n1549;
wire n1550;
wire n1551;
wire n1552;
wire n1553;
wire n1554;
wire n1555;
wire n1556;
wire n1557;
wire n1558;
wire n1559;
wire n1560;
wire n1561;
wire n1562;
wire n1563;
wire n1564;
wire n1565;
wire n1566;
wire n1567;
wire n1568;
wire n1569;
wire n1570;
wire n1571;
wire n1572;
wire n1573;
wire n1574;
wire n1575;
wire n1576;
wire n1577;
wire n1578;
wire n1579;
wire n1580;
wire n1581;
wire n1582;
wire n1583;
wire n1584;
wire n1585;
wire n1586;
wire n1587;
wire n1588;
wire n1589;
wire n1590;
wire n1591;
wire n1592;
wire n1593;
wire n1594;
wire n1595;
wire n1596;
wire n1597;
wire n1598;
wire n1599;
wire n1600;
wire n1601;
wire n1602;
wire n1603;
wire n1604;
wire n1605;
wire n1606;
wire n1607;
wire n1608;
wire n1609;
wire n1610;
wire n1611;
wire n1612;
wire n1613;
wire n1614;
wire n1615;
wire n1616;
wire n1617;
wire n1618;
wire n1619;
wire n1620;
wire n1621;
wire n1622;
wire n1623;
wire n1624;
wire n1625;
wire n1626;
wire n1627;
wire n1628;
wire n1629;
wire n1630;
wire n1631;
wire n1632;
wire n1633;
wire n1634;
wire n1635;
wire n1636;
wire n1637;
wire n1638;
wire n1639;
wire n1640;
wire n1641;
wire n1642;
wire n1643;
wire n1644;
wire n1645;
wire n1646;
wire n1647;
wire n1648;
wire n1649;
wire n1650;
wire n1651;
wire n1652;
wire n1653;
wire n1654;
wire n1655;
wire n1656;
wire n1657;
wire n1658;
wire n1659;
wire n1660;
wire n1661;
wire n1662;
wire n1663;
wire n1664;
wire n1665;
wire n1666;
wire n1667;
wire n1668;
wire n1669;
wire n1670;
wire n1671;
wire n1672;
wire n1673;
wire n1674;
wire n1675;
wire n1676;
wire n1677;
wire n1678;
wire n1679;
wire n1680;
wire n1681;
wire n1682;
wire n1683;
wire n1684;
wire n1685;
wire n1686;
wire n1687;
wire n1688;
wire n1689;
wire n1690;
wire n1691;
wire n1692;
wire n1693;
wire n1694;
wire n1695;
wire n1696;
wire n1697;
wire n1698;
wire n1699;
wire n1700;
wire n1701;
wire n1702;
wire n1703;
wire n1704;
wire n1705;
wire n1706;
wire n1707;
wire n1708;
wire n1709;
wire n1710;
wire n1711;
wire n1712;
wire n1713;
wire n1714;
wire n1715;
wire n1716;
wire n1717;
wire n1718;
wire n1719;
wire n1720;
wire n1721;
wire n1722;
wire n1723;
wire n1724;
wire n1725;
wire n1726;
wire n1727;
wire n1728;
wire n1729;
wire n1730;
wire n1731;
wire n1732;
wire n1733;
wire n1734;
wire n1735;
wire n1736;
wire n1737;
wire n1738;
wire n1739;
wire n1740;
wire n1741;
wire n1742;
wire n1743;
wire n1744;
wire n1745;
wire n1746;
wire n1747;
wire n1748;
wire n1749;
wire n1750;
wire n1751;
wire n1752;
wire n1753;
wire n1754;
wire n1755;
wire n1756;
wire n1757;
wire n1758;
wire n1759;
wire n1760;
wire n1761;
wire n1762;
wire n1763;
wire n1764;
wire n1765;
wire n1766;
wire n1767;
wire n1768;
wire n1769;
wire n1770;
wire n1771;
wire n1772;
wire n1773;
wire n1774;
wire n1775;
wire n1776;
wire n1777;
wire n1778;
wire n1779;
wire n1780;
wire n1781;
wire n1782;
wire n1783;
wire n1784;
wire n1785;
wire n1786;
wire n1787;
wire n1788;
wire n1789;
wire n1790;
wire n1791;
wire n1792;
wire n1793;
wire n1794;
wire n1795;
wire n1796;
wire n1797;
wire n1798;
wire n1799;
wire n1800;
wire n1801;
wire n1802;
wire n1803;
wire n1804;
wire n1805;
wire n1806;
wire n1807;
wire n1808;
wire n1809;
wire n1810;
wire n1811;
wire n1812;
wire n1813;
wire n1814;
wire n1815;
wire n1816;
wire n1817;
wire n1818;
wire n1819;
wire n1820;
wire n1821;
wire n1822;
wire n1823;
wire n1824;
wire n1825;
wire n1826;
wire n1827;
wire n1828;
wire n1829;
wire n1830;
wire n1831;
wire n1832;
wire n1833;
wire n1834;
wire n1835;
wire n1836;
wire n1837;
wire n1838;
wire n1839;
wire n1840;
wire n1841;
wire n1842;
wire n1843;
wire n1844;
wire n1845;
wire n1846;
wire n1847;
wire n1848;
wire n1849;
wire n1850;
wire n1851;
wire n1852;
wire n1853;
wire n1854;
wire n1855;
wire n1856;
wire n1857;
wire n1858;
wire n1859;
wire n1860;
wire n1861;
wire n1862;
wire n1863;
wire n1864;
wire n1865;
wire n1866;
wire n1867;
wire n1868;
wire n1869;
wire n1870;
wire n1871;
wire n1872;
wire n1873;
wire n1874;
wire n1875;
wire n1876;
wire n1877;
wire n1878;
wire n1879;
wire n1880;
wire n1881;
wire n1882;
wire n1883;
wire n1884;
wire n1885;
wire n1886;
wire n1887;
wire n1888;
wire n1889;
wire n1890;
wire n1891;
wire n1892;
wire n1893;
wire n1894;
wire n1895;
wire n1896;
wire n1897;
wire n1898;
wire n1899;
wire n1900;
wire n1901;
wire n1902;
wire n1903;
wire n1904;
wire n1905;
wire n1906;
wire n1907;
wire n1908;
wire n1909;
wire n1910;
wire n1911;
wire n1912;
wire n1913;
wire n1914;
wire n1915;
wire n1916;
wire n1917;
wire n1918;
wire n1919;
wire n1920;
wire n1921;
wire n1922;
wire n1923;
wire n1924;
wire n1925;
wire n1926;
wire n1927;
wire n1928;
wire n1929;
wire n1930;
wire n1931;
wire n1932;
wire n1933;
wire n1934;
wire n1935;
wire n1936;
wire n1937;
wire n1938;
wire n1939;
wire n1940;
wire n1941;
wire n1942;
wire n1943;
wire n1944;
wire n1945;
wire n1946;
wire n1947;
wire n1948;
wire n1949;
wire n1950;
wire n1951;
wire n1952;
wire n1953;
wire n1954;
wire n1955;
wire n1956;
wire n1957;
wire n1958;
wire n1959;
wire n1960;
wire n1961;
wire n1962;
wire n1963;
wire n1964;
wire n1965;
wire n1966;
wire n1967;
wire n1968;
wire n1969;
wire n1970;
wire n1971;
wire n1972;
wire n1973;
wire n1974;
wire n1975;
wire n1976;
wire n1977;
wire n1978;
wire n1979;
wire n1980;
wire n1981;
wire n1982;
wire n1983;
wire n1984;
wire n1985;
wire n1986;
wire n1987;
wire n1988;
wire n1989;
wire n1990;
wire n1991;
wire n1992;
wire n1993;
wire n1994;
wire n1995;
wire n1996;
wire n1997;
wire n1998;
wire n1999;
wire n2000;
wire n2001;
wire n2002;
wire n2003;
wire n2004;
wire n2005;
wire n2006;
wire n2007;
wire n2008;
wire n2009;
wire n2010;
wire n2011;
wire n2012;
wire n2013;
wire n2014;
wire n2015;
wire n2016;
wire n2017;
wire n2018;
wire n2019;
wire n2020;
wire n2021;
wire n2022;
wire n2023;
wire n2024;
wire n2025;
wire n2026;
wire n2027;
wire n2028;
wire n2029;
wire n2030;
wire n2031;
wire n2032;
wire n2033;
wire n2034;
wire n2035;
wire n2036;
wire n2037;
wire n2038;
wire n2039;
wire n2040;
wire n2041;
wire n2042;
wire n2043;
wire n2044;
wire n2045;
wire n2046;
wire n2047;
wire n2048;
wire n2049;
wire n2050;
wire n2051;
wire n2052;
wire n2053;
wire n2054;
wire n2055;
wire n2056;
wire n2057;
wire n2058;
wire n2059;
wire n2060;
wire n2061;
wire n2062;
wire n2063;
wire n2064;
wire n2065;
wire n2066;
wire n2067;
wire n2068;
wire n2069;
wire n2070;
wire n2071;
wire n2072;
wire n2073;
wire n2074;
wire n2075;
wire n2076;
wire n2077;
wire n2078;
wire n2079;
wire n2080;
wire n2081;
wire n2082;
wire n2083;
wire n2084;
wire n2085;
wire n2086;
wire n2087;
wire n2088;
wire n2089;
wire n2090;
wire n2091;
wire n2092;
wire n2093;
wire n2094;
wire n2095;
wire n2096;
wire n2097;
wire n2098;
wire n2099;
wire n2100;
wire n2101;
wire n2102;
wire n2103;
wire n2104;
wire n2105;
wire n2106;
wire n2107;
wire n2108;
wire n2109;
wire n2110;
wire n2111;
wire n2112;
wire n2113;
wire n2114;
wire n2115;
wire n2116;
wire n2117;
wire n2118;
wire n2119;
wire n2120;
wire n2121;
wire n2122;
wire n2123;
wire n2124;
wire n2125;
wire n2126;
wire n2127;
wire n2128;
wire n2129;
wire n2130;
wire n2131;
wire n2132;
wire n2133;
wire n2134;
wire n2135;
wire n2136;
wire n2137;
wire n2138;
wire n2139;
wire n2140;
wire n2141;
wire n2142;
wire n2143;
wire n2144;
wire n2145;
wire n2146;
wire n2147;
wire n2148;
wire n2149;
wire n2150;
wire n2151;
wire n2152;
wire n2153;
wire n2154;
wire n2155;
wire n2156;
wire n2157;
wire n2158;
wire n2159;
wire n2160;
wire n2161;
wire n2162;
wire n2163;
wire n2164;
wire n2165;
wire n2166;
wire n2167;
wire n2168;
wire n2169;
wire n2170;
wire n2171;
wire n2172;
wire n2173;
wire n2174;
wire n2175;
wire n2176;
wire n2177;
wire n2178;
wire n2179;
wire n2180;
wire n2181;
wire n2182;
wire n2183;
wire n2184;
wire n2185;
wire n2186;
wire n2187;
wire n2188;
wire n2189;
wire n2190;
wire n2191;
wire n2192;
wire n2193;
wire n2194;
wire n2195;
wire n2196;
wire n2197;
wire n2198;
wire n2199;
wire n2200;
wire n2201;
wire n2202;
wire n2203;
wire n2204;
wire n2205;
wire n2206;
wire n2207;
wire n2208;
wire n2209;
wire n2210;
wire n2211;
wire n2212;
wire n2213;
wire n2214;
wire n2215;
wire n2216;
wire n2217;
wire n2218;
wire n2219;
wire n2220;
wire n2221;
wire n2222;
wire n2223;
wire n2224;
wire n2225;
wire n2226;
wire n2227;
wire n2228;
wire n2229;
wire n2230;
wire n2231;
wire n2232;
wire n2233;
wire n2234;
wire n2235;
wire n2236;
wire n2237;
wire n2238;
wire n2239;
wire n2240;
wire n2241;
wire n2242;
wire n2243;
wire n2244;
wire n2245;
wire n2246;
wire n2247;
wire n2248;
wire n2249;
wire n2250;
wire n2251;
wire n2252;
wire n2253;
wire n2254;
wire n2255;
wire n2256;
wire n2257;
wire n2258;
wire n2259;
wire n2260;
wire n2261;
wire n2262;
wire n2263;
wire n2264;
wire n2265;
wire n2266;
wire n2267;
wire n2268;
wire n2269;
wire n2270;
wire n2271;
wire n2272;
wire n2273;
wire n2274;
wire n2275;
wire n2276;
wire n2277;
wire n2278;
wire n2279;
wire n2280;
wire n2281;
wire n2282;
wire n2283;
wire n2284;
wire n2285;
wire n2286;
wire n2287;
wire n2288;
wire n2289;
wire n2290;
wire n2291;
wire n2292;
wire n2293;
wire n2294;
wire n2295;
wire n2296;
wire n2297;
wire n2298;
wire n2299;
wire n2300;
wire n2301;
wire n2302;
wire n2303;
wire n2304;
wire n2305;
wire n2306;
wire n2307;
wire n2308;
wire n2309;
wire n2310;
wire n2311;
wire n2312;
wire n2313;
wire n2314;
wire n2315;
wire n2316;
wire n2317;
wire n2318;
wire n2319;
wire n2320;
wire n2321;
wire n2322;
wire n2323;
wire n2324;
wire n2325;
wire n2326;
wire n2327;
wire n2328;
wire n2329;
wire n2330;
wire n2331;
wire n2332;
wire n2333;
wire n2334;
wire n2335;
wire n2336;
wire n2337;
wire n2338;
wire n2339;
wire n2340;
wire n2341;
wire n2342;
wire n2343;
wire n2344;
wire n2345;
wire n2346;
wire n2347;
wire n2348;
wire n2349;
wire n2350;
wire n2351;
wire n2352;
wire n2353;
wire n2354;
wire n2355;
wire n2356;
wire n2357;
wire n2358;
wire n2359;
wire n2360;
wire n2361;
wire n2362;
wire n2363;
wire n2364;
wire n2365;
wire n2366;
wire n2367;
wire n2368;
wire n2369;
wire n2370;
wire n2371;
wire n2372;
wire n2373;
wire n2374;
wire n2375;
wire n2376;
wire n2377;
wire n2378;
wire n2379;
wire n2380;
wire n2381;
wire n2382;
wire n2383;
wire n2384;
wire n2385;
wire n2386;
wire n2387;
wire n2388;
wire n2389;
wire n2390;
wire n2391;
wire n2392;
wire n2393;
wire n2394;
wire n2395;
wire n2396;
wire n2397;
wire n2398;
wire n2399;
wire n2400;
wire n2401;
wire n2402;
wire n2403;
wire n2404;
wire n2405;
wire n2406;
wire n2407;
wire n2408;
wire n2409;
wire n2410;
wire n2411;
wire n2412;
wire n2413;
wire n2414;
wire n2415;
wire n2416;
wire n2417;
wire n2418;
wire n2419;
wire n2420;
wire n2421;
wire n2422;
wire n2423;
wire n2424;
wire n2425;
wire n2426;
wire n2427;
wire n2428;
wire n2429;
wire n2430;
wire n2431;
wire n2432;
wire n2433;
wire n2434;
wire n2435;
wire n2436;
wire n2437;
wire n2438;
wire n2439;
wire n2440;
wire n2441;
wire n2442;
wire n2443;
wire n2444;
wire n2445;
wire n2446;
wire n2447;
wire n2448;
wire n2449;
wire n2450;
wire n2451;
wire n2452;
wire n2453;
wire n2454;
wire n2455;
wire n2456;
wire n2457;
wire n2458;
wire n2459;
wire n2460;
wire n2461;
wire n2462;
wire n2463;
wire n2464;
wire n2465;
wire n2466;
wire n2467;
wire n2468;
wire n2469;
wire n2470;
wire n2471;
wire n2472;
wire n2473;
wire n2474;
wire n2475;
wire n2476;
wire n2477;
wire n2478;
wire n2479;
wire n2480;
wire n2481;
wire n2482;
wire n2483;
wire n2484;
wire n2485;
wire n2486;
wire n2487;
wire n2488;
wire n2489;
wire n2490;
wire n2491;
wire n2492;
wire n2493;
wire n2494;
wire n2495;
wire n2496;
wire n2497;
wire n2498;
wire n2499;
wire n2500;
wire n2501;
wire n2502;
wire n2503;
wire n2504;
wire n2505;
wire n2506;
wire n2507;
wire n2508;
wire n2509;
wire n2510;
wire n2511;
wire n2512;
wire n2513;
wire n2514;
wire n2515;
wire n2516;
wire n2517;
wire n2518;
wire n2519;
wire n2520;
wire n2521;
wire n2522;
wire n2523;
wire n2524;
wire n2525;
wire n2526;
wire n2527;
wire n2528;
wire n2529;
wire n2530;
wire n2531;
wire n2532;
wire n2533;
wire n2534;
wire n2535;
wire n2536;
wire n2537;
wire n2538;
wire n2539;
wire n2540;
wire n2541;
wire n2542;
wire n2543;
wire n2544;
wire n2545;
wire n2546;
wire n2547;
wire n2548;
wire n2549;
wire n2550;
wire n2551;
wire n2552;
wire n2553;
wire n2554;
wire n2555;
wire n2556;
wire n2557;
wire n2558;
wire n2559;
wire n2560;
wire n2561;
wire n2562;
wire n2563;
wire n2564;
wire n2565;
wire n2566;
wire n2567;
wire n2568;
wire n2569;
wire n2570;
wire n2571;
wire n2572;
wire n2573;
wire n2574;
wire n2575;
wire n2576;
wire n2577;
wire n2578;
wire n2579;
wire n2580;
wire n2581;
wire n2582;
wire n2583;
wire n2584;
wire n2585;
wire n2586;
wire n2587;
wire n2588;
wire n2589;
wire n2590;
wire n2591;
wire n2592;
wire n2593;
wire n2594;
wire n2595;
wire n2596;
wire n2597;
wire n2598;
wire n2599;
wire n2600;
wire n2601;
wire n2602;
wire n2603;
wire n2604;
wire n2605;
wire n2606;
wire n2607;
wire n2608;
wire n2609;
wire n2610;
wire n2611;
wire n2612;
wire n2613;
wire n2614;
wire n2615;
wire n2616;
wire n2617;
wire n2618;
wire n2619;
wire n2620;
wire n2621;
wire n2622;
wire n2623;
wire n2624;
wire n2625;
wire n2626;
wire n2627;
wire n2628;
wire n2629;
wire n2630;
wire n2631;
wire n2632;
wire n2633;
wire n2634;
wire n2635;
wire n2636;
wire n2637;
wire n2638;
wire n2639;
wire n2640;
wire n2641;
wire n2642;
wire n2643;
wire n2644;
wire n2645;
wire n2646;
wire n2647;
wire n2648;
wire n2649;
wire n2650;
wire n2651;
wire n2652;
wire n2653;
wire n2654;
wire n2655;
wire n2656;
wire n2657;
wire n2658;
wire n2659;
wire n2660;
wire n2661;
wire n2662;
wire n2663;
wire n2664;
wire n2665;
wire n2666;
wire n2667;
wire n2668;
wire n2669;
wire n2670;
wire n2671;
wire n2672;
wire n2673;
wire n2674;
wire n2675;
wire n2676;
wire n2677;
wire n2678;
wire n2679;
wire n2680;
wire n2681;
wire n2682;
wire n2683;
wire n2684;
wire n2685;
wire n2686;
wire n2687;
wire n2688;
wire n2689;
wire n2690;
wire n2691;
wire n2692;
wire n2693;
wire n2694;
wire n2695;
wire n2696;
wire n2697;
wire n2698;
wire n2699;
wire n2700;
wire n2701;
wire n2702;
wire n2703;
wire n2704;
wire n2705;
wire n2706;
wire n2707;
wire n2708;
wire n2709;
wire n2710;
wire n2711;
wire n2712;
wire n2713;
wire n2714;
wire n2715;
wire n2716;
wire n2717;
wire n2718;
wire n2719;
wire n2720;
wire n2721;
wire n2722;
wire n2723;
wire n2724;
wire n2725;
wire n2726;
wire n2727;
wire n2728;
wire n2729;
wire n2730;
wire n2731;
wire n2732;
wire n2733;
wire n2734;
wire n2735;
wire n2736;
wire n2737;
wire n2738;
wire n2739;
wire n2740;
wire n2741;
wire n2742;
wire n2743;
wire n2744;
wire n2745;
wire n2746;
wire n2747;
wire n2748;
wire n2749;
wire n2750;
wire n2751;
wire n2752;
wire n2753;
wire n2754;
wire n2755;
wire n2756;
wire n2757;
wire n2758;
wire n2759;
wire n2760;
wire n2761;
wire n2762;
wire n2763;
wire n2764;
wire n2765;
wire n2766;
wire n2767;
wire n2768;
wire n2769;
wire n2770;
wire n2771;
wire n2772;
wire n2773;
wire n2774;
wire n2775;
wire n2776;
wire n2777;
wire n2778;
wire n2779;
wire n2780;
wire n2781;
wire n2782;
wire n2783;
wire n2784;
wire n2785;
wire n2786;
wire n2787;
wire n2788;
wire n2789;
wire n2790;
wire n2791;
wire n2792;
wire n2793;
wire n2794;
wire n2795;
wire n2796;
wire n2797;
wire n2798;
wire n2799;
wire n2800;
wire n2801;
wire n2802;
wire n2803;
wire n2804;
wire n2805;
wire n2806;
wire n2807;
wire n2808;
wire n2809;
wire n2810;
wire n2811;
wire n2812;
wire n2813;
wire n2814;
wire n2815;
wire n2816;
wire n2817;
wire n2818;
wire n2819;
wire n2820;
wire n2821;
wire n2822;
wire n2823;
wire n2824;
wire n2825;
wire n2826;
wire n2827;
wire n2828;
wire n2829;
wire n2830;
wire n2831;
wire n2832;
wire n2833;
wire n2834;
wire n2835;
wire n2836;
wire n2837;
wire n2838;
wire n2839;
wire n2840;
wire n2841;
wire n2842;
wire n2843;
wire n2844;
wire n2845;
wire n2846;
wire n2847;
wire n2848;
wire n2849;
wire n2850;
wire n2851;
wire n2852;
wire n2853;
wire n2854;
wire n2855;
wire n2856;
wire n2857;
wire n2858;
wire n2859;
wire n2860;
wire n2861;
wire n2862;
wire n2863;
wire n2864;
wire n2865;
wire n2866;
wire n2867;
wire n2868;
wire n2869;
wire n2870;
wire n2871;
wire n2872;
wire n2873;
wire n2874;
wire n2875;
wire n2876;
wire n2877;
wire n2878;
wire n2879;
wire n2880;
wire n2881;
wire n2882;
wire n2883;
wire n2884;
wire n2885;
wire n2886;
wire n2887;
wire n2888;
wire n2889;
wire n2890;
wire n2891;
wire n2892;
wire n2893;
wire n2894;
wire n2895;
wire n2896;
wire n2897;
wire n2898;
wire n2899;
wire n2900;
wire n2901;
wire n2902;
wire n2903;
wire n2904;
wire n2905;
wire n2906;
wire n2907;
wire n2908;
wire n2909;
wire n2910;
wire n2911;
wire n2912;
wire n2913;
wire n2914;
wire n2915;
wire n2916;
wire n2917;
wire n2918;
wire n2919;
wire n2920;
wire n2921;
wire n2922;
wire n2923;
wire n2924;
wire n2925;
wire n2926;
wire n2927;
wire n2928;
wire n2929;
wire n2930;
wire n2931;
wire n2932;
wire n2933;
wire n2934;
wire n2935;
wire n2936;
wire n2937;
wire n2938;
wire n2939;
wire n2940;
wire n2941;
wire n2942;
wire n2943;
wire n2944;
wire n2945;
wire n2946;
wire n2947;
wire n2948;
wire n2949;
wire n2950;
wire n2951;
wire n2952;
wire n2953;
wire n2954;
wire n2955;
wire n2956;
wire n2957;
wire n2958;
wire n2959;
wire n2960;
wire n2961;
wire n2962;
wire n2963;
wire n2964;
wire n2965;
wire n2966;
wire n2967;
wire n2968;
wire n2969;
wire n2970;
wire n2971;
wire n2972;
wire n2973;
wire n2974;
wire n2975;
wire n2976;
wire n2977;
wire n2978;
wire n2979;
wire n2980;
wire n2981;
wire n2982;
wire n2983;
wire n2984;
wire n2985;
wire n2986;
wire n2987;
wire n2988;
wire n2989;
wire n2990;
wire n2991;
wire n2992;
wire n2993;
wire n2994;
wire n2995;
wire n2996;
wire n2997;
wire n2998;
wire n2999;
wire n3000;
wire n3001;
wire n3002;
wire n3003;
wire n3004;
wire n3005;
wire n3006;
wire n3007;
wire n3008;
wire n3009;
wire n3010;
wire n3011;
wire n3012;
wire n3013;
wire n3014;
wire n3015;
wire n3016;
wire n3017;
wire n3018;
wire n3019;
wire n3020;
wire n3021;
wire n3022;
wire n3023;
wire n3024;
wire n3025;
wire n3026;
wire n3027;
wire n3028;
wire n3029;
wire n3030;
wire n3031;
wire n3032;
wire n3033;
wire n3034;
wire n3035;
wire n3036;
wire n3037;
wire n3038;
wire n3039;
wire n3040;
wire n3041;
wire n3042;
wire n3043;
wire n3044;
wire n3045;
wire n3046;
wire n3047;
wire n3048;
wire n3049;
wire n3050;
wire n3051;
wire n3052;
wire n3053;
wire n3054;
wire n3055;
wire n3056;
wire n3057;
wire n3058;
wire n3059;
wire n3060;
wire n3061;
wire n3062;
wire n3063;
wire n3064;
wire n3065;
wire n3066;
wire n3067;
wire n3068;
wire n3069;
wire n3070;
wire n3071;
wire n3072;
wire n3073;
wire n3074;
wire n3075;
wire n3076;
wire n3077;
wire n3078;
wire n3079;
wire n3080;
wire n3081;
wire n3082;
wire n3083;
wire n3084;
wire n3085;
wire n3086;
wire n3087;
wire n3088;
wire n3089;
wire n3090;
wire n3091;
wire n3092;
wire n3093;
wire n3094;
wire n3095;
wire n3096;
wire n3097;
wire n3098;
wire n3099;
wire n3100;
wire n3101;
wire n3102;
wire n3103;
wire n3104;
wire n3105;
wire n3106;
wire n3107;
wire n3108;
wire n3109;
wire n3110;
wire n3111;
wire n3112;
wire n3113;
wire n3114;
wire n3115;
wire n3116;
wire n3117;
wire n3118;
wire n3119;
wire n3120;
wire n3121;
wire n3122;
wire n3123;
wire n3124;
wire n3125;
wire n3126;
wire n3127;
wire n3128;
wire n3129;
wire n3130;
wire n3131;
wire n3132;
wire n3133;
wire n3134;
wire n3135;
wire n3136;
wire n3137;
wire n3138;
wire n3139;
xor (out,n0,n1758);
nand (n0,n1,n1757);
or (n1,n2,n276);
nand (n2,n3,n275);
or (n3,n4,n214);
xor (n4,n5,n177);
xor (n5,n6,n110);
or (n6,n7,n109);
and (n7,n8,n59);
xor (n8,n9,n33);
nand (n9,n10,n27);
or (n10,n11,n22);
nand (n11,n12,n19);
nor (n12,n13,n17);
and (n13,n14,n16);
not (n14,n15);
and (n17,n15,n18);
not (n18,n16);
xor (n19,n14,n20);
not (n20,n21);
nor (n22,n23,n25);
and (n23,n20,n24);
and (n25,n21,n26);
not (n26,n24);
or (n27,n12,n28);
nor (n28,n29,n31);
and (n29,n20,n30);
and (n31,n21,n32);
not (n32,n30);
not (n33,n34);
nand (n34,n35,n49);
or (n35,n36,n42);
not (n36,n37);
nand (n37,n38,n41);
or (n38,n16,n39);
not (n39,n40);
or (n41,n18,n40);
not (n42,n43);
nand (n43,n44,n48);
or (n44,n45,n47);
not (n45,n46);
nand (n48,n47,n45);
or (n49,n50,n54);
nand (n50,n42,n51);
nand (n51,n52,n53);
nand (n52,n45,n16);
nand (n53,n46,n18);
nor (n54,n55,n58);
and (n55,n56,n16);
not (n56,n57);
and (n58,n57,n18);
or (n59,n60,n108);
and (n60,n61,n93);
xor (n61,n62,n87);
nand (n62,n63,n81);
or (n63,n64,n72);
not (n64,n65);
nor (n65,n66,n71);
and (n66,n67,n69);
not (n67,n68);
not (n69,n70);
and (n71,n68,n70);
nand (n72,n73,n78);
not (n73,n74);
nand (n74,n75,n77);
or (n75,n20,n76);
nand (n77,n20,n76);
nand (n78,n79,n80);
or (n79,n76,n69);
nand (n80,n69,n76);
nand (n81,n74,n82);
nor (n82,n83,n86);
and (n83,n84,n69);
not (n84,n85);
and (n86,n85,n70);
nand (n87,n88,n92);
or (n88,n89,n50);
nor (n89,n90,n91);
and (n90,n18,n30);
and (n91,n16,n32);
or (n92,n42,n54);
nand (n93,n94,n104);
or (n94,n95,n97);
not (n95,n96);
not (n97,n98);
nor (n98,n99,n101);
not (n99,n100);
nand (n101,n102,n103);
or (n102,n69,n100);
nand (n103,n100,n69);
or (n104,n105,n106);
not (n105,n101);
not (n106,n107);
and (n108,n62,n87);
and (n109,n9,n33);
xor (n110,n111,n166);
xor (n111,n112,n150);
or (n112,n113,n149);
and (n113,n114,n127);
xor (n114,n115,n124);
nand (n115,n116,n118);
or (n116,n72,n117);
not (n117,n82);
or (n118,n73,n119);
nor (n119,n120,n122);
and (n120,n69,n121);
and (n122,n70,n123);
not (n123,n121);
nand (n124,n125,n126);
or (n125,n106,n97);
nand (n126,n101,n68);
nand (n127,n128,n147);
or (n128,n129,n142);
not (n129,n130);
nor (n130,n131,n137);
nor (n131,n132,n135);
and (n132,n133,n134);
not (n134,n47);
and (n135,n47,n136);
not (n136,n133);
nand (n137,n138,n141);
or (n138,n139,n133);
not (n139,n140);
nand (n141,n133,n139);
nor (n142,n143,n145);
and (n143,n134,n144);
and (n145,n47,n146);
not (n146,n144);
or (n147,n148,n134);
not (n148,n137);
and (n149,n115,n124);
xor (n150,n151,n160);
xor (n151,n152,n154);
nand (n152,n153,n47);
or (n153,n137,n130);
nand (n154,n155,n156);
or (n155,n50,n36);
or (n156,n42,n157);
nor (n157,n158,n159);
and (n158,n18,n144);
and (n159,n16,n146);
nand (n160,n161,n162);
or (n161,n72,n119);
or (n162,n73,n163);
nor (n163,n164,n165);
and (n164,n69,n24);
and (n165,n70,n26);
xor (n166,n167,n34);
xor (n167,n168,n171);
nand (n168,n169,n170);
or (n169,n97,n67);
or (n170,n105,n84);
nand (n171,n172,n173);
or (n172,n11,n28);
or (n173,n12,n174);
nor (n174,n175,n176);
and (n175,n20,n57);
and (n176,n21,n56);
or (n177,n178,n213);
and (n178,n179,n212);
xor (n179,n180,n211);
or (n180,n181,n210);
and (n181,n182,n204);
xor (n182,n183,n197);
nand (n183,n184,n140);
or (n184,n185,n192);
not (n185,n186);
nand (n186,n187,n191);
nand (n187,n188,n190);
or (n188,n189,n139);
nand (n190,n139,n189);
not (n191,n192);
nand (n192,n193,n196);
or (n193,n194,n189);
not (n194,n195);
nand (n196,n189,n194);
nand (n197,n198,n202);
or (n198,n199,n129);
nor (n199,n200,n201);
and (n200,n39,n47);
and (n201,n40,n134);
nand (n202,n203,n137);
not (n203,n142);
nand (n204,n205,n209);
or (n205,n206,n11);
nor (n206,n207,n208);
and (n207,n121,n20);
and (n208,n21,n123);
or (n209,n12,n22);
and (n210,n183,n197);
xor (n211,n114,n127);
xor (n212,n8,n59);
and (n213,n180,n211);
or (n214,n215,n274);
and (n215,n216,n252);
xor (n216,n217,n251);
or (n217,n218,n250);
and (n218,n219,n249);
xor (n219,n220,n226);
nand (n220,n221,n225);
or (n221,n129,n222);
nor (n222,n223,n224);
and (n223,n56,n47);
and (n224,n57,n134);
or (n225,n148,n199);
or (n226,n227,n248);
and (n227,n228,n242);
xor (n228,n229,n235);
nand (n229,n230,n234);
or (n230,n11,n231);
nor (n231,n232,n233);
and (n232,n85,n20);
and (n233,n21,n84);
or (n234,n206,n12);
nand (n235,n236,n237);
or (n236,n64,n73);
nand (n237,n238,n239);
not (n238,n72);
nor (n239,n240,n241);
and (n240,n106,n69);
and (n241,n107,n70);
nand (n242,n243,n247);
or (n243,n186,n244);
nor (n244,n245,n246);
and (n245,n139,n144);
and (n246,n140,n146);
or (n247,n191,n139);
and (n248,n229,n235);
xor (n249,n61,n93);
and (n250,n220,n226);
xor (n251,n179,n212);
or (n252,n253,n273);
and (n253,n254,n272);
xor (n254,n255,n256);
xor (n255,n182,n204);
or (n256,n257,n271);
and (n257,n258,n270);
xor (n258,n259,n264);
nand (n259,n260,n263);
or (n260,n97,n261);
not (n261,n262);
or (n263,n105,n95);
nand (n264,n265,n269);
or (n265,n266,n50);
nor (n266,n267,n268);
and (n267,n18,n24);
and (n268,n16,n26);
or (n269,n42,n89);
not (n270,n220);
and (n271,n259,n264);
xor (n272,n219,n249);
and (n273,n255,n256);
and (n274,n217,n251);
nand (n275,n214,n4);
nand (n276,n277,n1752);
or (n277,n278,n528);
not (n278,n279);
nor (n279,n280,n523);
nor (n280,n281,n514);
or (n281,n282,n513);
and (n282,n283,n418);
xor (n283,n284,n343);
xor (n284,n285,n342);
xor (n285,n286,n312);
or (n286,n287,n311);
and (n287,n288,n305);
xor (n288,n289,n298);
nand (n289,n290,n295);
or (n290,n291,n11);
not (n291,n292);
nand (n292,n293,n294);
or (n293,n67,n21);
or (n294,n68,n20);
nand (n295,n296,n297);
not (n296,n231);
not (n297,n12);
nand (n298,n299,n304);
or (n299,n300,n129);
not (n300,n301);
nor (n301,n302,n303);
and (n302,n32,n134);
and (n303,n30,n47);
or (n304,n148,n222);
nand (n305,n306,n309);
or (n306,n72,n307);
not (n307,n308);
xnor (n308,n95,n70);
or (n309,n73,n310);
not (n310,n239);
and (n311,n289,n298);
or (n312,n313,n341);
and (n313,n314,n335);
xor (n314,n315,n328);
nand (n315,n316,n195);
or (n316,n317,n323);
nand (n317,n318,n322);
or (n318,n319,n321);
not (n319,n320);
nand (n322,n321,n319);
nor (n323,n317,n324);
nor (n324,n325,n327);
and (n325,n326,n195);
not (n326,n321);
and (n327,n321,n194);
nand (n328,n329,n334);
or (n329,n186,n330);
not (n330,n331);
nor (n331,n332,n333);
and (n332,n39,n139);
and (n333,n40,n140);
or (n334,n191,n244);
nand (n335,n336,n340);
or (n336,n50,n337);
nor (n337,n338,n339);
and (n338,n123,n16);
and (n339,n121,n18);
or (n340,n42,n266);
and (n341,n315,n328);
xor (n342,n228,n242);
xor (n343,n344,n389);
xor (n344,n345,n346);
xor (n345,n258,n270);
or (n346,n347,n388);
and (n347,n348,n362);
xor (n348,n349,n354);
nand (n349,n350,n353);
or (n350,n97,n351);
not (n351,n352);
or (n353,n105,n261);
nand (n354,n355,n361);
or (n355,n356,n360);
not (n356,n357);
nor (n357,n358,n359);
and (n358,n144,n195);
and (n359,n146,n194);
not (n360,n323);
nand (n361,n317,n195);
or (n362,n363,n387);
and (n363,n364,n379);
xor (n364,n365,n372);
nand (n365,n366,n371);
or (n366,n367,n186);
not (n367,n368);
nor (n368,n369,n370);
and (n369,n57,n140);
and (n370,n56,n139);
nand (n371,n192,n331);
nand (n372,n373,n378);
or (n373,n374,n50);
not (n374,n375);
nor (n375,n376,n377);
and (n376,n84,n18);
and (n377,n85,n16);
or (n378,n42,n337);
nand (n379,n380,n381);
or (n380,n291,n12);
nand (n381,n382,n386);
not (n382,n383);
nor (n383,n384,n385);
and (n384,n20,n107);
and (n385,n106,n21);
not (n386,n11);
and (n387,n365,n372);
and (n388,n349,n354);
or (n389,n390,n417);
and (n390,n391,n416);
xor (n391,n392,n415);
or (n392,n393,n414);
and (n393,n394,n409);
xor (n394,n395,n402);
nand (n395,n396,n401);
or (n396,n397,n129);
not (n397,n398);
nor (n398,n399,n400);
and (n399,n26,n134);
and (n400,n24,n47);
nand (n401,n137,n301);
nand (n402,n403,n408);
or (n403,n404,n72);
not (n404,n405);
nand (n405,n406,n407);
or (n406,n70,n261);
or (n407,n69,n262);
nand (n408,n74,n308);
nand (n409,n410,n413);
or (n410,n411,n97);
not (n411,n412);
nand (n413,n101,n352);
and (n414,n395,n402);
xor (n415,n288,n305);
xor (n416,n314,n335);
and (n417,n392,n415);
or (n418,n419,n512);
and (n419,n420,n482);
xor (n420,n421,n422);
xor (n421,n348,n362);
or (n422,n423,n481);
and (n423,n424,n458);
xor (n424,n425,n426);
not (n425,n354);
or (n426,n427,n457);
and (n427,n428,n450);
xor (n428,n429,n443);
nand (n429,n430,n320);
or (n430,n431,n437);
nand (n431,n432,n436);
or (n432,n433,n435);
not (n433,n434);
nand (n436,n433,n435);
not (n437,n438);
nand (n438,n439,n440);
not (n439,n431);
nand (n440,n441,n442);
or (n441,n320,n433);
nand (n442,n433,n320);
nand (n443,n444,n449);
or (n444,n445,n360);
not (n445,n446);
nand (n446,n447,n448);
or (n447,n40,n194);
nand (n448,n194,n40);
nand (n449,n357,n317);
nand (n450,n451,n456);
or (n451,n452,n129);
not (n452,n453);
nand (n453,n454,n455);
or (n454,n47,n123);
or (n455,n134,n121);
nand (n456,n137,n398);
and (n457,n429,n443);
or (n458,n459,n480);
and (n459,n460,n473);
xor (n460,n461,n466);
nand (n461,n462,n465);
or (n462,n463,n97);
not (n463,n464);
nand (n465,n101,n412);
nand (n466,n467,n472);
or (n467,n468,n50);
not (n468,n469);
nor (n469,n470,n471);
and (n470,n67,n18);
and (n471,n68,n16);
nand (n472,n43,n375);
nand (n473,n474,n479);
or (n474,n186,n475);
not (n475,n476);
nor (n476,n477,n478);
and (n477,n32,n139);
and (n478,n30,n140);
or (n479,n191,n367);
and (n480,n461,n466);
and (n481,n425,n426);
or (n482,n483,n511);
and (n483,n484,n487);
xor (n484,n485,n486);
xor (n485,n394,n409);
xor (n486,n364,n379);
or (n487,n488,n510);
and (n488,n489,n503);
xor (n489,n490,n496);
nand (n490,n491,n495);
or (n491,n492,n11);
nor (n492,n493,n494);
and (n493,n21,n95);
and (n494,n20,n96);
nand (n495,n382,n297);
nand (n496,n497,n502);
or (n497,n498,n72);
not (n498,n499);
nor (n499,n500,n501);
and (n500,n351,n69);
and (n501,n352,n70);
nand (n502,n74,n405);
not (n503,n504);
nor (n504,n505,n509);
and (n505,n437,n506);
nor (n506,n507,n508);
and (n507,n146,n319);
and (n508,n144,n320);
nor (n509,n439,n319);
and (n510,n490,n496);
and (n511,n485,n486);
and (n512,n421,n422);
and (n513,n284,n343);
xor (n514,n515,n520);
xor (n515,n516,n519);
or (n516,n517,n518);
and (n517,n285,n342);
and (n518,n286,n312);
xor (n519,n254,n272);
or (n520,n521,n522);
and (n521,n344,n389);
and (n522,n345,n346);
nor (n523,n524,n525);
xor (n524,n216,n252);
or (n525,n526,n527);
and (n526,n515,n520);
and (n527,n516,n519);
not (n528,n529);
nand (n529,n530,n1233);
nor (n530,n531,n1219);
and (n531,n532,n894);
and (n532,n533,n877);
nor (n533,n534,n789);
nor (n534,n535,n709);
xor (n535,n536,n617);
xor (n536,n537,n564);
or (n537,n538,n563);
and (n538,n539,n542);
xor (n539,n540,n541);
xor (n540,n460,n473);
xor (n541,n489,n503);
or (n542,n543,n562);
and (n543,n544,n552);
xor (n544,n545,n504);
nand (n545,n546,n551);
or (n546,n547,n72);
not (n547,n548);
nor (n548,n549,n550);
and (n549,n411,n69);
and (n550,n412,n70);
nand (n551,n74,n499);
nand (n552,n553,n435);
nor (n553,n554,n558);
and (n554,n185,n555);
nor (n555,n556,n557);
and (n556,n123,n139);
and (n557,n121,n140);
and (n558,n192,n559);
nor (n559,n560,n561);
and (n560,n26,n139);
and (n561,n24,n140);
and (n562,n545,n504);
and (n563,n540,n541);
xor (n564,n565,n616);
xor (n565,n566,n567);
xor (n566,n424,n458);
or (n567,n568,n615);
and (n568,n569,n614);
xor (n569,n570,n591);
or (n570,n571,n590);
and (n571,n572,n584);
xor (n572,n573,n580);
nand (n573,n574,n579);
or (n574,n575,n50);
not (n575,n576);
nand (n576,n577,n578);
or (n577,n107,n18);
nand (n578,n18,n107);
nand (n579,n469,n43);
nand (n580,n581,n583);
or (n581,n582,n186);
not (n582,n559);
nand (n583,n192,n476);
nand (n584,n585,n589);
or (n585,n11,n586);
nor (n586,n587,n588);
and (n587,n262,n20);
and (n588,n21,n261);
or (n589,n492,n12);
and (n590,n573,n580);
or (n591,n592,n613);
and (n592,n593,n606);
xor (n593,n594,n601);
nand (n594,n595,n600);
or (n595,n596,n360);
not (n596,n597);
nor (n597,n598,n599);
and (n598,n56,n194);
and (n599,n57,n195);
nand (n600,n446,n317);
nand (n601,n602,n605);
or (n602,n603,n97);
not (n603,n604);
nand (n605,n101,n464);
nand (n606,n607,n612);
or (n607,n608,n129);
not (n608,n609);
nor (n609,n610,n611);
and (n610,n84,n134);
and (n611,n85,n47);
nand (n612,n137,n453);
and (n613,n594,n601);
xor (n614,n428,n450);
and (n615,n570,n591);
xor (n616,n484,n487);
or (n617,n618,n708);
and (n618,n619,n673);
xor (n619,n620,n621);
xor (n620,n569,n614);
or (n621,n622,n672);
and (n622,n623,n671);
xor (n623,n624,n648);
or (n624,n625,n647);
and (n625,n626,n639);
xor (n626,n627,n634);
nand (n627,n628,n633);
or (n628,n629,n72);
not (n629,n630);
nor (n630,n631,n632);
and (n631,n463,n69);
and (n632,n464,n70);
nand (n633,n548,n74);
nand (n634,n635,n638);
or (n635,n636,n97);
not (n636,n637);
nand (n638,n101,n604);
nand (n639,n640,n642);
or (n640,n641,n439);
not (n641,n506);
or (n642,n438,n643);
not (n643,n644);
or (n644,n645,n646);
and (n645,n39,n320);
and (n646,n40,n319);
and (n647,n627,n634);
or (n648,n649,n670);
and (n649,n650,n664);
xor (n650,n651,n658);
nand (n651,n652,n657);
or (n652,n653,n129);
not (n653,n654);
nor (n654,n655,n656);
and (n655,n67,n134);
and (n656,n68,n47);
nand (n657,n137,n609);
nand (n658,n659,n663);
or (n659,n660,n360);
nor (n660,n661,n662);
and (n661,n32,n195);
and (n662,n30,n194);
nand (n663,n597,n317);
nand (n664,n665,n669);
or (n665,n50,n666);
nor (n666,n667,n668);
and (n667,n18,n96);
and (n668,n16,n95);
or (n669,n42,n575);
and (n670,n651,n658);
xor (n671,n572,n584);
and (n672,n624,n648);
or (n673,n674,n707);
and (n674,n675,n678);
xor (n675,n676,n677);
xor (n676,n593,n606);
xor (n677,n544,n552);
and (n678,n679,n701);
or (n679,n680,n700);
and (n680,n681,n695);
xor (n681,n682,n688);
nand (n682,n683,n687);
or (n683,n684,n186);
nor (n684,n685,n686);
and (n685,n84,n140);
and (n686,n85,n139);
nand (n687,n555,n192);
nand (n688,n689,n694);
or (n689,n690,n72);
not (n690,n691);
nand (n691,n692,n693);
or (n692,n70,n603);
or (n693,n69,n604);
nand (n694,n74,n630);
nand (n695,n696,n699);
or (n696,n697,n97);
not (n697,n698);
nand (n699,n101,n637);
and (n700,n682,n688);
nand (n701,n702,n706);
or (n702,n11,n703);
nor (n703,n704,n705);
and (n704,n20,n352);
and (n705,n21,n351);
or (n706,n12,n586);
and (n707,n676,n677);
and (n708,n620,n621);
or (n709,n710,n788);
and (n710,n711,n714);
xor (n711,n712,n713);
xor (n712,n539,n542);
xor (n713,n619,n673);
or (n714,n715,n787);
and (n715,n716,n751);
xor (n716,n717,n718);
xor (n717,n623,n671);
or (n718,n719,n750);
and (n719,n720,n748);
xor (n720,n721,n747);
or (n721,n722,n746);
and (n722,n723,n738);
xor (n723,n724,n731);
nand (n724,n725,n730);
or (n725,n726,n438);
not (n726,n727);
nor (n727,n728,n729);
and (n728,n56,n319);
and (n729,n57,n320);
nand (n730,n431,n644);
nand (n731,n732,n737);
or (n732,n733,n129);
not (n733,n734);
nand (n734,n735,n736);
or (n735,n47,n106);
or (n736,n134,n107);
nand (n737,n137,n654);
nand (n738,n739,n744);
or (n739,n360,n740);
not (n740,n741);
nor (n741,n742,n743);
and (n742,n194,n26);
and (n743,n24,n195);
or (n744,n660,n745);
not (n745,n317);
and (n746,n724,n731);
xor (n747,n650,n664);
nand (n748,n749,n552);
or (n749,n435,n553);
and (n750,n721,n747);
or (n751,n752,n786);
and (n752,n753,n785);
xor (n753,n754,n755);
xor (n754,n626,n639);
or (n755,n756,n784);
and (n756,n757,n773);
xor (n757,n758,n766);
nand (n758,n759,n764);
or (n759,n760,n50);
not (n760,n761);
nor (n761,n762,n763);
and (n762,n261,n18);
and (n763,n262,n16);
nand (n764,n765,n43);
not (n765,n666);
nand (n766,n767,n772);
or (n767,n768,n11);
not (n768,n769);
nand (n769,n770,n771);
or (n770,n21,n411);
or (n771,n20,n412);
or (n772,n12,n703);
nand (n773,n774,n783);
or (n774,n775,n778);
nand (n775,n776,n435);
not (n776,n777);
not (n778,n779);
nor (n779,n780,n782);
and (n780,n146,n781);
not (n781,n435);
and (n782,n144,n435);
or (n783,n781,n776);
and (n784,n758,n766);
xor (n785,n679,n701);
and (n786,n754,n755);
and (n787,n717,n718);
and (n788,n712,n713);
nor (n789,n790,n791);
xor (n790,n711,n714);
or (n791,n792,n876);
and (n792,n793,n875);
xor (n793,n794,n795);
xor (n794,n675,n678);
or (n795,n796,n874);
and (n796,n797,n873);
xor (n797,n798,n866);
or (n798,n799,n865);
and (n799,n800,n842);
xor (n800,n801,n819);
or (n801,n802,n818);
and (n802,n803,n811);
xor (n803,n804,n805);
and (n804,n101,n698);
nand (n805,n806,n807);
or (n806,n776,n778);
or (n807,n808,n775);
nor (n808,n809,n810);
and (n809,n781,n40);
and (n810,n435,n39);
nand (n811,n812,n817);
or (n812,n438,n813);
not (n813,n814);
nor (n814,n815,n816);
and (n815,n32,n319);
and (n816,n30,n320);
nand (n817,n431,n727);
and (n818,n804,n805);
or (n819,n820,n841);
and (n820,n821,n835);
xor (n821,n822,n829);
nand (n822,n823,n828);
or (n823,n824,n360);
not (n824,n825);
nand (n825,n826,n827);
or (n826,n195,n123);
or (n827,n194,n121);
nand (n828,n741,n317);
nand (n829,n830,n834);
or (n830,n831,n50);
nor (n831,n832,n833);
and (n832,n351,n16);
and (n833,n352,n18);
nand (n834,n761,n43);
nand (n835,n836,n837);
or (n836,n768,n12);
or (n837,n11,n838);
nor (n838,n839,n840);
and (n839,n464,n20);
and (n840,n21,n463);
and (n841,n822,n829);
or (n842,n843,n864);
and (n843,n844,n858);
xor (n844,n845,n852);
nand (n845,n846,n851);
or (n846,n847,n72);
not (n847,n848);
nand (n848,n849,n850);
or (n849,n70,n636);
or (n850,n69,n637);
nand (n851,n691,n74);
nand (n852,n853,n857);
or (n853,n186,n854);
nor (n854,n855,n856);
and (n855,n67,n140);
and (n856,n68,n139);
or (n857,n191,n684);
nand (n858,n859,n863);
or (n859,n129,n860);
nor (n860,n861,n862);
and (n861,n95,n47);
and (n862,n96,n134);
or (n863,n148,n733);
and (n864,n845,n852);
and (n865,n801,n819);
or (n866,n867,n872);
and (n867,n868,n871);
xor (n868,n869,n870);
xor (n869,n681,n695);
xor (n870,n723,n738);
xor (n871,n757,n773);
and (n872,n869,n870);
xor (n873,n720,n748);
and (n874,n798,n866);
xor (n875,n716,n751);
and (n876,n794,n795);
nor (n877,n878,n889);
nor (n878,n879,n886);
xor (n879,n880,n883);
xor (n880,n881,n882);
xor (n881,n391,n416);
xor (n882,n420,n482);
or (n883,n884,n885);
and (n884,n565,n616);
and (n885,n566,n567);
or (n886,n887,n888);
and (n887,n536,n617);
and (n888,n537,n564);
nor (n889,n890,n891);
xor (n890,n283,n418);
or (n891,n892,n893);
and (n892,n880,n883);
and (n893,n881,n882);
nand (n894,n895,n1213);
or (n895,n896,n1195);
not (n896,n897);
nor (n897,n898,n1194);
and (n898,n899,n1135);
nand (n899,n900,n1043);
xor (n900,n901,n1030);
xor (n901,n902,n903);
xor (n902,n868,n871);
or (n903,n904,n1029);
and (n904,n905,n1000);
xor (n905,n906,n953);
or (n906,n907,n952);
and (n907,n908,n928);
xor (n908,n909,n915);
nand (n909,n910,n914);
or (n910,n11,n911);
nor (n911,n912,n913);
and (n912,n20,n604);
and (n913,n21,n603);
or (n914,n12,n838);
xor (n915,n916,n922);
nor (n916,n917,n69);
nor (n917,n918,n920);
and (n918,n919,n20);
nand (n919,n698,n76);
and (n920,n697,n921);
not (n921,n76);
nand (n922,n923,n927);
or (n923,n924,n775);
nor (n924,n925,n926);
and (n925,n56,n435);
and (n926,n57,n781);
or (n927,n808,n776);
or (n928,n929,n951);
and (n929,n930,n940);
xor (n930,n931,n932);
nor (n931,n73,n697);
nand (n932,n933,n938);
or (n933,n775,n934);
not (n934,n935);
nor (n935,n936,n937);
and (n936,n32,n781);
and (n937,n30,n435);
nand (n938,n939,n777);
not (n939,n924);
nand (n940,n941,n946);
or (n941,n438,n942);
not (n942,n943);
nand (n943,n944,n945);
or (n944,n320,n123);
or (n945,n319,n121);
or (n946,n439,n947);
not (n947,n948);
nand (n948,n949,n950);
or (n949,n320,n26);
or (n950,n319,n24);
and (n951,n931,n932);
and (n952,n909,n915);
xor (n953,n954,n977);
xor (n954,n955,n956);
and (n955,n916,n922);
or (n956,n957,n976);
and (n957,n958,n969);
xor (n958,n959,n962);
nand (n959,n960,n961);
or (n960,n947,n438);
nand (n961,n431,n814);
nand (n962,n963,n968);
or (n963,n964,n72);
not (n964,n965);
nand (n965,n966,n967);
or (n966,n69,n698);
or (n967,n70,n697);
nand (n968,n848,n74);
nand (n969,n970,n975);
or (n970,n186,n971);
not (n971,n972);
nor (n972,n973,n974);
and (n973,n106,n139);
and (n974,n107,n140);
or (n975,n191,n854);
and (n976,n959,n962);
or (n977,n978,n999);
and (n978,n979,n993);
xor (n979,n980,n987);
nand (n980,n981,n986);
or (n981,n982,n129);
not (n982,n983);
nor (n983,n984,n985);
and (n984,n261,n134);
and (n985,n262,n47);
or (n986,n860,n148);
nand (n987,n988,n992);
or (n988,n989,n360);
nor (n989,n990,n991);
and (n990,n194,n85);
and (n991,n195,n84);
nand (n992,n317,n825);
nand (n993,n994,n998);
or (n994,n50,n995);
nor (n995,n996,n997);
and (n996,n18,n412);
and (n997,n16,n411);
or (n998,n42,n831);
and (n999,n980,n987);
or (n1000,n1001,n1028);
and (n1001,n1002,n1027);
xor (n1002,n1003,n1026);
or (n1003,n1004,n1025);
and (n1004,n1005,n1019);
xor (n1005,n1006,n1013);
nand (n1006,n1007,n1012);
or (n1007,n1008,n186);
not (n1008,n1009);
nand (n1009,n1010,n1011);
or (n1010,n140,n95);
or (n1011,n139,n96);
nand (n1012,n192,n972);
nand (n1013,n1014,n1018);
or (n1014,n129,n1015);
nor (n1015,n1016,n1017);
and (n1016,n134,n352);
and (n1017,n47,n351);
nand (n1018,n137,n983);
nand (n1019,n1020,n1024);
or (n1020,n360,n1021);
nor (n1021,n1022,n1023);
and (n1022,n194,n68);
and (n1023,n195,n67);
or (n1024,n989,n745);
and (n1025,n1006,n1013);
xor (n1026,n979,n993);
xor (n1027,n958,n969);
and (n1028,n1003,n1026);
and (n1029,n906,n953);
xor (n1030,n1031,n1036);
xor (n1031,n1032,n1035);
or (n1032,n1033,n1034);
and (n1033,n954,n977);
and (n1034,n955,n956);
xor (n1035,n800,n842);
or (n1036,n1037,n1042);
and (n1037,n1038,n1041);
xor (n1038,n1039,n1040);
xor (n1039,n821,n835);
xor (n1040,n803,n811);
xor (n1041,n844,n858);
and (n1042,n1039,n1040);
or (n1043,n1044,n1134);
and (n1044,n1045,n1133);
xor (n1045,n1046,n1047);
xor (n1046,n1038,n1041);
or (n1047,n1048,n1132);
and (n1048,n1049,n1080);
xor (n1049,n1050,n1079);
or (n1050,n1051,n1078);
and (n1051,n1052,n1066);
xor (n1052,n1053,n1060);
nand (n1053,n1054,n1058);
or (n1054,n1055,n50);
nor (n1055,n1056,n1057);
and (n1056,n463,n16);
and (n1057,n464,n18);
nand (n1058,n1059,n43);
not (n1059,n995);
nand (n1060,n1061,n1065);
or (n1061,n1062,n11);
nor (n1062,n1063,n1064);
and (n1063,n20,n637);
and (n1064,n21,n636);
or (n1065,n12,n911);
and (n1066,n1067,n1072);
nor (n1067,n1068,n20);
nor (n1068,n1069,n1071);
and (n1069,n1070,n18);
nand (n1070,n698,n15);
and (n1071,n697,n14);
nand (n1072,n1073,n1074);
or (n1073,n776,n934);
or (n1074,n1075,n775);
nor (n1075,n1076,n1077);
and (n1076,n26,n435);
and (n1077,n24,n781);
and (n1078,n1053,n1060);
xor (n1079,n908,n928);
or (n1080,n1081,n1131);
and (n1081,n1082,n1130);
xor (n1082,n1083,n1108);
or (n1083,n1084,n1107);
and (n1084,n1085,n1100);
xor (n1085,n1086,n1093);
nand (n1086,n1087,n1092);
or (n1087,n1088,n438);
not (n1088,n1089);
nor (n1089,n1090,n1091);
and (n1090,n84,n319);
and (n1091,n85,n320);
nand (n1092,n943,n431);
nand (n1093,n1094,n1099);
or (n1094,n1095,n186);
not (n1095,n1096);
nand (n1096,n1097,n1098);
or (n1097,n140,n261);
or (n1098,n139,n262);
nand (n1099,n192,n1009);
nand (n1100,n1101,n1106);
or (n1101,n129,n1102);
not (n1102,n1103);
nand (n1103,n1104,n1105);
or (n1104,n47,n411);
or (n1105,n134,n412);
or (n1106,n148,n1015);
and (n1107,n1086,n1093);
or (n1108,n1109,n1129);
and (n1109,n1110,n1123);
xor (n1110,n1111,n1117);
nand (n1111,n1112,n1116);
or (n1112,n360,n1113);
nor (n1113,n1114,n1115);
and (n1114,n194,n107);
and (n1115,n195,n106);
or (n1116,n1021,n745);
nand (n1117,n1118,n1122);
or (n1118,n50,n1119);
nor (n1119,n1120,n1121);
and (n1120,n18,n604);
and (n1121,n16,n603);
or (n1122,n1055,n42);
nand (n1123,n1124,n1128);
or (n1124,n11,n1125);
nor (n1125,n1126,n1127);
and (n1126,n697,n21);
and (n1127,n698,n20);
or (n1128,n1062,n12);
and (n1129,n1111,n1117);
xor (n1130,n930,n940);
and (n1131,n1083,n1108);
and (n1132,n1050,n1079);
xor (n1133,n905,n1000);
and (n1134,n1046,n1047);
nand (n1135,n1136,n1137);
xor (n1136,n1045,n1133);
or (n1137,n1138,n1193);
and (n1138,n1139,n1192);
xor (n1139,n1140,n1141);
xor (n1140,n1002,n1027);
or (n1141,n1142,n1191);
and (n1142,n1143,n1146);
xor (n1143,n1144,n1145);
xor (n1144,n1005,n1019);
xor (n1145,n1052,n1066);
or (n1146,n1147,n1190);
and (n1147,n1148,n1168);
xor (n1148,n1149,n1150);
xor (n1149,n1067,n1072);
or (n1150,n1151,n1167);
and (n1151,n1152,n1161);
xor (n1152,n1153,n1154);
and (n1153,n297,n698);
nand (n1154,n1155,n1160);
or (n1155,n1156,n438);
not (n1156,n1157);
nand (n1157,n1158,n1159);
or (n1158,n320,n67);
or (n1159,n319,n68);
nand (n1160,n431,n1089);
nand (n1161,n1162,n1163);
or (n1162,n1095,n191);
or (n1163,n186,n1164);
nor (n1164,n1165,n1166);
and (n1165,n351,n140);
and (n1166,n352,n139);
and (n1167,n1153,n1154);
or (n1168,n1169,n1189);
and (n1169,n1170,n1183);
xor (n1170,n1171,n1177);
nand (n1171,n1172,n1176);
or (n1172,n1173,n129);
nor (n1173,n1174,n1175);
and (n1174,n463,n47);
and (n1175,n464,n134);
nand (n1176,n1103,n137);
nand (n1177,n1178,n1182);
or (n1178,n1179,n775);
nor (n1179,n1180,n1181);
and (n1180,n781,n121);
and (n1181,n435,n123);
or (n1182,n1075,n776);
nand (n1183,n1184,n1188);
or (n1184,n1185,n50);
nor (n1185,n1186,n1187);
and (n1186,n18,n637);
and (n1187,n16,n636);
or (n1188,n1119,n42);
and (n1189,n1171,n1177);
and (n1190,n1149,n1150);
and (n1191,n1144,n1145);
xor (n1192,n1049,n1080);
and (n1193,n1140,n1141);
nor (n1194,n900,n1043);
not (n1195,n1196);
nor (n1196,n1197,n1208);
nor (n1197,n1198,n1199);
xor (n1198,n793,n875);
or (n1199,n1200,n1207);
and (n1200,n1201,n1206);
xor (n1201,n1202,n1203);
xor (n1202,n753,n785);
or (n1203,n1204,n1205);
and (n1204,n1031,n1036);
and (n1205,n1032,n1035);
xor (n1206,n797,n873);
and (n1207,n1202,n1203);
nor (n1208,n1209,n1210);
xor (n1209,n1201,n1206);
or (n1210,n1211,n1212);
and (n1211,n901,n1030);
and (n1212,n902,n903);
nor (n1213,n1214,n1218);
and (n1214,n1215,n1216);
not (n1215,n1197);
not (n1216,n1217);
nand (n1217,n1209,n1210);
and (n1218,n1198,n1199);
nand (n1219,n1220,n1227);
or (n1220,n1221,n1222);
not (n1221,n877);
not (n1222,n1223);
nor (n1223,n1224,n534);
and (n1224,n1225,n1226);
nand (n1225,n709,n535);
nand (n1226,n790,n791);
nor (n1227,n1228,n1232);
and (n1228,n1229,n1230);
not (n1229,n889);
not (n1230,n1231);
nand (n1231,n879,n886);
and (n1232,n890,n891);
nand (n1233,n532,n1234,n1237);
and (n1234,n1196,n1235);
nor (n1235,n1194,n1236);
nor (n1236,n1136,n1137);
nand (n1237,n1238,n1739);
or (n1238,n1239,n1675);
not (n1239,n1240);
nand (n1240,n1241,n1664,n1674);
nand (n1241,n1242,n1420,n1524);
nand (n1242,n1243,n1384);
not (n1243,n1244);
xor (n1244,n1245,n1343);
xor (n1245,n1246,n1281);
xor (n1246,n1247,n1263);
xor (n1247,n1248,n1254);
nand (n1248,n1249,n1253);
or (n1249,n50,n1250);
nor (n1250,n1251,n1252);
and (n1251,n697,n16);
and (n1252,n18,n698);
or (n1253,n42,n1185);
nand (n1254,n1255,n1259);
or (n1255,n360,n1256);
nor (n1256,n1257,n1258);
and (n1257,n194,n262);
and (n1258,n195,n261);
or (n1259,n1260,n745);
nor (n1260,n1261,n1262);
and (n1261,n194,n96);
and (n1262,n195,n95);
nand (n1263,n1264,n1280);
or (n1264,n1265,n1272);
not (n1265,n1266);
nand (n1266,n1267,n16);
nand (n1267,n1268,n1269);
or (n1268,n698,n46);
nand (n1269,n1270,n134);
not (n1270,n1271);
and (n1271,n698,n46);
not (n1272,n1273);
nand (n1273,n1274,n1279);
or (n1274,n1275,n438);
not (n1275,n1276);
nand (n1276,n1277,n1278);
or (n1277,n320,n106);
or (n1278,n319,n107);
nand (n1279,n431,n1157);
or (n1280,n1273,n1266);
xor (n1281,n1282,n1332);
xor (n1282,n1283,n1304);
or (n1283,n1284,n1303);
and (n1284,n1285,n1293);
xor (n1285,n1286,n1287);
and (n1286,n43,n698);
nand (n1287,n1288,n1292);
or (n1288,n1289,n438);
nor (n1289,n1290,n1291);
and (n1290,n95,n320);
and (n1291,n96,n319);
nand (n1292,n431,n1276);
nand (n1293,n1294,n1299);
or (n1294,n186,n1295);
not (n1295,n1296);
nor (n1296,n1297,n1298);
and (n1297,n463,n139);
and (n1298,n464,n140);
or (n1299,n191,n1300);
nor (n1300,n1301,n1302);
and (n1301,n412,n139);
and (n1302,n411,n140);
and (n1303,n1286,n1287);
or (n1304,n1305,n1331);
and (n1305,n1306,n1325);
xor (n1306,n1307,n1316);
nand (n1307,n1308,n1312);
or (n1308,n129,n1309);
nor (n1309,n1310,n1311);
and (n1310,n636,n47);
and (n1311,n637,n134);
or (n1312,n148,n1313);
nor (n1313,n1314,n1315);
and (n1314,n604,n134);
and (n1315,n603,n47);
nand (n1316,n1317,n1321);
or (n1317,n1318,n775);
nor (n1318,n1319,n1320);
and (n1319,n781,n68);
and (n1320,n435,n67);
or (n1321,n1322,n776);
nor (n1322,n1323,n1324);
and (n1323,n781,n85);
and (n1324,n435,n84);
nand (n1325,n1326,n1330);
or (n1326,n360,n1327);
nor (n1327,n1328,n1329);
and (n1328,n194,n352);
and (n1329,n195,n351);
or (n1330,n1256,n745);
and (n1331,n1307,n1316);
xor (n1332,n1333,n1340);
xor (n1333,n1334,n1337);
nand (n1334,n1335,n1336);
or (n1335,n186,n1300);
or (n1336,n1164,n191);
nand (n1337,n1338,n1339);
or (n1338,n129,n1313);
or (n1339,n148,n1173);
nand (n1340,n1341,n1342);
or (n1341,n1322,n775);
or (n1342,n1179,n776);
or (n1343,n1344,n1383);
and (n1344,n1345,n1382);
xor (n1345,n1346,n1359);
and (n1346,n1347,n1353);
and (n1347,n1348,n47);
nand (n1348,n1349,n1350);
or (n1349,n698,n133);
nand (n1350,n1351,n139);
not (n1351,n1352);
and (n1352,n698,n133);
nand (n1353,n1354,n1358);
or (n1354,n438,n1355);
nor (n1355,n1356,n1357);
and (n1356,n319,n262);
and (n1357,n320,n261);
or (n1358,n439,n1289);
or (n1359,n1360,n1381);
and (n1360,n1361,n1375);
xor (n1361,n1362,n1369);
nand (n1362,n1363,n1368);
or (n1363,n1364,n186);
not (n1364,n1365);
nor (n1365,n1366,n1367);
and (n1366,n604,n140);
and (n1367,n603,n139);
nand (n1368,n192,n1296);
nand (n1369,n1370,n1374);
or (n1370,n129,n1371);
nor (n1371,n1372,n1373);
and (n1372,n47,n697);
and (n1373,n134,n698);
or (n1374,n148,n1309);
nand (n1375,n1376,n1380);
or (n1376,n775,n1377);
nor (n1377,n1378,n1379);
and (n1378,n781,n107);
and (n1379,n435,n106);
or (n1380,n1318,n776);
and (n1381,n1362,n1369);
xor (n1382,n1285,n1293);
and (n1383,n1346,n1359);
not (n1384,n1385);
or (n1385,n1386,n1419);
and (n1386,n1387,n1418);
xor (n1387,n1388,n1389);
xor (n1388,n1306,n1325);
or (n1389,n1390,n1417);
and (n1390,n1391,n1399);
xor (n1391,n1392,n1398);
nand (n1392,n1393,n1397);
or (n1393,n360,n1394);
nor (n1394,n1395,n1396);
and (n1395,n194,n412);
and (n1396,n195,n411);
or (n1397,n1327,n745);
xor (n1398,n1347,n1353);
or (n1399,n1400,n1416);
and (n1400,n1401,n1409);
xor (n1401,n1402,n1403);
and (n1402,n137,n698);
nand (n1403,n1404,n1408);
or (n1404,n1405,n775);
nor (n1405,n1406,n1407);
and (n1406,n781,n96);
and (n1407,n435,n95);
or (n1408,n1377,n776);
nand (n1409,n1410,n1415);
or (n1410,n186,n1411);
not (n1411,n1412);
nand (n1412,n1413,n1414);
or (n1413,n140,n636);
or (n1414,n139,n637);
or (n1415,n191,n1364);
and (n1416,n1402,n1403);
and (n1417,n1392,n1398);
xor (n1418,n1345,n1382);
and (n1419,n1388,n1389);
nor (n1420,n1421,n1461);
not (n1421,n1422);
or (n1422,n1423,n1424);
xor (n1423,n1387,n1418);
or (n1424,n1425,n1460);
and (n1425,n1426,n1459);
xor (n1426,n1427,n1428);
xor (n1427,n1361,n1375);
or (n1428,n1429,n1458);
and (n1429,n1430,n1443);
xor (n1430,n1431,n1437);
nand (n1431,n1432,n1436);
or (n1432,n438,n1433);
nor (n1433,n1434,n1435);
and (n1434,n319,n352);
and (n1435,n320,n351);
or (n1436,n439,n1355);
nand (n1437,n1438,n1442);
or (n1438,n360,n1439);
nor (n1439,n1440,n1441);
and (n1440,n194,n464);
and (n1441,n195,n463);
or (n1442,n1394,n745);
and (n1443,n1444,n1451);
nor (n1444,n1445,n139);
nor (n1445,n1446,n1449);
and (n1446,n1447,n194);
not (n1447,n1448);
and (n1448,n698,n189);
and (n1449,n697,n1450);
not (n1450,n189);
nand (n1451,n1452,n1457);
or (n1452,n775,n1453);
not (n1453,n1454);
nor (n1454,n1455,n1456);
and (n1455,n262,n435);
and (n1456,n261,n781);
or (n1457,n1405,n776);
and (n1458,n1431,n1437);
xor (n1459,n1391,n1399);
and (n1460,n1427,n1428);
nand (n1461,n1462,n1518);
not (n1462,n1463);
nor (n1463,n1464,n1493);
xor (n1464,n1465,n1492);
xor (n1465,n1466,n1491);
or (n1466,n1467,n1490);
and (n1467,n1468,n1484);
xor (n1468,n1469,n1476);
nand (n1469,n1470,n1475);
or (n1470,n1471,n186);
not (n1471,n1472);
nand (n1472,n1473,n1474);
or (n1473,n139,n698);
or (n1474,n140,n697);
nand (n1475,n192,n1412);
nand (n1476,n1477,n1482);
or (n1477,n1478,n438);
not (n1478,n1479);
nand (n1479,n1480,n1481);
or (n1480,n320,n411);
or (n1481,n319,n412);
nand (n1482,n1483,n431);
not (n1483,n1433);
nand (n1484,n1485,n1489);
or (n1485,n360,n1486);
nor (n1486,n1487,n1488);
and (n1487,n194,n604);
and (n1488,n195,n603);
or (n1489,n1439,n745);
and (n1490,n1469,n1476);
xor (n1491,n1401,n1409);
xor (n1492,n1430,n1443);
or (n1493,n1494,n1517);
and (n1494,n1495,n1516);
xor (n1495,n1496,n1497);
xor (n1496,n1444,n1451);
or (n1497,n1498,n1515);
and (n1498,n1499,n1508);
xor (n1499,n1500,n1501);
and (n1500,n192,n698);
nand (n1501,n1502,n1503);
or (n1502,n776,n1453);
or (n1503,n1504,n775);
not (n1504,n1505);
nand (n1505,n1506,n1507);
or (n1506,n352,n781);
nand (n1507,n781,n352);
nand (n1508,n1509,n1514);
or (n1509,n1510,n438);
not (n1510,n1511);
nand (n1511,n1512,n1513);
or (n1512,n320,n463);
or (n1513,n319,n464);
nand (n1514,n431,n1479);
and (n1515,n1500,n1501);
xor (n1516,n1468,n1484);
and (n1517,n1496,n1497);
not (n1518,n1519);
nor (n1519,n1520,n1521);
xor (n1520,n1426,n1459);
or (n1521,n1522,n1523);
and (n1522,n1465,n1492);
and (n1523,n1466,n1491);
or (n1524,n1525,n1663);
and (n1525,n1526,n1553);
xor (n1526,n1527,n1552);
or (n1527,n1528,n1551);
and (n1528,n1529,n1550);
xor (n1529,n1530,n1536);
nand (n1530,n1531,n1535);
or (n1531,n360,n1532);
nor (n1532,n1533,n1534);
and (n1533,n194,n637);
and (n1534,n195,n636);
or (n1535,n1486,n745);
nor (n1536,n1537,n1545);
not (n1537,n1538);
nand (n1538,n1539,n1544);
or (n1539,n775,n1540);
not (n1540,n1541);
nor (n1541,n1542,n1543);
and (n1542,n412,n435);
and (n1543,n411,n781);
nand (n1544,n1505,n777);
nand (n1545,n1546,n195);
nand (n1546,n1547,n1549);
or (n1547,n1548,n320);
and (n1548,n698,n321);
or (n1549,n698,n321);
xor (n1550,n1499,n1508);
and (n1551,n1530,n1536);
xor (n1552,n1495,n1516);
or (n1553,n1554,n1662);
and (n1554,n1555,n1579);
xor (n1555,n1556,n1578);
or (n1556,n1557,n1577);
and (n1557,n1558,n1573);
xor (n1558,n1559,n1566);
nand (n1559,n1560,n1565);
or (n1560,n1561,n438);
not (n1561,n1562);
nor (n1562,n1563,n1564);
and (n1563,n603,n319);
and (n1564,n604,n320);
nand (n1565,n431,n1511);
nand (n1566,n1567,n1572);
or (n1567,n1568,n360);
not (n1568,n1569);
nand (n1569,n1570,n1571);
or (n1570,n194,n698);
or (n1571,n697,n195);
or (n1572,n1532,n745);
nand (n1573,n1574,n1576);
or (n1574,n1575,n1537);
not (n1575,n1545);
or (n1576,n1538,n1545);
and (n1577,n1559,n1566);
xor (n1578,n1529,n1550);
or (n1579,n1580,n1661);
and (n1580,n1581,n1602);
xor (n1581,n1582,n1601);
or (n1582,n1583,n1600);
and (n1583,n1584,n1593);
xor (n1584,n1585,n1586);
and (n1585,n317,n698);
nand (n1586,n1587,n1592);
or (n1587,n1588,n438);
not (n1588,n1589);
nor (n1589,n1590,n1591);
and (n1590,n636,n319);
and (n1591,n637,n320);
nand (n1592,n431,n1562);
nand (n1593,n1594,n1595);
or (n1594,n776,n1540);
or (n1595,n775,n1596);
not (n1596,n1597);
nor (n1597,n1598,n1599);
and (n1598,n463,n781);
and (n1599,n464,n435);
and (n1600,n1585,n1586);
xor (n1601,n1558,n1573);
nand (n1602,n1603,n1660);
or (n1603,n1604,n1620);
nor (n1604,n1605,n1606);
xor (n1605,n1584,n1593);
and (n1606,n1607,n1614);
nand (n1607,n1608,n1609);
nand (n1608,n1597,n777);
nand (n1609,n1610,n1613);
nor (n1610,n1611,n1612);
and (n1611,n603,n781);
and (n1612,n604,n435);
not (n1613,n775);
not (n1614,n1615);
nand (n1615,n1616,n320);
nand (n1616,n1617,n1619);
or (n1617,n1618,n435);
and (n1618,n698,n434);
or (n1619,n698,n434);
nor (n1620,n1621,n1659);
and (n1621,n1622,n1633);
nand (n1622,n1623,n1627);
nor (n1623,n1624,n1626);
and (n1624,n1625,n1614);
not (n1625,n1607);
and (n1626,n1607,n1615);
nor (n1627,n1628,n1629);
and (n1628,n431,n1589);
and (n1629,n437,n1630);
nand (n1630,n1631,n1632);
or (n1631,n319,n698);
or (n1632,n697,n320);
nand (n1633,n1634,n1657);
or (n1634,n1635,n1649);
not (n1635,n1636);
and (n1636,n1637,n1647);
nand (n1637,n1638,n1643);
or (n1638,n776,n1639);
not (n1639,n1640);
nor (n1640,n1641,n1642);
and (n1641,n636,n781);
and (n1642,n637,n435);
nand (n1643,n1644,n1613);
nand (n1644,n1645,n1646);
or (n1645,n781,n698);
or (n1646,n435,n697);
nor (n1647,n1648,n781);
and (n1648,n698,n777);
not (n1649,n1650);
nand (n1650,n1651,n1656);
not (n1651,n1652);
nand (n1652,n1653,n1655);
or (n1653,n776,n1654);
not (n1654,n1610);
nand (n1655,n1640,n1613);
nand (n1656,n431,n698);
nand (n1657,n1658,n1652);
not (n1658,n1656);
nor (n1659,n1623,n1627);
nand (n1660,n1605,n1606);
and (n1661,n1582,n1601);
and (n1662,n1556,n1578);
and (n1663,n1527,n1552);
nand (n1664,n1665,n1242);
or (n1665,n1666,n1668);
not (n1666,n1667);
nand (n1667,n1423,n1424);
not (n1668,n1669);
nand (n1669,n1422,n1670);
nand (n1670,n1671,n1673);
or (n1671,n1519,n1672);
nand (n1672,n1464,n1493);
nand (n1673,n1520,n1521);
nand (n1674,n1244,n1385);
not (n1675,n1676);
nor (n1676,n1677,n1702);
nor (n1677,n1678,n1679);
xor (n1678,n1139,n1192);
or (n1679,n1680,n1701);
and (n1680,n1681,n1684);
xor (n1681,n1682,n1683);
xor (n1682,n1082,n1130);
xor (n1683,n1143,n1146);
or (n1684,n1685,n1700);
and (n1685,n1686,n1689);
xor (n1686,n1687,n1688);
xor (n1687,n1110,n1123);
xor (n1688,n1085,n1100);
or (n1689,n1690,n1699);
and (n1690,n1691,n1696);
xor (n1691,n1692,n1695);
nand (n1692,n1693,n1694);
or (n1693,n360,n1260);
or (n1694,n1113,n745);
and (n1695,n1273,n1265);
or (n1696,n1697,n1698);
and (n1697,n1333,n1340);
and (n1698,n1334,n1337);
and (n1699,n1692,n1695);
and (n1700,n1687,n1688);
and (n1701,n1682,n1683);
nand (n1702,n1703,n1732);
nor (n1703,n1704,n1727);
nor (n1704,n1705,n1718);
xor (n1705,n1706,n1717);
xor (n1706,n1707,n1708);
xor (n1707,n1148,n1168);
or (n1708,n1709,n1716);
and (n1709,n1710,n1713);
xor (n1710,n1711,n1712);
xor (n1711,n1170,n1183);
xor (n1712,n1152,n1161);
or (n1713,n1714,n1715);
and (n1714,n1247,n1263);
and (n1715,n1248,n1254);
and (n1716,n1711,n1712);
xor (n1717,n1686,n1689);
or (n1718,n1719,n1726);
and (n1719,n1720,n1725);
xor (n1720,n1721,n1722);
xor (n1721,n1691,n1696);
or (n1722,n1723,n1724);
and (n1723,n1282,n1332);
and (n1724,n1283,n1304);
xor (n1725,n1710,n1713);
and (n1726,n1721,n1722);
nor (n1727,n1728,n1731);
or (n1728,n1729,n1730);
and (n1729,n1245,n1343);
and (n1730,n1246,n1281);
xor (n1731,n1720,n1725);
nand (n1732,n1733,n1735);
not (n1733,n1734);
xor (n1734,n1681,n1684);
not (n1735,n1736);
or (n1736,n1737,n1738);
and (n1737,n1706,n1717);
and (n1738,n1707,n1708);
nor (n1739,n1740,n1751);
and (n1740,n1741,n1742);
not (n1741,n1677);
nand (n1742,n1743,n1750);
or (n1743,n1744,n1745);
not (n1744,n1732);
not (n1745,n1746);
nand (n1746,n1747,n1749);
or (n1747,n1704,n1748);
nand (n1748,n1728,n1731);
nand (n1749,n1705,n1718);
nand (n1750,n1734,n1736);
and (n1751,n1678,n1679);
not (n1752,n1753);
nand (n1753,n1754,n1756);
or (n1754,n1755,n523);
nand (n1755,n281,n514);
nand (n1756,n524,n525);
nand (n1757,n276,n2);
xor (n1758,n1759,n3083);
xor (n1759,n1760,n3082);
xor (n1760,n1761,n3025);
xor (n1761,n1762,n3024);
xor (n1762,n1763,n2955);
xor (n1763,n1764,n2954);
xor (n1764,n1765,n2879);
xor (n1765,n1766,n2878);
xor (n1766,n1767,n2797);
xor (n1767,n1768,n2796);
xor (n1768,n1769,n2712);
xor (n1769,n1770,n2711);
xor (n1770,n1771,n2619);
xor (n1771,n1772,n2618);
or (n1772,n1773,n2528);
and (n1773,n1774,n2527);
or (n1774,n1775,n2433);
and (n1775,n1776,n2432);
or (n1776,n1777,n2345);
and (n1777,n1778,n2344);
or (n1778,n1779,n2250);
and (n1779,n1780,n2249);
or (n1780,n1781,n2156);
and (n1781,n1782,n358);
or (n1782,n1783,n2062);
and (n1783,n1784,n2061);
or (n1784,n1785,n1971);
and (n1785,n1786,n508);
or (n1786,n1787,n1877);
and (n1787,n1788,n1876);
and (n1788,n782,n1789);
or (n1789,n1790,n1793);
and (n1790,n1791,n1792);
and (n1791,n144,n777);
and (n1792,n40,n435);
and (n1793,n1794,n1795);
xor (n1794,n1791,n1792);
or (n1795,n1796,n1799);
and (n1796,n1797,n1798);
and (n1797,n40,n777);
and (n1798,n57,n435);
and (n1799,n1800,n1801);
xor (n1800,n1797,n1798);
or (n1801,n1802,n1804);
and (n1802,n1803,n937);
and (n1803,n57,n777);
and (n1804,n1805,n1806);
xor (n1805,n1803,n937);
or (n1806,n1807,n1810);
and (n1807,n1808,n1809);
and (n1808,n30,n777);
and (n1809,n24,n435);
and (n1810,n1811,n1812);
xor (n1811,n1808,n1809);
or (n1812,n1813,n1816);
and (n1813,n1814,n1815);
and (n1814,n24,n777);
and (n1815,n121,n435);
and (n1816,n1817,n1818);
xor (n1817,n1814,n1815);
or (n1818,n1819,n1822);
and (n1819,n1820,n1821);
and (n1820,n121,n777);
and (n1821,n85,n435);
and (n1822,n1823,n1824);
xor (n1823,n1820,n1821);
or (n1824,n1825,n1828);
and (n1825,n1826,n1827);
and (n1826,n85,n777);
and (n1827,n68,n435);
and (n1828,n1829,n1830);
xor (n1829,n1826,n1827);
or (n1830,n1831,n1834);
and (n1831,n1832,n1833);
and (n1832,n68,n777);
and (n1833,n107,n435);
and (n1834,n1835,n1836);
xor (n1835,n1832,n1833);
or (n1836,n1837,n1840);
and (n1837,n1838,n1839);
and (n1838,n107,n777);
and (n1839,n96,n435);
and (n1840,n1841,n1842);
xor (n1841,n1838,n1839);
or (n1842,n1843,n1845);
and (n1843,n1844,n1455);
and (n1844,n96,n777);
and (n1845,n1846,n1847);
xor (n1846,n1844,n1455);
or (n1847,n1848,n1851);
and (n1848,n1849,n1850);
and (n1849,n262,n777);
and (n1850,n352,n435);
and (n1851,n1852,n1853);
xor (n1852,n1849,n1850);
or (n1853,n1854,n1856);
and (n1854,n1855,n1542);
and (n1855,n352,n777);
and (n1856,n1857,n1858);
xor (n1857,n1855,n1542);
or (n1858,n1859,n1861);
and (n1859,n1860,n1599);
and (n1860,n412,n777);
and (n1861,n1862,n1863);
xor (n1862,n1860,n1599);
or (n1863,n1864,n1866);
and (n1864,n1865,n1612);
and (n1865,n464,n777);
and (n1866,n1867,n1868);
xor (n1867,n1865,n1612);
or (n1868,n1869,n1871);
and (n1869,n1870,n1642);
and (n1870,n604,n777);
and (n1871,n1872,n1873);
xor (n1872,n1870,n1642);
and (n1873,n1874,n1875);
and (n1874,n637,n777);
and (n1875,n698,n435);
and (n1876,n144,n434);
and (n1877,n1878,n1879);
xor (n1878,n1788,n1876);
or (n1879,n1880,n1883);
and (n1880,n1881,n1882);
xor (n1881,n782,n1789);
and (n1882,n40,n434);
and (n1883,n1884,n1885);
xor (n1884,n1881,n1882);
or (n1885,n1886,n1889);
and (n1886,n1887,n1888);
xor (n1887,n1794,n1795);
and (n1888,n57,n434);
and (n1889,n1890,n1891);
xor (n1890,n1887,n1888);
or (n1891,n1892,n1895);
and (n1892,n1893,n1894);
xor (n1893,n1800,n1801);
and (n1894,n30,n434);
and (n1895,n1896,n1897);
xor (n1896,n1893,n1894);
or (n1897,n1898,n1901);
and (n1898,n1899,n1900);
xor (n1899,n1805,n1806);
and (n1900,n24,n434);
and (n1901,n1902,n1903);
xor (n1902,n1899,n1900);
or (n1903,n1904,n1907);
and (n1904,n1905,n1906);
xor (n1905,n1811,n1812);
and (n1906,n121,n434);
and (n1907,n1908,n1909);
xor (n1908,n1905,n1906);
or (n1909,n1910,n1913);
and (n1910,n1911,n1912);
xor (n1911,n1817,n1818);
and (n1912,n85,n434);
and (n1913,n1914,n1915);
xor (n1914,n1911,n1912);
or (n1915,n1916,n1919);
and (n1916,n1917,n1918);
xor (n1917,n1823,n1824);
and (n1918,n68,n434);
and (n1919,n1920,n1921);
xor (n1920,n1917,n1918);
or (n1921,n1922,n1925);
and (n1922,n1923,n1924);
xor (n1923,n1829,n1830);
and (n1924,n107,n434);
and (n1925,n1926,n1927);
xor (n1926,n1923,n1924);
or (n1927,n1928,n1931);
and (n1928,n1929,n1930);
xor (n1929,n1835,n1836);
and (n1930,n96,n434);
and (n1931,n1932,n1933);
xor (n1932,n1929,n1930);
or (n1933,n1934,n1937);
and (n1934,n1935,n1936);
xor (n1935,n1841,n1842);
and (n1936,n262,n434);
and (n1937,n1938,n1939);
xor (n1938,n1935,n1936);
or (n1939,n1940,n1943);
and (n1940,n1941,n1942);
xor (n1941,n1846,n1847);
and (n1942,n352,n434);
and (n1943,n1944,n1945);
xor (n1944,n1941,n1942);
or (n1945,n1946,n1949);
and (n1946,n1947,n1948);
xor (n1947,n1852,n1853);
and (n1948,n412,n434);
and (n1949,n1950,n1951);
xor (n1950,n1947,n1948);
or (n1951,n1952,n1955);
and (n1952,n1953,n1954);
xor (n1953,n1857,n1858);
and (n1954,n464,n434);
and (n1955,n1956,n1957);
xor (n1956,n1953,n1954);
or (n1957,n1958,n1961);
and (n1958,n1959,n1960);
xor (n1959,n1862,n1863);
and (n1960,n604,n434);
and (n1961,n1962,n1963);
xor (n1962,n1959,n1960);
or (n1963,n1964,n1967);
and (n1964,n1965,n1966);
xor (n1965,n1867,n1868);
and (n1966,n637,n434);
and (n1967,n1968,n1969);
xor (n1968,n1965,n1966);
and (n1969,n1970,n1618);
xor (n1970,n1872,n1873);
and (n1971,n1972,n1973);
xor (n1972,n1786,n508);
or (n1973,n1974,n1977);
and (n1974,n1975,n1976);
xor (n1975,n1878,n1879);
and (n1976,n40,n320);
and (n1977,n1978,n1979);
xor (n1978,n1975,n1976);
or (n1979,n1980,n1982);
and (n1980,n1981,n729);
xor (n1981,n1884,n1885);
and (n1982,n1983,n1984);
xor (n1983,n1981,n729);
or (n1984,n1985,n1987);
and (n1985,n1986,n816);
xor (n1986,n1890,n1891);
and (n1987,n1988,n1989);
xor (n1988,n1986,n816);
or (n1989,n1990,n1993);
and (n1990,n1991,n1992);
xor (n1991,n1896,n1897);
and (n1992,n24,n320);
and (n1993,n1994,n1995);
xor (n1994,n1991,n1992);
or (n1995,n1996,n1999);
and (n1996,n1997,n1998);
xor (n1997,n1902,n1903);
and (n1998,n121,n320);
and (n1999,n2000,n2001);
xor (n2000,n1997,n1998);
or (n2001,n2002,n2004);
and (n2002,n2003,n1091);
xor (n2003,n1908,n1909);
and (n2004,n2005,n2006);
xor (n2005,n2003,n1091);
or (n2006,n2007,n2010);
and (n2007,n2008,n2009);
xor (n2008,n1914,n1915);
and (n2009,n68,n320);
and (n2010,n2011,n2012);
xor (n2011,n2008,n2009);
or (n2012,n2013,n2016);
and (n2013,n2014,n2015);
xor (n2014,n1920,n1921);
and (n2015,n107,n320);
and (n2016,n2017,n2018);
xor (n2017,n2014,n2015);
or (n2018,n2019,n2022);
and (n2019,n2020,n2021);
xor (n2020,n1926,n1927);
and (n2021,n96,n320);
and (n2022,n2023,n2024);
xor (n2023,n2020,n2021);
or (n2024,n2025,n2028);
and (n2025,n2026,n2027);
xor (n2026,n1932,n1933);
and (n2027,n262,n320);
and (n2028,n2029,n2030);
xor (n2029,n2026,n2027);
or (n2030,n2031,n2034);
and (n2031,n2032,n2033);
xor (n2032,n1938,n1939);
and (n2033,n352,n320);
and (n2034,n2035,n2036);
xor (n2035,n2032,n2033);
or (n2036,n2037,n2040);
and (n2037,n2038,n2039);
xor (n2038,n1944,n1945);
and (n2039,n412,n320);
and (n2040,n2041,n2042);
xor (n2041,n2038,n2039);
or (n2042,n2043,n2046);
and (n2043,n2044,n2045);
xor (n2044,n1950,n1951);
and (n2045,n464,n320);
and (n2046,n2047,n2048);
xor (n2047,n2044,n2045);
or (n2048,n2049,n2051);
and (n2049,n2050,n1564);
xor (n2050,n1956,n1957);
and (n2051,n2052,n2053);
xor (n2052,n2050,n1564);
or (n2053,n2054,n2056);
and (n2054,n2055,n1591);
xor (n2055,n1962,n1963);
and (n2056,n2057,n2058);
xor (n2057,n2055,n1591);
and (n2058,n2059,n2060);
xor (n2059,n1968,n1969);
and (n2060,n698,n320);
and (n2061,n144,n321);
and (n2062,n2063,n2064);
xor (n2063,n1784,n2061);
or (n2064,n2065,n2068);
and (n2065,n2066,n2067);
xor (n2066,n1972,n1973);
and (n2067,n40,n321);
and (n2068,n2069,n2070);
xor (n2069,n2066,n2067);
or (n2070,n2071,n2074);
and (n2071,n2072,n2073);
xor (n2072,n1978,n1979);
and (n2073,n57,n321);
and (n2074,n2075,n2076);
xor (n2075,n2072,n2073);
or (n2076,n2077,n2080);
and (n2077,n2078,n2079);
xor (n2078,n1983,n1984);
and (n2079,n30,n321);
and (n2080,n2081,n2082);
xor (n2081,n2078,n2079);
or (n2082,n2083,n2086);
and (n2083,n2084,n2085);
xor (n2084,n1988,n1989);
and (n2085,n24,n321);
and (n2086,n2087,n2088);
xor (n2087,n2084,n2085);
or (n2088,n2089,n2092);
and (n2089,n2090,n2091);
xor (n2090,n1994,n1995);
and (n2091,n121,n321);
and (n2092,n2093,n2094);
xor (n2093,n2090,n2091);
or (n2094,n2095,n2098);
and (n2095,n2096,n2097);
xor (n2096,n2000,n2001);
and (n2097,n85,n321);
and (n2098,n2099,n2100);
xor (n2099,n2096,n2097);
or (n2100,n2101,n2104);
and (n2101,n2102,n2103);
xor (n2102,n2005,n2006);
and (n2103,n68,n321);
and (n2104,n2105,n2106);
xor (n2105,n2102,n2103);
or (n2106,n2107,n2110);
and (n2107,n2108,n2109);
xor (n2108,n2011,n2012);
and (n2109,n107,n321);
and (n2110,n2111,n2112);
xor (n2111,n2108,n2109);
or (n2112,n2113,n2116);
and (n2113,n2114,n2115);
xor (n2114,n2017,n2018);
and (n2115,n96,n321);
and (n2116,n2117,n2118);
xor (n2117,n2114,n2115);
or (n2118,n2119,n2122);
and (n2119,n2120,n2121);
xor (n2120,n2023,n2024);
and (n2121,n262,n321);
and (n2122,n2123,n2124);
xor (n2123,n2120,n2121);
or (n2124,n2125,n2128);
and (n2125,n2126,n2127);
xor (n2126,n2029,n2030);
and (n2127,n352,n321);
and (n2128,n2129,n2130);
xor (n2129,n2126,n2127);
or (n2130,n2131,n2134);
and (n2131,n2132,n2133);
xor (n2132,n2035,n2036);
and (n2133,n412,n321);
and (n2134,n2135,n2136);
xor (n2135,n2132,n2133);
or (n2136,n2137,n2140);
and (n2137,n2138,n2139);
xor (n2138,n2041,n2042);
and (n2139,n464,n321);
and (n2140,n2141,n2142);
xor (n2141,n2138,n2139);
or (n2142,n2143,n2146);
and (n2143,n2144,n2145);
xor (n2144,n2047,n2048);
and (n2145,n604,n321);
and (n2146,n2147,n2148);
xor (n2147,n2144,n2145);
or (n2148,n2149,n2152);
and (n2149,n2150,n2151);
xor (n2150,n2052,n2053);
and (n2151,n637,n321);
and (n2152,n2153,n2154);
xor (n2153,n2150,n2151);
and (n2154,n2155,n1548);
xor (n2155,n2057,n2058);
and (n2156,n2157,n2158);
xor (n2157,n1782,n358);
or (n2158,n2159,n2162);
and (n2159,n2160,n2161);
xor (n2160,n2063,n2064);
and (n2161,n40,n195);
and (n2162,n2163,n2164);
xor (n2163,n2160,n2161);
or (n2164,n2165,n2167);
and (n2165,n2166,n599);
xor (n2166,n2069,n2070);
and (n2167,n2168,n2169);
xor (n2168,n2166,n599);
or (n2169,n2170,n2173);
and (n2170,n2171,n2172);
xor (n2171,n2075,n2076);
and (n2172,n30,n195);
and (n2173,n2174,n2175);
xor (n2174,n2171,n2172);
or (n2175,n2176,n2178);
and (n2176,n2177,n743);
xor (n2177,n2081,n2082);
and (n2178,n2179,n2180);
xor (n2179,n2177,n743);
or (n2180,n2181,n2184);
and (n2181,n2182,n2183);
xor (n2182,n2087,n2088);
and (n2183,n121,n195);
and (n2184,n2185,n2186);
xor (n2185,n2182,n2183);
or (n2186,n2187,n2190);
and (n2187,n2188,n2189);
xor (n2188,n2093,n2094);
and (n2189,n85,n195);
and (n2190,n2191,n2192);
xor (n2191,n2188,n2189);
or (n2192,n2193,n2196);
and (n2193,n2194,n2195);
xor (n2194,n2099,n2100);
and (n2195,n68,n195);
and (n2196,n2197,n2198);
xor (n2197,n2194,n2195);
or (n2198,n2199,n2202);
and (n2199,n2200,n2201);
xor (n2200,n2105,n2106);
and (n2201,n107,n195);
and (n2202,n2203,n2204);
xor (n2203,n2200,n2201);
or (n2204,n2205,n2208);
and (n2205,n2206,n2207);
xor (n2206,n2111,n2112);
and (n2207,n96,n195);
and (n2208,n2209,n2210);
xor (n2209,n2206,n2207);
or (n2210,n2211,n2214);
and (n2211,n2212,n2213);
xor (n2212,n2117,n2118);
and (n2213,n262,n195);
and (n2214,n2215,n2216);
xor (n2215,n2212,n2213);
or (n2216,n2217,n2220);
and (n2217,n2218,n2219);
xor (n2218,n2123,n2124);
and (n2219,n352,n195);
and (n2220,n2221,n2222);
xor (n2221,n2218,n2219);
or (n2222,n2223,n2226);
and (n2223,n2224,n2225);
xor (n2224,n2129,n2130);
and (n2225,n412,n195);
and (n2226,n2227,n2228);
xor (n2227,n2224,n2225);
or (n2228,n2229,n2232);
and (n2229,n2230,n2231);
xor (n2230,n2135,n2136);
and (n2231,n464,n195);
and (n2232,n2233,n2234);
xor (n2233,n2230,n2231);
or (n2234,n2235,n2238);
and (n2235,n2236,n2237);
xor (n2236,n2141,n2142);
and (n2237,n604,n195);
and (n2238,n2239,n2240);
xor (n2239,n2236,n2237);
or (n2240,n2241,n2244);
and (n2241,n2242,n2243);
xor (n2242,n2147,n2148);
and (n2243,n637,n195);
and (n2244,n2245,n2246);
xor (n2245,n2242,n2243);
and (n2246,n2247,n2248);
xor (n2247,n2153,n2154);
and (n2248,n698,n195);
and (n2249,n144,n189);
and (n2250,n2251,n2252);
xor (n2251,n1780,n2249);
or (n2252,n2253,n2256);
and (n2253,n2254,n2255);
xor (n2254,n2157,n2158);
and (n2255,n40,n189);
and (n2256,n2257,n2258);
xor (n2257,n2254,n2255);
or (n2258,n2259,n2262);
and (n2259,n2260,n2261);
xor (n2260,n2163,n2164);
and (n2261,n57,n189);
and (n2262,n2263,n2264);
xor (n2263,n2260,n2261);
or (n2264,n2265,n2268);
and (n2265,n2266,n2267);
xor (n2266,n2168,n2169);
and (n2267,n30,n189);
and (n2268,n2269,n2270);
xor (n2269,n2266,n2267);
or (n2270,n2271,n2274);
and (n2271,n2272,n2273);
xor (n2272,n2174,n2175);
and (n2273,n24,n189);
and (n2274,n2275,n2276);
xor (n2275,n2272,n2273);
or (n2276,n2277,n2280);
and (n2277,n2278,n2279);
xor (n2278,n2179,n2180);
and (n2279,n121,n189);
and (n2280,n2281,n2282);
xor (n2281,n2278,n2279);
or (n2282,n2283,n2286);
and (n2283,n2284,n2285);
xor (n2284,n2185,n2186);
and (n2285,n85,n189);
and (n2286,n2287,n2288);
xor (n2287,n2284,n2285);
or (n2288,n2289,n2292);
and (n2289,n2290,n2291);
xor (n2290,n2191,n2192);
and (n2291,n68,n189);
and (n2292,n2293,n2294);
xor (n2293,n2290,n2291);
or (n2294,n2295,n2298);
and (n2295,n2296,n2297);
xor (n2296,n2197,n2198);
and (n2297,n107,n189);
and (n2298,n2299,n2300);
xor (n2299,n2296,n2297);
or (n2300,n2301,n2304);
and (n2301,n2302,n2303);
xor (n2302,n2203,n2204);
and (n2303,n96,n189);
and (n2304,n2305,n2306);
xor (n2305,n2302,n2303);
or (n2306,n2307,n2310);
and (n2307,n2308,n2309);
xor (n2308,n2209,n2210);
and (n2309,n262,n189);
and (n2310,n2311,n2312);
xor (n2311,n2308,n2309);
or (n2312,n2313,n2316);
and (n2313,n2314,n2315);
xor (n2314,n2215,n2216);
and (n2315,n352,n189);
and (n2316,n2317,n2318);
xor (n2317,n2314,n2315);
or (n2318,n2319,n2322);
and (n2319,n2320,n2321);
xor (n2320,n2221,n2222);
and (n2321,n412,n189);
and (n2322,n2323,n2324);
xor (n2323,n2320,n2321);
or (n2324,n2325,n2328);
and (n2325,n2326,n2327);
xor (n2326,n2227,n2228);
and (n2327,n464,n189);
and (n2328,n2329,n2330);
xor (n2329,n2326,n2327);
or (n2330,n2331,n2334);
and (n2331,n2332,n2333);
xor (n2332,n2233,n2234);
and (n2333,n604,n189);
and (n2334,n2335,n2336);
xor (n2335,n2332,n2333);
or (n2336,n2337,n2340);
and (n2337,n2338,n2339);
xor (n2338,n2239,n2240);
and (n2339,n637,n189);
and (n2340,n2341,n2342);
xor (n2341,n2338,n2339);
and (n2342,n2343,n1448);
xor (n2343,n2245,n2246);
and (n2344,n144,n140);
and (n2345,n2346,n2347);
xor (n2346,n1778,n2344);
or (n2347,n2348,n2350);
and (n2348,n2349,n333);
xor (n2349,n2251,n2252);
and (n2350,n2351,n2352);
xor (n2351,n2349,n333);
or (n2352,n2353,n2355);
and (n2353,n2354,n369);
xor (n2354,n2257,n2258);
and (n2355,n2356,n2357);
xor (n2356,n2354,n369);
or (n2357,n2358,n2360);
and (n2358,n2359,n478);
xor (n2359,n2263,n2264);
and (n2360,n2361,n2362);
xor (n2361,n2359,n478);
or (n2362,n2363,n2365);
and (n2363,n2364,n561);
xor (n2364,n2269,n2270);
and (n2365,n2366,n2367);
xor (n2366,n2364,n561);
or (n2367,n2368,n2370);
and (n2368,n2369,n557);
xor (n2369,n2275,n2276);
and (n2370,n2371,n2372);
xor (n2371,n2369,n557);
or (n2372,n2373,n2376);
and (n2373,n2374,n2375);
xor (n2374,n2281,n2282);
and (n2375,n85,n140);
and (n2376,n2377,n2378);
xor (n2377,n2374,n2375);
or (n2378,n2379,n2382);
and (n2379,n2380,n2381);
xor (n2380,n2287,n2288);
and (n2381,n68,n140);
and (n2382,n2383,n2384);
xor (n2383,n2380,n2381);
or (n2384,n2385,n2387);
and (n2385,n2386,n974);
xor (n2386,n2293,n2294);
and (n2387,n2388,n2389);
xor (n2388,n2386,n974);
or (n2389,n2390,n2393);
and (n2390,n2391,n2392);
xor (n2391,n2299,n2300);
and (n2392,n96,n140);
and (n2393,n2394,n2395);
xor (n2394,n2391,n2392);
or (n2395,n2396,n2399);
and (n2396,n2397,n2398);
xor (n2397,n2305,n2306);
and (n2398,n262,n140);
and (n2399,n2400,n2401);
xor (n2400,n2397,n2398);
or (n2401,n2402,n2405);
and (n2402,n2403,n2404);
xor (n2403,n2311,n2312);
and (n2404,n352,n140);
and (n2405,n2406,n2407);
xor (n2406,n2403,n2404);
or (n2407,n2408,n2411);
and (n2408,n2409,n2410);
xor (n2409,n2317,n2318);
and (n2410,n412,n140);
and (n2411,n2412,n2413);
xor (n2412,n2409,n2410);
or (n2413,n2414,n2416);
and (n2414,n2415,n1298);
xor (n2415,n2323,n2324);
and (n2416,n2417,n2418);
xor (n2417,n2415,n1298);
or (n2418,n2419,n2421);
and (n2419,n2420,n1366);
xor (n2420,n2329,n2330);
and (n2421,n2422,n2423);
xor (n2422,n2420,n1366);
or (n2423,n2424,n2427);
and (n2424,n2425,n2426);
xor (n2425,n2335,n2336);
and (n2426,n637,n140);
and (n2427,n2428,n2429);
xor (n2428,n2425,n2426);
and (n2429,n2430,n2431);
xor (n2430,n2341,n2342);
and (n2431,n698,n140);
and (n2432,n144,n133);
and (n2433,n2434,n2435);
xor (n2434,n1776,n2432);
or (n2435,n2436,n2439);
and (n2436,n2437,n2438);
xor (n2437,n2346,n2347);
and (n2438,n40,n133);
and (n2439,n2440,n2441);
xor (n2440,n2437,n2438);
or (n2441,n2442,n2445);
and (n2442,n2443,n2444);
xor (n2443,n2351,n2352);
and (n2444,n57,n133);
and (n2445,n2446,n2447);
xor (n2446,n2443,n2444);
or (n2447,n2448,n2451);
and (n2448,n2449,n2450);
xor (n2449,n2356,n2357);
and (n2450,n30,n133);
and (n2451,n2452,n2453);
xor (n2452,n2449,n2450);
or (n2453,n2454,n2457);
and (n2454,n2455,n2456);
xor (n2455,n2361,n2362);
and (n2456,n24,n133);
and (n2457,n2458,n2459);
xor (n2458,n2455,n2456);
or (n2459,n2460,n2463);
and (n2460,n2461,n2462);
xor (n2461,n2366,n2367);
and (n2462,n121,n133);
and (n2463,n2464,n2465);
xor (n2464,n2461,n2462);
or (n2465,n2466,n2469);
and (n2466,n2467,n2468);
xor (n2467,n2371,n2372);
and (n2468,n85,n133);
and (n2469,n2470,n2471);
xor (n2470,n2467,n2468);
or (n2471,n2472,n2475);
and (n2472,n2473,n2474);
xor (n2473,n2377,n2378);
and (n2474,n68,n133);
and (n2475,n2476,n2477);
xor (n2476,n2473,n2474);
or (n2477,n2478,n2481);
and (n2478,n2479,n2480);
xor (n2479,n2383,n2384);
and (n2480,n107,n133);
and (n2481,n2482,n2483);
xor (n2482,n2479,n2480);
or (n2483,n2484,n2487);
and (n2484,n2485,n2486);
xor (n2485,n2388,n2389);
and (n2486,n96,n133);
and (n2487,n2488,n2489);
xor (n2488,n2485,n2486);
or (n2489,n2490,n2493);
and (n2490,n2491,n2492);
xor (n2491,n2394,n2395);
and (n2492,n262,n133);
and (n2493,n2494,n2495);
xor (n2494,n2491,n2492);
or (n2495,n2496,n2499);
and (n2496,n2497,n2498);
xor (n2497,n2400,n2401);
and (n2498,n352,n133);
and (n2499,n2500,n2501);
xor (n2500,n2497,n2498);
or (n2501,n2502,n2505);
and (n2502,n2503,n2504);
xor (n2503,n2406,n2407);
and (n2504,n412,n133);
and (n2505,n2506,n2507);
xor (n2506,n2503,n2504);
or (n2507,n2508,n2511);
and (n2508,n2509,n2510);
xor (n2509,n2412,n2413);
and (n2510,n464,n133);
and (n2511,n2512,n2513);
xor (n2512,n2509,n2510);
or (n2513,n2514,n2517);
and (n2514,n2515,n2516);
xor (n2515,n2417,n2418);
and (n2516,n604,n133);
and (n2517,n2518,n2519);
xor (n2518,n2515,n2516);
or (n2519,n2520,n2523);
and (n2520,n2521,n2522);
xor (n2521,n2422,n2423);
and (n2522,n637,n133);
and (n2523,n2524,n2525);
xor (n2524,n2521,n2522);
and (n2525,n2526,n1352);
xor (n2526,n2428,n2429);
and (n2527,n144,n47);
and (n2528,n2529,n2530);
xor (n2529,n1774,n2527);
or (n2530,n2531,n2534);
and (n2531,n2532,n2533);
xor (n2532,n2434,n2435);
and (n2533,n40,n47);
and (n2534,n2535,n2536);
xor (n2535,n2532,n2533);
or (n2536,n2537,n2540);
and (n2537,n2538,n2539);
xor (n2538,n2440,n2441);
and (n2539,n57,n47);
and (n2540,n2541,n2542);
xor (n2541,n2538,n2539);
or (n2542,n2543,n2545);
and (n2543,n2544,n303);
xor (n2544,n2446,n2447);
and (n2545,n2546,n2547);
xor (n2546,n2544,n303);
or (n2547,n2548,n2550);
and (n2548,n2549,n400);
xor (n2549,n2452,n2453);
and (n2550,n2551,n2552);
xor (n2551,n2549,n400);
or (n2552,n2553,n2556);
and (n2553,n2554,n2555);
xor (n2554,n2458,n2459);
and (n2555,n121,n47);
and (n2556,n2557,n2558);
xor (n2557,n2554,n2555);
or (n2558,n2559,n2561);
and (n2559,n2560,n611);
xor (n2560,n2464,n2465);
and (n2561,n2562,n2563);
xor (n2562,n2560,n611);
or (n2563,n2564,n2566);
and (n2564,n2565,n656);
xor (n2565,n2470,n2471);
and (n2566,n2567,n2568);
xor (n2567,n2565,n656);
or (n2568,n2569,n2572);
and (n2569,n2570,n2571);
xor (n2570,n2476,n2477);
and (n2571,n107,n47);
and (n2572,n2573,n2574);
xor (n2573,n2570,n2571);
or (n2574,n2575,n2578);
and (n2575,n2576,n2577);
xor (n2576,n2482,n2483);
and (n2577,n96,n47);
and (n2578,n2579,n2580);
xor (n2579,n2576,n2577);
or (n2580,n2581,n2583);
and (n2581,n2582,n985);
xor (n2582,n2488,n2489);
and (n2583,n2584,n2585);
xor (n2584,n2582,n985);
or (n2585,n2586,n2589);
and (n2586,n2587,n2588);
xor (n2587,n2494,n2495);
and (n2588,n352,n47);
and (n2589,n2590,n2591);
xor (n2590,n2587,n2588);
or (n2591,n2592,n2595);
and (n2592,n2593,n2594);
xor (n2593,n2500,n2501);
and (n2594,n412,n47);
and (n2595,n2596,n2597);
xor (n2596,n2593,n2594);
or (n2597,n2598,n2601);
and (n2598,n2599,n2600);
xor (n2599,n2506,n2507);
and (n2600,n464,n47);
and (n2601,n2602,n2603);
xor (n2602,n2599,n2600);
or (n2603,n2604,n2607);
and (n2604,n2605,n2606);
xor (n2605,n2512,n2513);
and (n2606,n604,n47);
and (n2607,n2608,n2609);
xor (n2608,n2605,n2606);
or (n2609,n2610,n2613);
and (n2610,n2611,n2612);
xor (n2611,n2518,n2519);
and (n2612,n637,n47);
and (n2613,n2614,n2615);
xor (n2614,n2611,n2612);
and (n2615,n2616,n2617);
xor (n2616,n2524,n2525);
and (n2617,n698,n47);
and (n2618,n144,n46);
or (n2619,n2620,n2623);
and (n2620,n2621,n2622);
xor (n2621,n2529,n2530);
and (n2622,n40,n46);
and (n2623,n2624,n2625);
xor (n2624,n2621,n2622);
or (n2625,n2626,n2629);
and (n2626,n2627,n2628);
xor (n2627,n2535,n2536);
and (n2628,n57,n46);
and (n2629,n2630,n2631);
xor (n2630,n2627,n2628);
or (n2631,n2632,n2635);
and (n2632,n2633,n2634);
xor (n2633,n2541,n2542);
and (n2634,n30,n46);
and (n2635,n2636,n2637);
xor (n2636,n2633,n2634);
or (n2637,n2638,n2641);
and (n2638,n2639,n2640);
xor (n2639,n2546,n2547);
and (n2640,n24,n46);
and (n2641,n2642,n2643);
xor (n2642,n2639,n2640);
or (n2643,n2644,n2647);
and (n2644,n2645,n2646);
xor (n2645,n2551,n2552);
and (n2646,n121,n46);
and (n2647,n2648,n2649);
xor (n2648,n2645,n2646);
or (n2649,n2650,n2653);
and (n2650,n2651,n2652);
xor (n2651,n2557,n2558);
and (n2652,n85,n46);
and (n2653,n2654,n2655);
xor (n2654,n2651,n2652);
or (n2655,n2656,n2659);
and (n2656,n2657,n2658);
xor (n2657,n2562,n2563);
and (n2658,n68,n46);
and (n2659,n2660,n2661);
xor (n2660,n2657,n2658);
or (n2661,n2662,n2665);
and (n2662,n2663,n2664);
xor (n2663,n2567,n2568);
and (n2664,n107,n46);
and (n2665,n2666,n2667);
xor (n2666,n2663,n2664);
or (n2667,n2668,n2671);
and (n2668,n2669,n2670);
xor (n2669,n2573,n2574);
and (n2670,n96,n46);
and (n2671,n2672,n2673);
xor (n2672,n2669,n2670);
or (n2673,n2674,n2677);
and (n2674,n2675,n2676);
xor (n2675,n2579,n2580);
and (n2676,n262,n46);
and (n2677,n2678,n2679);
xor (n2678,n2675,n2676);
or (n2679,n2680,n2683);
and (n2680,n2681,n2682);
xor (n2681,n2584,n2585);
and (n2682,n352,n46);
and (n2683,n2684,n2685);
xor (n2684,n2681,n2682);
or (n2685,n2686,n2689);
and (n2686,n2687,n2688);
xor (n2687,n2590,n2591);
and (n2688,n412,n46);
and (n2689,n2690,n2691);
xor (n2690,n2687,n2688);
or (n2691,n2692,n2695);
and (n2692,n2693,n2694);
xor (n2693,n2596,n2597);
and (n2694,n464,n46);
and (n2695,n2696,n2697);
xor (n2696,n2693,n2694);
or (n2697,n2698,n2701);
and (n2698,n2699,n2700);
xor (n2699,n2602,n2603);
and (n2700,n604,n46);
and (n2701,n2702,n2703);
xor (n2702,n2699,n2700);
or (n2703,n2704,n2707);
and (n2704,n2705,n2706);
xor (n2705,n2608,n2609);
and (n2706,n637,n46);
and (n2707,n2708,n2709);
xor (n2708,n2705,n2706);
and (n2709,n2710,n1271);
xor (n2710,n2614,n2615);
and (n2711,n40,n16);
or (n2712,n2713,n2716);
and (n2713,n2714,n2715);
xor (n2714,n2624,n2625);
and (n2715,n57,n16);
and (n2716,n2717,n2718);
xor (n2717,n2714,n2715);
or (n2718,n2719,n2722);
and (n2719,n2720,n2721);
xor (n2720,n2630,n2631);
and (n2721,n30,n16);
and (n2722,n2723,n2724);
xor (n2723,n2720,n2721);
or (n2724,n2725,n2728);
and (n2725,n2726,n2727);
xor (n2726,n2636,n2637);
and (n2727,n24,n16);
and (n2728,n2729,n2730);
xor (n2729,n2726,n2727);
or (n2730,n2731,n2734);
and (n2731,n2732,n2733);
xor (n2732,n2642,n2643);
and (n2733,n121,n16);
and (n2734,n2735,n2736);
xor (n2735,n2732,n2733);
or (n2736,n2737,n2739);
and (n2737,n2738,n377);
xor (n2738,n2648,n2649);
and (n2739,n2740,n2741);
xor (n2740,n2738,n377);
or (n2741,n2742,n2744);
and (n2742,n2743,n471);
xor (n2743,n2654,n2655);
and (n2744,n2745,n2746);
xor (n2745,n2743,n471);
or (n2746,n2747,n2750);
and (n2747,n2748,n2749);
xor (n2748,n2660,n2661);
and (n2749,n107,n16);
and (n2750,n2751,n2752);
xor (n2751,n2748,n2749);
or (n2752,n2753,n2756);
and (n2753,n2754,n2755);
xor (n2754,n2666,n2667);
and (n2755,n96,n16);
and (n2756,n2757,n2758);
xor (n2757,n2754,n2755);
or (n2758,n2759,n2761);
and (n2759,n2760,n763);
xor (n2760,n2672,n2673);
and (n2761,n2762,n2763);
xor (n2762,n2760,n763);
or (n2763,n2764,n2767);
and (n2764,n2765,n2766);
xor (n2765,n2678,n2679);
and (n2766,n352,n16);
and (n2767,n2768,n2769);
xor (n2768,n2765,n2766);
or (n2769,n2770,n2773);
and (n2770,n2771,n2772);
xor (n2771,n2684,n2685);
and (n2772,n412,n16);
and (n2773,n2774,n2775);
xor (n2774,n2771,n2772);
or (n2775,n2776,n2779);
and (n2776,n2777,n2778);
xor (n2777,n2690,n2691);
and (n2778,n464,n16);
and (n2779,n2780,n2781);
xor (n2780,n2777,n2778);
or (n2781,n2782,n2785);
and (n2782,n2783,n2784);
xor (n2783,n2696,n2697);
and (n2784,n604,n16);
and (n2785,n2786,n2787);
xor (n2786,n2783,n2784);
or (n2787,n2788,n2791);
and (n2788,n2789,n2790);
xor (n2789,n2702,n2703);
and (n2790,n637,n16);
and (n2791,n2792,n2793);
xor (n2792,n2789,n2790);
and (n2793,n2794,n2795);
xor (n2794,n2708,n2709);
and (n2795,n698,n16);
and (n2796,n57,n15);
or (n2797,n2798,n2801);
and (n2798,n2799,n2800);
xor (n2799,n2717,n2718);
and (n2800,n30,n15);
and (n2801,n2802,n2803);
xor (n2802,n2799,n2800);
or (n2803,n2804,n2807);
and (n2804,n2805,n2806);
xor (n2805,n2723,n2724);
and (n2806,n24,n15);
and (n2807,n2808,n2809);
xor (n2808,n2805,n2806);
or (n2809,n2810,n2813);
and (n2810,n2811,n2812);
xor (n2811,n2729,n2730);
and (n2812,n121,n15);
and (n2813,n2814,n2815);
xor (n2814,n2811,n2812);
or (n2815,n2816,n2819);
and (n2816,n2817,n2818);
xor (n2817,n2735,n2736);
and (n2818,n85,n15);
and (n2819,n2820,n2821);
xor (n2820,n2817,n2818);
or (n2821,n2822,n2825);
and (n2822,n2823,n2824);
xor (n2823,n2740,n2741);
and (n2824,n68,n15);
and (n2825,n2826,n2827);
xor (n2826,n2823,n2824);
or (n2827,n2828,n2831);
and (n2828,n2829,n2830);
xor (n2829,n2745,n2746);
and (n2830,n107,n15);
and (n2831,n2832,n2833);
xor (n2832,n2829,n2830);
or (n2833,n2834,n2837);
and (n2834,n2835,n2836);
xor (n2835,n2751,n2752);
and (n2836,n96,n15);
and (n2837,n2838,n2839);
xor (n2838,n2835,n2836);
or (n2839,n2840,n2843);
and (n2840,n2841,n2842);
xor (n2841,n2757,n2758);
and (n2842,n262,n15);
and (n2843,n2844,n2845);
xor (n2844,n2841,n2842);
or (n2845,n2846,n2849);
and (n2846,n2847,n2848);
xor (n2847,n2762,n2763);
and (n2848,n352,n15);
and (n2849,n2850,n2851);
xor (n2850,n2847,n2848);
or (n2851,n2852,n2855);
and (n2852,n2853,n2854);
xor (n2853,n2768,n2769);
and (n2854,n412,n15);
and (n2855,n2856,n2857);
xor (n2856,n2853,n2854);
or (n2857,n2858,n2861);
and (n2858,n2859,n2860);
xor (n2859,n2774,n2775);
and (n2860,n464,n15);
and (n2861,n2862,n2863);
xor (n2862,n2859,n2860);
or (n2863,n2864,n2867);
and (n2864,n2865,n2866);
xor (n2865,n2780,n2781);
and (n2866,n604,n15);
and (n2867,n2868,n2869);
xor (n2868,n2865,n2866);
or (n2869,n2870,n2873);
and (n2870,n2871,n2872);
xor (n2871,n2786,n2787);
and (n2872,n637,n15);
and (n2873,n2874,n2875);
xor (n2874,n2871,n2872);
and (n2875,n2876,n2877);
xor (n2876,n2792,n2793);
not (n2877,n1070);
and (n2878,n30,n21);
or (n2879,n2880,n2883);
and (n2880,n2881,n2882);
xor (n2881,n2802,n2803);
and (n2882,n24,n21);
and (n2883,n2884,n2885);
xor (n2884,n2881,n2882);
or (n2885,n2886,n2889);
and (n2886,n2887,n2888);
xor (n2887,n2808,n2809);
and (n2888,n121,n21);
and (n2889,n2890,n2891);
xor (n2890,n2887,n2888);
or (n2891,n2892,n2895);
and (n2892,n2893,n2894);
xor (n2893,n2814,n2815);
and (n2894,n85,n21);
and (n2895,n2896,n2897);
xor (n2896,n2893,n2894);
or (n2897,n2898,n2901);
and (n2898,n2899,n2900);
xor (n2899,n2820,n2821);
and (n2900,n68,n21);
and (n2901,n2902,n2903);
xor (n2902,n2899,n2900);
or (n2903,n2904,n2907);
and (n2904,n2905,n2906);
xor (n2905,n2826,n2827);
and (n2906,n107,n21);
and (n2907,n2908,n2909);
xor (n2908,n2905,n2906);
or (n2909,n2910,n2913);
and (n2910,n2911,n2912);
xor (n2911,n2832,n2833);
and (n2912,n96,n21);
and (n2913,n2914,n2915);
xor (n2914,n2911,n2912);
or (n2915,n2916,n2919);
and (n2916,n2917,n2918);
xor (n2917,n2838,n2839);
and (n2918,n262,n21);
and (n2919,n2920,n2921);
xor (n2920,n2917,n2918);
or (n2921,n2922,n2925);
and (n2922,n2923,n2924);
xor (n2923,n2844,n2845);
and (n2924,n352,n21);
and (n2925,n2926,n2927);
xor (n2926,n2923,n2924);
or (n2927,n2928,n2931);
and (n2928,n2929,n2930);
xor (n2929,n2850,n2851);
and (n2930,n412,n21);
and (n2931,n2932,n2933);
xor (n2932,n2929,n2930);
or (n2933,n2934,n2937);
and (n2934,n2935,n2936);
xor (n2935,n2856,n2857);
and (n2936,n464,n21);
and (n2937,n2938,n2939);
xor (n2938,n2935,n2936);
or (n2939,n2940,n2943);
and (n2940,n2941,n2942);
xor (n2941,n2862,n2863);
and (n2942,n604,n21);
and (n2943,n2944,n2945);
xor (n2944,n2941,n2942);
or (n2945,n2946,n2949);
and (n2946,n2947,n2948);
xor (n2947,n2868,n2869);
and (n2948,n637,n21);
and (n2949,n2950,n2951);
xor (n2950,n2947,n2948);
and (n2951,n2952,n2953);
xor (n2952,n2874,n2875);
and (n2953,n698,n21);
and (n2954,n24,n76);
or (n2955,n2956,n2959);
and (n2956,n2957,n2958);
xor (n2957,n2884,n2885);
and (n2958,n121,n76);
and (n2959,n2960,n2961);
xor (n2960,n2957,n2958);
or (n2961,n2962,n2965);
and (n2962,n2963,n2964);
xor (n2963,n2890,n2891);
and (n2964,n85,n76);
and (n2965,n2966,n2967);
xor (n2966,n2963,n2964);
or (n2967,n2968,n2971);
and (n2968,n2969,n2970);
xor (n2969,n2896,n2897);
and (n2970,n68,n76);
and (n2971,n2972,n2973);
xor (n2972,n2969,n2970);
or (n2973,n2974,n2977);
and (n2974,n2975,n2976);
xor (n2975,n2902,n2903);
and (n2976,n107,n76);
and (n2977,n2978,n2979);
xor (n2978,n2975,n2976);
or (n2979,n2980,n2983);
and (n2980,n2981,n2982);
xor (n2981,n2908,n2909);
and (n2982,n96,n76);
and (n2983,n2984,n2985);
xor (n2984,n2981,n2982);
or (n2985,n2986,n2989);
and (n2986,n2987,n2988);
xor (n2987,n2914,n2915);
and (n2988,n262,n76);
and (n2989,n2990,n2991);
xor (n2990,n2987,n2988);
or (n2991,n2992,n2995);
and (n2992,n2993,n2994);
xor (n2993,n2920,n2921);
and (n2994,n352,n76);
and (n2995,n2996,n2997);
xor (n2996,n2993,n2994);
or (n2997,n2998,n3001);
and (n2998,n2999,n3000);
xor (n2999,n2926,n2927);
and (n3000,n412,n76);
and (n3001,n3002,n3003);
xor (n3002,n2999,n3000);
or (n3003,n3004,n3007);
and (n3004,n3005,n3006);
xor (n3005,n2932,n2933);
and (n3006,n464,n76);
and (n3007,n3008,n3009);
xor (n3008,n3005,n3006);
or (n3009,n3010,n3013);
and (n3010,n3011,n3012);
xor (n3011,n2938,n2939);
and (n3012,n604,n76);
and (n3013,n3014,n3015);
xor (n3014,n3011,n3012);
or (n3015,n3016,n3019);
and (n3016,n3017,n3018);
xor (n3017,n2944,n2945);
and (n3018,n637,n76);
and (n3019,n3020,n3021);
xor (n3020,n3017,n3018);
and (n3021,n3022,n3023);
xor (n3022,n2950,n2951);
not (n3023,n919);
and (n3024,n121,n70);
or (n3025,n3026,n3028);
and (n3026,n3027,n86);
xor (n3027,n2960,n2961);
and (n3028,n3029,n3030);
xor (n3029,n3027,n86);
or (n3030,n3031,n3033);
and (n3031,n3032,n71);
xor (n3032,n2966,n2967);
and (n3033,n3034,n3035);
xor (n3034,n3032,n71);
or (n3035,n3036,n3038);
and (n3036,n3037,n241);
xor (n3037,n2972,n2973);
and (n3038,n3039,n3040);
xor (n3039,n3037,n241);
or (n3040,n3041,n3044);
and (n3041,n3042,n3043);
xor (n3042,n2978,n2979);
and (n3043,n96,n70);
and (n3044,n3045,n3046);
xor (n3045,n3042,n3043);
or (n3046,n3047,n3050);
and (n3047,n3048,n3049);
xor (n3048,n2984,n2985);
and (n3049,n262,n70);
and (n3050,n3051,n3052);
xor (n3051,n3048,n3049);
or (n3052,n3053,n3055);
and (n3053,n3054,n501);
xor (n3054,n2990,n2991);
and (n3055,n3056,n3057);
xor (n3056,n3054,n501);
or (n3057,n3058,n3060);
and (n3058,n3059,n550);
xor (n3059,n2996,n2997);
and (n3060,n3061,n3062);
xor (n3061,n3059,n550);
or (n3062,n3063,n3065);
and (n3063,n3064,n632);
xor (n3064,n3002,n3003);
and (n3065,n3066,n3067);
xor (n3066,n3064,n632);
or (n3067,n3068,n3071);
and (n3068,n3069,n3070);
xor (n3069,n3008,n3009);
and (n3070,n604,n70);
and (n3071,n3072,n3073);
xor (n3072,n3069,n3070);
or (n3073,n3074,n3077);
and (n3074,n3075,n3076);
xor (n3075,n3014,n3015);
and (n3076,n637,n70);
and (n3077,n3078,n3079);
xor (n3078,n3075,n3076);
and (n3079,n3080,n3081);
xor (n3080,n3020,n3021);
and (n3081,n698,n70);
and (n3082,n85,n100);
or (n3083,n3084,n3087);
and (n3084,n3085,n3086);
xor (n3085,n3029,n3030);
and (n3086,n68,n100);
and (n3087,n3088,n3089);
xor (n3088,n3085,n3086);
or (n3089,n3090,n3093);
and (n3090,n3091,n3092);
xor (n3091,n3034,n3035);
and (n3092,n107,n100);
and (n3093,n3094,n3095);
xor (n3094,n3091,n3092);
or (n3095,n3096,n3099);
and (n3096,n3097,n3098);
xor (n3097,n3039,n3040);
and (n3098,n96,n100);
and (n3099,n3100,n3101);
xor (n3100,n3097,n3098);
or (n3101,n3102,n3105);
and (n3102,n3103,n3104);
xor (n3103,n3045,n3046);
and (n3104,n262,n100);
and (n3105,n3106,n3107);
xor (n3106,n3103,n3104);
or (n3107,n3108,n3111);
and (n3108,n3109,n3110);
xor (n3109,n3051,n3052);
and (n3110,n352,n100);
and (n3111,n3112,n3113);
xor (n3112,n3109,n3110);
or (n3113,n3114,n3117);
and (n3114,n3115,n3116);
xor (n3115,n3056,n3057);
and (n3116,n412,n100);
and (n3117,n3118,n3119);
xor (n3118,n3115,n3116);
or (n3119,n3120,n3123);
and (n3120,n3121,n3122);
xor (n3121,n3061,n3062);
and (n3122,n464,n100);
and (n3123,n3124,n3125);
xor (n3124,n3121,n3122);
or (n3125,n3126,n3129);
and (n3126,n3127,n3128);
xor (n3127,n3066,n3067);
and (n3128,n604,n100);
and (n3129,n3130,n3131);
xor (n3130,n3127,n3128);
or (n3131,n3132,n3135);
and (n3132,n3133,n3134);
xor (n3133,n3072,n3073);
and (n3134,n637,n100);
and (n3135,n3136,n3137);
xor (n3136,n3133,n3134);
and (n3137,n3138,n3139);
xor (n3138,n3078,n3079);
and (n3139,n698,n100);
endmodule
