module top (out,n19,n20,n24,n26,n28,n29,n30,n33,n34
        ,n38,n40,n42,n43,n46,n48,n50,n52,n53,n54
        ,n55,n56,n57,n58,n59,n60,n61,n62,n63,n64
        ,n65,n66,n67,n68,n69,n70,n71,n72,n73,n74
        ,n75,n76,n77,n78,n79,n80,n88,n89,n90,n97
        ,n98,n99,n106,n107,n108,n117,n118,n119,n123,n124
        ,n125,n133,n134,n135,n143,n144,n145,n159,n160,n161
        ,n164,n165,n166,n176,n177,n178,n185,n186,n187,n194
        ,n195,n196,n209,n210,n211,n230,n231,n232,n248,n249
        ,n250,n269,n270,n271,n279,n280,n281,n309,n310,n311
        ,n333,n334,n335,n353,n354,n355,n623,n624,n628,n630
        ,n632,n635,n636,n640,n642,n644,n645,n648,n650,n652
        ,n654,n655,n656,n657,n658,n659,n660,n661,n662,n663
        ,n664,n665,n666,n667,n668,n669,n670,n671,n672,n673
        ,n674,n675,n676,n677,n678,n679,n680,n681,n682,n685
        ,n686,n689,n690,n691);
output out;
input n19;
input n20;
input n24;
input n26;
input n28;
input n29;
input n30;
input n33;
input n34;
input n38;
input n40;
input n42;
input n43;
input n46;
input n48;
input n50;
input n52;
input n53;
input n54;
input n55;
input n56;
input n57;
input n58;
input n59;
input n60;
input n61;
input n62;
input n63;
input n64;
input n65;
input n66;
input n67;
input n68;
input n69;
input n70;
input n71;
input n72;
input n73;
input n74;
input n75;
input n76;
input n77;
input n78;
input n79;
input n80;
input n88;
input n89;
input n90;
input n97;
input n98;
input n99;
input n106;
input n107;
input n108;
input n117;
input n118;
input n119;
input n123;
input n124;
input n125;
input n133;
input n134;
input n135;
input n143;
input n144;
input n145;
input n159;
input n160;
input n161;
input n164;
input n165;
input n166;
input n176;
input n177;
input n178;
input n185;
input n186;
input n187;
input n194;
input n195;
input n196;
input n209;
input n210;
input n211;
input n230;
input n231;
input n232;
input n248;
input n249;
input n250;
input n269;
input n270;
input n271;
input n279;
input n280;
input n281;
input n309;
input n310;
input n311;
input n333;
input n334;
input n335;
input n353;
input n354;
input n355;
input n623;
input n624;
input n628;
input n630;
input n632;
input n635;
input n636;
input n640;
input n642;
input n644;
input n645;
input n648;
input n650;
input n652;
input n654;
input n655;
input n656;
input n657;
input n658;
input n659;
input n660;
input n661;
input n662;
input n663;
input n664;
input n665;
input n666;
input n667;
input n668;
input n669;
input n670;
input n671;
input n672;
input n673;
input n674;
input n675;
input n676;
input n677;
input n678;
input n679;
input n680;
input n681;
input n682;
input n685;
input n686;
input n689;
input n690;
input n691;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n21;
wire n22;
wire n23;
wire n25;
wire n27;
wire n31;
wire n32;
wire n35;
wire n36;
wire n37;
wire n39;
wire n41;
wire n44;
wire n45;
wire n47;
wire n49;
wire n51;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n120;
wire n121;
wire n122;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n162;
wire n163;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n173;
wire n174;
wire n175;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n625;
wire n626;
wire n627;
wire n629;
wire n631;
wire n633;
wire n634;
wire n637;
wire n638;
wire n639;
wire n641;
wire n643;
wire n646;
wire n647;
wire n649;
wire n651;
wire n653;
wire n683;
wire n684;
wire n687;
wire n688;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
xor (out,n0,n696);
and (n0,n1,n614);
nand (n1,n2,n613);
or (n2,n3,n396);
not (n3,n4);
nand (n4,n5,n395);
not (n5,n6);
nor (n6,n7,n357);
xor (n7,n8,n294);
xor (n8,n9,n198);
xor (n9,n10,n152);
xor (n10,n11,n110);
nand (n11,n12,n101);
or (n12,n13,n82);
not (n13,n14);
nand (n14,n15,n81);
or (n15,n16,n31);
not (n16,n17);
wire s0n17,s1n17,notn17;
or (n17,s0n17,s1n17);
not(notn17,n30);
and (s0n17,notn17,n18);
and (s1n17,n30,n29);
wire s0n18,s1n18,notn18;
or (n18,s0n18,s1n18);
not(notn18,n21);
and (s0n18,notn18,n19);
and (s1n18,n21,n20);
and (n21,n22,n27);
and (n22,n23,n25);
not (n23,n24);
not (n25,n26);
not (n27,n28);
wire s0n31,s1n31,notn31;
or (n31,s0n31,s1n31);
not(notn31,n44);
and (s0n31,notn31,n32);
and (s1n31,n44,n43);
wire s0n32,s1n32,notn32;
or (n32,s0n32,s1n32);
not(notn32,n35);
and (s0n32,notn32,n33);
and (s1n32,n35,n34);
and (n35,n36,n41);
and (n36,n37,n39);
not (n37,n38);
not (n39,n40);
not (n41,n42);
and (n44,n45,n47);
not (n45,n46);
or (n47,n48,n49);
and (n49,n50,n51);
or (n51,n52,n53,n54,n55,n56,n57,n58,n59,n60,n61,n62,n63,n64,n65,n66,n67,n68,n69,n70,n71,n72,n73,n74,n75,n76,n77,n78,n79,n80);
nand (n81,n16,n31);
not (n82,n83);
nor (n83,n84,n93);
nor (n84,n85,n91);
and (n85,n16,n86);
wire s0n86,s1n86,notn86;
or (n86,s0n86,s1n86);
not(notn86,n30);
and (s0n86,notn86,n87);
and (s1n86,n30,n90);
wire s0n87,s1n87,notn87;
or (n87,s0n87,s1n87);
not(notn87,n21);
and (s0n87,notn87,n88);
and (s1n87,n21,n89);
and (n91,n17,n92);
not (n92,n86);
nand (n93,n94,n100);
or (n94,n92,n95);
wire s0n95,s1n95,notn95;
or (n95,s0n95,s1n95);
not(notn95,n30);
and (s0n95,notn95,n96);
and (s1n95,n30,n99);
wire s0n96,s1n96,notn96;
or (n96,s0n96,s1n96);
not(notn96,n21);
and (s0n96,notn96,n97);
and (s1n96,n21,n98);
nand (n100,n95,n92);
nand (n101,n102,n93);
nand (n102,n103,n109);
or (n103,n16,n104);
wire s0n104,s1n104,notn104;
or (n104,s0n104,s1n104);
not(notn104,n44);
and (s0n104,notn104,n105);
and (s1n104,n44,n108);
wire s0n105,s1n105,notn105;
or (n105,s0n105,s1n105);
not(notn105,n35);
and (s0n105,notn105,n106);
and (s1n105,n35,n107);
nand (n109,n16,n104);
nand (n110,n111,n137);
or (n111,n112,n127);
not (n112,n113);
nand (n113,n114,n126);
or (n114,n115,n120);
wire s0n115,s1n115,notn115;
or (n115,s0n115,s1n115);
not(notn115,n30);
and (s0n115,notn115,n116);
and (s1n115,n30,n119);
wire s0n116,s1n116,notn116;
or (n116,s0n116,s1n116);
not(notn116,n21);
and (s0n116,notn116,n117);
and (s1n116,n21,n118);
not (n120,n121);
wire s0n121,s1n121,notn121;
or (n121,s0n121,s1n121);
not(notn121,n30);
and (s0n121,notn121,n122);
and (s1n121,n30,n125);
wire s0n122,s1n122,notn122;
or (n122,s0n122,s1n122);
not(notn122,n21);
and (s0n122,notn122,n123);
and (s1n122,n21,n124);
nand (n126,n120,n115);
not (n127,n128);
nand (n128,n129,n136);
or (n129,n130,n131);
not (n130,n95);
wire s0n131,s1n131,notn131;
or (n131,s0n131,s1n131);
not(notn131,n44);
and (s0n131,notn131,n132);
and (s1n131,n44,n135);
wire s0n132,s1n132,notn132;
or (n132,s0n132,s1n132);
not(notn132,n35);
and (s0n132,notn132,n133);
and (s1n132,n35,n134);
nand (n136,n131,n130);
nand (n137,n138,n147);
nand (n138,n139,n146);
or (n139,n95,n140);
not (n140,n141);
wire s0n141,s1n141,notn141;
or (n141,s0n141,s1n141);
not(notn141,n44);
and (s0n141,notn141,n142);
and (s1n141,n44,n145);
wire s0n142,s1n142,notn142;
or (n142,s0n142,s1n142);
not(notn142,n35);
and (s0n142,notn142,n143);
and (s1n142,n35,n144);
nand (n146,n140,n95);
not (n147,n148);
nand (n148,n112,n149);
nand (n149,n150,n151);
or (n150,n120,n95);
nand (n151,n95,n120);
nand (n152,n153,n189);
or (n153,n154,n170);
not (n154,n155);
nor (n155,n156,n167);
and (n156,n157,n162);
wire s0n157,s1n157,notn157;
or (n157,s0n157,s1n157);
not(notn157,n44);
and (s0n157,notn157,n158);
and (s1n157,n44,n161);
wire s0n158,s1n158,notn158;
or (n158,s0n158,s1n158);
not(notn158,n35);
and (s0n158,notn158,n159);
and (s1n158,n35,n160);
wire s0n162,s1n162,notn162;
or (n162,s0n162,s1n162);
not(notn162,n30);
and (s0n162,notn162,n163);
and (s1n162,n30,n166);
wire s0n163,s1n163,notn163;
or (n163,s0n163,s1n163);
not(notn163,n21);
and (s0n163,notn163,n164);
and (s1n163,n21,n165);
and (n167,n168,n169);
not (n168,n162);
not (n169,n157);
not (n170,n171);
nor (n171,n172,n181);
nor (n172,n173,n179);
and (n173,n168,n174);
wire s0n174,s1n174,notn174;
or (n174,s0n174,s1n174);
not(notn174,n30);
and (s0n174,notn174,n175);
and (s1n174,n30,n178);
wire s0n175,s1n175,notn175;
or (n175,s0n175,s1n175);
not(notn175,n21);
and (s0n175,notn175,n176);
and (s1n175,n21,n177);
and (n179,n162,n180);
not (n180,n174);
nand (n181,n182,n188);
or (n182,n183,n180);
wire s0n183,s1n183,notn183;
or (n183,s0n183,s1n183);
not(notn183,n30);
and (s0n183,notn183,n184);
and (s1n183,n30,n187);
wire s0n184,s1n184,notn184;
or (n184,s0n184,s1n184);
not(notn184,n21);
and (s0n184,notn184,n185);
and (s1n184,n21,n186);
nand (n188,n180,n183);
nand (n189,n190,n181);
nand (n190,n191,n197);
or (n191,n168,n192);
wire s0n192,s1n192,notn192;
or (n192,s0n192,s1n192);
not(notn192,n44);
and (s0n192,notn192,n193);
and (s1n192,n44,n196);
wire s0n193,s1n193,notn193;
or (n193,s0n193,s1n193);
not(notn193,n35);
and (s0n193,notn193,n194);
and (s1n193,n35,n195);
nand (n197,n192,n168);
or (n198,n199,n293);
and (n199,n200,n252);
xor (n200,n201,n214);
nand (n201,n202,n213);
or (n202,n82,n203);
not (n203,n204);
nor (n204,n205,n212);
and (n205,n16,n206);
not (n206,n207);
wire s0n207,s1n207,notn207;
or (n207,s0n207,s1n207);
not(notn207,n44);
and (s0n207,notn207,n208);
and (s1n207,n44,n211);
wire s0n208,s1n208,notn208;
or (n208,s0n208,s1n208);
not(notn208,n35);
and (s0n208,notn208,n209);
and (s1n208,n35,n210);
and (n212,n207,n17);
nand (n213,n93,n14);
xor (n214,n215,n221);
nor (n215,n216,n16);
and (n216,n217,n220);
nand (n217,n218,n130);
not (n218,n219);
and (n219,n207,n86);
nand (n220,n206,n92);
nand (n221,n222,n243);
or (n222,n223,n238);
not (n223,n224);
nor (n224,n225,n234);
nand (n225,n226,n233);
or (n226,n227,n162);
not (n227,n228);
wire s0n228,s1n228,notn228;
or (n228,s0n228,s1n228);
not(notn228,n30);
and (s0n228,notn228,n229);
and (s1n228,n30,n232);
wire s0n229,s1n229,notn229;
or (n229,s0n229,s1n229);
not(notn229,n21);
and (s0n229,notn229,n230);
and (s1n229,n21,n231);
nand (n233,n162,n227);
not (n234,n235);
nand (n235,n236,n237);
or (n236,n115,n227);
nand (n237,n227,n115);
not (n238,n239);
nand (n239,n240,n242);
or (n240,n241,n131);
not (n241,n115);
nand (n242,n131,n241);
nand (n243,n244,n225);
nand (n244,n245,n251);
or (n245,n241,n246);
wire s0n246,s1n246,notn246;
or (n246,s0n246,s1n246);
not(notn246,n44);
and (s0n246,notn246,n247);
and (s1n246,n44,n250);
wire s0n247,s1n247,notn247;
or (n247,s0n247,s1n247);
not(notn247,n35);
and (s0n247,notn247,n248);
and (s1n247,n35,n249);
nand (n251,n246,n241);
or (n252,n253,n292);
and (n253,n254,n273);
xor (n254,n255,n256);
and (n255,n93,n207);
nand (n256,n257,n263);
or (n257,n258,n170);
not (n258,n259);
nand (n259,n260,n262);
or (n260,n162,n261);
not (n261,n246);
nand (n262,n261,n162);
nand (n263,n264,n181);
nand (n264,n265,n272);
or (n265,n162,n266);
not (n266,n267);
wire s0n267,s1n267,notn267;
or (n267,s0n267,s1n267);
not(notn267,n44);
and (s0n267,notn267,n268);
and (s1n267,n44,n271);
wire s0n268,s1n268,notn268;
or (n268,s0n268,s1n268);
not(notn268,n35);
and (s0n268,notn268,n269);
and (s1n268,n35,n270);
nand (n272,n266,n162);
nand (n273,n274,n287);
or (n274,n275,n283);
not (n275,n276);
nor (n276,n277,n282);
wire s0n277,s1n277,notn277;
or (n277,s0n277,s1n277);
not(notn277,n30);
and (s0n277,notn277,n278);
and (s1n277,n30,n281);
wire s0n278,s1n278,notn278;
or (n278,s0n278,s1n278);
not(notn278,n21);
and (s0n278,notn278,n279);
and (s1n278,n21,n280);
not (n282,n183);
not (n283,n284);
nand (n284,n285,n286);
or (n285,n183,n169);
nand (n286,n169,n183);
nand (n287,n288,n277);
nand (n288,n289,n291);
or (n289,n183,n290);
not (n290,n192);
nand (n291,n290,n183);
and (n292,n255,n256);
and (n293,n201,n214);
xor (n294,n295,n325);
xor (n295,n296,n297);
and (n296,n215,n221);
or (n297,n298,n324);
and (n298,n299,n317);
xor (n299,n300,n313);
nand (n300,n301,n303);
or (n301,n275,n302);
not (n302,n288);
nand (n303,n304,n277);
nand (n304,n305,n312);
or (n305,n183,n306);
not (n306,n307);
wire s0n307,s1n307,notn307;
or (n307,s0n307,s1n307);
not(notn307,n44);
and (s0n307,notn307,n308);
and (s1n307,n44,n311);
wire s0n308,s1n308,notn308;
or (n308,s0n308,s1n308);
not(notn308,n35);
and (s0n308,notn308,n309);
and (s1n308,n35,n310);
nand (n312,n306,n183);
nand (n313,n314,n316);
or (n314,n315,n170);
not (n315,n264);
nand (n316,n155,n181);
nand (n317,n318,n323);
or (n318,n319,n148);
not (n319,n320);
nand (n320,n321,n322);
or (n321,n130,n104);
nand (n322,n104,n130);
nand (n323,n138,n113);
and (n324,n300,n313);
xor (n325,n326,n344);
xor (n326,n327,n337);
nor (n327,n206,n328);
nor (n328,n329,n336);
and (n329,n17,n330);
not (n330,n331);
wire s0n331,s1n331,notn331;
or (n331,s0n331,s1n331);
not(notn331,n30);
and (s0n331,notn331,n332);
and (s1n331,n30,n335);
wire s0n332,s1n332,notn332;
or (n332,s0n332,s1n332);
not(notn332,n21);
and (s0n332,notn332,n333);
and (s1n332,n21,n334);
and (n336,n16,n331);
nand (n337,n338,n340);
or (n338,n223,n339);
not (n339,n244);
nand (n340,n341,n225);
nand (n341,n342,n343);
or (n342,n115,n266);
nand (n343,n266,n115);
nand (n344,n345,n347);
or (n345,n346,n275);
not (n346,n304);
nand (n347,n348,n277);
nand (n348,n349,n356);
or (n349,n183,n350);
not (n350,n351);
wire s0n351,s1n351,notn351;
or (n351,s0n351,s1n351);
not(notn351,n44);
and (s0n351,notn351,n352);
and (s1n351,n44,n355);
wire s0n352,s1n352,notn352;
or (n352,s0n352,s1n352);
not(notn352,n35);
and (s0n352,notn352,n353);
and (s1n352,n35,n354);
nand (n356,n350,n183);
or (n357,n358,n394);
and (n358,n359,n393);
xor (n359,n360,n361);
xor (n360,n299,n317);
or (n361,n362,n392);
and (n362,n363,n378);
xor (n363,n364,n371);
nand (n364,n365,n370);
or (n365,n366,n148);
not (n366,n367);
nand (n367,n368,n369);
or (n368,n130,n31);
nand (n369,n31,n130);
nand (n370,n320,n113);
nand (n371,n372,n377);
or (n372,n373,n223);
not (n373,n374);
nand (n374,n375,n376);
or (n375,n241,n141);
nand (n376,n141,n241);
nand (n377,n239,n225);
and (n378,n379,n386);
nand (n379,n380,n385);
or (n380,n381,n170);
not (n381,n382);
nand (n382,n383,n384);
or (n383,n168,n131);
nand (n384,n131,n168);
nand (n385,n259,n181);
nor (n386,n387,n130);
and (n387,n388,n391);
nand (n388,n389,n241);
not (n389,n390);
and (n390,n207,n121);
nand (n391,n206,n120);
and (n392,n364,n371);
xor (n393,n200,n252);
and (n394,n360,n361);
nand (n395,n7,n357);
not (n396,n397);
nand (n397,n398,n608);
or (n398,n399,n464);
not (n399,n400);
nor (n400,n401,n434);
nor (n401,n402,n403);
xor (n402,n359,n393);
or (n403,n404,n433);
and (n404,n405,n432);
xor (n405,n406,n431);
or (n406,n407,n430);
and (n407,n408,n423);
xor (n408,n409,n416);
nand (n409,n410,n415);
or (n410,n275,n411);
not (n411,n412);
nand (n412,n413,n414);
or (n413,n183,n266);
nand (n414,n266,n183);
nand (n415,n284,n277);
nand (n416,n417,n422);
or (n417,n418,n148);
not (n418,n419);
nand (n419,n420,n421);
or (n420,n95,n206);
or (n421,n207,n130);
nand (n422,n367,n113);
nand (n423,n424,n429);
or (n424,n425,n223);
not (n425,n426);
nand (n426,n427,n428);
or (n427,n241,n104);
nand (n428,n104,n241);
nand (n429,n374,n225);
and (n430,n409,n416);
xor (n431,n254,n273);
xor (n432,n363,n378);
and (n433,n406,n431);
nor (n434,n435,n436);
xor (n435,n405,n432);
or (n436,n437,n463);
and (n437,n438,n462);
xor (n438,n439,n443);
nand (n439,n440,n442);
or (n440,n386,n441);
not (n441,n379);
nand (n442,n441,n386);
or (n443,n444,n461);
and (n444,n445,n454);
xor (n445,n446,n447);
and (n446,n113,n207);
nand (n447,n448,n453);
or (n448,n449,n170);
not (n449,n450);
nand (n450,n451,n452);
or (n451,n162,n140);
nand (n452,n140,n162);
nand (n453,n382,n181);
nand (n454,n455,n460);
or (n455,n456,n223);
not (n456,n457);
nand (n457,n458,n459);
or (n458,n241,n31);
nand (n459,n31,n241);
nand (n460,n426,n225);
and (n461,n446,n447);
xor (n462,n408,n423);
and (n463,n439,n443);
not (n464,n465);
nand (n465,n466,n607);
or (n466,n467,n498);
not (n467,n468);
nand (n468,n469,n471);
not (n469,n470);
xor (n470,n438,n462);
not (n471,n472);
or (n472,n473,n497);
and (n473,n474,n496);
xor (n474,n475,n482);
nand (n475,n476,n481);
or (n476,n275,n477);
not (n477,n478);
nand (n478,n479,n480);
or (n479,n282,n246);
nand (n480,n246,n282);
nand (n481,n412,n277);
and (n482,n483,n489);
nor (n483,n484,n241);
and (n484,n485,n488);
nand (n485,n486,n168);
not (n486,n487);
and (n487,n207,n228);
nand (n488,n206,n227);
nand (n489,n490,n495);
or (n490,n491,n170);
not (n491,n492);
nand (n492,n493,n494);
or (n493,n168,n104);
nand (n494,n104,n168);
nand (n495,n450,n181);
xor (n496,n445,n454);
and (n497,n475,n482);
not (n498,n499);
nand (n499,n500,n606);
or (n500,n501,n601);
nor (n501,n502,n600);
and (n502,n503,n543);
nand (n503,n504,n523);
not (n504,n505);
xor (n505,n506,n522);
xor (n506,n507,n514);
nand (n507,n508,n513);
or (n508,n509,n223);
not (n509,n510);
nor (n510,n511,n512);
and (n511,n207,n115);
and (n512,n241,n206);
nand (n513,n225,n457);
nand (n514,n515,n517);
or (n515,n516,n477);
not (n516,n277);
nand (n517,n518,n276);
nand (n518,n519,n521);
or (n519,n183,n520);
not (n520,n131);
nand (n521,n183,n520);
xor (n522,n483,n489);
not (n523,n524);
or (n524,n525,n542);
and (n525,n526,n535);
xor (n526,n527,n528);
and (n527,n225,n207);
nand (n528,n529,n531);
or (n529,n516,n530);
not (n530,n518);
nand (n531,n532,n276);
nand (n532,n533,n534);
or (n533,n183,n140);
nand (n534,n140,n183);
nand (n535,n536,n541);
or (n536,n537,n170);
not (n537,n538);
nand (n538,n539,n540);
or (n539,n168,n31);
nand (n540,n31,n168);
nand (n541,n492,n181);
and (n542,n527,n528);
nand (n543,n544,n598);
or (n544,n545,n563);
not (n545,n546);
nand (n546,n547,n549);
not (n547,n548);
xor (n548,n526,n535);
nand (n549,n550,n557);
nand (n550,n551,n553);
or (n551,n516,n552);
not (n552,n532);
nand (n553,n554,n276);
nand (n554,n555,n556);
or (n555,n282,n104);
nand (n556,n104,n282);
nor (n557,n558,n168);
and (n558,n559,n562);
nand (n559,n560,n282);
not (n560,n561);
and (n561,n207,n174);
nand (n562,n206,n180);
not (n563,n564);
or (n564,n565,n597);
and (n565,n566,n578);
xor (n566,n567,n574);
nand (n567,n568,n573);
or (n568,n569,n170);
not (n569,n570);
nor (n570,n571,n572);
and (n571,n207,n162);
and (n572,n168,n206);
nand (n573,n181,n538);
nand (n574,n575,n577);
or (n575,n576,n550);
not (n576,n557);
nand (n577,n550,n576);
or (n578,n579,n596);
and (n579,n580,n589);
xor (n580,n581,n582);
and (n581,n207,n181);
nand (n582,n583,n585);
or (n583,n516,n584);
not (n584,n554);
nand (n585,n586,n276);
nand (n586,n587,n588);
or (n587,n282,n31);
nand (n588,n31,n282);
nor (n589,n590,n593);
nor (n590,n591,n592);
and (n591,n276,n206);
and (n592,n586,n277);
nand (n593,n594,n183);
not (n594,n595);
and (n595,n207,n277);
and (n596,n581,n582);
and (n597,n567,n574);
nand (n598,n548,n599);
not (n599,n549);
and (n600,n505,n524);
nor (n601,n602,n603);
xor (n602,n474,n496);
or (n603,n604,n605);
and (n604,n506,n522);
and (n605,n507,n514);
nand (n606,n602,n603);
nand (n607,n470,n472);
not (n608,n609);
nand (n609,n610,n612);
or (n610,n401,n611);
nand (n611,n435,n436);
nand (n612,n402,n403);
nand (n613,n396,n3);
xor (n614,n615,n692);
xor (n615,n616,n619);
xor (n616,n617,n618);
and (n617,n184,n207);
and (n618,n278,n31);
not (n619,n620);
xor (n620,n621,n683);
and (n621,n622,n633);
wire s0n622,s1n622,notn622;
or (n622,s0n622,s1n622);
not(notn622,n625);
and (s0n622,notn622,n623);
and (s1n622,n625,n624);
and (n625,n626,n631);
and (n626,n627,n629);
not (n627,n628);
not (n629,n630);
not (n631,n632);
wire s0n633,s1n633,notn633;
or (n633,s0n633,s1n633);
not(notn633,n646);
and (s0n633,notn633,n634);
and (s1n633,n646,n645);
wire s0n634,s1n634,notn634;
or (n634,s0n634,s1n634);
not(notn634,n637);
and (s0n634,notn634,n635);
and (s1n634,n637,n636);
and (n637,n638,n643);
and (n638,n639,n641);
not (n639,n640);
not (n641,n642);
not (n643,n644);
and (n646,n647,n649);
not (n647,n648);
or (n649,n650,n651);
and (n651,n652,n653);
or (n653,n654,n655,n656,n657,n658,n659,n660,n661,n662,n663,n664,n665,n666,n667,n668,n669,n670,n671,n672,n673,n674,n675,n676,n677,n678,n679,n680,n681,n682);
and (n683,n684,n687);
wire s0n684,s1n684,notn684;
or (n684,s0n684,s1n684);
not(notn684,n625);
and (s0n684,notn684,n685);
and (s1n684,n625,n686);
wire s0n687,s1n687,notn687;
or (n687,s0n687,s1n687);
not(notn687,n646);
and (s0n687,notn687,n688);
and (s1n687,n646,n691);
wire s0n688,s1n688,notn688;
or (n688,s0n688,s1n688);
not(notn688,n637);
and (s0n688,notn688,n689);
and (s1n688,n637,n690);
or (n692,n693,n694);
and (n693,n278,n207);
not (n694,n695);
and (n695,n684,n633);
and (n696,n614,n697);
xor (n697,n698,n961);
xor (n698,n699,n959);
xor (n699,n700,n958);
xor (n700,n701,n950);
xor (n701,n702,n949);
xor (n702,n703,n934);
xor (n703,n704,n933);
xor (n704,n705,n913);
xor (n705,n706,n912);
xor (n706,n707,n886);
xor (n707,n708,n885);
xor (n708,n709,n853);
xor (n709,n710,n852);
xor (n710,n711,n814);
xor (n711,n712,n156);
xor (n712,n713,n770);
xor (n713,n714,n769);
xor (n714,n715,n718);
xor (n715,n716,n717);
and (n716,n351,n277);
and (n717,n307,n183);
or (n718,n719,n722);
and (n719,n720,n721);
and (n720,n307,n277);
and (n721,n192,n183);
and (n722,n723,n724);
xor (n723,n720,n721);
or (n724,n725,n728);
and (n725,n726,n727);
and (n726,n192,n277);
and (n727,n157,n183);
and (n728,n729,n730);
xor (n729,n726,n727);
or (n730,n731,n734);
and (n731,n732,n733);
and (n732,n157,n277);
and (n733,n267,n183);
and (n734,n735,n736);
xor (n735,n732,n733);
or (n736,n737,n740);
and (n737,n738,n739);
and (n738,n267,n277);
and (n739,n246,n183);
and (n740,n741,n742);
xor (n741,n738,n739);
or (n742,n743,n746);
and (n743,n744,n745);
and (n744,n246,n277);
and (n745,n131,n183);
and (n746,n747,n748);
xor (n747,n744,n745);
or (n748,n749,n752);
and (n749,n750,n751);
and (n750,n131,n277);
and (n751,n141,n183);
and (n752,n753,n754);
xor (n753,n750,n751);
or (n754,n755,n758);
and (n755,n756,n757);
and (n756,n141,n277);
and (n757,n104,n183);
and (n758,n759,n760);
xor (n759,n756,n757);
or (n760,n761,n764);
and (n761,n762,n763);
and (n762,n104,n277);
and (n763,n31,n183);
and (n764,n765,n766);
xor (n765,n762,n763);
and (n766,n767,n768);
and (n767,n31,n277);
and (n768,n207,n183);
and (n769,n192,n174);
or (n770,n771,n774);
and (n771,n772,n773);
xor (n772,n723,n724);
and (n773,n157,n174);
and (n774,n775,n776);
xor (n775,n772,n773);
or (n776,n777,n780);
and (n777,n778,n779);
xor (n778,n729,n730);
and (n779,n267,n174);
and (n780,n781,n782);
xor (n781,n778,n779);
or (n782,n783,n786);
and (n783,n784,n785);
xor (n784,n735,n736);
and (n785,n246,n174);
and (n786,n787,n788);
xor (n787,n784,n785);
or (n788,n789,n792);
and (n789,n790,n791);
xor (n790,n741,n742);
and (n791,n131,n174);
and (n792,n793,n794);
xor (n793,n790,n791);
or (n794,n795,n798);
and (n795,n796,n797);
xor (n796,n747,n748);
and (n797,n141,n174);
and (n798,n799,n800);
xor (n799,n796,n797);
or (n800,n801,n804);
and (n801,n802,n803);
xor (n802,n753,n754);
and (n803,n104,n174);
and (n804,n805,n806);
xor (n805,n802,n803);
or (n806,n807,n810);
and (n807,n808,n809);
xor (n808,n759,n760);
and (n809,n31,n174);
and (n810,n811,n812);
xor (n811,n808,n809);
and (n812,n813,n561);
xor (n813,n765,n766);
or (n814,n815,n818);
and (n815,n816,n817);
xor (n816,n775,n776);
and (n817,n267,n162);
and (n818,n819,n820);
xor (n819,n816,n817);
or (n820,n821,n824);
and (n821,n822,n823);
xor (n822,n781,n782);
and (n823,n246,n162);
and (n824,n825,n826);
xor (n825,n822,n823);
or (n826,n827,n830);
and (n827,n828,n829);
xor (n828,n787,n788);
and (n829,n131,n162);
and (n830,n831,n832);
xor (n831,n828,n829);
or (n832,n833,n836);
and (n833,n834,n835);
xor (n834,n793,n794);
and (n835,n141,n162);
and (n836,n837,n838);
xor (n837,n834,n835);
or (n838,n839,n842);
and (n839,n840,n841);
xor (n840,n799,n800);
and (n841,n104,n162);
and (n842,n843,n844);
xor (n843,n840,n841);
or (n844,n845,n848);
and (n845,n846,n847);
xor (n846,n805,n806);
and (n847,n31,n162);
and (n848,n849,n850);
xor (n849,n846,n847);
and (n850,n851,n571);
xor (n851,n811,n812);
and (n852,n267,n228);
or (n853,n854,n857);
and (n854,n855,n856);
xor (n855,n819,n820);
and (n856,n246,n228);
and (n857,n858,n859);
xor (n858,n855,n856);
or (n859,n860,n863);
and (n860,n861,n862);
xor (n861,n825,n826);
and (n862,n131,n228);
and (n863,n864,n865);
xor (n864,n861,n862);
or (n865,n866,n869);
and (n866,n867,n868);
xor (n867,n831,n832);
and (n868,n141,n228);
and (n869,n870,n871);
xor (n870,n867,n868);
or (n871,n872,n875);
and (n872,n873,n874);
xor (n873,n837,n838);
and (n874,n104,n228);
and (n875,n876,n877);
xor (n876,n873,n874);
or (n877,n878,n881);
and (n878,n879,n880);
xor (n879,n843,n844);
and (n880,n31,n228);
and (n881,n882,n883);
xor (n882,n879,n880);
and (n883,n884,n487);
xor (n884,n849,n850);
and (n885,n246,n115);
or (n886,n887,n890);
and (n887,n888,n889);
xor (n888,n858,n859);
and (n889,n131,n115);
and (n890,n891,n892);
xor (n891,n888,n889);
or (n892,n893,n896);
and (n893,n894,n895);
xor (n894,n864,n865);
and (n895,n141,n115);
and (n896,n897,n898);
xor (n897,n894,n895);
or (n898,n899,n902);
and (n899,n900,n901);
xor (n900,n870,n871);
and (n901,n104,n115);
and (n902,n903,n904);
xor (n903,n900,n901);
or (n904,n905,n908);
and (n905,n906,n907);
xor (n906,n876,n877);
and (n907,n31,n115);
and (n908,n909,n910);
xor (n909,n906,n907);
and (n910,n911,n511);
xor (n911,n882,n883);
and (n912,n131,n121);
or (n913,n914,n917);
and (n914,n915,n916);
xor (n915,n891,n892);
and (n916,n141,n121);
and (n917,n918,n919);
xor (n918,n915,n916);
or (n919,n920,n923);
and (n920,n921,n922);
xor (n921,n897,n898);
and (n922,n104,n121);
and (n923,n924,n925);
xor (n924,n921,n922);
or (n925,n926,n929);
and (n926,n927,n928);
xor (n927,n903,n904);
and (n928,n31,n121);
and (n929,n930,n931);
xor (n930,n927,n928);
and (n931,n932,n390);
xor (n932,n909,n910);
and (n933,n141,n95);
or (n934,n935,n938);
and (n935,n936,n937);
xor (n936,n918,n919);
and (n937,n104,n95);
and (n938,n939,n940);
xor (n939,n936,n937);
or (n940,n941,n944);
and (n941,n942,n943);
xor (n942,n924,n925);
and (n943,n31,n95);
and (n944,n945,n946);
xor (n945,n942,n943);
and (n946,n947,n948);
xor (n947,n930,n931);
and (n948,n207,n95);
and (n949,n104,n86);
or (n950,n951,n954);
and (n951,n952,n953);
xor (n952,n939,n940);
and (n953,n31,n86);
and (n954,n955,n956);
xor (n955,n952,n953);
and (n956,n957,n219);
xor (n957,n945,n946);
and (n958,n31,n17);
and (n959,n960,n212);
xor (n960,n955,n956);
and (n961,n207,n331);
endmodule
