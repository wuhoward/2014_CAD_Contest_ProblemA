module top (out,n4,n5,n6,n23,n24,n26,n31,n36,n37
        ,n42,n48,n65,n69,n73,n81,n89,n91,n97,n103
        ,n109,n120,n122,n129,n139,n148,n158,n165,n171,n195
        ,n208,n226);
output out;
input n4;
input n5;
input n6;
input n23;
input n24;
input n26;
input n31;
input n36;
input n37;
input n42;
input n48;
input n65;
input n69;
input n73;
input n81;
input n89;
input n91;
input n97;
input n103;
input n109;
input n120;
input n122;
input n129;
input n139;
input n148;
input n158;
input n165;
input n171;
input n195;
input n208;
input n226;
wire n0;
wire n1;
wire n2;
wire n3;
wire n7;
wire n8;
wire n9;
wire n10;
wire n11;
wire n12;
wire n13;
wire n14;
wire n15;
wire n16;
wire n17;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n25;
wire n27;
wire n28;
wire n29;
wire n30;
wire n32;
wire n33;
wire n34;
wire n35;
wire n38;
wire n39;
wire n40;
wire n41;
wire n43;
wire n44;
wire n45;
wire n46;
wire n47;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n63;
wire n64;
wire n66;
wire n67;
wire n68;
wire n70;
wire n71;
wire n72;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n90;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n121;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n172;
wire n173;
wire n174;
wire n175;
wire n176;
wire n177;
wire n178;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n185;
wire n186;
wire n187;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n194;
wire n196;
wire n197;
wire n198;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n219;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
wire n548;
wire n549;
wire n550;
wire n551;
wire n552;
wire n553;
wire n554;
wire n555;
wire n556;
wire n557;
wire n558;
wire n559;
wire n560;
wire n561;
wire n562;
wire n563;
wire n564;
wire n565;
wire n566;
wire n567;
wire n568;
wire n569;
wire n570;
wire n571;
wire n572;
wire n573;
wire n574;
wire n575;
wire n576;
wire n577;
wire n578;
wire n579;
wire n580;
wire n581;
wire n582;
wire n583;
wire n584;
wire n585;
wire n586;
wire n587;
wire n588;
wire n589;
wire n590;
wire n591;
wire n592;
wire n593;
wire n594;
wire n595;
wire n596;
wire n597;
wire n598;
wire n599;
wire n600;
wire n601;
wire n602;
wire n603;
wire n604;
wire n605;
wire n606;
wire n607;
wire n608;
wire n609;
wire n610;
wire n611;
wire n612;
wire n613;
wire n614;
wire n615;
wire n616;
wire n617;
wire n618;
wire n619;
wire n620;
wire n621;
wire n622;
wire n623;
wire n624;
wire n625;
wire n626;
wire n627;
wire n628;
wire n629;
wire n630;
wire n631;
wire n632;
wire n633;
wire n634;
wire n635;
wire n636;
wire n637;
wire n638;
wire n639;
wire n640;
wire n641;
wire n642;
wire n643;
wire n644;
wire n645;
wire n646;
wire n647;
wire n648;
wire n649;
wire n650;
wire n651;
wire n652;
wire n653;
wire n654;
wire n655;
wire n656;
wire n657;
wire n658;
wire n659;
wire n660;
wire n661;
wire n662;
wire n663;
wire n664;
wire n665;
wire n666;
wire n667;
wire n668;
wire n669;
wire n670;
wire n671;
wire n672;
wire n673;
wire n674;
wire n675;
wire n676;
wire n677;
wire n678;
wire n679;
wire n680;
wire n681;
wire n682;
wire n683;
wire n684;
wire n685;
wire n686;
wire n687;
wire n688;
wire n689;
wire n690;
wire n691;
wire n692;
wire n693;
wire n694;
wire n695;
wire n696;
wire n697;
wire n698;
wire n699;
wire n700;
wire n701;
wire n702;
wire n703;
wire n704;
wire n705;
wire n706;
wire n707;
wire n708;
wire n709;
wire n710;
wire n711;
wire n712;
wire n713;
wire n714;
wire n715;
wire n716;
wire n717;
wire n718;
wire n719;
wire n720;
wire n721;
wire n722;
wire n723;
wire n724;
wire n725;
wire n726;
wire n727;
wire n728;
wire n729;
wire n730;
wire n731;
wire n732;
wire n733;
wire n734;
wire n735;
wire n736;
wire n737;
wire n738;
wire n739;
wire n740;
wire n741;
wire n742;
wire n743;
wire n744;
wire n745;
wire n746;
wire n747;
wire n748;
wire n749;
wire n750;
wire n751;
wire n752;
wire n753;
wire n754;
wire n755;
wire n756;
wire n757;
wire n758;
wire n759;
wire n760;
wire n761;
wire n762;
wire n763;
wire n764;
wire n765;
wire n766;
wire n767;
wire n768;
wire n769;
wire n770;
wire n771;
wire n772;
wire n773;
wire n774;
wire n775;
wire n776;
wire n777;
wire n778;
wire n779;
wire n780;
wire n781;
wire n782;
wire n783;
wire n784;
wire n785;
wire n786;
wire n787;
wire n788;
wire n789;
wire n790;
wire n791;
wire n792;
wire n793;
wire n794;
wire n795;
wire n796;
wire n797;
wire n798;
wire n799;
wire n800;
wire n801;
wire n802;
wire n803;
wire n804;
wire n805;
wire n806;
wire n807;
wire n808;
wire n809;
wire n810;
wire n811;
wire n812;
wire n813;
wire n814;
wire n815;
wire n816;
wire n817;
wire n818;
wire n819;
wire n820;
wire n821;
wire n822;
wire n823;
wire n824;
wire n825;
wire n826;
wire n827;
wire n828;
wire n829;
wire n830;
wire n831;
wire n832;
wire n833;
wire n834;
wire n835;
wire n836;
wire n837;
wire n838;
wire n839;
wire n840;
wire n841;
wire n842;
wire n843;
wire n844;
wire n845;
wire n846;
wire n847;
wire n848;
wire n849;
wire n850;
wire n851;
wire n852;
wire n853;
wire n854;
wire n855;
wire n856;
wire n857;
wire n858;
wire n859;
wire n860;
wire n861;
wire n862;
wire n863;
wire n864;
wire n865;
wire n866;
wire n867;
wire n868;
wire n869;
wire n870;
wire n871;
wire n872;
wire n873;
wire n874;
wire n875;
wire n876;
wire n877;
wire n878;
wire n879;
wire n880;
wire n881;
wire n882;
wire n883;
wire n884;
wire n885;
wire n886;
wire n887;
wire n888;
wire n889;
wire n890;
wire n891;
wire n892;
wire n893;
wire n894;
wire n895;
wire n896;
wire n897;
wire n898;
wire n899;
wire n900;
wire n901;
wire n902;
wire n903;
wire n904;
wire n905;
wire n906;
wire n907;
wire n908;
wire n909;
wire n910;
wire n911;
wire n912;
wire n913;
wire n914;
wire n915;
wire n916;
wire n917;
wire n918;
wire n919;
wire n920;
wire n921;
wire n922;
wire n923;
wire n924;
wire n925;
wire n926;
wire n927;
wire n928;
wire n929;
wire n930;
wire n931;
wire n932;
wire n933;
wire n934;
wire n935;
wire n936;
wire n937;
wire n938;
wire n939;
wire n940;
wire n941;
wire n942;
wire n943;
wire n944;
wire n945;
wire n946;
wire n947;
wire n948;
wire n949;
wire n950;
wire n951;
wire n952;
wire n953;
wire n954;
wire n955;
wire n956;
wire n957;
wire n958;
wire n959;
wire n960;
wire n961;
wire n962;
wire n963;
wire n964;
wire n965;
wire n966;
wire n967;
wire n968;
wire n969;
wire n970;
wire n971;
wire n972;
wire n973;
wire n974;
wire n975;
wire n976;
wire n977;
wire n978;
wire n979;
wire n980;
wire n981;
wire n982;
wire n983;
wire n984;
wire n985;
wire n986;
wire n987;
wire n988;
wire n989;
wire n990;
wire n991;
wire n992;
wire n993;
wire n994;
wire n995;
wire n996;
wire n997;
wire n998;
wire n999;
wire n1000;
wire n1001;
wire n1002;
wire n1003;
wire n1004;
wire n1005;
wire n1006;
wire n1007;
wire n1008;
wire n1009;
wire n1010;
wire n1011;
wire n1012;
wire n1013;
wire n1014;
wire n1015;
wire n1016;
wire n1017;
wire n1018;
wire n1019;
wire n1020;
wire n1021;
wire n1022;
wire n1023;
wire n1024;
wire n1025;
wire n1026;
wire n1027;
wire n1028;
wire n1029;
wire n1030;
wire n1031;
wire n1032;
wire n1033;
wire n1034;
wire n1035;
wire n1036;
wire n1037;
wire n1038;
wire n1039;
wire n1040;
wire n1041;
wire n1042;
wire n1043;
wire n1044;
wire n1045;
wire n1046;
wire n1047;
wire n1048;
wire n1049;
wire n1050;
wire n1051;
wire n1052;
wire n1053;
wire n1054;
wire n1055;
wire n1056;
wire n1057;
wire n1058;
wire n1059;
wire n1060;
wire n1061;
wire n1062;
wire n1063;
wire n1064;
wire n1065;
wire n1066;
wire n1067;
wire n1068;
wire n1069;
wire n1070;
wire n1071;
wire n1072;
wire n1073;
wire n1074;
wire n1075;
wire n1076;
wire n1077;
wire n1078;
wire n1079;
wire n1080;
wire n1081;
wire n1082;
wire n1083;
wire n1084;
wire n1085;
wire n1086;
wire n1087;
wire n1088;
wire n1089;
wire n1090;
wire n1091;
wire n1092;
wire n1093;
wire n1094;
wire n1095;
wire n1096;
wire n1097;
wire n1098;
wire n1099;
wire n1100;
wire n1101;
wire n1102;
wire n1103;
wire n1104;
wire n1105;
wire n1106;
wire n1107;
wire n1108;
wire n1109;
wire n1110;
wire n1111;
wire n1112;
wire n1113;
wire n1114;
wire n1115;
wire n1116;
wire n1117;
wire n1118;
wire n1119;
wire n1120;
wire n1121;
wire n1122;
wire n1123;
wire n1124;
wire n1125;
wire n1126;
wire n1127;
wire n1128;
wire n1129;
wire n1130;
wire n1131;
wire n1132;
wire n1133;
wire n1134;
wire n1135;
wire n1136;
wire n1137;
wire n1138;
wire n1139;
wire n1140;
wire n1141;
wire n1142;
wire n1143;
wire n1144;
wire n1145;
wire n1146;
wire n1147;
wire n1148;
wire n1149;
wire n1150;
wire n1151;
wire n1152;
wire n1153;
wire n1154;
wire n1155;
wire n1156;
wire n1157;
wire n1158;
wire n1159;
wire n1160;
wire n1161;
wire n1162;
wire n1163;
wire n1164;
wire n1165;
wire n1166;
wire n1167;
wire n1168;
wire n1169;
wire n1170;
wire n1171;
wire n1172;
wire n1173;
wire n1174;
wire n1175;
wire n1176;
wire n1177;
wire n1178;
wire n1179;
wire n1180;
xor (out,n0,n722);
not (n0,n1);
nor (n1,n2,n7);
and (n2,n3,n6);
nor (n3,n4,n5);
and (n7,n8,n719);
nand (n8,n9,n718);
or (n9,n10,n371);
not (n10,n11);
nand (n11,n12,n370);
not (n12,n13);
nor (n13,n14,n318);
xor (n14,n15,n232);
xor (n15,n16,n175);
xor (n16,n17,n112);
xor (n17,n18,n51);
xor (n18,n19,n32);
nor (n19,n20,n30);
nor (n20,n21,n27);
and (n21,n22,n25);
nand (n22,n23,n24);
not (n25,n26);
and (n27,n28,n29);
not (n28,n23);
not (n29,n24);
not (n30,n31);
nand (n32,n33,n45);
or (n33,n34,n38);
nand (n34,n35,n37);
not (n35,n36);
not (n38,n39);
nor (n39,n40,n44);
and (n40,n41,n43);
not (n41,n42);
not (n43,n37);
and (n44,n42,n37);
or (n45,n35,n46);
nor (n46,n47,n49);
and (n47,n43,n48);
and (n49,n37,n50);
not (n50,n48);
or (n51,n52,n111);
and (n52,n53,n84);
xor (n53,n54,n58);
nor (n54,n55,n28);
nor (n55,n56,n57);
and (n56,n29,n26);
and (n57,n24,n25);
nand (n58,n59,n77);
or (n59,n60,n71);
nand (n60,n61,n67);
not (n61,n62);
nand (n62,n63,n66);
or (n63,n64,n37);
not (n64,n65);
nand (n66,n64,n37);
nand (n67,n68,n70);
or (n68,n69,n64);
nand (n70,n64,n69);
nor (n71,n72,n75);
and (n72,n73,n74);
not (n74,n69);
and (n75,n76,n69);
not (n76,n73);
nand (n77,n78,n62);
not (n78,n79);
nor (n79,n80,n82);
and (n80,n81,n74);
and (n82,n83,n69);
not (n83,n81);
nand (n84,n85,n105);
or (n85,n86,n99);
nand (n86,n87,n93);
nand (n87,n88,n92);
or (n88,n89,n90);
not (n90,n91);
nand (n92,n90,n89);
not (n93,n94);
nand (n94,n95,n98);
or (n95,n96,n89);
not (n96,n97);
nand (n98,n89,n96);
not (n99,n100);
nor (n100,n101,n104);
and (n101,n102,n90);
not (n102,n103);
and (n104,n103,n91);
or (n105,n93,n106);
nor (n106,n107,n110);
and (n107,n108,n91);
not (n108,n109);
and (n110,n109,n90);
and (n111,n54,n58);
or (n112,n113,n174);
and (n113,n114,n151);
xor (n114,n115,n142);
nand (n115,n116,n135);
or (n116,n117,n125);
not (n117,n118);
nand (n118,n119,n123);
or (n119,n120,n121);
not (n121,n122);
or (n123,n122,n124);
not (n124,n120);
not (n125,n126);
nor (n126,n127,n132);
nor (n127,n128,n130);
and (n128,n129,n124);
and (n130,n120,n131);
not (n131,n129);
nand (n132,n133,n134);
or (n133,n90,n129);
nand (n134,n129,n90);
nand (n135,n136,n132);
not (n136,n137);
nor (n137,n138,n140);
and (n138,n124,n139);
and (n140,n141,n120);
not (n141,n139);
nand (n142,n143,n150);
or (n143,n34,n144);
not (n144,n145);
nor (n145,n146,n149);
and (n146,n147,n43);
not (n147,n148);
and (n149,n148,n37);
nand (n150,n39,n36);
nand (n151,n152,n168);
or (n152,n153,n163);
nand (n153,n154,n160);
not (n154,n155);
nand (n155,n156,n159);
or (n156,n157,n120);
not (n157,n158);
nand (n159,n120,n157);
nand (n160,n161,n162);
nand (n161,n157,n26);
nand (n162,n158,n25);
nor (n163,n164,n166);
and (n164,n25,n165);
and (n166,n26,n167);
not (n167,n165);
or (n168,n154,n169);
nor (n169,n170,n172);
and (n170,n25,n171);
and (n172,n26,n173);
not (n173,n171);
and (n174,n115,n142);
or (n175,n176,n231);
and (n176,n177,n180);
xor (n177,n178,n179);
xor (n178,n114,n151);
xor (n179,n53,n84);
or (n180,n181,n230);
and (n181,n182,n211);
xor (n182,n183,n189);
nand (n183,n184,n188);
or (n184,n153,n185);
nor (n185,n186,n187);
and (n186,n28,n26);
and (n187,n23,n25);
or (n188,n154,n163);
nand (n189,n190,n204);
or (n190,n191,n201);
not (n191,n192);
nor (n192,n193,n197);
nand (n193,n194,n196);
or (n194,n74,n195);
nand (n196,n195,n74);
nor (n197,n198,n200);
and (n198,n199,n97);
not (n199,n195);
and (n200,n195,n96);
nor (n201,n202,n203);
and (n202,n96,n109);
and (n203,n97,n108);
or (n204,n205,n206);
not (n205,n193);
nor (n206,n207,n209);
and (n207,n96,n208);
and (n209,n97,n210);
not (n210,n208);
nand (n211,n212,n229);
or (n212,n213,n220);
not (n213,n214);
nand (n214,n215,n26);
nand (n215,n216,n217);
or (n216,n23,n158);
nand (n217,n218,n124);
not (n218,n219);
and (n219,n23,n158);
not (n220,n221);
nand (n221,n222,n223);
or (n222,n71,n61);
or (n223,n60,n224);
nor (n224,n225,n227);
and (n225,n226,n74);
and (n227,n228,n69);
not (n228,n226);
or (n229,n221,n214);
and (n230,n183,n189);
and (n231,n178,n179);
xor (n232,n233,n286);
xor (n233,n234,n263);
xor (n234,n235,n252);
xor (n235,n236,n246);
nand (n236,n237,n241);
or (n237,n238,n191);
nor (n238,n239,n240);
and (n239,n96,n226);
and (n240,n97,n228);
nand (n241,n242,n193);
not (n242,n243);
nor (n243,n244,n245);
and (n244,n96,n73);
and (n245,n97,n76);
nand (n246,n247,n248);
or (n247,n153,n169);
or (n248,n154,n249);
nor (n249,n250,n251);
and (n250,n25,n122);
and (n251,n26,n121);
nand (n252,n253,n259);
or (n253,n254,n256);
nand (n254,n55,n255);
xor (n255,n29,n30);
nor (n256,n257,n258);
and (n257,n28,n31);
and (n258,n23,n30);
or (n259,n260,n55);
nor (n260,n261,n262);
and (n261,n30,n165);
and (n262,n31,n167);
xor (n263,n264,n279);
xor (n264,n265,n272);
nand (n265,n266,n267);
or (n266,n60,n79);
nand (n267,n268,n62);
not (n268,n269);
nor (n269,n270,n271);
and (n270,n148,n74);
and (n271,n147,n69);
nand (n272,n273,n278);
or (n273,n274,n93);
not (n274,n275);
nor (n275,n276,n277);
and (n276,n208,n91);
and (n277,n210,n90);
or (n278,n86,n106);
nand (n279,n280,n281);
or (n280,n125,n137);
or (n281,n282,n283);
not (n282,n132);
nor (n283,n284,n285);
and (n284,n124,n103);
and (n285,n120,n102);
or (n286,n287,n317);
and (n287,n288,n293);
xor (n288,n289,n292);
nand (n289,n290,n291);
or (n290,n191,n206);
or (n291,n205,n238);
and (n292,n221,n213);
or (n293,n294,n316);
and (n294,n295,n310);
xor (n295,n296,n303);
nand (n296,n297,n302);
or (n297,n298,n86);
not (n298,n299);
nand (n299,n300,n301);
or (n300,n91,n141);
or (n301,n90,n139);
nand (n302,n94,n100);
nand (n303,n304,n309);
or (n304,n305,n125);
not (n305,n306);
nand (n306,n307,n308);
or (n307,n120,n173);
or (n308,n124,n171);
nand (n309,n132,n118);
nand (n310,n311,n312);
or (n311,n35,n144);
or (n312,n313,n34);
nor (n313,n314,n315);
and (n314,n43,n81);
and (n315,n37,n83);
and (n316,n296,n303);
and (n317,n289,n292);
or (n318,n319,n369);
and (n319,n320,n368);
xor (n320,n321,n322);
xor (n321,n288,n293);
or (n322,n323,n367);
and (n323,n324,n366);
xor (n324,n325,n343);
or (n325,n326,n342);
and (n326,n327,n336);
xor (n327,n328,n329);
nor (n328,n154,n28);
nand (n329,n330,n334);
or (n330,n331,n60);
nor (n331,n332,n333);
and (n332,n74,n208);
and (n333,n69,n210);
nand (n334,n335,n62);
not (n335,n224);
nand (n336,n337,n338);
or (n337,n298,n93);
or (n338,n86,n339);
nor (n339,n340,n341);
and (n340,n90,n122);
and (n341,n91,n121);
and (n342,n328,n329);
or (n343,n344,n365);
and (n344,n345,n359);
xor (n345,n346,n353);
nand (n346,n347,n352);
or (n347,n348,n125);
not (n348,n349);
nand (n349,n350,n351);
or (n350,n120,n167);
or (n351,n124,n165);
nand (n352,n132,n306);
nand (n353,n354,n358);
or (n354,n355,n34);
nor (n355,n356,n357);
and (n356,n43,n73);
and (n357,n37,n76);
or (n358,n313,n35);
nand (n359,n360,n364);
or (n360,n191,n361);
nor (n361,n362,n363);
and (n362,n96,n103);
and (n363,n97,n102);
or (n364,n205,n201);
and (n365,n346,n353);
xor (n366,n295,n310);
and (n367,n325,n343);
xor (n368,n177,n180);
and (n369,n321,n322);
nand (n370,n14,n318);
not (n371,n372);
nand (n372,n373,n717);
or (n373,n374,n711);
not (n374,n375);
nand (n375,n376,n710);
or (n376,n377,n459);
not (n377,n378);
or (n378,n379,n425);
xor (n379,n380,n383);
xor (n380,n381,n382);
xor (n381,n182,n211);
xor (n382,n324,n366);
or (n383,n384,n424);
and (n384,n385,n423);
xor (n385,n386,n399);
and (n386,n387,n393);
and (n387,n388,n120);
nand (n388,n389,n390);
or (n389,n23,n129);
nand (n390,n391,n90);
not (n391,n392);
and (n392,n23,n129);
nand (n393,n394,n398);
or (n394,n60,n395);
nor (n395,n396,n397);
and (n396,n74,n109);
and (n397,n69,n108);
or (n398,n61,n331);
or (n399,n400,n422);
and (n400,n401,n416);
xor (n401,n402,n409);
nand (n402,n403,n407);
or (n403,n404,n86);
nor (n404,n405,n406);
and (n405,n90,n171);
and (n406,n91,n173);
nand (n407,n408,n94);
not (n408,n339);
nand (n409,n410,n411);
or (n410,n348,n282);
nand (n411,n412,n126);
not (n412,n413);
nor (n413,n414,n415);
and (n414,n28,n120);
and (n415,n124,n23);
nand (n416,n417,n421);
or (n417,n34,n418);
nor (n418,n419,n420);
and (n419,n43,n226);
and (n420,n37,n228);
or (n421,n355,n35);
and (n422,n402,n409);
xor (n423,n327,n336);
and (n424,n386,n399);
or (n425,n426,n458);
and (n426,n427,n457);
xor (n427,n428,n429);
xor (n428,n345,n359);
or (n429,n430,n456);
and (n430,n431,n439);
xor (n431,n432,n438);
nand (n432,n433,n437);
or (n433,n191,n434);
nor (n434,n435,n436);
and (n435,n96,n139);
and (n436,n97,n141);
or (n437,n205,n361);
xor (n438,n387,n393);
or (n439,n440,n455);
and (n440,n441,n449);
xor (n441,n442,n443);
nor (n442,n282,n28);
nand (n443,n444,n448);
or (n444,n445,n34);
nor (n445,n446,n447);
and (n446,n210,n37);
and (n447,n208,n43);
or (n448,n418,n35);
nand (n449,n450,n454);
or (n450,n86,n451);
nor (n451,n452,n453);
and (n452,n90,n165);
and (n453,n91,n167);
or (n454,n93,n404);
and (n455,n442,n443);
and (n456,n432,n438);
xor (n457,n385,n423);
and (n458,n428,n429);
not (n459,n460);
or (n460,n461,n709);
and (n461,n462,n502);
xor (n462,n463,n501);
or (n463,n464,n500);
and (n464,n465,n499);
xor (n465,n466,n467);
xor (n466,n401,n416);
or (n467,n468,n498);
and (n468,n469,n484);
xor (n469,n470,n478);
nand (n470,n471,n476);
or (n471,n472,n60);
not (n472,n473);
nand (n473,n474,n475);
or (n474,n69,n102);
or (n475,n74,n103);
nand (n476,n477,n62);
not (n477,n395);
nand (n478,n479,n483);
or (n479,n191,n480);
nor (n480,n481,n482);
and (n481,n96,n122);
and (n482,n97,n121);
or (n483,n205,n434);
and (n484,n485,n491);
nor (n485,n486,n90);
nor (n486,n487,n489);
and (n487,n28,n488);
not (n488,n89);
nor (n489,n490,n97);
and (n490,n23,n89);
nand (n491,n492,n497);
or (n492,n34,n493);
not (n493,n494);
nor (n494,n495,n496);
and (n495,n108,n43);
and (n496,n109,n37);
or (n497,n445,n35);
and (n498,n470,n478);
xor (n499,n431,n439);
and (n500,n466,n467);
xor (n501,n427,n457);
nand (n502,n503,n706,n708);
nand (n503,n504,n539,n699);
nand (n504,n505,n507);
not (n505,n506);
xor (n506,n465,n499);
not (n507,n508);
or (n508,n509,n538);
and (n509,n510,n537);
xor (n510,n511,n536);
or (n511,n512,n535);
and (n512,n513,n529);
xor (n513,n514,n522);
nand (n514,n515,n520);
or (n515,n516,n86);
not (n516,n517);
nand (n517,n518,n519);
or (n518,n90,n23);
or (n519,n28,n91);
nand (n520,n521,n94);
not (n521,n451);
nand (n522,n523,n528);
or (n523,n524,n60);
not (n524,n525);
nand (n525,n526,n527);
or (n526,n69,n141);
or (n527,n74,n139);
nand (n528,n62,n473);
nand (n529,n530,n534);
or (n530,n191,n531);
nor (n531,n532,n533);
and (n532,n96,n171);
and (n533,n97,n173);
or (n534,n205,n480);
and (n535,n514,n522);
xor (n536,n441,n449);
xor (n537,n469,n484);
and (n538,n511,n536);
nand (n539,n540,n698);
or (n540,n541,n591);
not (n541,n542);
nand (n542,n543,n567);
not (n543,n544);
xor (n544,n545,n566);
xor (n545,n546,n547);
xor (n546,n485,n491);
or (n547,n548,n565);
and (n548,n549,n558);
xor (n549,n550,n551);
and (n550,n94,n23);
nand (n551,n552,n557);
or (n552,n34,n553);
not (n553,n554);
nor (n554,n555,n556);
and (n555,n102,n43);
and (n556,n103,n37);
nand (n557,n494,n36);
nand (n558,n559,n564);
or (n559,n560,n60);
not (n560,n561);
nor (n561,n562,n563);
and (n562,n121,n74);
and (n563,n122,n69);
nand (n564,n62,n525);
and (n565,n550,n551);
xor (n566,n513,n529);
not (n567,n568);
or (n568,n569,n590);
and (n569,n570,n589);
xor (n570,n571,n577);
nand (n571,n572,n576);
or (n572,n191,n573);
nor (n573,n574,n575);
and (n574,n167,n97);
and (n575,n165,n96);
or (n576,n205,n531);
and (n577,n578,n583);
and (n578,n579,n97);
nand (n579,n580,n582);
or (n580,n581,n69);
and (n581,n23,n195);
or (n582,n23,n195);
nand (n583,n584,n585);
or (n584,n35,n553);
or (n585,n586,n34);
nor (n586,n587,n588);
and (n587,n43,n139);
and (n588,n37,n141);
xor (n589,n549,n558);
and (n590,n571,n577);
not (n591,n592);
nand (n592,n593,n697);
or (n593,n594,n617);
not (n594,n595);
nand (n595,n596,n598);
not (n596,n597);
xor (n597,n570,n589);
not (n598,n599);
or (n599,n600,n616);
and (n600,n601,n615);
xor (n601,n602,n609);
nand (n602,n603,n608);
or (n603,n604,n60);
not (n604,n605);
nor (n605,n606,n607);
and (n606,n173,n74);
and (n607,n171,n69);
nand (n608,n561,n62);
nand (n609,n610,n611);
or (n610,n205,n573);
nand (n611,n192,n612);
nand (n612,n613,n614);
or (n613,n23,n96);
or (n614,n28,n97);
xor (n615,n578,n583);
and (n616,n602,n609);
not (n617,n618);
or (n618,n619,n696);
and (n619,n620,n641);
xor (n620,n621,n640);
or (n621,n622,n639);
and (n622,n623,n632);
xor (n623,n624,n625);
and (n624,n193,n23);
nand (n625,n626,n631);
or (n626,n627,n60);
not (n627,n628);
nor (n628,n629,n630);
and (n629,n167,n74);
and (n630,n165,n69);
nand (n631,n605,n62);
nand (n632,n633,n638);
or (n633,n34,n634);
not (n634,n635);
nor (n635,n636,n637);
and (n636,n121,n43);
and (n637,n122,n37);
or (n638,n586,n35);
and (n639,n624,n625);
xor (n640,n601,n615);
nand (n641,n642,n695);
or (n642,n643,n659);
nor (n643,n644,n645);
xor (n644,n623,n632);
nor (n645,n646,n654);
not (n646,n647);
nand (n647,n648,n649);
or (n648,n35,n634);
nand (n649,n650,n653);
nand (n650,n651,n652);
or (n651,n171,n43);
nand (n652,n43,n171);
not (n653,n34);
nand (n654,n655,n69);
nand (n655,n656,n658);
or (n656,n657,n37);
and (n657,n23,n65);
or (n658,n23,n65);
nor (n659,n660,n694);
and (n660,n661,n673);
nand (n661,n662,n669);
not (n662,n663);
nand (n663,n664,n668);
or (n664,n60,n665);
nor (n665,n666,n667);
and (n666,n69,n28);
and (n667,n23,n74);
or (n668,n61,n627);
nor (n669,n670,n671);
and (n670,n654,n647);
and (n671,n672,n646);
not (n672,n654);
or (n673,n674,n693);
and (n674,n675,n684);
xor (n675,n676,n677);
nor (n676,n61,n28);
nand (n677,n678,n683);
or (n678,n34,n679);
not (n679,n680);
nand (n680,n681,n682);
or (n681,n167,n37);
nand (n682,n37,n167);
nand (n683,n650,n36);
nor (n684,n685,n691);
nor (n685,n686,n687);
and (n686,n680,n36);
nor (n687,n688,n34);
nor (n688,n689,n690);
and (n689,n28,n37);
and (n690,n23,n43);
or (n691,n692,n43);
and (n692,n23,n36);
and (n693,n676,n677);
nor (n694,n662,n669);
nand (n695,n644,n645);
and (n696,n621,n640);
nand (n697,n597,n599);
nand (n698,n544,n568);
nand (n699,n700,n704);
not (n700,n701);
or (n701,n702,n703);
and (n702,n545,n566);
and (n703,n546,n547);
not (n704,n705);
xor (n705,n510,n537);
nand (n706,n504,n707);
and (n707,n705,n701);
nand (n708,n508,n506);
and (n709,n463,n501);
nand (n710,n379,n425);
not (n711,n712);
or (n712,n713,n716);
or (n713,n714,n715);
and (n714,n380,n383);
and (n715,n381,n382);
xor (n716,n320,n368);
nand (n717,n713,n716);
or (n718,n372,n11);
not (n719,n720);
nand (n720,n721,n4);
not (n721,n5);
wire s0n722,s1n722,notn722;
or (n722,s0n722,s1n722);
not(notn722,n5);
and (s0n722,notn722,n723);
and (s1n722,n5,1'b0);
wire s0n723,s1n723,notn723;
or (n723,s0n723,s1n723);
not(notn723,n4);
and (s0n723,notn723,n6);
and (s1n723,n4,n724);
xor (n724,n725,n1180);
xor (n725,n726,n1177);
xor (n726,n727,n1176);
xor (n727,n728,n1167);
xor (n728,n729,n1166);
xor (n729,n730,n1152);
xor (n730,n731,n1151);
xor (n731,n732,n1130);
xor (n732,n733,n1129);
xor (n733,n734,n1103);
xor (n734,n735,n1102);
xor (n735,n736,n1070);
xor (n736,n737,n1069);
xor (n737,n738,n1031);
xor (n738,n739,n1030);
xor (n739,n740,n985);
xor (n740,n741,n984);
xor (n741,n742,n934);
xor (n742,n743,n933);
xor (n743,n744,n879);
xor (n744,n745,n878);
xor (n745,n746,n816);
xor (n746,n747,n815);
xor (n747,n748,n750);
xor (n748,n749,n44);
and (n749,n48,n36);
or (n750,n751,n753);
and (n751,n752,n149);
and (n752,n42,n36);
and (n753,n754,n755);
xor (n754,n752,n149);
or (n755,n756,n759);
and (n756,n757,n758);
and (n757,n148,n36);
and (n758,n81,n37);
and (n759,n760,n761);
xor (n760,n757,n758);
or (n761,n762,n765);
and (n762,n763,n764);
and (n763,n81,n36);
and (n764,n73,n37);
and (n765,n766,n767);
xor (n766,n763,n764);
or (n767,n768,n771);
and (n768,n769,n770);
and (n769,n73,n36);
and (n770,n226,n37);
and (n771,n772,n773);
xor (n772,n769,n770);
or (n773,n774,n777);
and (n774,n775,n776);
and (n775,n226,n36);
and (n776,n208,n37);
and (n777,n778,n779);
xor (n778,n775,n776);
or (n779,n780,n782);
and (n780,n781,n496);
and (n781,n208,n36);
and (n782,n783,n784);
xor (n783,n781,n496);
or (n784,n785,n787);
and (n785,n786,n556);
and (n786,n109,n36);
and (n787,n788,n789);
xor (n788,n786,n556);
or (n789,n790,n793);
and (n790,n791,n792);
and (n791,n103,n36);
and (n792,n139,n37);
and (n793,n794,n795);
xor (n794,n791,n792);
or (n795,n796,n798);
and (n796,n797,n637);
and (n797,n139,n36);
and (n798,n799,n800);
xor (n799,n797,n637);
or (n800,n801,n804);
and (n801,n802,n803);
and (n802,n122,n36);
and (n803,n171,n37);
and (n804,n805,n806);
xor (n805,n802,n803);
or (n806,n807,n810);
and (n807,n808,n809);
and (n808,n171,n36);
and (n809,n165,n37);
and (n810,n811,n812);
xor (n811,n808,n809);
and (n812,n813,n814);
and (n813,n165,n36);
and (n814,n23,n37);
and (n815,n148,n65);
or (n816,n817,n820);
and (n817,n818,n819);
xor (n818,n754,n755);
and (n819,n81,n65);
and (n820,n821,n822);
xor (n821,n818,n819);
or (n822,n823,n826);
and (n823,n824,n825);
xor (n824,n760,n761);
and (n825,n73,n65);
and (n826,n827,n828);
xor (n827,n824,n825);
or (n828,n829,n832);
and (n829,n830,n831);
xor (n830,n766,n767);
and (n831,n226,n65);
and (n832,n833,n834);
xor (n833,n830,n831);
or (n834,n835,n838);
and (n835,n836,n837);
xor (n836,n772,n773);
and (n837,n208,n65);
and (n838,n839,n840);
xor (n839,n836,n837);
or (n840,n841,n844);
and (n841,n842,n843);
xor (n842,n778,n779);
and (n843,n109,n65);
and (n844,n845,n846);
xor (n845,n842,n843);
or (n846,n847,n850);
and (n847,n848,n849);
xor (n848,n783,n784);
and (n849,n103,n65);
and (n850,n851,n852);
xor (n851,n848,n849);
or (n852,n853,n856);
and (n853,n854,n855);
xor (n854,n788,n789);
and (n855,n139,n65);
and (n856,n857,n858);
xor (n857,n854,n855);
or (n858,n859,n862);
and (n859,n860,n861);
xor (n860,n794,n795);
and (n861,n122,n65);
and (n862,n863,n864);
xor (n863,n860,n861);
or (n864,n865,n868);
and (n865,n866,n867);
xor (n866,n799,n800);
and (n867,n171,n65);
and (n868,n869,n870);
xor (n869,n866,n867);
or (n870,n871,n874);
and (n871,n872,n873);
xor (n872,n805,n806);
and (n873,n165,n65);
and (n874,n875,n876);
xor (n875,n872,n873);
and (n876,n877,n657);
xor (n877,n811,n812);
and (n878,n81,n69);
or (n879,n880,n883);
and (n880,n881,n882);
xor (n881,n821,n822);
and (n882,n73,n69);
and (n883,n884,n885);
xor (n884,n881,n882);
or (n885,n886,n889);
and (n886,n887,n888);
xor (n887,n827,n828);
and (n888,n226,n69);
and (n889,n890,n891);
xor (n890,n887,n888);
or (n891,n892,n895);
and (n892,n893,n894);
xor (n893,n833,n834);
and (n894,n208,n69);
and (n895,n896,n897);
xor (n896,n893,n894);
or (n897,n898,n901);
and (n898,n899,n900);
xor (n899,n839,n840);
and (n900,n109,n69);
and (n901,n902,n903);
xor (n902,n899,n900);
or (n903,n904,n907);
and (n904,n905,n906);
xor (n905,n845,n846);
and (n906,n103,n69);
and (n907,n908,n909);
xor (n908,n905,n906);
or (n909,n910,n913);
and (n910,n911,n912);
xor (n911,n851,n852);
and (n912,n139,n69);
and (n913,n914,n915);
xor (n914,n911,n912);
or (n915,n916,n918);
and (n916,n917,n563);
xor (n917,n857,n858);
and (n918,n919,n920);
xor (n919,n917,n563);
or (n920,n921,n923);
and (n921,n922,n607);
xor (n922,n863,n864);
and (n923,n924,n925);
xor (n924,n922,n607);
or (n925,n926,n928);
and (n926,n927,n630);
xor (n927,n869,n870);
and (n928,n929,n930);
xor (n929,n927,n630);
and (n930,n931,n932);
xor (n931,n875,n876);
and (n932,n23,n69);
and (n933,n73,n195);
or (n934,n935,n938);
and (n935,n936,n937);
xor (n936,n884,n885);
and (n937,n226,n195);
and (n938,n939,n940);
xor (n939,n936,n937);
or (n940,n941,n944);
and (n941,n942,n943);
xor (n942,n890,n891);
and (n943,n208,n195);
and (n944,n945,n946);
xor (n945,n942,n943);
or (n946,n947,n950);
and (n947,n948,n949);
xor (n948,n896,n897);
and (n949,n109,n195);
and (n950,n951,n952);
xor (n951,n948,n949);
or (n952,n953,n956);
and (n953,n954,n955);
xor (n954,n902,n903);
and (n955,n103,n195);
and (n956,n957,n958);
xor (n957,n954,n955);
or (n958,n959,n962);
and (n959,n960,n961);
xor (n960,n908,n909);
and (n961,n139,n195);
and (n962,n963,n964);
xor (n963,n960,n961);
or (n964,n965,n968);
and (n965,n966,n967);
xor (n966,n914,n915);
and (n967,n122,n195);
and (n968,n969,n970);
xor (n969,n966,n967);
or (n970,n971,n974);
and (n971,n972,n973);
xor (n972,n919,n920);
and (n973,n171,n195);
and (n974,n975,n976);
xor (n975,n972,n973);
or (n976,n977,n980);
and (n977,n978,n979);
xor (n978,n924,n925);
and (n979,n165,n195);
and (n980,n981,n982);
xor (n981,n978,n979);
and (n982,n983,n581);
xor (n983,n929,n930);
and (n984,n226,n97);
or (n985,n986,n989);
and (n986,n987,n988);
xor (n987,n939,n940);
and (n988,n208,n97);
and (n989,n990,n991);
xor (n990,n987,n988);
or (n991,n992,n995);
and (n992,n993,n994);
xor (n993,n945,n946);
and (n994,n109,n97);
and (n995,n996,n997);
xor (n996,n993,n994);
or (n997,n998,n1001);
and (n998,n999,n1000);
xor (n999,n951,n952);
and (n1000,n103,n97);
and (n1001,n1002,n1003);
xor (n1002,n999,n1000);
or (n1003,n1004,n1007);
and (n1004,n1005,n1006);
xor (n1005,n957,n958);
and (n1006,n139,n97);
and (n1007,n1008,n1009);
xor (n1008,n1005,n1006);
or (n1009,n1010,n1013);
and (n1010,n1011,n1012);
xor (n1011,n963,n964);
and (n1012,n122,n97);
and (n1013,n1014,n1015);
xor (n1014,n1011,n1012);
or (n1015,n1016,n1019);
and (n1016,n1017,n1018);
xor (n1017,n969,n970);
and (n1018,n171,n97);
and (n1019,n1020,n1021);
xor (n1020,n1017,n1018);
or (n1021,n1022,n1025);
and (n1022,n1023,n1024);
xor (n1023,n975,n976);
and (n1024,n165,n97);
and (n1025,n1026,n1027);
xor (n1026,n1023,n1024);
and (n1027,n1028,n1029);
xor (n1028,n981,n982);
and (n1029,n23,n97);
and (n1030,n208,n89);
or (n1031,n1032,n1035);
and (n1032,n1033,n1034);
xor (n1033,n990,n991);
and (n1034,n109,n89);
and (n1035,n1036,n1037);
xor (n1036,n1033,n1034);
or (n1037,n1038,n1041);
and (n1038,n1039,n1040);
xor (n1039,n996,n997);
and (n1040,n103,n89);
and (n1041,n1042,n1043);
xor (n1042,n1039,n1040);
or (n1043,n1044,n1047);
and (n1044,n1045,n1046);
xor (n1045,n1002,n1003);
and (n1046,n139,n89);
and (n1047,n1048,n1049);
xor (n1048,n1045,n1046);
or (n1049,n1050,n1053);
and (n1050,n1051,n1052);
xor (n1051,n1008,n1009);
and (n1052,n122,n89);
and (n1053,n1054,n1055);
xor (n1054,n1051,n1052);
or (n1055,n1056,n1059);
and (n1056,n1057,n1058);
xor (n1057,n1014,n1015);
and (n1058,n171,n89);
and (n1059,n1060,n1061);
xor (n1060,n1057,n1058);
or (n1061,n1062,n1065);
and (n1062,n1063,n1064);
xor (n1063,n1020,n1021);
and (n1064,n165,n89);
and (n1065,n1066,n1067);
xor (n1066,n1063,n1064);
and (n1067,n1068,n490);
xor (n1068,n1026,n1027);
and (n1069,n109,n91);
or (n1070,n1071,n1073);
and (n1071,n1072,n104);
xor (n1072,n1036,n1037);
and (n1073,n1074,n1075);
xor (n1074,n1072,n104);
or (n1075,n1076,n1079);
and (n1076,n1077,n1078);
xor (n1077,n1042,n1043);
and (n1078,n139,n91);
and (n1079,n1080,n1081);
xor (n1080,n1077,n1078);
or (n1081,n1082,n1085);
and (n1082,n1083,n1084);
xor (n1083,n1048,n1049);
and (n1084,n122,n91);
and (n1085,n1086,n1087);
xor (n1086,n1083,n1084);
or (n1087,n1088,n1091);
and (n1088,n1089,n1090);
xor (n1089,n1054,n1055);
and (n1090,n171,n91);
and (n1091,n1092,n1093);
xor (n1092,n1089,n1090);
or (n1093,n1094,n1097);
and (n1094,n1095,n1096);
xor (n1095,n1060,n1061);
and (n1096,n165,n91);
and (n1097,n1098,n1099);
xor (n1098,n1095,n1096);
and (n1099,n1100,n1101);
xor (n1100,n1066,n1067);
and (n1101,n23,n91);
and (n1102,n103,n129);
or (n1103,n1104,n1107);
and (n1104,n1105,n1106);
xor (n1105,n1074,n1075);
and (n1106,n139,n129);
and (n1107,n1108,n1109);
xor (n1108,n1105,n1106);
or (n1109,n1110,n1113);
and (n1110,n1111,n1112);
xor (n1111,n1080,n1081);
and (n1112,n122,n129);
and (n1113,n1114,n1115);
xor (n1114,n1111,n1112);
or (n1115,n1116,n1119);
and (n1116,n1117,n1118);
xor (n1117,n1086,n1087);
and (n1118,n171,n129);
and (n1119,n1120,n1121);
xor (n1120,n1117,n1118);
or (n1121,n1122,n1125);
and (n1122,n1123,n1124);
xor (n1123,n1092,n1093);
and (n1124,n165,n129);
and (n1125,n1126,n1127);
xor (n1126,n1123,n1124);
and (n1127,n1128,n392);
xor (n1128,n1098,n1099);
and (n1129,n139,n120);
or (n1130,n1131,n1134);
and (n1131,n1132,n1133);
xor (n1132,n1108,n1109);
and (n1133,n122,n120);
and (n1134,n1135,n1136);
xor (n1135,n1132,n1133);
or (n1136,n1137,n1140);
and (n1137,n1138,n1139);
xor (n1138,n1114,n1115);
and (n1139,n171,n120);
and (n1140,n1141,n1142);
xor (n1141,n1138,n1139);
or (n1142,n1143,n1146);
and (n1143,n1144,n1145);
xor (n1144,n1120,n1121);
and (n1145,n165,n120);
and (n1146,n1147,n1148);
xor (n1147,n1144,n1145);
and (n1148,n1149,n1150);
xor (n1149,n1126,n1127);
and (n1150,n23,n120);
and (n1151,n122,n158);
or (n1152,n1153,n1156);
and (n1153,n1154,n1155);
xor (n1154,n1135,n1136);
and (n1155,n171,n158);
and (n1156,n1157,n1158);
xor (n1157,n1154,n1155);
or (n1158,n1159,n1162);
and (n1159,n1160,n1161);
xor (n1160,n1141,n1142);
and (n1161,n165,n158);
and (n1162,n1163,n1164);
xor (n1163,n1160,n1161);
and (n1164,n1165,n219);
xor (n1165,n1147,n1148);
and (n1166,n171,n26);
or (n1167,n1168,n1171);
and (n1168,n1169,n1170);
xor (n1169,n1157,n1158);
and (n1170,n165,n26);
and (n1171,n1172,n1173);
xor (n1172,n1169,n1170);
and (n1173,n1174,n1175);
xor (n1174,n1163,n1164);
and (n1175,n23,n26);
and (n1176,n165,n24);
and (n1177,n1178,n1179);
xor (n1178,n1172,n1173);
not (n1179,n22);
and (n1180,n23,n31);
endmodule
